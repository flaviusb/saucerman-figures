time,BARK_RESENS,PKA_RESENS,HYD,REASSOC,b1_AR_tot,b1_AR_d,b1_AR_p,Gs_agtp_tot,Gs_agdp,Gs_bg,cAMP_tot,PLB,Inhib1,Inhib1_DEPHOSPH,PLB_p,Inhib1p_tot,frac_PLB_p,frac_PLB,LCCa,LCCa_DEPHOSPH,LCCb,LCCb_DEPHOSPH,LCCa_p,LCCb_p,frac_LCCa_p,frac_LCCb_p,E_Na,E_K,E_Ca,Na_i,K_i,Ca_i,am,bm,ah,aj,bh,bj,m,h,j,I_Na,V_m,a_lcc,b_lcc,f_lcc,y_lcc_inf,tau_y_lcc,gamma,v_gamma,v_omega,v,w,x,y,z,i_bar_Ca,i_bar_K,f_avail,I_Ca,I_CaK,I_Ca_tot,r_toss,s_toss,tau_r_to,tau_s_to,tau_ss_to,r_to,s_to,ss_to,I_to,r_ss_inf,tau_r_ss,s_ss_inf,r_ss,s_ss,I_ss,a_Ki,b_Ki,Ki_ss,I_Ki,Kp,I_Kp,s4,s5,I_NCX,f_NaK,I_NaK,I_PCa,I_CaB,I_NaB,I_Na_tot,I_K_tot,I_Ca_tot,t_rel,ryr_on,ryr_off,g_rel,I_rel,Ca_jsr,trel,Km_up,I_up,I_leak,I_tr,B_jsr,Ca_nsr,SR_content,b_trpn,b_cmdn,b_indo,B_myo,I_app,V_clamp,I_pace
0.001 2.90118e-11 2.5388e-06 0.020175 0.0201691 0.01205 1.31872e-08 0.001154 0.0252187 0.000644604 0.0258587 0.8453 101.895 0.2474 0.699601 4.105 0.0526 0.0387264 0.961274 0.019897 0.00422319 0.019159 0.00406791 0.005103 0.005841 0.20412 0.23364 57.9406 -87.8925 124.761 16 145 0.00015794 0.267094 192.917 0.310688 0.0673859 0.00409497 0.000561604 0.00138259 0.989185 0.990114 -2.97382e-06 -85.6679 0.0929843 31195 300.011 0.983521 0.319147 0.819315 0.81931 9.99958 2.9809e-06 1.19243e-05 0.130395 0.960074 0.920046 -0.0132933 4.89107e-06 0.500034 -1.81349e-20 6.67248e-24 -1.81282e-20 0.00139513 0.997818 8.59296e-05 0.152554 2.85172 0.00139518 0.999986 0.613135 0.0010384 0.00187967 0.000859296 0.455648 0.06315 0.430012 0.00422877 1.02 0.887304 0.534786 0.285531 1.71633e-07 3.05458e-09 2399.65 3484.98 -0.0821782 0.482121 0.277787 0.276061 -0.589201 -0.169458 0.417364 -0.264775 -0.148784 0.903 1 8.24217e-197 272.41 4.31077e-194 1.92011 0.901 0.000299995 1.02001 0.601723 0.498071 0.381411 1.92039 122.313 79.7879 18.475 58.8514 0.00420341 0 -40 10
0.002 5.80234e-11 2.5388e-06 0.0203099 0.0203008 0.01205 2.63743e-08 0.001154 0.0253874 0.000644612 0.0260274 0.8453 101.895 0.2474 0.699601 4.105 0.0526 0.0387264 0.961274 0.019897 0.00422319 0.019159 0.00406791 0.005103 0.005841 0.20412 0.23364 57.9406 -87.8925 124.766 15.9999 145 0.000157881 0.267054 192.952 0.310777 0.0673969 0.00409434 0.000561464 0.00138213 0.988594 0.99022 -2.96945e-06 -85.6699 0.092966 31199.8 300.011 0.983525 0.319147 0.819007 0.819002 9.99958 2.97973e-06 1.19185e-05 0.130435 0.960147 0.920091 -0.0132936 4.88667e-06 0.500034 -1.81148e-20 6.65892e-24 -1.81081e-20 0.00139489 0.997819 8.59127e-05 0.152522 2.85153 0.0013949 0.999972 0.61327 0.00103728 0.00187936 0.000859127 0.455696 0.0210061 0.430024 0.00140545 1.02 0.88714 0.534832 0.285304 1.71576e-07 3.05089e-09 2399.57 3483.84 -0.0820954 0.482105 0.277777 0.275981 -0.589221 -0.16946 0.417582 -0.267808 -0.149048 0.904 1 4.99913e-197 272.49 2.6157e-194 1.92034 0.902 0.000299995 1.01941 0.601835 0.713458 0.381452 1.92075 122.331 79.8021 18.4759 58.8584 0.00420277 0 -40 10
0.003 8.7035e-11 2.5388e-06 0.0204447 0.0204326 0.01205 3.95614e-08 0.001154 0.0255558 0.000644622 0.0261958 0.845301 101.895 0.2474 0.699601 4.105 0.0526 0.0387264 0.961274 0.019897 0.00422319 0.019159 0.00406791 0.005103 0.005841 0.20412 0.23364 57.9407 -87.8925 124.771 15.9999 145 0.000157821 0.26705 192.955 0.310786 0.067398 0.00409428 0.000561451 0.00138209 0.988163 0.99032 -2.96818e-06 -85.67 0.0929643 31200.2 300.011 0.983526 0.319147 0.818699 0.818694 9.99958 2.9796e-06 1.19183e-05 0.130439 0.96022 0.920137 -0.0132936 4.88627e-06 0.500034 -1.81145e-20 6.65825e-24 -1.81078e-20 0.00139487 0.997819 8.59112e-05 0.152519 2.85151 0.00139487 0.999958 0.613405 0.00103718 0.00187933 0.000859112 0.4557 0.0078478 0.430037 0.000525043 1.02 0.887125 0.534836 0.285283 1.71571e-07 3.05055e-09 2399.55 3482.54 -0.0819988 0.482103 0.277776 0.275903 -0.589235 -0.169461 0.417868 -0.268707 -0.149335 0.905 1 3.03212e-197 272.576 1.58725e-194 1.92064 0.903 0.000299995 1.01881 0.601944 0.806082 0.381503 1.9211 122.349 79.8162 18.4767 58.8654 0.00420213 0 -40 10
0.004 1.16046e-10 2.5388e-06 0.0205793 0.0205643 0.0120499 5.27484e-08 0.001154 0.0257242 0.000644636 0.0263642 0.845301 101.895 0.2474 0.699601 4.105 0.0526 0.0387264 0.961274 0.019897 0.00422319 0.019159 0.00406791 0.00510301 0.00584101 0.20412 0.23364 57.9407 -87.8926 124.776 15.9999 145 0.000157762 0.267057 192.949 0.310771 0.0673962 0.00409438 0.000561473 0.00138216 0.987848 0.990413 -2.96798e-06 -85.6697 0.0929673 31199.4 300.011 0.983525 0.319147 0.818392 0.818387 9.99958 2.97976e-06 1.19189e-05 0.130439 0.960293 0.920182 -0.0132936 4.88698e-06 0.500034 -1.81206e-20 6.66149e-24 -1.81139e-20 0.00139491 0.997819 8.59139e-05 0.152524 2.85154 0.0013949 0.999944 0.613539 0.00103736 0.00187938 0.000859139 0.455692 0.00374245 0.430049 0.000250428 1.02 0.887152 0.534829 0.28532 1.7158e-07 3.05115e-09 2399.55 3481.21 -0.0818986 0.482106 0.277777 0.275824 -0.589248 -0.16946 0.418173 -0.268947 -0.149627 0.906 1 1.83908e-197 272.664 9.63184e-195 1.92095 0.904 0.000299995 1.01821 0.60205 0.845394 0.381558 1.92144 122.367 79.8303 18.4776 58.8723 0.0042015 0 -40 10
0.005 1.45058e-10 2.5388e-06 0.0207139 0.0206961 0.0120499 6.59354e-08 0.001154 0.0258924 0.000644652 0.0265324 0.845302 101.895 0.2474 0.699601 4.105 0.0526 0.0387265 0.961274 0.019897 0.00422319 0.019159 0.00406791 0.00510301 0.00584101 0.20412 0.23364 57.9408 -87.8926 124.781 15.9998 145 0.000157703 0.267065 192.942 0.310752 0.0673938 0.00409451 0.000561503 0.00138226 0.987618 0.9905 -2.96817e-06 -85.6693 0.0929712 31198.4 300.011 0.983524 0.319147 0.818086 0.818081 9.99958 2.97998e-06 1.19198e-05 0.130439 0.960366 0.920227 -0.0132935 4.88794e-06 0.500034 -1.81281e-20 6.66561e-24 -1.81215e-20 0.00139496 0.997819 8.59175e-05 0.152531 2.85158 0.00139496 0.99993 0.613674 0.0010376 0.00187944 0.000859175 0.455682 0.00246159 0.430061 0.000164754 1.02 0.887187 0.534819 0.285369 1.71592e-07 3.05195e-09 2399.55 3479.87 -0.0817979 0.482109 0.277779 0.275746 -0.589261 -0.16946 0.41848 -0.268986 -0.14992 0.907 1 1.11546e-197 272.753 5.84489e-195 1.92128 0.905 0.000299995 1.01762 0.602155 0.861565 0.381614 1.92177 122.385 79.8443 18.4784 58.8792 0.00420086 0 -40 10
0.006 1.74069e-10 2.5388e-06 0.0208483 0.0208278 0.0120499 7.91223e-08 0.001154 0.0260604 0.000644672 0.0267005 0.845302 101.895 0.2474 0.699601 4.105 0.0526 0.0387265 0.961274 0.019897 0.0042232 0.019159 0.00406791 0.00510301 0.00584101 0.20412 0.23364 57.9408 -87.8926 124.786 15.9998 145 0.000157645 0.267074 192.935 0.310733 0.0673915 0.00409465 0.000561533 0.00138236 0.987449 0.990581 -2.96851e-06 -85.6689 0.092975 31197.4 300.011 0.983523 0.319147 0.817782 0.817777 9.99958 2.9802e-06 1.19207e-05 0.130439 0.960438 0.920272 -0.0132934 4.88887e-06 0.500035 -1.81356e-20 6.66965e-24 -1.81289e-20 0.00139501 0.997818 8.5921e-05 0.152538 2.85163 0.00139501 0.999916 0.613809 0.00103783 0.00187951 0.00085921 0.455672 0.00206078 0.430073 0.000137956 1.02 0.887222 0.534809 0.285417 1.71604e-07 3.05273e-09 2399.55 3478.54 -0.0816976 0.482113 0.277781 0.275668 -0.589274 -0.169459 0.418787 -0.268968 -0.150211 0.908 1 6.76558e-198 272.841 3.54686e-195 1.92161 0.906 0.000299995 1.01702 0.602259 0.867697 0.381671 1.9221 122.403 79.8583 18.4793 58.8861 0.00420023 0 -40 10
0.007 2.0308e-10 2.5388e-06 0.0209827 0.0209595 0.0120499 9.23092e-08 0.001154 0.0262284 0.000644693 0.0268685 0.845303 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961274 0.019897 0.0042232 0.019159 0.00406791 0.00510301 0.00584101 0.20412 0.23364 57.9409 -87.8926 124.791 15.9998 145 0.000157586 0.267081 192.928 0.310716 0.0673894 0.00409477 0.000561559 0.00138244 0.987326 0.990657 -2.96891e-06 -85.6685 0.0929785 31196.6 300.011 0.983522 0.319147 0.817478 0.817473 9.99958 2.98039e-06 1.19214e-05 0.130439 0.96051 0.920316 -0.0132934 4.88971e-06 0.500035 -1.81425e-20 6.67337e-24 -1.81358e-20 0.00139505 0.997818 8.59242e-05 0.152544 2.85166 0.00139505 0.999902 0.613943 0.00103804 0.00187957 0.000859242 0.455663 0.00193596 0.430085 0.000129632 1.02 0.887253 0.5348 0.285461 1.71615e-07 3.05343e-09 2399.54 3477.22 -0.081598 0.482116 0.277782 0.27559 -0.589287 -0.169459 0.41909 -0.268936 -0.150501 0.909 1 4.10353e-198 272.928 2.15234e-195 1.92194 0.907 0.000299995 1.01643 0.602364 0.869468 0.381729 1.92244 122.421 79.8723 18.4801 58.893 0.0041996 0 -40 10
0.008 2.32091e-10 2.5388e-06 0.0211169 0.0210912 0.0120499 1.05496e-07 0.001154 0.0263962 0.000644718 0.0270363 0.845304 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961274 0.019897 0.0042232 0.019159 0.00406792 0.00510301 0.00584101 0.20412 0.23364 57.9409 -87.8926 124.796 15.9997 145 0.000157528 0.267088 192.923 0.310702 0.0673876 0.00409487 0.000561582 0.00138252 0.987236 0.990728 -2.96933e-06 -85.6682 0.0929815 31195.8 300.011 0.983522 0.319147 0.817175 0.81717 9.99958 2.98056e-06 1.19221e-05 0.130439 0.960582 0.920361 -0.0132933 4.89044e-06 0.500035 -1.81488e-20 6.67673e-24 -1.81422e-20 0.00139509 0.997818 8.5927e-05 0.152549 2.85169 0.00139509 0.999889 0.614078 0.00103823 0.00187962 0.00085927 0.455656 0.00189702 0.430098 0.000127047 1.02 0.88728 0.534793 0.285499 1.71624e-07 3.05405e-09 2399.54 3475.91 -0.081499 0.482118 0.277783 0.275512 -0.5893 -0.169459 0.419391 -0.268903 -0.150789 0.91 1 2.48892e-198 273.015 1.3061e-195 1.92227 0.908 0.000299995 1.01584 0.602468 0.869351 0.381787 1.92277 122.438 79.8862 18.481 58.8999 0.00419898 0 -40 10
0.009 2.61102e-10 2.5388e-06 0.0212511 0.0212229 0.0120499 1.18683e-07 0.001154 0.0265638 0.000644745 0.027204 0.845305 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961274 0.019897 0.0042232 0.019159 0.00406792 0.00510301 0.00584101 0.204121 0.233641 57.941 -87.8926 124.801 15.9997 145 0.00015747 0.267094 192.918 0.310689 0.067386 0.00409496 0.000561602 0.00138258 0.98717 0.990794 -2.96974e-06 -85.6679 0.0929841 31195.1 300.011 0.983521 0.319147 0.816874 0.816869 9.99958 2.98071e-06 1.19227e-05 0.130439 0.960654 0.920405 -0.0132933 4.89108e-06 0.500035 -1.81546e-20 6.67975e-24 -1.8148e-20 0.00139513 0.997818 8.59294e-05 0.152554 2.85172 0.00139513 0.999875 0.614213 0.00103839 0.00187966 0.000859294 0.455649 0.00188468 0.43011 0.000126234 1.02 0.887304 0.534786 0.285531 1.71632e-07 3.05458e-09 2399.53 3474.6 -0.0814008 0.48212 0.277784 0.275435 -0.589313 -0.169458 0.419689 -0.268872 -0.151076 0.911 1 1.50961e-198 273.102 7.92579e-196 1.9226 0.909 0.000299995 1.01525 0.602571 0.86842 0.381844 1.9231 122.456 79.9 18.4818 58.9067 0.00419835 0 -40 10
0.01 2.90113e-10 2.5388e-06 0.0213851 0.0213546 0.0120499 1.3187e-07 0.001154 0.0267314 0.000644774 0.0273715 0.845306 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961274 0.019897 0.0042232 0.019159 0.00406792 0.00510301 0.00584101 0.204121 0.233641 57.941 -87.8926 124.806 15.9997 145 0.000157412 0.267098 192.913 0.310678 0.0673847 0.00409504 0.000561619 0.00138264 0.987122 0.990856 -2.97013e-06 -85.6677 0.0929863 31194.5 300.011 0.983521 0.319147 0.816573 0.816568 9.99958 2.98084e-06 1.19232e-05 0.130439 0.960726 0.920449 -0.0132932 4.89163e-06 0.500035 -1.81599e-20 6.68246e-24 -1.81532e-20 0.00139516 0.997818 8.59314e-05 0.152558 2.85174 0.00139516 0.999862 0.614347 0.00103853 0.0018797 0.000859314 0.455643 0.00188129 0.430122 0.000126025 1.02 0.887324 0.53478 0.28556 1.71639e-07 3.05504e-09 2399.53 3473.3 -0.0813031 0.482122 0.277785 0.275358 -0.589326 -0.169458 0.419985 -0.268846 -0.151362 0.912 1 9.15622e-199 273.188 4.80958e-196 1.92294 0.91 0.000299995 1.01467 0.602675 0.867128 0.381902 1.92343 122.474 79.9139 18.4827 58.9136 0.00419773 0 -40 10
0.011 3.19124e-10 2.5388e-06 0.021519 0.0214863 0.0120499 1.45056e-07 0.001154 0.0268988 0.000644806 0.027539 0.845308 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961273 0.019897 0.0042232 0.019159 0.00406792 0.00510302 0.00584102 0.204121 0.233641 57.9411 -87.8926 124.811 15.9996 145 0.000157354 0.267103 192.91 0.310668 0.0673835 0.00409511 0.000561634 0.00138268 0.987086 0.990914 -2.9705e-06 -85.6675 0.0929882 31194 300.011 0.98352 0.319147 0.816273 0.816268 9.99958 2.98095e-06 1.19237e-05 0.130439 0.960797 0.920493 -0.0132932 4.8921e-06 0.500035 -1.81648e-20 6.6849e-24 -1.81581e-20 0.00139518 0.997818 8.59332e-05 0.152561 2.85176 0.00139518 0.999848 0.614482 0.00103865 0.00187973 0.000859332 0.455638 0.00188047 0.430134 0.000125987 1.02 0.887342 0.534775 0.285584 1.71645e-07 3.05543e-09 2399.52 3472.01 -0.0812061 0.482124 0.277786 0.275281 -0.589339 -0.169458 0.420278 -0.268823 -0.151646 0.913 1 5.55353e-199 273.274 2.91858e-196 1.92327 0.911 0.000299995 1.01408 0.602778 0.865685 0.381959 1.92376 122.491 79.9276 18.4835 58.9203 0.00419711 0 -40 10
0.012 3.48135e-10 2.5388e-06 0.0216528 0.021618 0.0120498 1.58243e-07 0.001154 0.027066 0.000644839 0.0277063 0.845309 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961273 0.019897 0.0042232 0.019159 0.00406792 0.00510302 0.00584102 0.204121 0.233641 57.9411 -87.8926 124.816 15.9996 145 0.000157296 0.267106 192.907 0.31066 0.0673825 0.00409516 0.000561647 0.00138272 0.98706 0.990968 -2.97084e-06 -85.6673 0.0929899 31193.6 300.011 0.98352 0.319147 0.815975 0.81597 9.99958 2.98104e-06 1.19241e-05 0.130439 0.960868 0.920536 -0.0132932 4.8925e-06 0.500035 -1.81692e-20 6.6871e-24 -1.81625e-20 0.0013952 0.997818 8.59347e-05 0.152564 2.85178 0.0013952 0.999835 0.614616 0.00103876 0.00187976 0.000859347 0.455634 0.00188 0.430146 0.000125969 1.02 0.887357 0.534771 0.285605 1.7165e-07 3.05577e-09 2399.51 3470.72 -0.0811096 0.482125 0.277786 0.275204 -0.589352 -0.169458 0.420569 -0.268803 -0.151929 0.914 1 3.36839e-199 273.359 1.77107e-196 1.9236 0.912 0.000299995 1.0135 0.602882 0.864193 0.382016 1.92409 122.509 79.9414 18.4844 58.9271 0.00419649 0 -40 10
0.013 3.77145e-10 2.5388e-06 0.0217865 0.0217496 0.0120498 1.7143e-07 0.001154 0.0272332 0.000644875 0.0278734 0.845311 101.895 0.2474 0.699601 4.10501 0.0526 0.0387265 0.961273 0.019897 0.0042232 0.019159 0.00406792 0.00510302 0.00584102 0.204121 0.233641 57.9412 -87.8926 124.82 15.9996 145 0.000157239 0.267109 192.904 0.310654 0.0673817 0.00409521 0.000561657 0.00138276 0.987041 0.991018 -2.97116e-06 -85.6671 0.0929913 31193.3 300.011 0.983519 0.319147 0.815677 0.815672 9.99958 2.98112e-06 1.19244e-05 0.130439 0.960939 0.92058 -0.0132932 4.89285e-06 0.500035 -1.81733e-20 6.6891e-24 -1.81666e-20 0.00139522 0.997818 8.5936e-05 0.152566 2.8518 0.00139522 0.999822 0.61475 0.00103885 0.00187979 0.00085936 0.45563 0.00187983 0.430158 0.000125968 1.02 0.88737 0.534767 0.285623 1.71654e-07 3.05606e-09 2399.5 3469.44 -0.0810136 0.482127 0.277787 0.275128 -0.589365 -0.169458 0.420859 -0.268786 -0.15221 0.915 1 2.04303e-199 273.445 1.07472e-196 1.92393 0.913 0.000299995 1.01292 0.602985 0.862671 0.382073 1.92442 122.527 79.9551 18.4852 58.9339 0.00419588 0 -40 10
0.014 4.06156e-10 2.5388e-06 0.0219201 0.0218812 0.0120498 1.84616e-07 0.001154 0.0274001 0.000644913 0.0280405 0.845313 101.895 0.2474 0.699602 4.10501 0.0526 0.0387265 0.961273 0.019897 0.00422321 0.019159 0.00406792 0.00510302 0.00584102 0.204121 0.233641 57.9412 -87.8926 124.825 15.9996 145 0.000157182 0.267112 192.902 0.310648 0.067381 0.00409525 0.000561666 0.00138279 0.987027 0.991065 -2.97144e-06 -85.667 0.0929924 31192.9 300.011 0.983519 0.319147 0.81538 0.815375 9.99958 2.98119e-06 1.19246e-05 0.130439 0.96101 0.920623 -0.0132931 4.89314e-06 0.500035 -1.81771e-20 6.6909e-24 -1.81704e-20 0.00139524 0.997818 8.59371e-05 0.152568 2.85181 0.00139524 0.999809 0.614885 0.00103892 0.00187981 0.000859371 0.455627 0.0018798 0.43017 0.000125977 1.02 0.887381 0.534764 0.285638 1.71658e-07 3.0563e-09 2399.49 3468.17 -0.0809181 0.482128 0.277787 0.275052 -0.589379 -0.169458 0.421146 -0.268771 -0.152491 0.916 1 1.23916e-199 273.529 6.52167e-197 1.92426 0.914 0.000299995 1.01234 0.603088 0.861141 0.38213 1.92475 122.544 79.9687 18.486 58.9406 0.00419526 0 -40 10
0.015 4.35166e-10 2.5388e-06 0.0220536 0.0220128 0.0120498 1.97803e-07 0.001154 0.027567 0.000644953 0.0282074 0.845314 101.895 0.2474 0.699602 4.10501 0.0526001 0.0387265 0.961273 0.019897 0.00422321 0.019159 0.00406792 0.00510302 0.00584102 0.204121 0.233641 57.9413 -87.8926 124.83 15.9995 145 0.000157125 0.267114 192.9 0.310643 0.0673804 0.00409529 0.000561674 0.00138281 0.987017 0.991109 -2.9717e-06 -85.6669 0.0929934 31192.7 300.012 0.983519 0.319147 0.815084 0.81508 9.99958 2.98125e-06 1.19249e-05 0.130439 0.96108 0.920666 -0.0132931 4.89339e-06 0.500035 -1.81806e-20 6.69255e-24 -1.81739e-20 0.00139525 0.997818 8.5938e-05 0.15257 2.85182 0.00139525 0.999796 0.615019 0.00103899 0.00187982 0.00085938 0.455625 0.00187982 0.430183 0.000125988 1.02 0.88739 0.534762 0.285651 1.71661e-07 3.0565e-09 2399.48 3466.9 -0.0808232 0.482128 0.277787 0.274976 -0.589392 -0.169458 0.421432 -0.268759 -0.15277 0.917 1 7.51588e-200 273.614 3.95749e-197 1.92459 0.915 0.000299995 1.01177 0.60319 0.859611 0.382187 1.92508 122.562 79.9823 18.4869 58.9473 0.00419465 0 -40 10
0.016 4.64177e-10 2.5388e-06 0.022187 0.0221444 0.0120498 2.10989e-07 0.001154 0.0277337 0.000644995 0.0283741 0.845316 101.895 0.2474 0.699602 4.10501 0.0526001 0.0387265 0.961273 0.019897 0.00422321 0.019159 0.00406792 0.00510302 0.00584102 0.204121 0.233641 57.9414 -87.8926 124.835 15.9995 145 0.000157068 0.267116 192.899 0.310639 0.0673799 0.00409532 0.00056168 0.00138283 0.987009 0.99115 -2.97193e-06 -85.6668 0.0929943 31192.5 300.012 0.983519 0.319147 0.81479 0.814785 9.99958 2.98129e-06 1.19251e-05 0.130439 0.96115 0.920709 -0.0132931 4.89359e-06 0.500035 -1.8184e-20 6.69406e-24 -1.81773e-20 0.00139526 0.997818 8.59388e-05 0.152572 2.85183 0.00139526 0.999783 0.615153 0.00103904 0.00187984 0.000859388 0.455622 0.00187984 0.430195 0.000125994 1.02 0.887398 0.53476 0.285661 1.71664e-07 3.05668e-09 2399.47 3465.64 -0.0807286 0.482129 0.277787 0.2749 -0.589405 -0.169458 0.421716 -0.268748 -0.153048 0.918 1 4.55861e-200 273.698 2.40149e-197 1.92491 0.916 0.000299995 1.01119 0.603293 0.858089 0.382244 1.9254 122.579 79.9959 18.4877 58.954 0.00419404 0 -40 10
0.017 4.93187e-10 2.5388e-06 0.0223203 0.022276 0.0120498 2.24176e-07 0.001154 0.0279003 0.000645038 0.0285408 0.845319 101.895 0.2474 0.699602 4.10501 0.0526001 0.0387266 0.961273 0.019897 0.00422321 0.019159 0.00406793 0.00510303 0.00584103 0.204121 0.233641 57.9414 -87.8926 124.84 15.9995 145 0.000157011 0.267117 192.897 0.310635 0.0673795 0.00409534 0.000561685 0.00138285 0.987003 0.991188 -2.97214e-06 -85.6667 0.0929949 31192.3 300.012 0.983519 0.319147 0.814496 0.814491 9.99958 2.98133e-06 1.19252e-05 0.130439 0.96122 0.920751 -0.0132931 4.89377e-06 0.500035 -1.81871e-20 6.69544e-24 -1.81804e-20 0.00139527 0.997818 8.59394e-05 0.152573 2.85184 0.00139527 0.99977 0.615287 0.00103909 0.00187985 0.000859394 0.455621 0.00187985 0.430207 0.000126004 1.02 0.887404 0.534758 0.28567 1.71666e-07 3.05682e-09 2399.46 3464.39 -0.0806345 0.48213 0.277787 0.274825 -0.589418 -0.169458 0.421998 -0.26874 -0.153325 0.919 1 2.76494e-200 273.782 1.45727e-197 1.92524 0.917 0.000299995 1.01062 0.603395 0.856564 0.382301 1.92573 122.597 80.0094 18.4885 58.9607 0.00419343 0 -40 10
0.018 5.22197e-10 2.5388e-06 0.0224534 0.0224075 0.0120498 2.37362e-07 0.001154 0.0280668 0.000645083 0.0287073 0.845321 101.895 0.2474 0.699603 4.10502 0.0526001 0.0387266 0.961273 0.019897 0.00422321 0.019159 0.00406793 0.00510303 0.00584103 0.204121 0.233641 57.9415 -87.8926 124.845 15.9994 145 0.000156955 0.267119 192.896 0.310633 0.0673792 0.00409536 0.00056169 0.00138286 0.986999 0.991224 -2.97232e-06 -85.6667 0.0929955 31192.2 300.012 0.983518 0.319147 0.814203 0.814198 9.99958 2.98136e-06 1.19253e-05 0.130439 0.96129 0.920794 -0.0132931 4.89391e-06 0.500035 -1.819e-20 6.69672e-24 -1.81833e-20 0.00139528 0.997818 8.59399e-05 0.152574 2.85184 0.00139528 0.999757 0.615421 0.00103913 0.00187986 0.000859399 0.455619 0.00187985 0.430219 0.000126014 1.02 0.887409 0.534756 0.285678 1.71667e-07 3.05694e-09 2399.44 3463.14 -0.0805408 0.48213 0.277787 0.27475 -0.589432 -0.169458 0.422279 -0.268732 -0.153601 0.92 1 1.67702e-200 273.865 8.84299e-198 1.92557 0.918 0.000299995 1.01005 0.603498 0.855043 0.382358 1.92606 122.614 80.0229 18.4893 58.9673 0.00419283 0 -40 10
0.019 5.51207e-10 2.5388e-06 0.0225865 0.022539 0.0120497 2.50549e-07 0.001154 0.0282331 0.00064513 0.0288736 0.845323 101.895 0.2474 0.699603 4.10502 0.0526002 0.0387266 0.961273 0.019897 0.00422321 0.019159 0.00406793 0.00510303 0.00584103 0.204121 0.233641 57.9415 -87.8926 124.849 15.9994 145 0.000156899 0.26712 192.895 0.310631 0.0673789 0.00409538 0.000561693 0.00138287 0.986996 0.991257 -2.97248e-06 -85.6666 0.0929959 31192 300.012 0.983518 0.319147 0.813911 0.813906 9.99958 2.98139e-06 1.19254e-05 0.130439 0.961359 0.920836 -0.0132931 4.89402e-06 0.500035 -1.81927e-20 6.6979e-24 -1.8186e-20 0.00139528 0.997818 8.59403e-05 0.152575 2.85185 0.00139528 0.999744 0.615555 0.00103916 0.00187987 0.000859403 0.455618 0.00187986 0.430231 0.000126021 1.02 0.887414 0.534755 0.285684 1.71669e-07 3.05703e-09 2399.43 3461.89 -0.0804476 0.482131 0.277787 0.274675 -0.589445 -0.169458 0.422559 -0.268726 -0.153875 0.921 1 1.01716e-200 273.949 5.36608e-198 1.9259 0.919 0.000299995 1.00948 0.6036 0.853528 0.382414 1.92638 122.632 80.0364 18.4902 58.974 0.00419222 0 -40 10
0.02 5.80217e-10 2.5388e-06 0.0227194 0.0226704 0.0120497 2.63735e-07 0.001154 0.0283993 0.000645178 0.0290399 0.845326 101.895 0.2474 0.699604 4.10502 0.0526002 0.0387266 0.961273 0.019897 0.00422321 0.019159 0.00406793 0.00510303 0.00584103 0.204121 0.233641 57.9416 -87.8926 124.854 15.9994 145 0.000156842 0.26712 192.895 0.310629 0.0673787 0.00409539 0.000561696 0.00138288 0.986994 0.991288 -2.97263e-06 -85.6666 0.0929963 31192 300.012 0.983518 0.319147 0.81362 0.813615 9.99958 2.98141e-06 1.19255e-05 0.130439 0.961429 0.920878 -0.0132931 4.89412e-06 0.500035 -1.81954e-20 6.69899e-24 -1.81887e-20 0.00139529 0.997818 8.59406e-05 0.152575 2.85185 0.00139529 0.999732 0.615689 0.00103919 0.00187987 0.000859406 0.455617 0.00187987 0.430243 0.000126028 1.02 0.887417 0.534754 0.285688 1.7167e-07 3.05711e-09 2399.42 3460.65 -0.0803547 0.482131 0.277787 0.2746 -0.589458 -0.169458 0.422837 -0.268721 -0.154149 0.922 1 6.16941e-201 274.032 3.25623e-198 1.92622 0.92 0.000299995 1.00892 0.603702 0.852019 0.382471 1.92671 122.649 80.0498 18.491 58.9806 0.00419162 0 -40 10
0.021 6.09227e-10 2.5388e-06 0.0228523 0.0228019 0.0120497 2.76921e-07 0.001154 0.0285654 0.000645228 0.029206 0.845328 101.895 0.2474 0.699604 4.10502 0.0526003 0.0387266 0.961273 0.019897 0.00422322 0.019159 0.00406793 0.00510303 0.00584103 0.204121 0.233641 57.9416 -87.8926 124.859 15.9993 145 0.000156787 0.267121 192.894 0.310628 0.0673785 0.0040954 0.000561698 0.00138289 0.986992 0.991318 -2.97275e-06 -85.6666 0.0929965 31191.9 300.012 0.983518 0.319147 0.81333 0.813326 9.99958 2.98142e-06 1.19256e-05 0.130439 0.961498 0.92092 -0.0132931 4.89419e-06 0.500035 -1.81979e-20 6.70002e-24 -1.81912e-20 0.00139529 0.997818 8.59409e-05 0.152576 2.85185 0.00139529 0.999719 0.615823 0.00103921 0.00187988 0.000859409 0.455617 0.00187987 0.430255 0.000126033 1.02 0.88742 0.534753 0.285692 1.71671e-07 3.05717e-09 2399.4 3459.41 -0.0802622 0.482131 0.277787 0.274525 -0.589472 -0.169458 0.423114 -0.268717 -0.154422 0.923 1 3.74194e-201 274.114 1.97593e-198 1.92655 0.921 0.000299995 1.00835 0.603803 0.850514 0.382527 1.92703 122.666 80.0631 18.4918 58.9872 0.00419102 0 -40 10
0.022 6.38237e-10 2.5388e-06 0.022985 0.0229333 0.0120497 2.90108e-07 0.001154 0.0287313 0.000645279 0.029372 0.845331 101.895 0.2474 0.699605 4.10502 0.0526003 0.0387266 0.961273 0.019897 0.00422322 0.019159 0.00406793 0.00510303 0.00584103 0.204121 0.233641 57.9417 -87.8926 124.864 15.9993 145 0.000156731 0.267121 192.894 0.310627 0.0673784 0.0040954 0.000561699 0.00138289 0.986991 0.991345 -2.97286e-06 -85.6666 0.0929967 31191.8 300.012 0.983518 0.319147 0.813041 0.813037 9.99958 2.98144e-06 1.19256e-05 0.130439 0.961567 0.920961 -0.0132931 4.89424e-06 0.500035 -1.82003e-20 6.70098e-24 -1.81936e-20 0.00139529 0.997818 8.59411e-05 0.152576 2.85185 0.00139529 0.999707 0.615957 0.00103923 0.00187988 0.000859411 0.455616 0.00187988 0.430267 0.000126039 1.02 0.887422 0.534753 0.285695 1.71671e-07 3.05721e-09 2399.39 3458.18 -0.0801701 0.482131 0.277787 0.274451 -0.589485 -0.169458 0.42339 -0.268714 -0.154694 0.924 1 2.2696e-201 274.197 1.19903e-198 1.92687 0.922 0.000299995 1.00779 0.603905 0.849014 0.382584 1.92736 122.684 80.0765 18.4926 58.9937 0.00419043 0 -40 10
0.023 6.67246e-10 2.5388e-06 0.0231177 0.0230646 0.0120497 3.03294e-07 0.001154 0.0288971 0.000645332 0.0295378 0.845334 101.895 0.2474 0.699606 4.10502 0.0526004 0.0387266 0.961273 0.019897 0.00422322 0.019159 0.00406793 0.00510304 0.00584104 0.204121 0.233641 57.9417 -87.8926 124.868 15.9993 145 0.000156675 0.267122 192.894 0.310626 0.0673783 0.00409541 0.0005617 0.0013829 0.98699 0.99137 -2.97296e-06 -85.6665 0.0929969 31191.8 300.012 0.983518 0.319147 0.812753 0.812748 9.99958 2.98144e-06 1.19257e-05 0.130439 0.961635 0.921003 -0.0132931 4.89428e-06 0.500035 -1.82026e-20 6.70188e-24 -1.81959e-20 0.0013953 0.997818 8.59412e-05 0.152576 2.85186 0.0013953 0.999695 0.616091 0.00103924 0.00187988 0.000859412 0.455616 0.00187988 0.430279 0.000126043 1.02 0.887423 0.534752 0.285697 1.71672e-07 3.05724e-09 2399.37 3456.96 -0.0800783 0.482131 0.277787 0.274377 -0.589498 -0.169458 0.423665 -0.268711 -0.154964 0.925 1 1.37658e-201 274.279 7.27587e-199 1.9272 0.923 0.000299995 1.00723 0.604006 0.847519 0.38264 1.92768 122.701 80.0897 18.4934 59.0003 0.00418983 0 -40 10
0.024 6.96256e-10 2.5388e-06 0.0232502 0.023196 0.0120497 3.1648e-07 0.001154 0.0290628 0.000645385 0.0297035 0.845337 101.895 0.2474 0.699606 4.10502 0.0526004 0.0387266 0.961273 0.019897 0.00422322 0.019159 0.00406793 0.00510304 0.00584104 0.204122 0.233642 57.9418 -87.8926 124.873 15.9992 145 0.00015662 0.267122 192.893 0.310626 0.0673783 0.00409541 0.000561701 0.0013829 0.986989 0.991394 -2.97304e-06 -85.6665 0.0929969 31191.8 300.012 0.983518 0.319147 0.812466 0.812461 9.99958 2.98145e-06 1.19257e-05 0.130439 0.961704 0.921044 -0.0132931 4.89431e-06 0.500036 -1.82048e-20 6.70274e-24 -1.81981e-20 0.0013953 0.997818 8.59412e-05 0.152576 2.85186 0.0013953 0.999682 0.616225 0.00103926 0.00187988 0.000859412 0.455615 0.00187988 0.430291 0.000126048 1.02 0.887424 0.534752 0.285698 1.71672e-07 3.05726e-09 2399.36 3455.74 -0.0799869 0.482132 0.277786 0.274303 -0.589511 -0.169458 0.423938 -0.268709 -0.155234 0.926 1 8.34939e-202 274.361 4.4151e-199 1.92752 0.924 0.000299995 1.00667 0.604108 0.846029 0.382696 1.928 122.718 80.103 18.4942 59.0068 0.00418924 0 -40 10
0.025 7.25265e-10 2.5388e-06 0.0233826 0.0233273 0.0120497 3.29666e-07 0.001154 0.0292283 0.00064544 0.0298691 0.84534 101.895 0.2474 0.699607 4.10502 0.0526005 0.0387266 0.961273 0.019897 0.00422322 0.019159 0.00406793 0.00510304 0.00584104 0.204122 0.233642 57.9418 -87.8926 124.878 15.9992 145.001 0.000156565 0.267122 192.893 0.310625 0.0673783 0.00409541 0.000561701 0.0013829 0.986989 0.991416 -2.97311e-06 -85.6665 0.092997 31191.8 300.012 0.983518 0.319147 0.81218 0.812175 9.99958 2.98145e-06 1.19257e-05 0.130439 0.961772 0.921085 -0.0132931 4.89433e-06 0.500036 -1.82069e-20 6.70355e-24 -1.82002e-20 0.0013953 0.997818 8.59413e-05 0.152576 2.85186 0.0013953 0.99967 0.616359 0.00103926 0.00187988 0.000859413 0.455615 0.00187988 0.430303 0.000126052 1.02 0.887425 0.534752 0.285699 1.71672e-07 3.05727e-09 2399.35 3454.52 -0.0798958 0.482132 0.277786 0.27423 -0.589524 -0.169458 0.42421 -0.268708 -0.155503 0.927 1 5.06416e-202 274.442 2.67914e-199 1.92784 0.925 0.000299995 1.00611 0.604209 0.844543 0.382752 1.92833 122.735 80.1162 18.495 59.0133 0.00418864 0 -40 10
0.026 7.54275e-10 2.5388e-06 0.0235149 0.0234585 0.0120497 3.42852e-07 0.001154 0.0293937 0.000645496 0.0300346 0.845344 101.895 0.247399 0.699608 4.10502 0.0526005 0.0387266 0.961273 0.019897 0.00422322 0.019159 0.00406794 0.00510304 0.00584104 0.204122 0.233642 57.9419 -87.8926 124.883 15.9992 145.001 0.00015651 0.267122 192.893 0.310626 0.0673783 0.00409541 0.000561701 0.0013829 0.986988 0.991437 -2.97317e-06 -85.6665 0.092997 31191.8 300.012 0.983518 0.319147 0.811895 0.81189 9.99958 2.98145e-06 1.19257e-05 0.130439 0.96184 0.921126 -0.0132931 4.89433e-06 0.500036 -1.8209e-20 6.70433e-24 -1.82023e-20 0.0013953 0.997818 8.59413e-05 0.152576 2.85186 0.0013953 0.999658 0.616493 0.00103927 0.00187988 0.000859413 0.455615 0.00187988 0.430315 0.000126055 1.02 0.887425 0.534752 0.285699 1.71672e-07 3.05728e-09 2399.33 3453.31 -0.0798051 0.482132 0.277786 0.274156 -0.589537 -0.169458 0.424482 -0.268707 -0.155771 0.928 1 3.07157e-202 274.524 1.62573e-199 1.92817 0.926 0.000299995 1.00556 0.60431 0.843063 0.382808 1.92865 122.753 80.1293 18.4958 59.0198 0.00418805 0 -40 10
0.027 7.83284e-10 2.5388e-06 0.0236472 0.0235897 0.0120496 3.56038e-07 0.001154 0.0295589 0.000645553 0.0301999 0.845347 101.895 0.247399 0.699609 4.10503 0.0526006 0.0387267 0.961273 0.019897 0.00422322 0.019159 0.00406794 0.00510304 0.00584104 0.204122 0.233642 57.9419 -87.8926 124.887 15.9991 145.001 0.000156455 0.267122 192.894 0.310626 0.0673783 0.00409541 0.000561701 0.0013829 0.986988 0.991456 -2.97322e-06 -85.6665 0.0929969 31191.8 300.012 0.983518 0.319147 0.811611 0.811606 9.99958 2.98145e-06 1.19257e-05 0.130439 0.961908 0.921167 -0.0132931 4.89433e-06 0.500036 -1.82111e-20 6.70507e-24 -1.82043e-20 0.0013953 0.997818 8.59412e-05 0.152576 2.85186 0.0013953 0.999646 0.616626 0.00103927 0.00187988 0.000859412 0.455616 0.00187988 0.430328 0.000126059 1.02 0.887425 0.534752 0.285699 1.71672e-07 3.05727e-09 2399.32 3452.1 -0.0797147 0.482131 0.277786 0.274083 -0.589551 -0.169458 0.424752 -0.268707 -0.156038 0.929 1 1.863e-202 274.605 9.86514e-200 1.92849 0.927 0.000299995 1.005 0.60441 0.841587 0.382864 1.92897 122.77 80.1425 18.4966 59.0263 0.00418747 0 -40 10
0.028 8.12293e-10 2.5388e-06 0.0237793 0.0237209 0.0120496 3.69224e-07 0.001154 0.0297241 0.000645611 0.0303651 0.845351 101.895 0.247399 0.69961 4.10503 0.0526007 0.0387267 0.961273 0.019897 0.00422323 0.019159 0.00406794 0.00510305 0.00584105 0.204122 0.233642 57.942 -87.8926 124.892 15.9991 145.001 0.0001564 0.267122 192.894 0.310626 0.0673783 0.00409541 0.0005617 0.0013829 0.986988 0.991475 -2.97326e-06 -85.6665 0.0929968 31191.8 300.012 0.983518 0.319147 0.811327 0.811322 9.99958 2.98144e-06 1.19257e-05 0.130439 0.961976 0.921208 -0.0132931 4.89432e-06 0.500036 -1.8213e-20 6.70578e-24 -1.82063e-20 0.0013953 0.997818 8.59411e-05 0.152576 2.85185 0.0013953 0.999634 0.61676 0.00103927 0.00187988 0.000859411 0.455616 0.00187988 0.43034 0.000126062 1.02 0.887425 0.534752 0.285699 1.71671e-07 3.05726e-09 2399.3 3450.89 -0.0796246 0.482131 0.277785 0.27401 -0.589564 -0.169458 0.425021 -0.268707 -0.156304 0.93 1 1.12997e-202 274.686 5.98627e-200 1.92881 0.928 0.000299995 1.00445 0.604511 0.840115 0.38292 1.92929 122.787 80.1556 18.4974 59.0327 0.00418688 0 -40 10
0.029 8.41302e-10 2.5388e-06 0.0239113 0.023852 0.0120496 3.8241e-07 0.001154 0.0298891 0.00064567 0.0305302 0.845354 101.895 0.247399 0.699611 4.10503 0.0526008 0.0387267 0.961273 0.019897 0.00422323 0.019159 0.00406794 0.00510305 0.00584105 0.204122 0.233642 57.9421 -87.8926 124.897 15.9991 145.001 0.000156346 0.267121 192.894 0.310627 0.0673784 0.0040954 0.000561699 0.00138289 0.986988 0.991492 -2.9733e-06 -85.6666 0.0929967 31191.8 300.012 0.983518 0.319147 0.811045 0.81104 9.99958 2.98143e-06 1.19256e-05 0.130439 0.962043 0.921248 -0.0132931 4.8943e-06 0.500036 -1.8215e-20 6.70647e-24 -1.82083e-20 0.00139529 0.997818 8.5941e-05 0.152576 2.85185 0.00139529 0.999622 0.616893 0.00103928 0.00187988 0.00085941 0.455616 0.00187988 0.430352 0.000126065 1.02 0.887424 0.534752 0.285698 1.71671e-07 3.05724e-09 2399.29 3449.69 -0.0795348 0.482131 0.277785 0.273938 -0.589577 -0.169458 0.425289 -0.268707 -0.156569 0.931 1 6.8536e-203 274.766 3.63253e-200 1.92913 0.929 0.000299995 1.0039 0.604612 0.838649 0.382975 1.92961 122.804 80.1686 18.4982 59.0391 0.0041863 0 -40 10
0.03 8.70311e-10 2.5388e-06 0.0240432 0.0239831 0.0120496 3.95596e-07 0.001154 0.0300539 0.000645729 0.0306951 0.845358 101.895 0.247399 0.699612 4.10503 0.0526009 0.0387267 0.961273 0.019897 0.00422323 0.019159 0.00406794 0.00510305 0.00584105 0.204122 0.233642 57.9421 -87.8927 124.901 15.999 145.001 0.000156292 0.267121 192.894 0.310627 0.0673785 0.0040954 0.000561698 0.00138289 0.986988 0.991507 -2.97332e-06 -85.6666 0.0929966 31191.9 300.012 0.983518 0.319147 0.810763 0.810759 9.99958 2.98143e-06 1.19256e-05 0.130439 0.96211 0.921288 -0.0132931 4.89428e-06 0.500036 -1.82169e-20 6.70713e-24 -1.82101e-20 0.00139529 0.997818 8.59409e-05 0.152576 2.85185 0.00139529 0.99961 0.617027 0.00103927 0.00187988 0.000859409 0.455616 0.00187988 0.430364 0.000126068 1.02 0.887423 0.534753 0.285696 1.71671e-07 3.05722e-09 2399.27 3448.5 -0.0794454 0.482131 0.277785 0.273865 -0.58959 -0.169458 0.425556 -0.268707 -0.156834 0.932 1 4.15692e-203 274.846 2.20425e-200 1.92945 0.93 0.000299995 1.00335 0.604712 0.837187 0.383031 1.92993 122.821 80.1816 18.499 59.0455 0.00418572 0 -40 10
0.031 8.9932e-10 2.5388e-06 0.0241749 0.0241141 0.0120496 4.08782e-07 0.001154 0.0302187 0.00064579 0.0308599 0.845362 101.895 0.247399 0.699613 4.10503 0.052601 0.0387267 0.961273 0.0198969 0.00422323 0.0191589 0.00406794 0.00510305 0.00584105 0.204122 0.233642 57.9422 -87.8927 124.906 15.999 145.001 0.000156238 0.267121 192.894 0.310628 0.0673786 0.00409539 0.000561697 0.00138289 0.986987 0.991522 -2.97335e-06 -85.6666 0.0929964 31191.9 300.012 0.983518 0.319147 0.810483 0.810478 9.99958 2.98142e-06 1.19256e-05 0.130439 0.962177 0.921328 -0.0132931 4.89425e-06 0.500036 -1.82187e-20 6.70777e-24 -1.8212e-20 0.00139529 0.997818 8.59408e-05 0.152575 2.85185 0.00139529 0.999599 0.61716 0.00103927 0.00187987 0.000859408 0.455617 0.00187988 0.430376 0.00012607 1.02 0.887422 0.534753 0.285695 1.7167e-07 3.0572e-09 2399.26 3447.3 -0.0793563 0.482131 0.277784 0.273793 -0.589603 -0.169458 0.425823 -0.268708 -0.157097 0.933 1 2.5213e-203 274.927 1.33756e-200 1.92977 0.931 0.000299995 1.00281 0.604812 0.83573 0.383086 1.93025 122.838 80.1946 18.4998 59.0519 0.00418514 0 -40 10
0.032 9.28329e-10 2.5388e-06 0.0243066 0.024245 0.0120496 4.21968e-07 0.001154 0.0303833 0.000645851 0.0310245 0.845366 101.895 0.247399 0.699614 4.10503 0.0526011 0.0387267 0.961273 0.0198969 0.00422323 0.0191589 0.00406794 0.00510305 0.00584105 0.204122 0.233642 57.9422 -87.8927 124.91 15.999 145.001 0.000156184 0.26712 192.895 0.310629 0.0673787 0.00409539 0.000561696 0.00138288 0.986987 0.991536 -2.97336e-06 -85.6666 0.0929963 31192 300.012 0.983518 0.319147 0.810203 0.810198 9.99958 2.98141e-06 1.19255e-05 0.130439 0.962244 0.921368 -0.0132931 4.89422e-06 0.500036 -1.82205e-20 6.7084e-24 -1.82138e-20 0.00139529 0.997818 8.59406e-05 0.152575 2.85185 0.00139529 0.999587 0.617294 0.00103927 0.00187987 0.000859406 0.455617 0.00187987 0.430388 0.000126073 1.02 0.887421 0.534753 0.285693 1.7167e-07 3.05717e-09 2399.24 3446.12 -0.0792675 0.482131 0.277784 0.273721 -0.589616 -0.169458 0.426088 -0.268709 -0.15736 0.934 1 1.52924e-203 275.006 8.11639e-201 1.93009 0.932 0.000299995 1.00226 0.604912 0.834277 0.383142 1.93057 122.855 80.2075 18.5006 59.0583 0.00418456 0 -40 10
0.033 9.57338e-10 2.5388e-06 0.0244382 0.024376 0.0120496 4.35153e-07 0.001154 0.0305478 0.000645913 0.0311891 0.84537 101.895 0.247399 0.699616 4.10503 0.0526012 0.0387267 0.961273 0.0198969 0.00422323 0.0191589 0.00406795 0.00510306 0.00584106 0.204122 0.233642 57.9423 -87.8927 124.915 15.9989 145.001 0.00015613 0.26712 192.895 0.31063 0.0673788 0.00409538 0.000561694 0.00138288 0.986987 0.991549 -2.97337e-06 -85.6666 0.0929961 31192 300.012 0.983518 0.319147 0.809925 0.80992 9.99958 2.9814e-06 1.19255e-05 0.130439 0.96231 0.921408 -0.0132931 4.89418e-06 0.500036 -1.82223e-20 6.70901e-24 -1.82156e-20 0.00139529 0.997818 8.59404e-05 0.152575 2.85185 0.00139529 0.999576 0.617427 0.00103927 0.00187987 0.000859404 0.455618 0.00187987 0.4304 0.000126075 1.02 0.887419 0.534754 0.285691 1.71669e-07 3.05713e-09 2399.23 3444.93 -0.079179 0.482131 0.277784 0.273649 -0.589629 -0.169459 0.426352 -0.26871 -0.157621 0.935 1 9.27534e-204 275.086 4.92508e-201 1.93041 0.933 0.000299995 1.00172 0.605012 0.83283 0.383197 1.93089 122.873 80.2204 18.5014 59.0646 0.00418398 0 -40 10
0.034 9.86346e-10 2.5388e-06 0.0245697 0.0245068 0.0120496 4.48339e-07 0.001154 0.0307121 0.000645975 0.0313535 0.845375 101.895 0.247399 0.699617 4.10503 0.0526013 0.0387267 0.961273 0.0198969 0.00422324 0.0191589 0.00406795 0.00510306 0.00584106 0.204122 0.233642 57.9423 -87.8927 124.92 15.9989 145.001 0.000156076 0.267119 192.895 0.310631 0.0673789 0.00409537 0.000561693 0.00138287 0.986987 0.991561 -2.97338e-06 -85.6666 0.0929959 31192.1 300.012 0.983518 0.319147 0.809647 0.809642 9.99958 2.98139e-06 1.19254e-05 0.130439 0.962377 0.921447 -0.0132931 4.89414e-06 0.500036 -1.82241e-20 6.70961e-24 -1.82174e-20 0.00139528 0.997818 8.59403e-05 0.152574 2.85185 0.00139528 0.999564 0.617561 0.00103926 0.00187986 0.000859403 0.455618 0.00187987 0.430412 0.000126078 1.02 0.887418 0.534754 0.285689 1.71669e-07 3.0571e-09 2399.21 3443.75 -0.0790908 0.482131 0.277783 0.273578 -0.589641 -0.169459 0.426615 -0.268712 -0.157882 0.936 1 5.62578e-204 275.165 2.98857e-201 1.93073 0.934 0.000299995 1.00118 0.605111 0.831386 0.383252 1.93121 122.89 80.2332 18.5022 59.071 0.00418341 0 -40 10
0.035 1.01535e-09 2.5388e-06 0.024701 0.0246376 0.0120495 4.61525e-07 0.001154 0.0308763 0.000646039 0.0315177 0.845379 101.895 0.247399 0.699619 4.10504 0.0526014 0.0387267 0.961273 0.0198969 0.00422324 0.0191589 0.00406795 0.00510306 0.00584106 0.204122 0.233642 57.9424 -87.8927 124.924 15.9989 145.001 0.000156023 0.267119 192.896 0.310632 0.067379 0.00409537 0.000561691 0.00138287 0.986987 0.991572 -2.97338e-06 -85.6667 0.0929957 31192.1 300.012 0.983518 0.319147 0.80937 0.809365 9.99958 2.98138e-06 1.19254e-05 0.130439 0.962443 0.921487 -0.0132931 4.8941e-06 0.500036 -1.82259e-20 6.7102e-24 -1.82192e-20 0.00139528 0.997818 8.59401e-05 0.152574 2.85184 0.00139528 0.999553 0.617694 0.00103926 0.00187986 0.000859401 0.455619 0.00187986 0.430424 0.00012608 1.02 0.887416 0.534754 0.285687 1.71668e-07 3.05706e-09 2399.19 3442.58 -0.0790029 0.48213 0.277783 0.273507 -0.589654 -0.169459 0.426878 -0.268713 -0.158142 0.937 1 3.41221e-204 275.244 1.81348e-201 1.93105 0.935 0.000299995 1.00064 0.605211 0.829948 0.383307 1.93152 122.906 80.246 18.5029 59.0773 0.00418284 0 -40 10
0.036 1.04436e-09 2.5388e-06 0.0248323 0.0247684 0.0120495 4.74711e-07 0.001154 0.0310404 0.000646102 0.0316819 0.845384 101.895 0.247398 0.69962 4.10504 0.0526015 0.0387268 0.961273 0.0198969 0.00422324 0.0191589 0.00406795 0.00510306 0.00584106 0.204122 0.233642 57.9424 -87.8927 124.929 15.9988 145.001 0.00015597 0.267118 192.896 0.310633 0.0673792 0.00409536 0.000561689 0.00138286 0.986988 0.991583 -2.97338e-06 -85.6667 0.0929954 31192.2 300.012 0.983518 0.319147 0.809094 0.809089 9.99958 2.98136e-06 1.19253e-05 0.130439 0.962509 0.921526 -0.0132931 4.89406e-06 0.500036 -1.82276e-20 6.71077e-24 -1.82209e-20 0.00139528 0.997818 8.59399e-05 0.152574 2.85184 0.00139528 0.999541 0.617827 0.00103925 0.00187986 0.000859399 0.455619 0.00187986 0.430436 0.000126082 1.02 0.887415 0.534755 0.285685 1.71667e-07 3.05702e-09 2399.18 3441.41 -0.0789153 0.48213 0.277782 0.273435 -0.589667 -0.169459 0.427139 -0.268714 -0.158401 0.938 1 2.06961e-204 275.323 1.10043e-201 1.93137 0.936 0.000299995 1.0001 0.60531 0.828514 0.383362 1.93184 122.923 80.2588 18.5037 59.0836 0.00418227 0 -40 10
0.037 1.07337e-09 2.5388e-06 0.0249635 0.0248991 0.0120495 4.87896e-07 0.001154 0.0312043 0.000646166 0.0318459 0.845388 101.895 0.247398 0.699622 4.10504 0.0526017 0.0387268 0.961273 0.0198969 0.00422324 0.0191589 0.00406795 0.00510306 0.00584106 0.204123 0.233643 57.9425 -87.8927 124.933 15.9988 145.001 0.000155917 0.267118 192.897 0.310634 0.0673793 0.00409535 0.000561688 0.00138286 0.986988 0.991593 -2.97337e-06 -85.6667 0.0929952 31192.2 300.012 0.983518 0.319147 0.808819 0.808814 9.99958 2.98135e-06 1.19253e-05 0.130439 0.962575 0.921565 -0.0132931 4.89401e-06 0.500036 -1.82293e-20 6.71134e-24 -1.82226e-20 0.00139527 0.997818 8.59397e-05 0.152573 2.85184 0.00139528 0.99953 0.61796 0.00103924 0.00187985 0.000859397 0.45562 0.00187986 0.430448 0.000126084 1.02 0.887413 0.534755 0.285683 1.71667e-07 3.05698e-09 2399.16 3440.24 -0.0788281 0.48213 0.277782 0.273365 -0.58968 -0.169459 0.4274 -0.268716 -0.158659 0.939 1 1.25528e-204 275.402 6.67743e-202 1.93169 0.937 0.000299995 0.999568 0.605409 0.827085 0.383417 1.93216 122.94 80.2715 18.5045 59.0898 0.0041817 0 -40 10
0.038 1.10238e-09 2.5388e-06 0.0250945 0.0250297 0.0120495 5.01082e-07 0.001154 0.0313681 0.000646231 0.0320098 0.845393 101.895 0.247398 0.699624 4.10504 0.0526018 0.0387268 0.961273 0.0198969 0.00422324 0.0191589 0.00406795 0.00510307 0.00584107 0.204123 0.233643 57.9425 -87.8927 124.938 15.9988 145.001 0.000155864 0.267117 192.897 0.310635 0.0673795 0.00409534 0.000561686 0.00138285 0.986988 0.991602 -2.97337e-06 -85.6667 0.092995 31192.3 300.012 0.983519 0.319147 0.808545 0.80854 9.99958 2.98134e-06 1.19252e-05 0.130439 0.96264 0.921604 -0.0132931 4.89396e-06 0.500037 -1.8231e-20 6.7119e-24 -1.82243e-20 0.00139527 0.997818 8.59394e-05 0.152573 2.85184 0.00139527 0.999519 0.618094 0.00103924 0.00187985 0.000859394 0.455621 0.00187985 0.43046 0.000126086 1.02 0.887411 0.534756 0.28568 1.71666e-07 3.05694e-09 2399.15 3439.07 -0.0787411 0.48213 0.277782 0.273294 -0.589693 -0.169459 0.42766 -0.268718 -0.158917 0.94 1 7.61366e-205 275.48 4.05188e-202 1.932 0.938 0.000299995 0.999034 0.605508 0.82566 0.383472 1.93247 122.957 80.2842 18.5053 59.0961 0.00418113 0 -40 10
0.039 1.13139e-09 2.5388e-06 0.0252255 0.0251603 0.0120495 5.14267e-07 0.001154 0.0315318 0.000646296 0.0321735 0.845398 101.895 0.247398 0.699626 4.10504 0.052602 0.0387268 0.961273 0.0198969 0.00422324 0.0191589 0.00406795 0.00510307 0.00584107 0.204123 0.233643 57.9426 -87.8927 124.942 15.9987 145.001 0.000155811 0.267117 192.898 0.310636 0.0673796 0.00409533 0.000561684 0.00138285 0.986988 0.99161 -2.97336e-06 -85.6668 0.0929948 31192.4 300.013 0.983519 0.319147 0.808272 0.808267 9.99958 2.98132e-06 1.19252e-05 0.13044 0.962705 0.921642 -0.0132931 4.89391e-06 0.500037 -1.82327e-20 6.71245e-24 -1.8226e-20 0.00139527 0.997818 8.59392e-05 0.152572 2.85183 0.00139527 0.999508 0.618227 0.00103923 0.00187985 0.000859392 0.455621 0.00187985 0.430472 0.000126088 1.02 0.887409 0.534756 0.285678 1.71665e-07 3.0569e-09 2399.13 3437.91 -0.0786544 0.48213 0.277781 0.273224 -0.589705 -0.169459 0.427918 -0.268719 -0.159173 0.941 1 4.61792e-205 275.559 2.45869e-202 1.93232 0.939 0.000299994 0.998503 0.605607 0.82424 0.383527 1.93279 122.974 80.2969 18.506 59.1023 0.00418057 0 -40 10
0.04 1.1604e-09 2.5388e-06 0.0253563 0.0252908 0.0120495 5.27453e-07 0.001154 0.0316954 0.000646361 0.0323371 0.845403 101.895 0.247398 0.699628 4.10504 0.0526021 0.0387268 0.961273 0.0198969 0.00422325 0.0191589 0.00406796 0.00510307 0.00584107 0.204123 0.233643 57.9427 -87.8927 124.947 15.9987 145.001 0.000155759 0.267116 192.898 0.310638 0.0673797 0.00409533 0.000561682 0.00138284 0.986988 0.991618 -2.97334e-06 -85.6668 0.0929945 31192.4 300.013 0.983519 0.319147 0.807999 0.807994 9.99958 2.98131e-06 1.19251e-05 0.13044 0.962771 0.921681 -0.0132931 4.89386e-06 0.500037 -1.82344e-20 6.71299e-24 -1.82276e-20 0.00139527 0.997818 8.5939e-05 0.152572 2.85183 0.00139527 0.999497 0.61836 0.00103922 0.00187984 0.00085939 0.455622 0.00187984 0.430484 0.00012609 1.02 0.887408 0.534757 0.285675 1.71664e-07 3.05685e-09 2399.12 3436.76 -0.078568 0.482129 0.277781 0.273153 -0.589718 -0.169459 0.428176 -0.268721 -0.159429 0.942 1 2.80091e-205 275.636 1.49194e-202 1.93264 0.94 0.000299994 0.997973 0.605706 0.822824 0.383582 1.9331 122.991 80.3095 18.5068 59.1085 0.00418 0 -40 10
0.041 1.1894e-09 2.5388e-06 0.025487 0.0254212 0.0120495 5.40638e-07 0.001154 0.0318588 0.000646427 0.0325006 0.845408 101.895 0.247398 0.69963 4.10504 0.0526023 0.0387268 0.961273 0.0198969 0.00422325 0.0191589 0.00406796 0.00510307 0.00584107 0.204123 0.233643 57.9427 -87.8927 124.951 15.9987 145.001 0.000155707 0.267116 192.898 0.310639 0.0673799 0.00409532 0.00056168 0.00138283 0.986988 0.991626 -2.97333e-06 -85.6668 0.0929943 31192.5 300.013 0.983519 0.319147 0.807728 0.807723 9.99958 2.9813e-06 1.19251e-05 0.13044 0.962835 0.921719 -0.0132931 4.89381e-06 0.500037 -1.8236e-20 6.71353e-24 -1.82293e-20 0.00139526 0.997818 8.59388e-05 0.152572 2.85183 0.00139526 0.999486 0.618493 0.00103922 0.00187984 0.000859388 0.455622 0.00187984 0.430496 0.000126092 1.02 0.887406 0.534757 0.285672 1.71664e-07 3.05681e-09 2399.1 3435.61 -0.0784819 0.482129 0.27778 0.273083 -0.589731 -0.169459 0.428433 -0.268723 -0.159684 0.943 1 1.69884e-205 275.714 9.05309e-203 1.93295 0.941 0.000299994 0.997445 0.605805 0.821413 0.383636 1.93342 123.008 80.322 18.5076 59.1147 0.00417944 0 -40 10
0.042 1.21841e-09 2.5388e-06 0.0256177 0.0255516 0.0120494 5.53823e-07 0.001154 0.0320221 0.000646493 0.032664 0.845414 101.895 0.247398 0.699632 4.10505 0.0526024 0.0387268 0.961273 0.0198969 0.00422325 0.0191589 0.00406796 0.00510308 0.00584108 0.204123 0.233643 57.9428 -87.8927 124.956 15.9986 145.001 0.000155654 0.267115 192.899 0.31064 0.06738 0.00409531 0.000561678 0.00138283 0.986988 0.991633 -2.97331e-06 -85.6668 0.092994 31192.5 300.013 0.983519 0.319147 0.807457 0.807452 9.99958 2.98128e-06 1.1925e-05 0.13044 0.9629 0.921758 -0.0132931 4.89376e-06 0.500037 -1.82377e-20 6.71406e-24 -1.8231e-20 0.00139526 0.997818 8.59385e-05 0.152571 2.85183 0.00139526 0.999475 0.618626 0.00103921 0.00187983 0.000859385 0.455623 0.00187984 0.430508 0.000126094 1.02 0.887404 0.534758 0.28567 1.71663e-07 3.05676e-09 2399.09 3434.46 -0.0783961 0.482129 0.27778 0.273014 -0.589743 -0.169459 0.428689 -0.268725 -0.159938 0.944 1 1.0304e-205 275.792 5.49341e-203 1.93327 0.942 0.000299994 0.996918 0.605903 0.820006 0.383691 1.93373 123.025 80.3346 18.5083 59.1209 0.00417888 0 -40 10
0.043 1.24742e-09 2.5388e-06 0.0257482 0.0256819 0.0120494 5.67009e-07 0.001154 0.0321853 0.000646559 0.0328272 0.845419 101.895 0.247397 0.699634 4.10505 0.0526026 0.0387269 0.961273 0.0198969 0.00422325 0.0191589 0.00406796 0.00510308 0.00584108 0.204123 0.233643 57.9428 -87.8927 124.96 15.9986 145.001 0.000155602 0.267115 192.899 0.310641 0.0673802 0.0040953 0.000561676 0.00138282 0.986988 0.99164 -2.97329e-06 -85.6669 0.0929938 31192.6 300.013 0.983519 0.319147 0.807187 0.807183 9.99958 2.98127e-06 1.1925e-05 0.13044 0.962965 0.921796 -0.0132931 4.89371e-06 0.500037 -1.82393e-20 6.71459e-24 -1.82326e-20 0.00139526 0.997818 8.59383e-05 0.152571 2.85182 0.00139526 0.999464 0.618759 0.0010392 0.00187983 0.000859383 0.455624 0.00187983 0.430519 0.000126096 1.02 0.887402 0.534759 0.285667 1.71662e-07 3.05672e-09 2399.07 3433.31 -0.0783106 0.482129 0.27778 0.272944 -0.589756 -0.169459 0.428945 -0.268727 -0.160191 0.945 1 6.24967e-206 275.869 3.3334e-203 1.93358 0.943 0.000299994 0.996394 0.606001 0.818604 0.383745 1.93405 123.041 80.3471 18.5091 59.127 0.00417833 0 -40 10
0.044 1.27643e-09 2.5388e-06 0.0258786 0.0258122 0.0120494 5.80194e-07 0.001154 0.0323483 0.000646626 0.0329903 0.845425 101.895 0.247397 0.699636 4.10505 0.0526028 0.0387269 0.961273 0.0198969 0.00422326 0.0191589 0.00406796 0.00510308 0.00584108 0.204123 0.233643 57.9429 -87.8927 124.965 15.9986 145.001 0.000155551 0.267114 192.9 0.310642 0.0673803 0.00409529 0.000561675 0.00138282 0.986988 0.991646 -2.97327e-06 -85.6669 0.0929935 31192.7 300.013 0.983519 0.319147 0.806919 0.806914 9.99958 2.98125e-06 1.19249e-05 0.13044 0.963029 0.921833 -0.0132931 4.89366e-06 0.500037 -1.82409e-20 6.71512e-24 -1.82342e-20 0.00139525 0.997818 8.59381e-05 0.15257 2.85182 0.00139525 0.999453 0.618892 0.00103919 0.00187982 0.000859381 0.455624 0.00187983 0.430531 0.000126098 1.02 0.8874 0.534759 0.285664 1.71661e-07 3.05667e-09 2399.06 3432.17 -0.0782253 0.482129 0.277779 0.272875 -0.589768 -0.16946 0.429199 -0.268729 -0.160443 0.946 1 3.79062e-206 275.946 2.0227e-203 1.93389 0.944 0.000299994 0.995871 0.606099 0.817207 0.383799 1.93436 123.058 80.3595 18.5098 59.1331 0.00417777 0 -40 10
0.045 1.30543e-09 2.5388e-06 0.0260089 0.0259423 0.0120494 5.93379e-07 0.001154 0.0325112 0.000646692 0.0331533 0.84543 101.895 0.247397 0.699639 4.10505 0.052603 0.0387269 0.961273 0.0198969 0.00422326 0.0191589 0.00406797 0.00510308 0.00584108 0.204123 0.233643 57.9429 -87.8927 124.969 15.9985 145.001 0.000155499 0.267114 192.9 0.310644 0.0673805 0.00409528 0.000561673 0.00138281 0.986988 0.991651 -2.97325e-06 -85.6669 0.0929933 31192.7 300.013 0.983519 0.319147 0.806651 0.806646 9.99958 2.98124e-06 1.19248e-05 0.13044 0.963093 0.921871 -0.0132931 4.8936e-06 0.500037 -1.82426e-20 6.71564e-24 -1.82358e-20 0.00139525 0.997818 8.59378e-05 0.15257 2.85182 0.00139525 0.999443 0.619025 0.00103919 0.00187982 0.000859378 0.455625 0.00187982 0.430543 0.0001261 1.02 0.887398 0.53476 0.285662 1.7166e-07 3.05663e-09 2399.04 3431.03 -0.0781404 0.482128 0.277779 0.272806 -0.589781 -0.16946 0.429453 -0.268731 -0.160695 0.947 1 2.29913e-206 276.023 1.22737e-203 1.93421 0.945 0.000299994 0.995349 0.606197 0.815813 0.383854 1.93467 123.075 80.372 18.5106 59.1392 0.00417722 0 -40 10
0.046 1.33444e-09 2.5388e-06 0.0261392 0.0260725 0.0120494 6.06565e-07 0.001154 0.0326739 0.000646759 0.0333161 0.845436 101.895 0.247397 0.699641 4.10505 0.0526032 0.0387269 0.961273 0.0198969 0.00422326 0.0191589 0.00406797 0.00510309 0.00584109 0.204123 0.233643 57.943 -87.8927 124.974 15.9985 145.001 0.000155447 0.267113 192.901 0.310645 0.0673807 0.00409527 0.000561671 0.0013828 0.986988 0.991657 -2.97323e-06 -85.667 0.092993 31192.8 300.013 0.983519 0.319147 0.806384 0.806379 9.99958 2.98122e-06 1.19248e-05 0.13044 0.963157 0.921909 -0.0132931 4.89355e-06 0.500037 -1.82442e-20 6.71616e-24 -1.82374e-20 0.00139525 0.997818 8.59376e-05 0.152569 2.85181 0.00139525 0.999432 0.619157 0.00103918 0.00187982 0.000859376 0.455626 0.00187982 0.430555 0.000126102 1.02 0.887396 0.53476 0.285659 1.7166e-07 3.05658e-09 2399.02 3429.9 -0.0780557 0.482128 0.277778 0.272737 -0.589793 -0.16946 0.429705 -0.268733 -0.160945 0.948 1 1.39449e-206 276.099 7.44765e-204 1.93452 0.946 0.000299994 0.99483 0.606295 0.814425 0.383908 1.93498 123.092 80.3843 18.5113 59.1453 0.00417667 0 -40 10
0.047 1.36345e-09 2.5388e-06 0.0262693 0.0262025 0.0120494 6.1975e-07 0.001154 0.0328366 0.000646825 0.0334788 0.845442 101.895 0.247397 0.699644 4.10505 0.0526034 0.0387269 0.961273 0.0198969 0.00422326 0.0191589 0.00406797 0.00510309 0.00584109 0.204124 0.233644 57.943 -87.8927 124.978 15.9985 145.001 0.000155396 0.267113 192.901 0.310646 0.0673808 0.00409526 0.000561669 0.0013828 0.986988 0.991662 -2.9732e-06 -85.667 0.0929927 31192.9 300.013 0.983519 0.319147 0.806118 0.806113 9.99958 2.98121e-06 1.19247e-05 0.13044 0.963221 0.921946 -0.0132931 4.8935e-06 0.500037 -1.82458e-20 6.71668e-24 -1.82391e-20 0.00139524 0.997818 8.59374e-05 0.152569 2.85181 0.00139524 0.999421 0.61929 0.00103917 0.00187981 0.000859374 0.455626 0.00187981 0.430567 0.000126103 1.02 0.887394 0.534761 0.285656 1.71659e-07 3.05653e-09 2399.01 3428.77 -0.0779713 0.482128 0.277778 0.272668 -0.589806 -0.16946 0.429957 -0.268734 -0.161195 0.949 1 8.45801e-207 276.175 4.5192e-204 1.93483 0.947 0.000299994 0.994312 0.606393 0.81304 0.383962 1.9353 123.108 80.3967 18.5121 59.1514 0.00417612 0 -40 10
0.048 1.39246e-09 2.5388e-06 0.0263993 0.0263324 0.0120494 6.32935e-07 0.001154 0.0329991 0.000646892 0.0336414 0.845448 101.895 0.247396 0.699647 4.10506 0.0526036 0.0387269 0.961273 0.0198969 0.00422326 0.0191589 0.00406797 0.00510309 0.00584109 0.204124 0.233644 57.9431 -87.8927 124.982 15.9984 145.001 0.000155345 0.267112 192.902 0.310647 0.067381 0.00409526 0.000561667 0.00138279 0.986988 0.991667 -2.97318e-06 -85.667 0.0929925 31192.9 300.013 0.983519 0.319147 0.805852 0.805847 9.99958 2.9812e-06 1.19247e-05 0.13044 0.963284 0.921983 -0.0132931 4.89345e-06 0.500037 -1.82474e-20 6.71719e-24 -1.82406e-20 0.00139524 0.997818 8.59371e-05 0.152568 2.85181 0.00139524 0.999411 0.619423 0.00103917 0.00187981 0.000859371 0.455627 0.00187981 0.430579 0.000126105 1.02 0.887392 0.534761 0.285653 1.71658e-07 3.05649e-09 2398.99 3427.64 -0.0778872 0.482128 0.277778 0.2726 -0.589818 -0.16946 0.430208 -0.268736 -0.161444 0.95 1 5.13004e-207 276.252 2.74223e-204 1.93514 0.948 0.000299994 0.993796 0.60649 0.81166 0.384016 1.93561 123.125 80.409 18.5128 59.1575 0.00417557 0 -40 10
0.049 1.42146e-09 2.5388e-06 0.0265292 0.0264623 0.0120494 6.4612e-07 0.001154 0.0331615 0.000646959 0.0338038 0.845454 101.895 0.247396 0.69965 4.10506 0.0526038 0.038727 0.961273 0.0198969 0.00422327 0.0191589 0.00406797 0.0051031 0.0058411 0.204124 0.233644 57.9431 -87.8927 124.987 15.9984 145.001 0.000155294 0.267111 192.902 0.310649 0.0673811 0.00409525 0.000561665 0.00138278 0.986988 0.991671 -2.97315e-06 -85.667 0.0929922 31193 300.013 0.983519 0.319147 0.805588 0.805583 9.99958 2.98118e-06 1.19246e-05 0.13044 0.963347 0.92202 -0.0132931 4.89339e-06 0.500038 -1.8249e-20 6.7177e-24 -1.82422e-20 0.00139524 0.997818 8.59369e-05 0.152568 2.85181 0.00139524 0.999401 0.619556 0.00103916 0.0018798 0.000859369 0.455628 0.00187981 0.430591 0.000126107 1.02 0.88739 0.534762 0.285651 1.71657e-07 3.05644e-09 2398.98 3426.52 -0.0778034 0.482127 0.277777 0.272531 -0.589831 -0.16946 0.430458 -0.268738 -0.161692 0.951 1 3.11153e-207 276.327 1.66397e-204 1.93546 0.949 0.000299994 0.993282 0.606588 0.810285 0.38407 1.93592 123.141 80.4213 18.5136 59.1635 0.00417502 0 -40 10
0.05 1.45047e-09 2.5388e-06 0.026659 0.0265921 0.0120493 6.59305e-07 0.001154 0.0333237 0.000647026 0.0339661 0.845461 101.895 0.247396 0.699652 4.10506 0.0526041 0.038727 0.961273 0.0198969 0.00422327 0.0191589 0.00406797 0.0051031 0.0058411 0.204124 0.233644 57.9432 -87.8927 124.991 15.9984 145.001 0.000155243 0.267111 192.903 0.31065 0.0673813 0.00409524 0.000561663 0.00138278 0.986988 0.991675 -2.97313e-06 -85.6671 0.092992 31193.1 300.013 0.983519 0.319147 0.805324 0.80532 9.99958 2.98117e-06 1.19246e-05 0.13044 0.963411 0.922057 -0.0132931 4.89334e-06 0.500038 -1.82505e-20 6.71821e-24 -1.82438e-20 0.00139523 0.997818 8.59367e-05 0.152568 2.8518 0.00139523 0.99939 0.619688 0.00103915 0.0018798 0.000859367 0.455628 0.0018798 0.430603 0.000126109 1.02 0.887388 0.534762 0.285648 1.71657e-07 3.05639e-09 2398.96 3425.4 -0.0777199 0.482127 0.277777 0.272463 -0.589843 -0.16946 0.430707 -0.26874 -0.16194 0.952 1 1.88724e-207 276.403 1.00969e-204 1.93577 0.95 0.000299994 0.99277 0.606685 0.808914 0.384123 1.93623 123.158 80.4335 18.5143 59.1695 0.00417448 0 -40 10
0.051 1.47948e-09 2.5388e-06 0.0267887 0.0267219 0.0120493 6.7249e-07 0.001154 0.0334858 0.000647093 0.0341283 0.845467 101.895 0.247396 0.699656 4.10506 0.0526043 0.038727 0.961273 0.0198969 0.00422327 0.0191589 0.00406798 0.0051031 0.0058411 0.204124 0.233644 57.9433 -87.8927 124.995 15.9983 145.001 0.000155193 0.26711 192.903 0.310651 0.0673814 0.00409523 0.000561661 0.00138277 0.986989 0.991679 -2.9731e-06 -85.6671 0.0929917 31193.1 300.013 0.983519 0.319147 0.805062 0.805057 9.99958 2.98115e-06 1.19245e-05 0.13044 0.963473 0.922094 -0.0132931 4.89329e-06 0.500038 -1.82521e-20 6.71872e-24 -1.82454e-20 0.00139523 0.997818 8.59364e-05 0.152567 2.8518 0.00139523 0.99938 0.619821 0.00103914 0.00187979 0.000859364 0.455629 0.0018798 0.430615 0.000126111 1.02 0.887386 0.534763 0.285645 1.71656e-07 3.05635e-09 2398.95 3424.29 -0.0776366 0.482127 0.277776 0.272395 -0.589855 -0.16946 0.430956 -0.268742 -0.162186 0.953 1 1.14467e-207 276.478 6.12673e-205 1.93608 0.951 0.000299994 0.992259 0.606782 0.807547 0.384177 1.93654 123.175 80.4457 18.5151 59.1755 0.00417394 0 -40 10
0.052 1.50848e-09 2.5388e-06 0.0269183 0.0268515 0.0120493 6.85675e-07 0.001154 0.0336478 0.00064716 0.0342904 0.845473 101.895 0.247395 0.699659 4.10506 0.0526046 0.038727 0.961273 0.0198969 0.00422327 0.0191589 0.00406798 0.0051031 0.0058411 0.204124 0.233644 57.9433 -87.8927 125 15.9983 145.001 0.000155142 0.26711 192.904 0.310652 0.0673816 0.00409522 0.000561659 0.00138276 0.986989 0.991682 -2.97307e-06 -85.6671 0.0929915 31193.2 300.013 0.983519 0.319147 0.8048 0.804795 9.99958 2.98114e-06 1.19244e-05 0.13044 0.963536 0.922131 -0.0132932 4.89324e-06 0.500038 -1.82537e-20 6.71922e-24 -1.8247e-20 0.00139523 0.997818 8.59362e-05 0.152567 2.8518 0.00139523 0.99937 0.619953 0.00103914 0.00187979 0.000859362 0.45563 0.00187979 0.430627 0.000126113 1.02 0.887384 0.534764 0.285642 1.71655e-07 3.0563e-09 2398.93 3423.18 -0.0775536 0.482127 0.277776 0.272328 -0.589867 -0.16946 0.431204 -0.268744 -0.162432 0.954 1 6.94276e-208 276.554 3.71765e-205 1.93639 0.952 0.000299994 0.99175 0.606879 0.806184 0.384231 1.93685 123.191 80.4578 18.5158 59.1815 0.0041734 0 -40 10
0.053 1.53749e-09 2.5388e-06 0.0270477 0.0269811 0.0120493 6.9886e-07 0.001154 0.0338097 0.000647226 0.0344523 0.84548 101.895 0.247395 0.699662 4.10507 0.0526048 0.038727 0.961273 0.0198969 0.00422328 0.0191589 0.00406798 0.00510311 0.00584111 0.204124 0.233644 57.9434 -87.8927 125.004 15.9983 145.001 0.000155092 0.267109 192.904 0.310654 0.0673817 0.00409521 0.000561657 0.00138276 0.986989 0.991686 -2.97304e-06 -85.6671 0.0929912 31193.3 300.013 0.983519 0.319147 0.804539 0.804534 9.99958 2.98112e-06 1.19244e-05 0.13044 0.963599 0.922167 -0.0132932 4.89318e-06 0.500038 -1.82553e-20 6.71972e-24 -1.82485e-20 0.00139522 0.997818 8.5936e-05 0.152566 2.8518 0.00139522 0.99936 0.620086 0.00103913 0.00187978 0.00085936 0.45563 0.00187979 0.430639 0.000126115 1.02 0.887382 0.534764 0.28564 1.71654e-07 3.05625e-09 2398.91 3422.07 -0.0774709 0.482127 0.277775 0.27226 -0.58988 -0.16946 0.43145 -0.268746 -0.162677 0.955 1 4.211e-208 276.629 2.25584e-205 1.9367 0.953 0.000299994 0.991242 0.606975 0.804826 0.384284 1.93716 123.208 80.47 18.5165 59.1875 0.00417286 0 -40 10
0.054 1.5665e-09 2.5388e-06 0.0271771 0.0271106 0.0120493 7.12045e-07 0.001154 0.0339714 0.000647293 0.0346141 0.845487 101.895 0.247395 0.699665 4.10507 0.0526051 0.0387271 0.961273 0.0198969 0.00422328 0.0191589 0.00406798 0.00510311 0.00584111 0.204124 0.233644 57.9434 -87.8927 125.008 15.9982 145.001 0.000155042 0.267109 192.905 0.310655 0.0673819 0.0040952 0.000561655 0.00138275 0.986989 0.991689 -2.97301e-06 -85.6672 0.092991 31193.3 300.013 0.983519 0.319147 0.804279 0.804274 9.99958 2.98111e-06 1.19243e-05 0.13044 0.963661 0.922204 -0.0132932 4.89313e-06 0.500038 -1.82568e-20 6.72023e-24 -1.82501e-20 0.00139522 0.997818 8.59357e-05 0.152566 2.85179 0.00139522 0.99935 0.620218 0.00103912 0.00187978 0.000859357 0.455631 0.00187978 0.430651 0.000126116 1.02 0.88738 0.534765 0.285637 1.71653e-07 3.05621e-09 2398.9 3420.96 -0.0773885 0.482126 0.277775 0.272193 -0.589892 -0.169461 0.431696 -0.268748 -0.162921 0.956 1 2.5541e-208 276.703 1.36883e-205 1.93701 0.954 0.000299994 0.990737 0.607072 0.803472 0.384338 1.93746 123.224 80.482 18.5173 59.1934 0.00417232 0 -40 10
0.055 1.5955e-09 2.5388e-06 0.0273064 0.02724 0.0120493 7.25229e-07 0.001154 0.034133 0.000647359 0.0347758 0.845494 101.895 0.247395 0.699669 4.10507 0.0526054 0.0387271 0.961273 0.0198969 0.00422328 0.0191589 0.00406799 0.00510311 0.00584111 0.204125 0.233645 57.9435 -87.8927 125.013 15.9982 145.001 0.000154992 0.267108 192.905 0.310656 0.067382 0.00409519 0.000561653 0.00138275 0.986989 0.991692 -2.97298e-06 -85.6672 0.0929907 31193.4 300.014 0.98352 0.319147 0.80402 0.804015 9.99958 2.98109e-06 1.19243e-05 0.13044 0.963723 0.92224 -0.0132932 4.89308e-06 0.500038 -1.82584e-20 6.72073e-24 -1.82517e-20 0.00139522 0.997818 8.59355e-05 0.152565 2.85179 0.00139522 0.99934 0.620351 0.00103912 0.00187978 0.000859355 0.455632 0.00187978 0.430663 0.000126118 1.02 0.887378 0.534765 0.285634 1.71653e-07 3.05616e-09 2398.88 3419.86 -0.0773063 0.482126 0.277775 0.272126 -0.589904 -0.169461 0.431941 -0.26875 -0.163165 0.957 1 1.54914e-208 276.778 8.30591e-206 1.93731 0.955 0.000299994 0.990233 0.607169 0.802123 0.384391 1.93777 123.241 80.4941 18.518 59.1993 0.00417179 0 -40 10
0.056 1.62451e-09 2.5388e-06 0.0274356 0.0273693 0.0120493 7.38414e-07 0.001154 0.0342945 0.000647426 0.0349373 0.845501 101.895 0.247394 0.699672 4.10507 0.0526057 0.0387271 0.961273 0.0198969 0.00422328 0.0191589 0.00406799 0.00510312 0.00584112 0.204125 0.233645 57.9435 -87.8927 125.017 15.9982 145.001 0.000154942 0.267108 192.906 0.310657 0.0673822 0.00409519 0.000561651 0.00138274 0.986989 0.991695 -2.97295e-06 -85.6672 0.0929905 31193.5 300.014 0.98352 0.319147 0.803761 0.803756 9.99958 2.98108e-06 1.19242e-05 0.13044 0.963785 0.922276 -0.0132932 4.89303e-06 0.500038 -1.82599e-20 6.72123e-24 -1.82532e-20 0.00139521 0.997818 8.59353e-05 0.152565 2.85179 0.00139521 0.99933 0.620483 0.00103911 0.00187977 0.000859353 0.455632 0.00187978 0.430674 0.00012612 1.02 0.887376 0.534766 0.285632 1.71652e-07 3.05612e-09 2398.87 3418.77 -0.0772244 0.482126 0.277774 0.27206 -0.589916 -0.169461 0.432186 -0.268752 -0.163408 0.958 1 9.396e-209 276.852 5.03994e-206 1.93762 0.956 0.000299994 0.98973 0.607265 0.800777 0.384444 1.93808 123.257 80.5061 18.5187 59.2052 0.00417125 0 -40 10
0.057 1.65352e-09 2.5388e-06 0.0275646 0.0274986 0.0120492 7.51599e-07 0.001154 0.0344558 0.000647492 0.0350987 0.845508 101.895 0.247394 0.699676 4.10507 0.0526059 0.0387271 0.961273 0.0198969 0.00422329 0.0191589 0.00406799 0.00510312 0.00584112 0.204125 0.233645 57.9436 -87.8928 125.021 15.9981 145.001 0.000154892 0.267107 192.906 0.310659 0.0673823 0.00409518 0.000561649 0.00138273 0.986989 0.991697 -2.97292e-06 -85.6673 0.0929902 31193.5 300.014 0.98352 0.319147 0.803504 0.803499 9.99958 2.98107e-06 1.19242e-05 0.13044 0.963847 0.922312 -0.0132932 4.89298e-06 0.500038 -1.82615e-20 6.72172e-24 -1.82548e-20 0.00139521 0.997818 8.5935e-05 0.152564 2.85179 0.00139521 0.99932 0.620615 0.00103911 0.00187977 0.00085935 0.455633 0.00187977 0.430686 0.000126122 1.02 0.887374 0.534766 0.285629 1.71651e-07 3.05607e-09 2398.85 3417.67 -0.0771428 0.482126 0.277774 0.271993 -0.589928 -0.169461 0.432429 -0.268753 -0.163649 0.959 1 5.69896e-209 276.926 3.05818e-206 1.93793 0.957 0.000299994 0.98923 0.607361 0.799436 0.384497 1.93839 123.273 80.5181 18.5194 59.2111 0.00417072 0 -40 10
0.058 1.68252e-09 2.5388e-06 0.0276936 0.0276278 0.0120492 7.64784e-07 0.001154 0.034617 0.000647558 0.03526 0.845515 101.895 0.247394 0.69968 4.10508 0.0526063 0.0387271 0.961273 0.0198969 0.00422329 0.0191589 0.00406799 0.00510312 0.00584112 0.204125 0.233645 57.9436 -87.8928 125.026 15.9981 145.001 0.000154843 0.267107 192.907 0.31066 0.0673825 0.00409517 0.000561647 0.00138273 0.986989 0.9917 -2.97289e-06 -85.6673 0.09299 31193.6 300.014 0.98352 0.319147 0.803247 0.803242 9.99958 2.98105e-06 1.19241e-05 0.13044 0.963908 0.922347 -0.0132932 4.89293e-06 0.500038 -1.8263e-20 6.72222e-24 -1.82563e-20 0.00139521 0.997818 8.59348e-05 0.152564 2.85178 0.00139521 0.99931 0.620747 0.0010391 0.00187976 0.000859348 0.455634 0.00187977 0.430698 0.000126124 1.02 0.887373 0.534767 0.285626 1.7165e-07 3.05603e-09 2398.84 3416.58 -0.0770615 0.482126 0.277773 0.271927 -0.58994 -0.169461 0.432672 -0.268755 -0.16389 0.96 1 3.4566e-209 277 1.85567e-206 1.93824 0.958 0.000299994 0.988731 0.607457 0.7981 0.384551 1.93869 123.29 80.53 18.5202 59.217 0.00417019 0 -40 10
0.059 1.71153e-09 2.5388e-06 0.0278225 0.0277568 0.0120492 7.77968e-07 0.001154 0.0347781 0.000647623 0.0354211 0.845523 101.895 0.247393 0.699684 4.10508 0.0526066 0.0387272 0.961273 0.0198969 0.00422329 0.0191589 0.00406799 0.00510313 0.00584113 0.204125 0.233645 57.9437 -87.8928 125.03 15.9981 145.001 0.000154793 0.267106 192.907 0.310661 0.0673826 0.00409516 0.000561646 0.00138272 0.986989 0.991702 -2.97286e-06 -85.6673 0.0929897 31193.6 300.014 0.98352 0.319147 0.802991 0.802986 9.99958 2.98104e-06 1.1924e-05 0.13044 0.96397 0.922383 -0.0132932 4.89288e-06 0.500039 -1.82646e-20 6.72272e-24 -1.82578e-20 0.0013952 0.997818 8.59346e-05 0.152564 2.85178 0.0013952 0.9993 0.62088 0.00103909 0.00187976 0.000859346 0.455634 0.00187976 0.43071 0.000126126 1.02 0.887371 0.534767 0.285624 1.7165e-07 3.05598e-09 2398.82 3415.5 -0.0769804 0.482125 0.277773 0.27186 -0.589952 -0.169461 0.432914 -0.268757 -0.164131 0.961 1 2.09653e-209 277.074 1.126e-206 1.93854 0.959 0.000299994 0.988233 0.607553 0.796767 0.384604 1.939 123.306 80.5419 18.5209 59.2228 0.00416966 0 -40 10
0.06 1.74054e-09 2.5388e-06 0.0279512 0.0278858 0.0120492 7.91153e-07 0.001154 0.034939 0.000647689 0.0355821 0.84553 101.895 0.247393 0.699688 4.10508 0.0526069 0.0387272 0.961273 0.0198969 0.0042233 0.0191589 0.004068 0.00510313 0.00584113 0.204125 0.233645 57.9438 -87.8928 125.034 15.998 145.001 0.000154744 0.267105 192.907 0.310662 0.0673828 0.00409515 0.000561644 0.00138272 0.986989 0.991704 -2.97283e-06 -85.6673 0.0929895 31193.7 300.014 0.98352 0.319147 0.802736 0.802731 9.99958 2.98102e-06 1.1924e-05 0.13044 0.964031 0.922418 -0.0132932 4.89283e-06 0.500039 -1.82661e-20 6.72321e-24 -1.82594e-20 0.0013952 0.997818 8.59344e-05 0.152563 2.85178 0.0013952 0.99929 0.621012 0.00103909 0.00187976 0.000859344 0.455635 0.00187976 0.430722 0.000126128 1.02 0.887369 0.534768 0.285621 1.71649e-07 3.05594e-09 2398.8 3414.42 -0.0768996 0.482125 0.277773 0.271795 -0.589964 -0.169461 0.433155 -0.268759 -0.16437 0.962 1 1.27161e-209 277.147 6.83241e-207 1.93885 0.96 0.000299994 0.987738 0.607649 0.795439 0.384656 1.9393 123.323 80.5538 18.5216 59.2287 0.00416914 0 -40 10
0.061 1.76954e-09 2.5388e-06 0.0280799 0.0280148 0.0120492 8.04337e-07 0.001154 0.0350999 0.000647754 0.035743 0.845538 101.895 0.247393 0.699692 4.10508 0.0526072 0.0387272 0.961273 0.0198969 0.0042233 0.0191589 0.004068 0.00510314 0.00584113 0.204125 0.233645 57.9438 -87.8928 125.038 15.998 145.001 0.000154695 0.267105 192.908 0.310663 0.0673829 0.00409514 0.000561642 0.00138271 0.986989 0.991706 -2.9728e-06 -85.6674 0.0929892 31193.8 300.014 0.98352 0.319147 0.802482 0.802477 9.99958 2.98101e-06 1.19239e-05 0.13044 0.964092 0.922453 -0.0132932 4.89278e-06 0.500039 -1.82676e-20 6.72371e-24 -1.82609e-20 0.0013952 0.997818 8.59341e-05 0.152563 2.85178 0.0013952 0.999281 0.621144 0.00103908 0.00187975 0.000859341 0.455635 0.00187975 0.430734 0.00012613 1.02 0.887367 0.534768 0.285619 1.71648e-07 3.0559e-09 2398.79 3413.34 -0.0768191 0.482125 0.277772 0.271729 -0.589976 -0.169461 0.433395 -0.268761 -0.164609 0.963 1 7.71271e-210 277.22 4.14582e-207 1.93916 0.961 0.000299994 0.987244 0.607744 0.794115 0.384709 1.93961 123.339 80.5656 18.5223 59.2345 0.00416861 0 -40 10
0.062 1.79855e-09 2.5388e-06 0.0282085 0.0281436 0.0120492 8.17522e-07 0.001154 0.0352606 0.000647819 0.0359038 0.845546 101.895 0.247392 0.699696 4.10509 0.0526076 0.0387272 0.961273 0.0198969 0.0042233 0.0191589 0.004068 0.00510314 0.00584114 0.204126 0.233646 57.9439 -87.8928 125.043 15.998 145.001 0.000154646 0.267104 192.908 0.310665 0.0673831 0.00409513 0.00056164 0.0013827 0.986989 0.991708 -2.97277e-06 -85.6674 0.092989 31193.8 300.014 0.98352 0.319147 0.802228 0.802224 9.99958 2.981e-06 1.19239e-05 0.13044 0.964153 0.922489 -0.0132932 4.89273e-06 0.500039 -1.82692e-20 6.7242e-24 -1.82624e-20 0.00139519 0.997818 8.59339e-05 0.152562 2.85177 0.00139519 0.999271 0.621276 0.00103908 0.00187975 0.000859339 0.455636 0.00187975 0.430746 0.000126132 1.02 0.887365 0.534769 0.285616 1.71647e-07 3.05585e-09 2398.77 3412.26 -0.0767388 0.482125 0.277772 0.271663 -0.589988 -0.169461 0.433635 -0.268762 -0.164847 0.964 1 4.67799e-210 277.293 2.51562e-207 1.93946 0.962 0.000299994 0.986751 0.60784 0.792795 0.384762 1.93991 123.355 80.5774 18.523 59.2403 0.00416809 0 -40 10
0.063 1.82755e-09 2.5388e-06 0.0283369 0.0282723 0.0120492 8.30706e-07 0.001154 0.0354211 0.000647884 0.0360644 0.845554 101.895 0.247392 0.699701 4.10509 0.0526079 0.0387273 0.961273 0.0198969 0.00422331 0.0191589 0.004068 0.00510314 0.00584114 0.204126 0.233646 57.9439 -87.8928 125.047 15.9979 145.001 0.000154598 0.267104 192.909 0.310666 0.0673832 0.00409513 0.000561638 0.0013827 0.986989 0.991709 -2.97274e-06 -85.6674 0.0929888 31193.9 300.014 0.98352 0.319147 0.801976 0.801971 9.99958 2.98098e-06 1.19238e-05 0.13044 0.964213 0.922524 -0.0132932 4.89268e-06 0.500039 -1.82707e-20 6.72469e-24 -1.8264e-20 0.00139519 0.997818 8.59337e-05 0.152562 2.85177 0.00139519 0.999262 0.621408 0.00103907 0.00187974 0.000859337 0.455637 0.00187975 0.430757 0.000126134 1.02 0.887363 0.534769 0.285614 1.71647e-07 3.05581e-09 2398.76 3411.19 -0.0766588 0.482124 0.277771 0.271598 -0.59 -0.169461 0.433873 -0.268764 -0.165084 0.965 1 2.83735e-210 277.366 1.52644e-207 1.93977 0.963 0.000299994 0.98626 0.607935 0.791479 0.384815 1.94022 123.371 80.5891 18.5237 59.246 0.00416757 0 -40 10
0.064 1.85656e-09 2.5388e-06 0.0284653 0.028401 0.0120492 8.43891e-07 0.001154 0.0355816 0.000647948 0.0362249 0.845562 101.895 0.247392 0.699705 4.10509 0.0526083 0.0387273 0.961273 0.0198969 0.00422331 0.0191589 0.00406801 0.00510315 0.00584115 0.204126 0.233646 57.944 -87.8928 125.051 15.9979 145.001 0.000154549 0.267103 192.909 0.310667 0.0673834 0.00409512 0.000561636 0.00138269 0.98699 0.991711 -2.97271e-06 -85.6674 0.0929885 31194 300.014 0.98352 0.319147 0.801724 0.801719 9.99958 2.98097e-06 1.19238e-05 0.13044 0.964274 0.922558 -0.0132932 4.89263e-06 0.500039 -1.82722e-20 6.72518e-24 -1.82655e-20 0.00139519 0.997818 8.59335e-05 0.152562 2.85177 0.00139519 0.999252 0.62154 0.00103907 0.00187974 0.000859335 0.455637 0.00187974 0.430769 0.000126136 1.02 0.887361 0.53477 0.285611 1.71646e-07 3.05577e-09 2398.74 3410.12 -0.0765791 0.482124 0.277771 0.271533 -0.590011 -0.169461 0.434111 -0.268766 -0.16532 0.966 1 1.72094e-210 277.438 9.26221e-208 1.94007 0.964 0.000299994 0.985771 0.60803 0.790168 0.384867 1.94052 123.388 80.6009 18.5245 59.2518 0.00416705 0 -40 10
0.065 1.88557e-09 2.5388e-06 0.0285935 0.0285295 0.0120491 8.57075e-07 0.001154 0.0357419 0.000648012 0.0363853 0.84557 101.895 0.247391 0.69971 4.10509 0.0526086 0.0387273 0.961273 0.0198968 0.00422331 0.0191589 0.00406801 0.00510315 0.00584115 0.204126 0.233646 57.944 -87.8928 125.055 15.9979 145.001 0.000154501 0.267103 192.91 0.310668 0.0673835 0.00409511 0.000561635 0.00138269 0.98699 0.991713 -2.97268e-06 -85.6675 0.0929883 31194 300.014 0.98352 0.319147 0.801473 0.801469 9.99958 2.98096e-06 1.19237e-05 0.13044 0.964334 0.922593 -0.0132932 4.89258e-06 0.500039 -1.82737e-20 6.72567e-24 -1.8267e-20 0.00139518 0.997818 8.59333e-05 0.152561 2.85177 0.00139518 0.999243 0.621672 0.00103906 0.00187974 0.000859333 0.455638 0.00187974 0.430781 0.000126138 1.02 0.88736 0.53477 0.285609 1.71645e-07 3.05573e-09 2398.73 3409.06 -0.0764996 0.482124 0.277771 0.271468 -0.590023 -0.169462 0.434348 -0.268767 -0.165556 0.967 1 1.0438e-210 277.511 5.62016e-208 1.94037 0.965 0.000299994 0.985284 0.608125 0.78886 0.38492 1.94082 123.404 80.6125 18.5252 59.2575 0.00416653 0 -40 10
0.066 1.91457e-09 2.5388e-06 0.0287216 0.028658 0.0120491 8.7026e-07 0.001154 0.0359021 0.000648076 0.0365455 0.845578 101.895 0.247391 0.699715 4.1051 0.052609 0.0387273 0.961273 0.0198968 0.00422332 0.0191588 0.00406801 0.00510316 0.00584115 0.204126 0.233646 57.9441 -87.8928 125.059 15.9979 145.001 0.000154453 0.267102 192.91 0.310669 0.0673836 0.0040951 0.000561633 0.00138268 0.98699 0.991714 -2.97265e-06 -85.6675 0.0929881 31194.1 300.014 0.98352 0.319147 0.801223 0.801219 9.99958 2.98094e-06 1.19237e-05 0.13044 0.964394 0.922628 -0.0132932 4.89254e-06 0.50004 -1.82752e-20 6.72616e-24 -1.82685e-20 0.00139518 0.997818 8.59331e-05 0.152561 2.85176 0.00139518 0.999234 0.621804 0.00103906 0.00187973 0.000859331 0.455638 0.00187973 0.430793 0.00012614 1.02 0.887358 0.534771 0.285606 1.71644e-07 3.05568e-09 2398.71 3407.99 -0.0764204 0.482124 0.27777 0.271403 -0.590035 -0.169462 0.434585 -0.268769 -0.165791 0.968 1 6.33098e-211 277.583 3.41022e-208 1.94068 0.966 0.000299994 0.984798 0.60822 0.787557 0.384972 1.94113 123.42 80.6242 18.5259 59.2633 0.00416602 0 -40 10
0.067 1.94358e-09 2.5388e-06 0.0288497 0.0287864 0.0120491 8.83444e-07 0.001154 0.0360621 0.00064814 0.0367056 0.845586 101.895 0.247391 0.69972 4.1051 0.0526094 0.0387274 0.961273 0.0198968 0.00422332 0.0191588 0.00406802 0.00510316 0.00584116 0.204126 0.233646 57.9441 -87.8928 125.063 15.9978 145.001 0.000154405 0.267102 192.911 0.31067 0.0673838 0.00409509 0.000561631 0.00138267 0.98699 0.991715 -2.97262e-06 -85.6675 0.0929878 31194.1 300.015 0.98352 0.319147 0.800974 0.800969 9.99958 2.98093e-06 1.19236e-05 0.13044 0.964454 0.922662 -0.0132932 4.89249e-06 0.50004 -1.82768e-20 6.72665e-24 -1.827e-20 0.00139518 0.997818 8.59328e-05 0.15256 2.85176 0.00139518 0.999224 0.621936 0.00103905 0.00187973 0.000859328 0.455639 0.00187973 0.430805 0.000126142 1.02 0.887356 0.534771 0.285604 1.71644e-07 3.05564e-09 2398.69 3406.94 -0.0763415 0.482124 0.27777 0.271339 -0.590047 -0.169462 0.43482 -0.268771 -0.166025 0.969 1 3.83993e-211 277.655 2.06926e-208 1.94098 0.967 0.000299994 0.984314 0.608314 0.786258 0.385025 1.94143 123.436 80.6358 18.5266 59.269 0.0041655 0 -40 10
0.068 1.97258e-09 2.5388e-06 0.0289776 0.0289147 0.0120491 8.96628e-07 0.001154 0.036222 0.000648203 0.0368656 0.845595 101.895 0.24739 0.699725 4.1051 0.0526098 0.0387274 0.961273 0.0198968 0.00422332 0.0191588 0.00406802 0.00510316 0.00584116 0.204127 0.233646 57.9442 -87.8928 125.068 15.9978 145.001 0.000154357 0.267101 192.911 0.310671 0.0673839 0.00409509 0.000561629 0.00138267 0.98699 0.991716 -2.97259e-06 -85.6675 0.0929876 31194.2 300.015 0.98352 0.319147 0.800726 0.800721 9.99958 2.98092e-06 1.19236e-05 0.13044 0.964513 0.922696 -0.0132932 4.89244e-06 0.50004 -1.82783e-20 6.72714e-24 -1.82715e-20 0.00139517 0.997818 8.59326e-05 0.15256 2.85176 0.00139518 0.999215 0.622067 0.00103905 0.00187972 0.000859326 0.45564 0.00187973 0.430817 0.000126144 1.02 0.887354 0.534772 0.285601 1.71643e-07 3.0556e-09 2398.68 3405.88 -0.0762628 0.482123 0.277769 0.271274 -0.590058 -0.169462 0.435055 -0.268772 -0.166258 0.97 1 2.32904e-211 277.726 1.25559e-208 1.94128 0.968 0.000299994 0.983831 0.608409 0.784963 0.385077 1.94173 123.452 80.6474 18.5273 59.2746 0.00416499 0 -40 10
0.069 2.00159e-09 2.5388e-06 0.0291055 0.0290429 0.0120491 9.09812e-07 0.001154 0.0363818 0.000648266 0.0370255 0.845603 101.895 0.24739 0.69973 4.10511 0.0526102 0.0387274 0.961273 0.0198968 0.00422333 0.0191588 0.00406802 0.00510317 0.00584117 0.204127 0.233647 57.9443 -87.8928 125.072 15.9978 145.001 0.000154309 0.267101 192.911 0.310673 0.067384 0.00409508 0.000561627 0.00138266 0.98699 0.991718 -2.97255e-06 -85.6676 0.0929874 31194.3 300.015 0.98352 0.319147 0.800478 0.800473 9.99958 2.98091e-06 1.19235e-05 0.13044 0.964573 0.92273 -0.0132932 4.8924e-06 0.50004 -1.82798e-20 6.72763e-24 -1.8273e-20 0.00139517 0.997818 8.59324e-05 0.152559 2.85176 0.00139517 0.999206 0.622199 0.00103904 0.00187972 0.000859324 0.45564 0.00187972 0.430828 0.000126146 1.02 0.887353 0.534772 0.285599 1.71642e-07 3.05556e-09 2398.66 3404.83 -0.0761844 0.482123 0.277769 0.27121 -0.59007 -0.169462 0.435289 -0.268774 -0.166491 0.971 1 1.41263e-211 277.798 7.61868e-209 1.94159 0.969 0.000299994 0.98335 0.608503 0.783672 0.385129 1.94203 123.468 80.6589 18.528 59.2803 0.00416448 0 -40 10
0.07 2.03059e-09 2.5388e-06 0.0292332 0.029171 0.0120491 9.22997e-07 0.001154 0.0365415 0.000648328 0.0371852 0.845612 101.895 0.247389 0.699735 4.10511 0.0526106 0.0387274 0.961273 0.0198968 0.00422333 0.0191588 0.00406802 0.00510317 0.00584117 0.204127 0.233647 57.9443 -87.8928 125.076 15.9977 145.001 0.000154261 0.2671 192.912 0.310674 0.0673842 0.00409507 0.000561626 0.00138266 0.98699 0.991719 -2.97252e-06 -85.6676 0.0929872 31194.3 300.015 0.98352 0.319147 0.800231 0.800227 9.99958 2.98089e-06 1.19235e-05 0.13044 0.964632 0.922764 -0.0132932 4.89235e-06 0.50004 -1.82813e-20 6.72812e-24 -1.82745e-20 0.00139517 0.997818 8.59322e-05 0.152559 2.85175 0.00139517 0.999197 0.622331 0.00103904 0.00187972 0.000859322 0.455641 0.00187972 0.43084 0.000126148 1.02 0.887351 0.534773 0.285597 1.71642e-07 3.05552e-09 2398.65 3403.78 -0.0761062 0.482123 0.277769 0.271146 -0.590082 -0.169462 0.435522 -0.268775 -0.166723 0.972 1 8.56805e-212 277.869 4.62287e-209 1.94189 0.97 0.000299994 0.982871 0.608598 0.782385 0.385181 1.94233 123.485 80.6704 18.5287 59.286 0.00416397 0 -40 10
0.071 2.0596e-09 2.5388e-06 0.0293608 0.029299 0.0120491 9.36181e-07 0.001154 0.036701 0.00064839 0.0373448 0.845621 101.895 0.247389 0.699741 4.10511 0.0526111 0.0387275 0.961273 0.0198968 0.00422333 0.0191588 0.00406803 0.00510318 0.00584118 0.204127 0.233647 57.9444 -87.8928 125.08 15.9977 145.001 0.000154214 0.2671 192.912 0.310675 0.0673843 0.00409506 0.000561624 0.00138265 0.98699 0.99172 -2.97249e-06 -85.6676 0.0929869 31194.4 300.015 0.98352 0.319147 0.799985 0.799981 9.99958 2.98088e-06 1.19234e-05 0.13044 0.964691 0.922798 -0.0132932 4.89231e-06 0.50004 -1.82828e-20 6.7286e-24 -1.8276e-20 0.00139517 0.997818 8.5932e-05 0.152559 2.85175 0.00139517 0.999188 0.622462 0.00103903 0.00187971 0.00085932 0.455641 0.00187972 0.430852 0.00012615 1.02 0.887349 0.534773 0.285594 1.71641e-07 3.05548e-09 2398.63 3402.74 -0.0760283 0.482123 0.277768 0.271083 -0.590093 -0.169462 0.435755 -0.268777 -0.166954 0.973 1 5.19678e-212 277.94 2.80506e-209 1.94219 0.971 0.000299994 0.982393 0.608692 0.781102 0.385233 1.94263 123.501 80.6819 18.5294 59.2916 0.00416346 0 -40 10
0.072 2.0886e-09 2.5388e-06 0.0294884 0.0294269 0.012049 9.49365e-07 0.001154 0.0368604 0.000648452 0.0375043 0.84563 101.895 0.247388 0.699746 4.10512 0.0526115 0.0387275 0.961272 0.0198968 0.00422334 0.0191588 0.00406803 0.00510318 0.00584118 0.204127 0.233647 57.9444 -87.8928 125.084 15.9977 145.001 0.000154167 0.267099 192.913 0.310676 0.0673845 0.00409505 0.000561622 0.00138265 0.98699 0.991721 -2.97246e-06 -85.6676 0.0929867 31194.4 300.015 0.98352 0.319147 0.79974 0.799735 9.99958 2.98087e-06 1.19234e-05 0.13044 0.96475 0.922832 -0.0132932 4.89226e-06 0.50004 -1.82842e-20 6.72909e-24 -1.82775e-20 0.00139516 0.997818 8.59318e-05 0.152558 2.85175 0.00139516 0.999179 0.622594 0.00103903 0.00187971 0.000859318 0.455642 0.00187971 0.430864 0.000126152 1.02 0.887348 0.534774 0.285592 1.7164e-07 3.05544e-09 2398.62 3401.7 -0.0759507 0.482123 0.277768 0.271019 -0.590105 -0.169462 0.435986 -0.268779 -0.167184 0.974 1 3.15201e-212 278.011 1.70205e-209 1.94249 0.972 0.000299994 0.981917 0.608786 0.779823 0.385285 1.94293 123.517 80.6933 18.53 59.2972 0.00416296 0 -40 10
0.073 2.11761e-09 2.5388e-06 0.0296158 0.0295547 0.012049 9.62549e-07 0.001154 0.0370197 0.000648513 0.0376636 0.845639 101.895 0.247388 0.699752 4.10512 0.052612 0.0387275 0.961272 0.0198968 0.00422334 0.0191588 0.00406803 0.00510319 0.00584118 0.204127 0.233647 57.9445 -87.8928 125.088 15.9976 145.001 0.00015412 0.267099 192.913 0.310677 0.0673846 0.00409505 0.000561621 0.00138264 0.98699 0.991722 -2.97243e-06 -85.6677 0.0929865 31194.5 300.015 0.98352 0.319147 0.799496 0.799491 9.99958 2.98085e-06 1.19233e-05 0.13044 0.964809 0.922865 -0.0132932 4.89222e-06 0.500041 -1.82857e-20 6.72957e-24 -1.8279e-20 0.00139516 0.997818 8.59316e-05 0.152558 2.85175 0.00139516 0.99917 0.622726 0.00103903 0.0018797 0.000859316 0.455643 0.00187971 0.430876 0.000126154 1.02 0.887346 0.534774 0.28559 1.7164e-07 3.0554e-09 2398.6 3400.66 -0.0758733 0.482123 0.277767 0.270956 -0.590116 -0.169462 0.436217 -0.26878 -0.167414 0.975 1 1.91179e-212 278.081 1.03277e-209 1.94279 0.973 0.000299994 0.981442 0.60888 0.778548 0.385337 1.94323 123.533 80.7047 18.5307 59.3028 0.00416245 0 -40 10
0.074 2.14661e-09 2.5388e-06 0.0297431 0.0296824 0.012049 9.75733e-07 0.001154 0.0371789 0.000648574 0.0378229 0.845648 101.895 0.247388 0.699758 4.10512 0.0526124 0.0387276 0.961272 0.0198968 0.00422334 0.0191588 0.00406804 0.00510319 0.00584119 0.204128 0.233648 57.9445 -87.8928 125.092 15.9976 145.002 0.000154073 0.267098 192.914 0.310678 0.0673847 0.00409504 0.000561619 0.00138264 0.98699 0.991722 -2.9724e-06 -85.6677 0.0929863 31194.5 300.015 0.983521 0.319147 0.799252 0.799248 9.99958 2.98084e-06 1.19233e-05 0.130441 0.964867 0.922899 -0.0132932 4.89217e-06 0.500041 -1.82872e-20 6.73006e-24 -1.82805e-20 0.00139516 0.997818 8.59314e-05 0.152558 2.85174 0.00139516 0.999161 0.622857 0.00103902 0.0018797 0.000859314 0.455643 0.0018797 0.430887 0.000126156 1.02 0.887344 0.534775 0.285587 1.71639e-07 3.05536e-09 2398.58 3399.63 -0.0757962 0.482122 0.277767 0.270893 -0.590128 -0.169462 0.436447 -0.268781 -0.167642 0.976 1 1.15956e-212 278.152 6.26661e-210 1.94309 0.974 0.000299994 0.980969 0.608973 0.777278 0.385389 1.94353 123.549 80.7161 18.5314 59.3084 0.00416195 0 -40 10
0.075 2.17562e-09 2.5388e-06 0.0298703 0.02981 0.012049 9.88917e-07 0.001154 0.0373379 0.000648635 0.0379819 0.845658 101.895 0.247387 0.699764 4.10512 0.0526129 0.0387276 0.961272 0.0198968 0.00422335 0.0191588 0.00406804 0.0051032 0.00584119 0.204128 0.233648 57.9446 -87.8928 125.096 15.9976 145.002 0.000154026 0.267098 192.914 0.310679 0.0673848 0.00409503 0.000561617 0.00138263 0.98699 0.991723 -2.97237e-06 -85.6677 0.0929861 31194.6 300.015 0.983521 0.319147 0.79901 0.799005 9.99958 2.98083e-06 1.19232e-05 0.130441 0.964926 0.922932 -0.0132932 4.89213e-06 0.500041 -1.82887e-20 6.73054e-24 -1.8282e-20 0.00139515 0.997818 8.59312e-05 0.152557 2.85174 0.00139515 0.999153 0.622989 0.00103902 0.0018797 0.000859312 0.455644 0.0018797 0.430899 0.000126158 1.02 0.887343 0.534775 0.285585 1.71638e-07 3.05532e-09 2398.57 3398.6 -0.0757193 0.482122 0.277767 0.27083 -0.590139 -0.169463 0.436677 -0.268783 -0.16787 0.977 1 7.03308e-213 278.222 3.80244e-210 1.94339 0.975 0.000299994 0.980497 0.609067 0.776011 0.38544 1.94383 123.565 80.7274 18.5321 59.3139 0.00416145 0 -40 10
0.076 2.20462e-09 2.5388e-06 0.0299975 0.0299376 0.012049 1.0021e-06 0.001154 0.0374968 0.000648695 0.0381409 0.845667 101.895 0.247387 0.69977 4.10513 0.0526134 0.0387276 0.961272 0.0198968 0.00422335 0.0191588 0.00406804 0.0051032 0.0058412 0.204128 0.233648 57.9446 -87.8928 125.1 15.9975 145.002 0.000153979 0.267097 192.914 0.31068 0.067385 0.00409502 0.000561616 0.00138262 0.98699 0.991724 -2.97234e-06 -85.6677 0.0929858 31194.6 300.015 0.983521 0.319147 0.798768 0.798763 9.99958 2.98082e-06 1.19232e-05 0.130441 0.964984 0.922965 -0.0132932 4.89209e-06 0.500041 -1.82902e-20 6.73103e-24 -1.82835e-20 0.00139515 0.997818 8.5931e-05 0.152557 2.85174 0.00139515 0.999144 0.62312 0.00103902 0.00187969 0.00085931 0.455644 0.0018797 0.430911 0.00012616 1.02 0.887341 0.534776 0.285583 1.71638e-07 3.05529e-09 2398.55 3397.57 -0.0756427 0.482122 0.277766 0.270767 -0.59015 -0.169463 0.436905 -0.268784 -0.168098 0.978 1 4.26578e-213 278.292 2.30723e-210 1.94369 0.976 0.000299994 0.980027 0.60916 0.774748 0.385492 1.94413 123.581 80.7387 18.5328 59.3195 0.00416095 0 -40 10
0.077 2.23363e-09 2.5388e-06 0.0301245 0.030065 0.012049 1.01528e-06 0.001154 0.0376556 0.000648754 0.0382997 0.845677 101.895 0.247386 0.699776 4.10513 0.0526139 0.0387277 0.961272 0.0198968 0.00422336 0.0191588 0.00406805 0.00510321 0.0058412 0.204128 0.233648 57.9447 -87.8928 125.104 15.9975 145.002 0.000153933 0.267097 192.915 0.310681 0.0673851 0.00409502 0.000561614 0.00138262 0.98699 0.991725 -2.97231e-06 -85.6677 0.0929856 31194.7 300.016 0.983521 0.319147 0.798526 0.798522 9.99958 2.98081e-06 1.19231e-05 0.130441 0.965042 0.922998 -0.0132932 4.89204e-06 0.500041 -1.82917e-20 6.73151e-24 -1.82849e-20 0.00139515 0.997818 8.59308e-05 0.152556 2.85174 0.00139515 0.999135 0.623251 0.00103901 0.00187969 0.000859308 0.455645 0.00187969 0.430923 0.000126162 1.02 0.88734 0.534776 0.285581 1.71637e-07 3.05525e-09 2398.54 3396.54 -0.0755663 0.482122 0.277766 0.270705 -0.590162 -0.169463 0.437133 -0.268786 -0.168324 0.979 1 2.58733e-213 278.362 1.39997e-210 1.94399 0.977 0.000299994 0.979559 0.609254 0.773489 0.385544 1.94443 123.597 80.75 18.5335 59.325 0.00416045 0 -40 10
0.078 2.26263e-09 2.5388e-06 0.0302514 0.0301924 0.012049 1.02847e-06 0.001154 0.0378142 0.000648813 0.0384584 0.845686 101.895 0.247386 0.699783 4.10514 0.0526144 0.0387277 0.961272 0.0198968 0.00422336 0.0191588 0.00406805 0.00510321 0.00584121 0.204128 0.233648 57.9448 -87.8928 125.108 15.9975 145.002 0.000153886 0.267097 192.915 0.310682 0.0673852 0.00409501 0.000561612 0.00138261 0.986991 0.991725 -2.97228e-06 -85.6678 0.0929854 31194.8 300.016 0.983521 0.319147 0.798286 0.798281 9.99958 2.98079e-06 1.19231e-05 0.130441 0.9651 0.923031 -0.0132933 4.892e-06 0.500041 -1.82931e-20 6.73199e-24 -1.82864e-20 0.00139515 0.997818 8.59306e-05 0.152556 2.85173 0.00139515 0.999127 0.623383 0.00103901 0.00187969 0.000859306 0.455645 0.00187969 0.430935 0.000126165 1.02 0.887338 0.534776 0.285579 1.71636e-07 3.05521e-09 2398.52 3395.52 -0.0754902 0.482122 0.277765 0.270642 -0.590173 -0.169463 0.43736 -0.268787 -0.16855 0.98 1 1.56929e-213 278.431 8.49468e-211 1.94428 0.978 0.000299994 0.979092 0.609347 0.772234 0.385595 1.94472 123.612 80.7612 18.5341 59.3305 0.00415996 0 -40 10
0.079 2.29163e-09 2.5388e-06 0.0303782 0.0303196 0.012049 1.04165e-06 0.001154 0.0379728 0.000648872 0.038617 0.845696 101.895 0.247385 0.699789 4.10514 0.0526149 0.0387277 0.961272 0.0198968 0.00422336 0.0191588 0.00406805 0.00510322 0.00584121 0.204129 0.233649 57.9448 -87.8928 125.112 15.9974 145.002 0.00015384 0.267096 192.916 0.310683 0.0673854 0.004095 0.000561611 0.00138261 0.986991 0.991726 -2.97225e-06 -85.6678 0.0929852 31194.8 300.016 0.983521 0.319147 0.798046 0.798042 9.99958 2.98078e-06 1.1923e-05 0.130441 0.965157 0.923064 -0.0132933 4.89196e-06 0.500042 -1.82946e-20 6.73247e-24 -1.82879e-20 0.00139514 0.997818 8.59304e-05 0.152556 2.85173 0.00139514 0.999118 0.623514 0.00103901 0.00187968 0.000859304 0.455646 0.00187969 0.430946 0.000126167 1.02 0.887336 0.534777 0.285576 1.71636e-07 3.05517e-09 2398.51 3394.51 -0.0754144 0.482121 0.277765 0.27058 -0.590184 -0.169463 0.437586 -0.268789 -0.168775 0.981 1 9.51824e-214 278.501 5.15435e-211 1.94458 0.979 0.000299994 0.978627 0.60944 0.770983 0.385646 1.94502 123.628 80.7724 18.5348 59.336 0.00415946 0 -40 10
0.08 2.32064e-09 2.5388e-06 0.0305049 0.0304467 0.0120489 1.05484e-06 0.001154 0.0381311 0.000648931 0.0387755 0.845706 101.895 0.247385 0.699796 4.10514 0.0526154 0.0387278 0.961272 0.0198968 0.00422337 0.0191588 0.00406806 0.00510322 0.00584122 0.204129 0.233649 57.9449 -87.8928 125.116 15.9974 145.002 0.000153794 0.267096 192.916 0.310684 0.0673855 0.004095 0.000561609 0.0013826 0.986991 0.991726 -2.97222e-06 -85.6678 0.092985 31194.9 300.016 0.983521 0.319147 0.797808 0.797803 9.99958 2.98077e-06 1.1923e-05 0.130441 0.965215 0.923097 -0.0132933 4.89192e-06 0.500042 -1.82961e-20 6.73295e-24 -1.82893e-20 0.00139514 0.997818 8.59302e-05 0.152555 2.85173 0.00139514 0.99911 0.623645 0.00103901 0.00187968 0.000859302 0.455646 0.00187968 0.430958 0.000126169 1.02 0.887335 0.534777 0.285574 1.71635e-07 3.05514e-09 2398.49 3393.49 -0.0753388 0.482121 0.277765 0.270518 -0.590196 -0.169463 0.437812 -0.26879 -0.169 0.982 1 5.7731e-214 278.57 3.12753e-211 1.94488 0.98 0.000299994 0.978163 0.609533 0.769736 0.385698 1.94532 123.644 80.7836 18.5355 59.3415 0.00415897 0 -40 10
0.081 2.34964e-09 2.5388e-06 0.0306315 0.0305738 0.0120489 1.06802e-06 0.001154 0.0382894 0.000648989 0.0389338 0.845716 101.895 0.247384 0.699803 4.10515 0.0526159 0.0387278 0.961272 0.0198968 0.00422337 0.0191588 0.00406806 0.00510323 0.00584122 0.204129 0.233649 57.9449 -87.8928 125.12 15.9973 145.002 0.000153748 0.267095 192.916 0.310685 0.0673856 0.00409499 0.000561608 0.0013826 0.986991 0.991727 -2.97219e-06 -85.6678 0.0929848 31194.9 300.016 0.983521 0.319147 0.79757 0.797565 9.99958 2.98076e-06 1.19229e-05 0.130441 0.965272 0.923129 -0.0132933 4.89188e-06 0.500042 -1.82975e-20 6.73343e-24 -1.82908e-20 0.00139514 0.997818 8.593e-05 0.152555 2.85173 0.00139514 0.999101 0.623776 0.001039 0.00187968 0.0008593 0.455647 0.00187968 0.43097 0.000126171 1.02 0.887333 0.534778 0.285572 1.71634e-07 3.0551e-09 2398.47 3392.48 -0.0752634 0.482121 0.277764 0.270457 -0.590207 -0.169463 0.438037 -0.268791 -0.169223 0.983 1 3.50156e-214 278.639 1.8977e-211 1.94517 0.981 0.000299994 0.977701 0.609625 0.768493 0.385749 1.94561 123.66 80.7947 18.5362 59.347 0.00415848 0 -40 10
0.082 2.37865e-09 2.5388e-06 0.030758 0.0307007 0.0120489 1.0812e-06 0.001154 0.0384476 0.000649046 0.039092 0.845726 101.895 0.247384 0.699809 4.10515 0.0526165 0.0387278 0.961272 0.0198968 0.00422338 0.0191588 0.00406806 0.00510323 0.00584123 0.204129 0.233649 57.945 -87.8928 125.124 15.9973 145.002 0.000153703 0.267095 192.917 0.310686 0.0673857 0.00409498 0.000561606 0.00138259 0.986991 0.991728 -2.97216e-06 -85.6679 0.0929846 31195 300.016 0.983521 0.319147 0.797332 0.797328 9.99958 2.98075e-06 1.19229e-05 0.130441 0.965329 0.923161 -0.0132933 4.89184e-06 0.500042 -1.8299e-20 6.73391e-24 -1.82923e-20 0.00139514 0.997818 8.59299e-05 0.152555 2.85173 0.00139514 0.999093 0.623907 0.001039 0.00187967 0.000859299 0.455647 0.00187967 0.430982 0.000126173 1.02 0.887332 0.534778 0.28557 1.71634e-07 3.05506e-09 2398.46 3391.47 -0.0751883 0.482121 0.277764 0.270395 -0.590218 -0.169463 0.438261 -0.268793 -0.169446 0.984 1 2.12381e-214 278.707 1.15147e-211 1.94547 0.982 0.000299994 0.977241 0.609718 0.767254 0.3858 1.94591 123.676 80.8058 18.5368 59.3524 0.00415799 0 -40 10
0.083 2.40765e-09 2.5388e-06 0.0308845 0.0308276 0.0120489 1.09439e-06 0.001154 0.0386056 0.000649103 0.0392501 0.845736 101.895 0.247383 0.699816 4.10515 0.0526171 0.0387279 0.961272 0.0198968 0.00422338 0.0191588 0.00406807 0.00510324 0.00584123 0.20413 0.233649 57.945 -87.8929 125.128 15.9973 145.002 0.000153657 0.267094 192.917 0.310687 0.0673858 0.00409497 0.000561605 0.00138259 0.986991 0.991728 -2.97213e-06 -85.6679 0.0929844 31195 300.016 0.983521 0.319147 0.797096 0.797091 9.99958 2.98074e-06 1.19228e-05 0.130441 0.965386 0.923194 -0.0132933 4.8918e-06 0.500042 -1.83004e-20 6.73439e-24 -1.82937e-20 0.00139513 0.997818 8.59297e-05 0.152554 2.85172 0.00139513 0.999084 0.624039 0.001039 0.00187967 0.000859297 0.455648 0.00187967 0.430993 0.000126175 1.02 0.88733 0.534779 0.285568 1.71633e-07 3.05503e-09 2398.44 3390.47 -0.0751135 0.482121 0.277764 0.270334 -0.590229 -0.169463 0.438484 -0.268794 -0.169668 0.985 1 1.28815e-214 278.776 6.98681e-212 1.94577 0.983 0.000299994 0.976781 0.60981 0.766019 0.385851 1.9462 123.692 80.8168 18.5375 59.3578 0.0041575 0 -40 10
0.084 2.43665e-09 2.5388e-06 0.0310108 0.0309543 0.0120489 1.10757e-06 0.001154 0.0387635 0.00064916 0.039408 0.845747 101.895 0.247382 0.699824 4.10516 0.0526176 0.0387279 0.961272 0.0198968 0.00422339 0.0191588 0.00406807 0.00510324 0.00584124 0.20413 0.23365 57.9451 -87.8929 125.132 15.9972 145.002 0.000153612 0.267094 192.917 0.310688 0.067386 0.00409497 0.000561603 0.00138258 0.986991 0.991728 -2.97211e-06 -85.6679 0.0929842 31195.1 300.016 0.983521 0.319147 0.79686 0.796855 9.99958 2.98072e-06 1.19228e-05 0.130441 0.965443 0.923226 -0.0132933 4.89176e-06 0.500042 -1.83019e-20 6.73487e-24 -1.82952e-20 0.00139513 0.997818 8.59295e-05 0.152554 2.85172 0.00139513 0.999076 0.62417 0.001039 0.00187967 0.000859295 0.455648 0.00187967 0.431005 0.000126178 1.02 0.887329 0.534779 0.285566 1.71633e-07 3.05499e-09 2398.43 3389.47 -0.0750389 0.482121 0.277763 0.270273 -0.59024 -0.169463 0.438706 -0.268795 -0.16989 0.986 1 7.81305e-215 278.844 4.2394e-212 1.94606 0.984 0.000299994 0.976324 0.609903 0.764787 0.385902 1.9465 123.707 80.8278 18.5382 59.3632 0.00415702 0 -40 10
0.085 2.46566e-09 2.5388e-06 0.031137 0.031081 0.0120489 1.12075e-06 0.001154 0.0389212 0.000649216 0.0395658 0.845757 101.895 0.247382 0.699831 4.10516 0.0526182 0.0387279 0.961272 0.0198968 0.00422339 0.0191588 0.00406808 0.00510325 0.00584125 0.20413 0.23365 57.9451 -87.8929 125.136 15.9972 145.002 0.000153566 0.267093 192.918 0.310689 0.0673861 0.00409496 0.000561602 0.00138258 0.986991 0.991729 -2.97208e-06 -85.6679 0.092984 31195.1 300.017 0.983521 0.319147 0.796625 0.79662 9.99958 2.98071e-06 1.19227e-05 0.130441 0.965499 0.923258 -0.0132933 4.89172e-06 0.500043 -1.83033e-20 6.73535e-24 -1.82966e-20 0.00139513 0.997818 8.59293e-05 0.152554 2.85172 0.00139513 0.999068 0.624301 0.001039 0.00187966 0.000859293 0.455649 0.00187966 0.431017 0.00012618 1.02 0.887327 0.534779 0.285564 1.71632e-07 3.05496e-09 2398.41 3388.47 -0.0749645 0.48212 0.277763 0.270212 -0.590251 -0.169463 0.438928 -0.268796 -0.170111 0.987 1 4.73885e-215 278.912 2.57234e-212 1.94636 0.985 0.000299994 0.975868 0.609995 0.76356 0.385953 1.94679 123.723 80.8388 18.5388 59.3686 0.00415653 0 -40 10
0.086 2.49466e-09 2.5388e-06 0.0312631 0.0312075 0.0120489 1.13394e-06 0.001154 0.0390788 0.000649272 0.0397235 0.845768 101.895 0.247381 0.699838 4.10517 0.0526188 0.038728 0.961272 0.0198967 0.0042234 0.0191587 0.00406808 0.00510326 0.00584125 0.20413 0.23365 57.9452 -87.8929 125.14 15.9972 145.002 0.000153521 0.267093 192.918 0.31069 0.0673862 0.00409495 0.0005616 0.00138257 0.986991 0.991729 -2.97205e-06 -85.6679 0.0929838 31195.2 300.017 0.983521 0.319147 0.796391 0.796386 9.99958 2.9807e-06 1.19227e-05 0.130441 0.965556 0.92329 -0.0132933 4.89168e-06 0.500043 -1.83048e-20 6.73583e-24 -1.82981e-20 0.00139512 0.997818 8.59291e-05 0.152553 2.85172 0.00139513 0.99906 0.624432 0.00103899 0.00187966 0.000859291 0.45565 0.00187966 0.431029 0.000126182 1.02 0.887326 0.53478 0.285562 1.71631e-07 3.05492e-09 2398.4 3387.48 -0.0748904 0.48212 0.277762 0.270151 -0.590262 -0.169464 0.439149 -0.268798 -0.170331 0.988 1 2.87426e-215 278.98 1.56082e-212 1.94665 0.986 0.000299994 0.975413 0.610087 0.762336 0.386004 1.94709 123.739 80.8498 18.5395 59.374 0.00415605 0 -40 10
0.087 2.52367e-09 2.5388e-06 0.0313891 0.031334 0.0120489 1.14712e-06 0.001154 0.0392364 0.000649327 0.0398811 0.845779 101.895 0.247381 0.699846 4.10517 0.0526194 0.038728 0.961272 0.0198967 0.0042234 0.0191587 0.00406808 0.00510326 0.00584126 0.20413 0.23365 57.9453 -87.8929 125.144 15.9971 145.002 0.000153476 0.267093 192.919 0.310691 0.0673863 0.00409495 0.000561599 0.00138257 0.986991 0.99173 -2.97202e-06 -85.668 0.0929836 31195.2 300.017 0.983521 0.319147 0.796158 0.796153 9.99958 2.98069e-06 1.19227e-05 0.130441 0.965612 0.923321 -0.0132933 4.89164e-06 0.500043 -1.83062e-20 6.7363e-24 -1.82995e-20 0.00139512 0.997818 8.59289e-05 0.152553 2.85172 0.00139512 0.999052 0.624562 0.00103899 0.00187966 0.000859289 0.45565 0.00187966 0.43104 0.000126184 1.02 0.887325 0.53478 0.28556 1.71631e-07 3.05489e-09 2398.38 3386.49 -0.0748166 0.48212 0.277762 0.27009 -0.590273 -0.169464 0.43937 -0.268799 -0.17055 0.989 1 1.74333e-215 279.048 9.47058e-213 1.94695 0.987 0.000299994 0.97496 0.610179 0.761116 0.386055 1.94738 123.754 80.8607 18.5402 59.3793 0.00415557 0 -40 10
0.088 2.55267e-09 2.5388e-06 0.031515 0.0314604 0.0120488 1.1603e-06 0.001154 0.0393937 0.000649382 0.0400385 0.84579 101.895 0.24738 0.699854 4.10517 0.05262 0.0387281 0.961272 0.0198967 0.00422341 0.0191587 0.00406809 0.00510327 0.00584126 0.204131 0.233651 57.9453 -87.8929 125.148 15.9971 145.002 0.000153431 0.267092 192.919 0.310692 0.0673864 0.00409494 0.000561597 0.00138256 0.986991 0.99173 -2.97199e-06 -85.668 0.0929834 31195.3 300.017 0.983521 0.319147 0.795925 0.79592 9.99958 2.98068e-06 1.19226e-05 0.130441 0.965668 0.923353 -0.0132933 4.89161e-06 0.500043 -1.83077e-20 6.73678e-24 -1.83009e-20 0.00139512 0.997818 8.59288e-05 0.152553 2.85171 0.00139512 0.999044 0.624693 0.00103899 0.00187965 0.000859288 0.455651 0.00187965 0.431052 0.000126187 1.02 0.887323 0.534781 0.285558 1.7163e-07 3.05486e-09 2398.36 3385.5 -0.0747429 0.48212 0.277762 0.27003 -0.590284 -0.169464 0.439589 -0.2688 -0.170769 0.99 1 1.05738e-215 279.115 5.74645e-213 1.94724 0.988 0.000299994 0.974509 0.610271 0.7599 0.386105 1.94767 123.77 80.8716 18.5408 59.3847 0.00415509 0 -40 10
0.089 2.58167e-09 2.5388e-06 0.0316408 0.0315866 0.0120488 1.17349e-06 0.001154 0.039551 0.000649436 0.0401958 0.845801 101.895 0.247379 0.699862 4.10518 0.0526206 0.0387281 0.961272 0.0198967 0.00422341 0.0191587 0.00406809 0.00510327 0.00584127 0.204131 0.233651 57.9454 -87.8929 125.152 15.9971 145.002 0.000153387 0.267092 192.919 0.310693 0.0673866 0.00409493 0.000561596 0.00138256 0.986991 0.99173 -2.97196e-06 -85.668 0.0929832 31195.3 300.017 0.983521 0.319147 0.795693 0.795688 9.99958 2.98067e-06 1.19226e-05 0.130441 0.965724 0.923384 -0.0132933 4.89157e-06 0.500043 -1.83091e-20 6.73725e-24 -1.83024e-20 0.00139512 0.997818 8.59286e-05 0.152552 2.85171 0.00139512 0.999036 0.624824 0.00103899 0.00187965 0.000859286 0.455651 0.00187965 0.431064 0.000126189 1.02 0.887322 0.534781 0.285556 1.7163e-07 3.05482e-09 2398.35 3384.51 -0.0746696 0.48212 0.277761 0.26997 -0.590295 -0.169464 0.439808 -0.268801 -0.170987 0.991 1 6.41334e-216 279.182 3.48677e-213 1.94753 0.989 0.000299994 0.974059 0.610362 0.758687 0.386156 1.94796 123.786 80.8824 18.5415 59.39 0.00415461 0 -40 10
0.09 2.61068e-09 2.5388e-06 0.0317665 0.0317128 0.0120488 1.18667e-06 0.001154 0.0397081 0.00064949 0.040353 0.845812 101.895 0.247379 0.69987 4.10518 0.0526213 0.0387281 0.961272 0.0198967 0.00422342 0.0191587 0.0040681 0.00510328 0.00584128 0.204131 0.233651 57.9454 -87.8929 125.156 15.997 145.002 0.000153342 0.267091 192.92 0.310694 0.0673867 0.00409493 0.000561594 0.00138256 0.986991 0.991731 -2.97194e-06 -85.668 0.092983 31195.4 300.017 0.983521 0.319147 0.795462 0.795457 9.99958 2.98066e-06 1.19225e-05 0.130441 0.965779 0.923416 -0.0132933 4.89153e-06 0.500044 -1.83105e-20 6.73773e-24 -1.83038e-20 0.00139511 0.997818 8.59284e-05 0.152552 2.85171 0.00139512 0.999028 0.624955 0.00103899 0.00187965 0.000859284 0.455651 0.00187965 0.431075 0.000126191 1.02 0.88732 0.534781 0.285554 1.71629e-07 3.05479e-09 2398.33 3383.53 -0.0745964 0.48212 0.277761 0.26991 -0.590306 -0.169464 0.440026 -0.268802 -0.171204 0.992 1 3.88989e-216 279.249 2.11566e-213 1.94783 0.99 0.000299994 0.97361 0.610454 0.757479 0.386206 1.94826 123.801 80.8933 18.5421 59.3953 0.00415414 0 -40 10
0.091 2.63968e-09 2.5388e-06 0.0318921 0.0318388 0.0120488 1.19985e-06 0.001154 0.0398651 0.000649544 0.0405101 0.845823 101.895 0.247378 0.699878 4.10519 0.0526219 0.0387282 0.961272 0.0198967 0.00422342 0.0191587 0.0040681 0.00510329 0.00584128 0.204131 0.233651 57.9455 -87.8929 125.16 15.997 145.002 0.000153298 0.267091 192.92 0.310695 0.0673868 0.00409492 0.000561593 0.00138255 0.986991 0.991731 -2.97191e-06 -85.668 0.0929829 31195.4 300.017 0.983521 0.319147 0.795232 0.795227 9.99958 2.98065e-06 1.19225e-05 0.130441 0.965835 0.923447 -0.0132933 4.8915e-06 0.500044 -1.8312e-20 6.7382e-24 -1.83052e-20 0.00139511 0.997818 8.59282e-05 0.152552 2.85171 0.00139511 0.99902 0.625086 0.00103899 0.00187964 0.000859282 0.455652 0.00187964 0.431087 0.000126193 1.02 0.887319 0.534782 0.285552 1.71628e-07 3.05476e-09 2398.32 3382.56 -0.0745236 0.482119 0.27776 0.26985 -0.590317 -0.169464 0.440244 -0.268803 -0.17142 0.993 1 2.35934e-216 279.316 1.28371e-213 1.94812 0.991 0.000299994 0.973163 0.610545 0.756274 0.386257 1.94855 123.817 80.904 18.5428 59.4006 0.00415366 0 -40 10
0.092 2.66868e-09 2.5388e-06 0.0320176 0.0319648 0.0120488 1.21304e-06 0.001154 0.040022 0.000649597 0.040667 0.845834 101.895 0.247377 0.699886 4.10519 0.0526226 0.0387282 0.961272 0.0198967 0.00422343 0.0191587 0.0040681 0.00510329 0.00584129 0.204132 0.233652 57.9455 -87.8929 125.163 15.997 145.002 0.000153253 0.267091 192.92 0.310696 0.0673869 0.00409491 0.000561591 0.00138255 0.986991 0.991731 -2.97188e-06 -85.6681 0.0929827 31195.5 300.017 0.983521 0.319147 0.795002 0.794997 9.99958 2.98064e-06 1.19224e-05 0.130441 0.96589 0.923478 -0.0132933 4.89146e-06 0.500044 -1.83134e-20 6.73868e-24 -1.83067e-20 0.00139511 0.997818 8.59281e-05 0.152551 2.85171 0.00139511 0.999012 0.625216 0.00103899 0.00187964 0.000859281 0.455652 0.00187964 0.431099 0.000126196 1.02 0.887318 0.534782 0.28555 1.71628e-07 3.05473e-09 2398.3 3381.58 -0.0744509 0.482119 0.27776 0.26979 -0.590328 -0.169464 0.44046 -0.268805 -0.171636 0.994 1 1.43101e-216 279.383 7.78912e-214 1.94841 0.992 0.000299994 0.972718 0.610636 0.755073 0.386307 1.94884 123.833 80.9148 18.5434 59.4059 0.00415319 0 -40 10
0.093 2.69768e-09 2.5388e-06 0.032143 0.0320906 0.0120488 1.22622e-06 0.001154 0.0401787 0.00064965 0.0408238 0.845846 101.895 0.247377 0.699895 4.1052 0.0526233 0.0387283 0.961272 0.0198967 0.00422343 0.0191587 0.00406811 0.0051033 0.0058413 0.204132 0.233652 57.9456 -87.8929 125.167 15.9969 145.002 0.000153209 0.26709 192.921 0.310697 0.067387 0.00409491 0.00056159 0.00138254 0.986991 0.991731 -2.97186e-06 -85.6681 0.0929825 31195.5 300.018 0.983521 0.319147 0.794773 0.794768 9.99958 2.98063e-06 1.19224e-05 0.130441 0.965945 0.923509 -0.0132933 4.89142e-06 0.500044 -1.83148e-20 6.73915e-24 -1.83081e-20 0.00139511 0.997818 8.59279e-05 0.152551 2.8517 0.00139511 0.999004 0.625347 0.00103899 0.00187964 0.000859279 0.455653 0.00187964 0.431111 0.000126198 1.02 0.887316 0.534783 0.285549 1.71627e-07 3.05469e-09 2398.28 3380.61 -0.0743785 0.482119 0.27776 0.269731 -0.590339 -0.169464 0.440676 -0.268806 -0.171851 0.995 1 8.67951e-217 279.449 4.72617e-214 1.9487 0.993 0.000299994 0.972274 0.610728 0.753876 0.386357 1.94913 123.848 80.9255 18.5441 59.4111 0.00415272 0 -40 10
0.094 2.72669e-09 2.5388e-06 0.0322683 0.0322164 0.0120488 1.2394e-06 0.001154 0.0403354 0.000649702 0.0409805 0.845857 101.895 0.247376 0.699903 4.1052 0.0526239 0.0387283 0.961272 0.0198967 0.00422344 0.0191587 0.00406811 0.00510331 0.0058413 0.204132 0.233652 57.9457 -87.8929 125.171 15.9969 145.002 0.000153165 0.26709 192.921 0.310698 0.0673871 0.0040949 0.000561589 0.00138254 0.986992 0.991732 -2.97183e-06 -85.6681 0.0929823 31195.6 300.018 0.983521 0.319147 0.794545 0.79454 9.99958 2.98062e-06 1.19224e-05 0.130441 0.966 0.92354 -0.0132933 4.89139e-06 0.500045 -1.83162e-20 6.73962e-24 -1.83095e-20 0.00139511 0.997818 8.59277e-05 0.152551 2.8517 0.00139511 0.998996 0.625478 0.00103899 0.00187963 0.000859277 0.455653 0.00187964 0.431122 0.0001262 1.02 0.887315 0.534783 0.285547 1.71627e-07 3.05466e-09 2398.27 3379.64 -0.0743064 0.482119 0.277759 0.269672 -0.59035 -0.169464 0.440892 -0.268807 -0.172065 0.996 1 5.26439e-217 279.516 2.86768e-214 1.94899 0.994 0.000299994 0.971831 0.610819 0.752682 0.386408 1.94942 123.864 80.9362 18.5447 59.4164 0.00415225 0 -40 10
0.095 2.75569e-09 2.5388e-06 0.0323935 0.032342 0.0120487 1.25259e-06 0.001154 0.0404919 0.000649753 0.041137 0.845869 101.895 0.247375 0.699912 4.10521 0.0526246 0.0387284 0.961272 0.0198967 0.00422344 0.0191587 0.00406812 0.00510331 0.00584131 0.204133 0.233652 57.9457 -87.8929 125.175 15.9969 145.002 0.000153122 0.267089 192.921 0.310698 0.0673872 0.0040949 0.000561587 0.00138253 0.986992 0.991732 -2.9718e-06 -85.6681 0.0929821 31195.6 300.018 0.983522 0.319147 0.794318 0.794313 9.99958 2.98061e-06 1.19223e-05 0.130442 0.966055 0.92357 -0.0132933 4.89135e-06 0.500045 -1.83177e-20 6.7401e-24 -1.83109e-20 0.0013951 0.997818 8.59276e-05 0.15255 2.8517 0.0013951 0.998989 0.625608 0.00103899 0.00187963 0.000859276 0.455654 0.00187963 0.431134 0.000126203 1.02 0.887314 0.534783 0.285545 1.71626e-07 3.05463e-09 2398.25 3378.67 -0.0742344 0.482119 0.277759 0.269613 -0.59036 -0.169464 0.441106 -0.268808 -0.172279 0.997 1 3.19301e-217 279.582 1.74e-214 1.94928 0.995 0.000299994 0.97139 0.610909 0.751493 0.386458 1.94971 123.879 80.9469 18.5453 59.4216 0.00415178 0 -40 10
0.096 2.78469e-09 2.5388e-06 0.0325186 0.0324675 0.0120487 1.26577e-06 0.001154 0.0406483 0.000649805 0.0412935 0.845881 101.895 0.247375 0.699921 4.10521 0.0526253 0.0387284 0.961272 0.0198967 0.00422345 0.0191587 0.00406812 0.00510332 0.00584132 0.204133 0.233653 57.9458 -87.8929 125.179 15.9968 145.002 0.000153078 0.267089 192.922 0.310699 0.0673873 0.00409489 0.000561586 0.00138253 0.986992 0.991732 -2.97178e-06 -85.6681 0.0929819 31195.7 300.018 0.983522 0.319147 0.794091 0.794086 9.99958 2.9806e-06 1.19223e-05 0.130442 0.96611 0.923601 -0.0132933 4.89132e-06 0.500045 -1.83191e-20 6.74057e-24 -1.83123e-20 0.0013951 0.997818 8.59274e-05 0.15255 2.8517 0.0013951 0.998981 0.625739 0.00103899 0.00187963 0.000859274 0.455654 0.00187963 0.431146 0.000126205 1.02 0.887312 0.534784 0.285543 1.71626e-07 3.0546e-09 2398.24 3377.71 -0.0741627 0.482119 0.277759 0.269554 -0.590371 -0.169464 0.44132 -0.268809 -0.172492 0.998 1 1.93666e-217 279.648 1.05577e-214 1.94957 0.996 0.000299994 0.97095 0.611 0.750307 0.386508 1.95 123.895 80.9575 18.546 59.4268 0.00415131 0 -40 10
0.097 2.8137e-09 2.5388e-06 0.0326436 0.032593 0.0120487 1.27895e-06 0.001154 0.0408045 0.000649856 0.0414498 0.845892 101.895 0.247374 0.69993 4.10522 0.0526261 0.0387285 0.961272 0.0198967 0.00422346 0.0191587 0.00406813 0.00510333 0.00584132 0.204133 0.233653 57.9458 -87.8929 125.183 15.9968 145.002 0.000153034 0.267089 192.922 0.3107 0.0673874 0.00409488 0.000561584 0.00138252 0.986992 0.991732 -2.97175e-06 -85.6682 0.0929818 31195.7 300.018 0.983522 0.319147 0.793865 0.793861 9.99958 2.98059e-06 1.19222e-05 0.130442 0.966164 0.923632 -0.0132933 4.89129e-06 0.500045 -1.83205e-20 6.74104e-24 -1.83137e-20 0.0013951 0.997818 8.59272e-05 0.15255 2.8517 0.0013951 0.998973 0.625869 0.00103899 0.00187962 0.000859272 0.455655 0.00187963 0.431157 0.000126207 1.02 0.887311 0.534784 0.285541 1.71625e-07 3.05457e-09 2398.22 3376.75 -0.0740913 0.482118 0.277758 0.269495 -0.590382 -0.169465 0.441533 -0.26881 -0.172704 0.999 1 1.17464e-217 279.713 6.40604e-215 1.94986 0.997 0.000299994 0.970512 0.611091 0.749124 0.386558 1.95029 123.91 80.9681 18.5466 59.432 0.00415085 0 -40 10
0.098 2.8427e-09 2.5388e-06 0.0327685 0.0327183 0.0120487 1.29214e-06 0.001154 0.0409606 0.000649906 0.0416059 0.845904 101.895 0.247373 0.699939 4.10522 0.0526268 0.0387285 0.961271 0.0198967 0.00422346 0.0191587 0.00406813 0.00510333 0.00584133 0.204133 0.233653 57.9459 -87.8929 125.186 15.9968 145.002 0.000152991 0.267088 192.922 0.310701 0.0673875 0.00409488 0.000561583 0.00138252 0.986992 0.991732 -2.97172e-06 -85.6682 0.0929816 31195.7 300.018 0.983522 0.319147 0.79364 0.793635 9.99958 2.98058e-06 1.19222e-05 0.130442 0.966219 0.923662 -0.0132933 4.89125e-06 0.500046 -1.83219e-20 6.74151e-24 -1.83152e-20 0.0013951 0.997818 8.59271e-05 0.152549 2.85169 0.0013951 0.998966 0.625999 0.00103899 0.00187962 0.000859271 0.455655 0.00187962 0.431169 0.00012621 1.02 0.88731 0.534784 0.28554 1.71624e-07 3.05454e-09 2398.21 3375.8 -0.0740201 0.482118 0.277758 0.269436 -0.590393 -0.169465 0.441745 -0.268811 -0.172916 1 1 7.12458e-218 279.779 3.88694e-215 1.95015 0.998 0.000299994 0.970076 0.611181 0.747945 0.386608 1.95058 123.926 80.9786 18.5473 59.4372 0.00415038 0 -40 10
0.099 2.8717e-09 2.5388e-06 0.0328933 0.0328436 0.0120487 1.30532e-06 0.001154 0.0411166 0.000649956 0.041762 0.845917 101.895 0.247372 0.699949 4.10523 0.0526275 0.0387286 0.961271 0.0198967 0.00422347 0.0191587 0.00406814 0.00510334 0.00584134 0.204134 0.233653 57.9459 -87.8929 125.19 15.9967 145.002 0.000152948 0.267088 192.923 0.310702 0.0673876 0.00409487 0.000561582 0.00138251 0.986992 0.991733 -2.9717e-06 -85.6682 0.0929814 31195.8 300.019 0.983522 0.319147 0.793416 0.793411 9.99958 2.98057e-06 1.19222e-05 0.130442 0.966273 0.923692 -0.0132933 4.89122e-06 0.500046 -1.83233e-20 6.74198e-24 -1.83166e-20 0.00139509 0.997818 8.59269e-05 0.152549 2.85169 0.00139509 0.998958 0.62613 0.00103899 0.00187962 0.000859269 0.455656 0.00187962 0.431181 0.000126212 1.02 0.887309 0.534785 0.285538 1.71624e-07 3.05451e-09 2398.19 3374.84 -0.0739491 0.482118 0.277757 0.269378 -0.590403 -0.169465 0.441957 -0.268812 -0.173127 1.001 1 4.32127e-218 279.844 2.35845e-215 1.95044 0.999 0.000299994 0.96964 0.611271 0.74677 0.386657 1.95087 123.941 80.9891 18.5479 59.4423 0.00414992 0 -40 10
0.1 2.9007e-09 2.5388e-06 0.033018 0.0329687 0.0120487 1.3185e-06 0.001154 0.0412725 0.000650005 0.0419179 0.845929 101.895 0.247372 0.699958 4.10523 0.0526283 0.0387286 0.961271 0.0198967 0.00422347 0.0191587 0.00406814 0.00510335 0.00584134 0.204134 0.233654 57.946 -87.8929 125.194 15.9967 145.002 0.000152905 0.267087 192.923 0.310703 0.0673877 0.00409486 0.00056158 0.00138251 0.986992 0.991733 -2.97167e-06 -85.6682 0.0929812 31195.8 300.019 0.983522 0.319147 0.793192 0.793187 9.99958 2.98056e-06 1.19221e-05 0.130442 0.966327 0.923722 -0.0132933 4.89119e-06 0.500046 -1.83247e-20 6.74245e-24 -1.8318e-20 0.00139509 0.997818 8.59268e-05 0.152549 2.85169 0.00139509 0.998951 0.62626 0.00103899 0.00187961 0.000859268 0.455656 0.00187962 0.431192 0.000126214 1.02 0.887307 0.534785 0.285536 1.71623e-07 3.05448e-09 2398.17 3373.89 -0.0738784 0.482118 0.277757 0.26932 -0.590414 -0.169465 0.442168 -0.268813 -0.173337 1.002 1 2.62099e-218 279.909 1.43102e-215 1.95073 1 0.000299994 0.969207 0.611362 0.745599 0.386707 1.95115 123.956 80.9996 18.5485 59.4475 0.00414946 0 -40 10
0.101 2.92971e-09 2.5388e-06 0.0331426 0.0330937 0.0120487 1.33168e-06 0.001154 0.0414283 0.000650054 0.0420737 0.845941 101.895 0.247371 0.699968 4.10524 0.052629 0.0387287 0.961271 0.0198966 0.00422348 0.0191586 0.00406815 0.00510336 0.00584135 0.204134 0.233654 57.946 -87.8929 125.198 15.9967 145.002 0.000152862 0.267087 192.923 0.310704 0.0673879 0.00409486 0.000561579 0.00138251 0.986992 0.991733 -2.97165e-06 -85.6682 0.0929811 31195.9 300.019 0.983522 0.319147 0.792969 0.792965 9.99958 2.98055e-06 1.19221e-05 0.130442 0.966381 0.923752 -0.0132933 4.89115e-06 0.500046 -1.83261e-20 6.74292e-24 -1.83194e-20 0.00139509 0.997818 8.59266e-05 0.152548 2.85169 0.00139509 0.998943 0.62639 0.00103899 0.00187961 0.000859266 0.455657 0.00187961 0.431204 0.000126217 1.02 0.887306 0.534785 0.285534 1.71623e-07 3.05445e-09 2398.16 3372.95 -0.0738079 0.482118 0.277757 0.269262 -0.590424 -0.169465 0.442378 -0.268814 -0.173547 1.003 1 1.58971e-218 279.974 8.68285e-216 1.95102 1.001 0.000299994 0.968774 0.611452 0.744431 0.386757 1.95144 123.972 81.0101 18.5492 59.4526 0.004149 0 -40 10
0.102 2.95871e-09 2.5388e-06 0.0332671 0.0332187 0.0120487 1.34487e-06 0.001154 0.0415839 0.000650103 0.0422294 0.845954 101.895 0.24737 0.699978 4.10524 0.0526298 0.0387287 0.961271 0.0198966 0.00422349 0.0191586 0.00406815 0.00510336 0.00584136 0.204135 0.233654 57.9461 -87.8929 125.201 15.9966 145.002 0.000152819 0.267087 192.924 0.310704 0.067388 0.00409485 0.000561578 0.0013825 0.986992 0.991733 -2.97162e-06 -85.6683 0.0929809 31195.9 300.019 0.983522 0.319147 0.792747 0.792742 9.99958 2.98054e-06 1.1922e-05 0.130442 0.966434 0.923782 -0.0132933 4.89112e-06 0.500047 -1.83275e-20 6.74339e-24 -1.83208e-20 0.00139509 0.997818 8.59265e-05 0.152548 2.85169 0.00139509 0.998936 0.626521 0.00103899 0.00187961 0.000859265 0.455657 0.00187961 0.431215 0.000126219 1.02 0.887305 0.534786 0.285533 1.71622e-07 3.05442e-09 2398.14 3372 -0.0737376 0.482118 0.277756 0.269204 -0.590435 -0.169465 0.442588 -0.268815 -0.173755 1.004 1 9.64207e-219 280.039 5.26841e-216 1.95131 1.002 0.000299994 0.968343 0.611542 0.743267 0.386807 1.95173 123.987 81.0205 18.5498 59.4577 0.00414854 0 -40 10
0.103 2.98771e-09 2.5388e-06 0.0333915 0.0333435 0.0120486 1.35805e-06 0.001154 0.0417394 0.000650151 0.0423849 0.845966 101.895 0.247369 0.699988 4.10525 0.0526306 0.0387288 0.961271 0.0198966 0.00422349 0.0191586 0.00406816 0.00510337 0.00584137 0.204135 0.233655 57.9462 -87.8929 125.205 15.9966 145.002 0.000152776 0.267086 192.924 0.310705 0.0673881 0.00409485 0.000561577 0.0013825 0.986992 0.991733 -2.9716e-06 -85.6683 0.0929807 31196 300.019 0.983522 0.319147 0.792526 0.792521 9.99958 2.98053e-06 1.1922e-05 0.130442 0.966488 0.923812 -0.0132933 4.89109e-06 0.500047 -1.83289e-20 6.74385e-24 -1.83221e-20 0.00139508 0.997818 8.59263e-05 0.152548 2.85169 0.00139508 0.998929 0.626651 0.00103899 0.00187961 0.000859263 0.455657 0.00187961 0.431227 0.000126222 1.02 0.887304 0.534786 0.285531 1.71622e-07 3.05439e-09 2398.13 3371.06 -0.0736676 0.482118 0.277756 0.269147 -0.590445 -0.169465 0.442797 -0.268815 -0.173964 1.005 1 5.84821e-219 280.103 3.19666e-216 1.95159 1.003 0.000299994 0.967914 0.611632 0.742107 0.386856 1.95202 124.002 81.0309 18.5504 59.4628 0.00414809 0 -40 10
0.104 3.01671e-09 2.5388e-06 0.0335158 0.0334682 0.0120486 1.37123e-06 0.001154 0.0418948 0.000650199 0.0425404 0.845979 101.895 0.247369 0.699998 4.10525 0.0526314 0.0387288 0.961271 0.0198966 0.0042235 0.0191586 0.00406816 0.00510338 0.00584137 0.204135 0.233655 57.9462 -87.8929 125.209 15.9966 145.002 0.000152733 0.267086 192.924 0.310706 0.0673882 0.00409484 0.000561575 0.00138249 0.986992 0.991733 -2.97157e-06 -85.6683 0.0929806 31196 300.019 0.983522 0.319147 0.792305 0.7923 9.99958 2.98052e-06 1.1922e-05 0.130442 0.966541 0.923842 -0.0132933 4.89106e-06 0.500047 -1.83303e-20 6.74432e-24 -1.83235e-20 0.00139508 0.997818 8.59261e-05 0.152548 2.85168 0.00139508 0.998922 0.626781 0.00103899 0.0018796 0.000859261 0.455658 0.00187961 0.431239 0.000126224 1.02 0.887303 0.534786 0.28553 1.71621e-07 3.05436e-09 2398.11 3370.13 -0.0735978 0.482117 0.277756 0.269089 -0.590456 -0.169465 0.443005 -0.268816 -0.174171 1.006 1 3.54712e-219 280.167 1.9396e-216 1.95188 1.004 0.000299994 0.967486 0.611721 0.74095 0.386906 1.9523 124.018 81.0413 18.551 59.4679 0.00414763 0 -40 10
0.105 3.04571e-09 2.5388e-06 0.03364 0.0335929 0.0120486 1.38441e-06 0.001154 0.04205 0.000650246 0.0426956 0.845992 101.895 0.247368 0.700008 4.10526 0.0526322 0.0387289 0.961271 0.0198966 0.0042235 0.0191586 0.00406817 0.00510339 0.00584138 0.204136 0.233655 57.9463 -87.8929 125.212 15.9965 145.002 0.000152691 0.267086 192.925 0.310707 0.0673883 0.00409484 0.000561574 0.00138249 0.986992 0.991734 -2.97155e-06 -85.6683 0.0929804 31196.1 300.02 0.983522 0.319147 0.792085 0.79208 9.99958 2.98051e-06 1.19219e-05 0.130442 0.966594 0.923871 -0.0132933 4.89103e-06 0.500047 -1.83317e-20 6.74479e-24 -1.83249e-20 0.00139508 0.997818 8.5926e-05 0.152547 2.85168 0.00139508 0.998914 0.626911 0.00103899 0.0018796 0.00085926 0.455658 0.0018796 0.43125 0.000126226 1.02 0.887301 0.534787 0.285528 1.71621e-07 3.05434e-09 2398.1 3369.19 -0.0735282 0.482117 0.277755 0.269032 -0.590466 -0.169465 0.443213 -0.268817 -0.174378 1.007 1 2.15144e-219 280.231 1.17687e-216 1.95217 1.005 0.000299994 0.967059 0.611811 0.739797 0.386955 1.95259 124.033 81.0516 18.5516 59.4729 0.00414718 0 -40 10
0.106 3.07471e-09 2.5388e-06 0.0337641 0.0337174 0.0120486 1.3976e-06 0.001154 0.0422051 0.000650293 0.0428508 0.846005 101.895 0.247367 0.700019 4.10526 0.052633 0.0387289 0.961271 0.0198966 0.00422351 0.0191586 0.00406817 0.0051034 0.00584139 0.204136 0.233656 57.9463 -87.8929 125.216 15.9965 145.002 0.000152649 0.267085 192.925 0.310708 0.0673883 0.00409483 0.000561573 0.00138249 0.986992 0.991734 -2.97153e-06 -85.6683 0.0929802 31196.1 300.02 0.983522 0.319147 0.791866 0.791861 9.99958 2.9805e-06 1.19219e-05 0.130442 0.966647 0.9239 -0.0132933 4.891e-06 0.500048 -1.83331e-20 6.74525e-24 -1.83263e-20 0.00139508 0.997818 8.59258e-05 0.152547 2.85168 0.00139508 0.998907 0.627041 0.00103899 0.0018796 0.000859258 0.455659 0.0018796 0.431262 0.000126229 1.02 0.8873 0.534787 0.285526 1.7162e-07 3.05431e-09 2398.08 3368.26 -0.0734589 0.482117 0.277755 0.268975 -0.590477 -0.169465 0.443419 -0.268818 -0.174584 1.008 1 1.30491e-219 280.295 7.14074e-217 1.95245 1.006 0.000299994 0.966634 0.6119 0.738647 0.387004 1.95287 124.048 81.0619 18.5523 59.478 0.00414673 0 -40 10
0.107 3.10372e-09 2.5388e-06 0.0338881 0.0338418 0.0120486 1.41078e-06 0.001154 0.0423601 0.00065034 0.0430059 0.846018 101.895 0.247366 0.700029 4.10527 0.0526339 0.038729 0.961271 0.0198966 0.00422352 0.0191586 0.00406818 0.00510341 0.0058414 0.204136 0.233656 57.9464 -87.8929 125.22 15.9965 145.002 0.000152607 0.267085 192.925 0.310708 0.0673884 0.00409482 0.000561572 0.00138248 0.986992 0.991734 -2.9715e-06 -85.6683 0.0929801 31196.1 300.02 0.983522 0.319147 0.791647 0.791642 9.99958 2.98049e-06 1.19219e-05 0.130442 0.9667 0.92393 -0.0132933 4.89097e-06 0.500048 -1.83344e-20 6.74572e-24 -1.83277e-20 0.00139508 0.997818 8.59257e-05 0.152547 2.85168 0.00139508 0.9989 0.627171 0.00103899 0.00187959 0.000859257 0.455659 0.0018796 0.431274 0.000126231 1.02 0.887299 0.534787 0.285525 1.7162e-07 3.05428e-09 2398.06 3367.33 -0.0733898 0.482117 0.277754 0.268918 -0.590487 -0.169465 0.443625 -0.268819 -0.174789 1.009 1 7.91469e-220 280.359 4.3327e-217 1.95274 1.007 0.000299994 0.96621 0.611989 0.737501 0.387053 1.95316 124.064 81.0722 18.5529 59.483 0.00414628 0 -40 10
0.108 3.13272e-09 2.5388e-06 0.034012 0.0339661 0.0120486 1.42396e-06 0.001154 0.042515 0.000650386 0.0431608 0.846031 101.895 0.247365 0.70004 4.10528 0.0526347 0.038729 0.961271 0.0198966 0.00422353 0.0191586 0.00406819 0.00510341 0.00584141 0.204137 0.233656 57.9464 -87.8929 125.224 15.9964 145.002 0.000152565 0.267085 192.926 0.310709 0.0673885 0.00409482 0.00056157 0.00138248 0.986992 0.991734 -2.97148e-06 -85.6684 0.0929799 31196.2 300.02 0.983522 0.319147 0.791429 0.791424 9.99958 2.98048e-06 1.19218e-05 0.130442 0.966752 0.923959 -0.0132933 4.89094e-06 0.500048 -1.83358e-20 6.74618e-24 -1.83291e-20 0.00139507 0.997818 8.59255e-05 0.152546 2.85168 0.00139507 0.998893 0.627301 0.001039 0.00187959 0.000859255 0.45566 0.00187959 0.431285 0.000126234 1.02 0.887298 0.534788 0.285523 1.71619e-07 3.05425e-09 2398.05 3366.41 -0.0733209 0.482117 0.277754 0.268861 -0.590497 -0.169465 0.443831 -0.26882 -0.174994 1.01 1 4.8005e-220 280.423 2.62889e-217 1.95302 1.008 0.000299994 0.965788 0.612079 0.736358 0.387103 1.95344 124.079 81.0824 18.5535 59.488 0.00414583 0 -40 10
0.109 3.16172e-09 2.5388e-06 0.0341358 0.0340903 0.0120486 1.43715e-06 0.001154 0.0426698 0.000650432 0.0433156 0.846044 101.895 0.247364 0.700051 4.10528 0.0526356 0.0387291 0.961271 0.0198966 0.00422353 0.0191586 0.00406819 0.00510342 0.00584141 0.204137 0.233657 57.9465 -87.8929 125.227 15.9964 145.002 0.000152523 0.267084 192.926 0.31071 0.0673886 0.00409481 0.000561569 0.00138247 0.986992 0.991734 -2.97146e-06 -85.6684 0.0929798 31196.2 300.02 0.983522 0.319147 0.791212 0.791207 9.99958 2.98047e-06 1.19218e-05 0.130442 0.966805 0.923988 -0.0132933 4.89091e-06 0.500048 -1.83372e-20 6.74665e-24 -1.83304e-20 0.00139507 0.997818 8.59254e-05 0.152546 2.85168 0.00139507 0.998886 0.627431 0.001039 0.00187959 0.000859254 0.45566 0.00187959 0.431297 0.000126236 1.02 0.887297 0.534788 0.285522 1.71619e-07 3.05423e-09 2398.03 3365.48 -0.0732523 0.482117 0.277754 0.268805 -0.590508 -0.169466 0.444036 -0.26882 -0.175198 1.011 1 2.91165e-220 280.486 1.5951e-217 1.95331 1.009 0.000299994 0.965367 0.612168 0.735219 0.387152 1.95373 124.094 81.0926 18.5541 59.493 0.00414538 0 -40 10
0.11 3.19072e-09 2.5388e-06 0.0342595 0.0342145 0.0120485 1.45033e-06 0.001154 0.0428244 0.000650477 0.0434703 0.846057 101.895 0.247364 0.700062 4.10529 0.0526365 0.0387291 0.961271 0.0198966 0.00422354 0.0191586 0.0040682 0.00510343 0.00584142 0.204137 0.233657 57.9466 -87.893 125.231 15.9964 145.002 0.000152481 0.267084 192.926 0.310711 0.0673887 0.00409481 0.000561568 0.00138247 0.986992 0.991734 -2.97143e-06 -85.6684 0.0929796 31196.3 300.021 0.983522 0.319147 0.790996 0.790991 9.99958 2.98046e-06 1.19218e-05 0.130443 0.966857 0.924017 -0.0132933 4.89088e-06 0.500049 -1.83386e-20 6.74711e-24 -1.83318e-20 0.00139507 0.997818 8.59253e-05 0.152546 2.85167 0.00139507 0.998879 0.627561 0.001039 0.00187959 0.000859253 0.45566 0.00187959 0.431308 0.000126239 1.02 0.887296 0.534788 0.28552 1.71618e-07 3.0542e-09 2398.02 3364.57 -0.0731838 0.482117 0.277753 0.268748 -0.590518 -0.169466 0.44424 -0.268821 -0.175402 1.012 1 1.76601e-220 280.549 9.67834e-218 1.95359 1.01 0.000299994 0.964947 0.612257 0.734084 0.387201 1.95401 124.109 81.1028 18.5547 59.498 0.00414494 0 -40 10
0.111 3.21972e-09 2.5388e-06 0.0343831 0.0343385 0.0120485 1.46351e-06 0.001154 0.0429789 0.000650522 0.0436248 0.846071 101.895 0.247363 0.700073 4.1053 0.0526374 0.0387292 0.961271 0.0198966 0.00422355 0.0191586 0.0040682 0.00510344 0.00584143 0.204138 0.233657 57.9466 -87.893 125.235 15.9963 145.002 0.000152439 0.267083 192.926 0.310711 0.0673888 0.0040948 0.000561567 0.00138247 0.986992 0.991734 -2.97141e-06 -85.6684 0.0929795 31196.3 300.021 0.983522 0.319147 0.79078 0.790775 9.99958 2.98046e-06 1.19217e-05 0.130443 0.966909 0.924046 -0.0132933 4.89085e-06 0.500049 -1.83399e-20 6.74758e-24 -1.83332e-20 0.00139507 0.997818 8.59251e-05 0.152546 2.85167 0.00139507 0.998872 0.627691 0.001039 0.00187958 0.000859251 0.455661 0.00187959 0.43132 0.000126241 1.02 0.887295 0.534789 0.285519 1.71618e-07 3.05417e-09 2398 3363.65 -0.0731157 0.482116 0.277753 0.268692 -0.590528 -0.169466 0.444443 -0.268822 -0.175605 1.013 1 1.07114e-220 280.612 5.87238e-218 1.95388 1.011 0.000299994 0.964529 0.612345 0.732952 0.38725 1.95429 124.124 81.1129 18.5553 59.503 0.00414449 0 -40 10
0.112 3.24872e-09 2.5388e-06 0.0345066 0.0344624 0.0120485 1.47669e-06 0.001154 0.0431333 0.000650566 0.0437793 0.846085 101.895 0.247362 0.700084 4.1053 0.0526383 0.0387293 0.961271 0.0198966 0.00422355 0.0191586 0.00406821 0.00510345 0.00584144 0.204138 0.233658 57.9467 -87.893 125.238 15.9963 145.002 0.000152398 0.267083 192.927 0.310712 0.0673889 0.0040948 0.000561566 0.00138246 0.986993 0.991734 -2.97139e-06 -85.6684 0.0929793 31196.3 300.021 0.983522 0.319147 0.790565 0.79056 9.99958 2.98045e-06 1.19217e-05 0.130443 0.966961 0.924075 -0.0132934 4.89082e-06 0.500049 -1.83413e-20 6.74804e-24 -1.83346e-20 0.00139507 0.997818 8.5925e-05 0.152545 2.85167 0.00139507 0.998865 0.62782 0.001039 0.00187958 0.00085925 0.455661 0.00187958 0.431332 0.000126244 1.02 0.887294 0.534789 0.285517 1.71617e-07 3.05415e-09 2397.98 3362.74 -0.0730477 0.482116 0.277753 0.268636 -0.590538 -0.169466 0.444646 -0.268823 -0.175807 1.014 1 6.49677e-221 280.675 3.56309e-218 1.95416 1.012 0.000299994 0.964112 0.612434 0.731823 0.387299 1.95458 124.139 81.123 18.5559 59.5079 0.00414405 0 -40 10
0.113 3.27772e-09 2.5388e-06 0.03463 0.0345862 0.0120485 1.48987e-06 0.001154 0.0432875 0.00065061 0.0439336 0.846098 101.895 0.247361 0.700096 4.10531 0.0526392 0.0387293 0.961271 0.0198965 0.00422356 0.0191586 0.00406821 0.00510346 0.00584145 0.204138 0.233658 57.9467 -87.893 125.242 15.9963 145.002 0.000152357 0.267083 192.927 0.310713 0.067389 0.00409479 0.000561564 0.00138246 0.986993 0.991734 -2.97137e-06 -85.6684 0.0929792 31196.4 300.021 0.983522 0.319147 0.790351 0.790346 9.99958 2.98044e-06 1.19216e-05 0.130443 0.967013 0.924103 -0.0132934 4.89079e-06 0.50005 -1.83427e-20 6.7485e-24 -1.83359e-20 0.00139506 0.997818 8.59248e-05 0.152545 2.85167 0.00139506 0.998858 0.62795 0.001039 0.00187958 0.000859248 0.455662 0.00187958 0.431343 0.000126246 1.02 0.887293 0.534789 0.285516 1.71617e-07 3.05412e-09 2397.97 3361.83 -0.0729799 0.482116 0.277752 0.26858 -0.590549 -0.169466 0.444848 -0.268823 -0.176008 1.015 1 3.94049e-221 280.737 2.16192e-218 1.95444 1.013 0.000299994 0.963697 0.612523 0.730698 0.387347 1.95486 124.155 81.1331 18.5565 59.5129 0.00414361 0 -40 10
0.114 3.30673e-09 2.5388e-06 0.0347533 0.0347099 0.0120485 1.50306e-06 0.001154 0.0434417 0.000650654 0.0440877 0.846112 101.895 0.24736 0.700107 4.10531 0.0526401 0.0387294 0.961271 0.0198965 0.00422357 0.0191585 0.00406822 0.00510347 0.00584146 0.204139 0.233658 57.9468 -87.893 125.245 15.9962 145.002 0.000152316 0.267082 192.927 0.310714 0.0673891 0.00409479 0.000561563 0.00138246 0.986993 0.991735 -2.97134e-06 -85.6685 0.092979 31196.4 300.021 0.983522 0.319147 0.790137 0.790132 9.99958 2.98043e-06 1.19216e-05 0.130443 0.967065 0.924132 -0.0132934 4.89077e-06 0.50005 -1.8344e-20 6.74896e-24 -1.83373e-20 0.00139506 0.997818 8.59247e-05 0.152545 2.85167 0.00139506 0.998852 0.62808 0.00103901 0.00187958 0.000859247 0.455662 0.00187958 0.431355 0.000126249 1.02 0.887292 0.534789 0.285514 1.71616e-07 3.0541e-09 2397.95 3360.92 -0.0729124 0.482116 0.277752 0.268525 -0.590559 -0.169466 0.445049 -0.268824 -0.176209 1.016 1 2.39003e-221 280.8 1.31175e-218 1.95473 1.014 0.000299994 0.963283 0.612611 0.729576 0.387396 1.95514 124.17 81.1431 18.5572 59.5178 0.00414317 0 -40 10
0.115 3.33573e-09 2.5388e-06 0.0348766 0.0348335 0.0120485 1.51624e-06 0.001154 0.0435957 0.000650697 0.0442418 0.846126 101.895 0.247359 0.700119 4.10532 0.052641 0.0387294 0.961271 0.0198965 0.00422358 0.0191585 0.00406823 0.00510348 0.00584147 0.204139 0.233659 57.9468 -87.893 125.249 15.9962 145.002 0.000152275 0.267082 192.928 0.310714 0.0673892 0.00409478 0.000561562 0.00138245 0.986993 0.991735 -2.97132e-06 -85.6685 0.0929789 31196.5 300.022 0.983522 0.319147 0.789924 0.789919 9.99958 2.98042e-06 1.19216e-05 0.130443 0.967116 0.92416 -0.0132934 4.89074e-06 0.50005 -1.83454e-20 6.74942e-24 -1.83386e-20 0.00139506 0.997818 8.59246e-05 0.152544 2.85167 0.00139506 0.998845 0.628209 0.00103901 0.00187957 0.000859246 0.455662 0.00187958 0.431366 0.000126251 1.02 0.887291 0.53479 0.285513 1.71616e-07 3.05407e-09 2397.94 3360.01 -0.0728451 0.482116 0.277751 0.268469 -0.590569 -0.169466 0.44525 -0.268825 -0.176409 1.017 1 1.44963e-221 280.862 7.95909e-219 1.95501 1.015 0.000299994 0.96287 0.612699 0.728458 0.387445 1.95542 124.185 81.1532 18.5578 59.5227 0.00414273 0 -40 10
0.116 3.36473e-09 2.5388e-06 0.0349997 0.034957 0.0120485 1.52942e-06 0.001154 0.0437496 0.00065074 0.0443957 0.84614 101.895 0.247358 0.700131 4.10533 0.052642 0.0387295 0.96127 0.0198965 0.00422358 0.0191585 0.00406823 0.00510349 0.00584148 0.204139 0.233659 57.9469 -87.893 125.253 15.9962 145.002 0.000152234 0.267082 192.928 0.310715 0.0673893 0.00409478 0.000561561 0.00138245 0.986993 0.991735 -2.9713e-06 -85.6685 0.0929787 31196.5 300.022 0.983522 0.319147 0.789712 0.789707 9.99958 2.98041e-06 1.19215e-05 0.130443 0.967168 0.924188 -0.0132934 4.89071e-06 0.500051 -1.83467e-20 6.74988e-24 -1.834e-20 0.00139506 0.997818 8.59244e-05 0.152544 2.85166 0.00139506 0.998838 0.628339 0.00103901 0.00187957 0.000859244 0.455663 0.00187957 0.431378 0.000126254 1.02 0.88729 0.53479 0.285512 1.71616e-07 3.05405e-09 2397.92 3359.11 -0.0727781 0.482116 0.277751 0.268414 -0.590579 -0.169466 0.44545 -0.268825 -0.176609 1.018 1 8.79243e-222 280.924 4.82919e-219 1.95529 1.016 0.000299994 0.962459 0.612788 0.727344 0.387493 1.9557 124.2 81.1631 18.5584 59.5276 0.00414229 0 -40 10
0.117 3.39373e-09 2.5388e-06 0.0351227 0.0350804 0.0120485 1.5426e-06 0.001154 0.0439033 0.000650783 0.0445495 0.846154 101.895 0.247357 0.700143 4.10533 0.0526429 0.0387296 0.96127 0.0198965 0.00422359 0.0191585 0.00406824 0.0051035 0.00584149 0.20414 0.233659 57.947 -87.893 125.256 15.9961 145.002 0.000152193 0.267082 192.928 0.310716 0.0673894 0.00409477 0.00056156 0.00138244 0.986993 0.991735 -2.97128e-06 -85.6685 0.0929786 31196.5 300.022 0.983522 0.319147 0.7895 0.789496 9.99958 2.98041e-06 1.19215e-05 0.130443 0.967219 0.924217 -0.0132934 4.89069e-06 0.500051 -1.83481e-20 6.75034e-24 -1.83413e-20 0.00139506 0.997818 8.59243e-05 0.152544 2.85166 0.00139506 0.998831 0.628469 0.00103901 0.00187957 0.000859243 0.455663 0.00187957 0.431389 0.000126256 1.02 0.887289 0.53479 0.28551 1.71615e-07 3.05402e-09 2397.91 3358.21 -0.0727112 0.482116 0.277751 0.268359 -0.590589 -0.169466 0.445649 -0.268826 -0.176808 1.019 1 5.33288e-222 280.986 2.93012e-219 1.95557 1.017 0.000299994 0.962049 0.612876 0.726233 0.387542 1.95599 124.215 81.1731 18.559 59.5324 0.00414186 0 -40 10
0.118 3.42273e-09 2.5388e-06 0.0352456 0.0352037 0.0120484 1.55579e-06 0.001154 0.044057 0.000650825 0.0447032 0.846169 101.895 0.247356 0.700156 4.10534 0.0526439 0.0387296 0.96127 0.0198965 0.0042236 0.0191585 0.00406825 0.0051035 0.00584149 0.20414 0.23366 57.947 -87.893 125.26 15.9961 145.002 0.000152152 0.267081 192.928 0.310717 0.0673895 0.00409477 0.000561559 0.00138244 0.986993 0.991735 -2.97126e-06 -85.6685 0.0929784 31196.6 300.022 0.983522 0.319147 0.789289 0.789285 9.99958 2.9804e-06 1.19215e-05 0.130443 0.96727 0.924245 -0.0132934 4.89066e-06 0.500051 -1.83494e-20 6.7508e-24 -1.83427e-20 0.00139505 0.997818 8.59242e-05 0.152544 2.85166 0.00139505 0.998825 0.628598 0.00103902 0.00187957 0.000859242 0.455663 0.00187957 0.431401 0.000126259 1.02 0.887288 0.534791 0.285509 1.71615e-07 3.054e-09 2397.89 3357.32 -0.0726446 0.482116 0.27775 0.268304 -0.590599 -0.169466 0.445848 -0.268827 -0.177006 1.02 1 3.23455e-222 281.047 1.77785e-219 1.95585 1.018 0.000299994 0.96164 0.612964 0.725125 0.38759 1.95627 124.23 81.183 18.5595 59.5373 0.00414142 0 -40 10
0.119 3.45173e-09 2.5388e-06 0.0353684 0.0353269 0.0120484 1.56897e-06 0.001154 0.0442105 0.000650866 0.0448568 0.846183 101.895 0.247355 0.700168 4.10535 0.0526449 0.0387297 0.96127 0.0198965 0.00422361 0.0191585 0.00406825 0.00510351 0.0058415 0.204141 0.23366 57.9471 -87.893 125.263 15.9961 145.002 0.000152112 0.267081 192.929 0.310717 0.0673895 0.00409476 0.000561558 0.00138244 0.986993 0.991735 -2.97124e-06 -85.6685 0.0929783 31196.6 300.022 0.983522 0.319147 0.789079 0.789075 9.99958 2.98039e-06 1.19215e-05 0.130443 0.967321 0.924273 -0.0132934 4.89064e-06 0.500052 -1.83508e-20 6.75126e-24 -1.8344e-20 0.00139505 0.997818 8.5924e-05 0.152543 2.85166 0.00139505 0.998818 0.628728 0.00103902 0.00187956 0.00085924 0.455664 0.00187957 0.431413 0.000126261 1.02 0.887287 0.534791 0.285507 1.71614e-07 3.05398e-09 2397.87 3356.43 -0.0725782 0.482115 0.27775 0.268249 -0.590609 -0.169466 0.446046 -0.268827 -0.177203 1.021 1 1.96186e-222 281.109 1.07871e-219 1.95613 1.019 0.000299994 0.961233 0.613051 0.724021 0.387639 1.95655 124.245 81.1929 18.5601 59.5421 0.00414099 0 -40 10
0.12 3.48073e-09 2.5388e-06 0.0354911 0.03545 0.0120484 1.58215e-06 0.001154 0.0443639 0.000650908 0.0450102 0.846197 101.895 0.247354 0.700181 4.10536 0.0526459 0.0387298 0.96127 0.0198965 0.00422362 0.0191585 0.00406826 0.00510352 0.00584151 0.204141 0.233661 57.9471 -87.893 125.267 15.996 145.002 0.000152071 0.267081 192.929 0.310718 0.0673896 0.00409476 0.000561557 0.00138243 0.986993 0.991735 -2.97122e-06 -85.6686 0.0929781 31196.6 300.023 0.983522 0.319147 0.78887 0.788865 9.99958 2.98038e-06 1.19214e-05 0.130443 0.967371 0.924301 -0.0132934 4.89061e-06 0.500052 -1.83521e-20 6.75172e-24 -1.83454e-20 0.00139505 0.997818 8.59239e-05 0.152543 2.85166 0.00139505 0.998812 0.628857 0.00103902 0.00187956 0.000859239 0.455664 0.00187956 0.431424 0.000126264 1.02 0.887286 0.534791 0.285506 1.71614e-07 3.05395e-09 2397.86 3355.54 -0.072512 0.482115 0.27775 0.268195 -0.590619 -0.169466 0.446243 -0.268828 -0.1774 1.022 1 1.18993e-222 281.17 6.54509e-220 1.95641 1.02 0.000299994 0.960827 0.613139 0.72292 0.387687 1.95683 124.26 81.2028 18.5607 59.547 0.00414056 0 -40 10
0.121 3.50973e-09 2.5388e-06 0.0356137 0.035573 0.0120484 1.59533e-06 0.001154 0.0445172 0.000650949 0.0451635 0.846212 101.895 0.247353 0.700193 4.10536 0.0526469 0.0387298 0.96127 0.0198965 0.00422362 0.0191585 0.00406827 0.00510353 0.00584152 0.204141 0.233661 57.9472 -87.893 125.27 15.996 145.002 0.000152031 0.26708 192.929 0.310719 0.0673897 0.00409475 0.000561556 0.00138243 0.986993 0.991735 -2.9712e-06 -85.6686 0.092978 31196.7 300.023 0.983522 0.319147 0.788661 0.788656 9.99958 2.98037e-06 1.19214e-05 0.130443 0.967422 0.924328 -0.0132934 4.89058e-06 0.500052 -1.83535e-20 6.75218e-24 -1.83467e-20 0.00139505 0.997818 8.59238e-05 0.152543 2.85166 0.00139505 0.998805 0.628986 0.00103903 0.00187956 0.000859238 0.455665 0.00187956 0.431436 0.000126267 1.02 0.887285 0.534791 0.285505 1.71613e-07 3.05393e-09 2397.84 3354.65 -0.0724461 0.482115 0.277749 0.26814 -0.590629 -0.169467 0.44644 -0.268828 -0.177597 1.023 1 7.21726e-223 281.231 3.97123e-220 1.95669 1.021 0.000299994 0.960423 0.613227 0.721822 0.387735 1.95711 124.275 81.2126 18.5613 59.5518 0.00414013 0 -40 10
0.122 3.53873e-09 2.5388e-06 0.0357363 0.0356958 0.0120484 1.60851e-06 0.001154 0.0446703 0.000650989 0.0453167 0.846227 101.895 0.247352 0.700206 4.10537 0.0526479 0.0387299 0.96127 0.0198965 0.00422363 0.0191585 0.00406827 0.00510354 0.00584153 0.204142 0.233661 57.9472 -87.893 125.274 15.996 145.003 0.000151991 0.26708 192.929 0.310719 0.0673898 0.00409475 0.000561554 0.00138243 0.986993 0.991735 -2.97117e-06 -85.6686 0.0929779 31196.7 300.023 0.983522 0.319147 0.788453 0.788448 9.99958 2.98037e-06 1.19214e-05 0.130443 0.967472 0.924356 -0.0132934 4.89056e-06 0.500053 -1.83548e-20 6.75264e-24 -1.83481e-20 0.00139505 0.997818 8.59236e-05 0.152543 2.85165 0.00139505 0.998799 0.629116 0.00103903 0.00187956 0.000859236 0.455665 0.00187956 0.431447 0.000126269 1.02 0.887284 0.534792 0.285504 1.71613e-07 3.05391e-09 2397.83 3353.77 -0.0723804 0.482115 0.277749 0.268086 -0.590639 -0.169467 0.446636 -0.268829 -0.177792 1.024 1 4.37749e-223 281.292 2.40954e-220 1.95697 1.022 0.000299994 0.960019 0.613314 0.720728 0.387783 1.95739 124.29 81.2224 18.5619 59.5566 0.0041397 0 -40 10
0.123 3.56773e-09 2.5388e-06 0.0358587 0.0358186 0.0120484 1.6217e-06 0.001154 0.0448234 0.00065103 0.0454698 0.846242 101.895 0.247351 0.700219 4.10538 0.0526489 0.03873 0.96127 0.0198964 0.00422364 0.0191585 0.00406828 0.00510356 0.00584154 0.204142 0.233662 57.9473 -87.893 125.277 15.9959 145.003 0.000151951 0.26708 192.93 0.31072 0.0673899 0.00409474 0.000561553 0.00138242 0.986993 0.991735 -2.97115e-06 -85.6686 0.0929777 31196.7 300.023 0.983523 0.319147 0.788246 0.788241 9.99958 2.98036e-06 1.19213e-05 0.130444 0.967522 0.924384 -0.0132934 4.89054e-06 0.500053 -1.83562e-20 6.75309e-24 -1.83494e-20 0.00139505 0.997818 8.59235e-05 0.152542 2.85165 0.00139505 0.998792 0.629245 0.00103903 0.00187955 0.000859235 0.455665 0.00187956 0.431459 0.000126272 1.02 0.887283 0.534792 0.285502 1.71613e-07 3.05388e-09 2397.81 3352.88 -0.0723148 0.482115 0.277749 0.268032 -0.590649 -0.169467 0.446831 -0.268829 -0.177987 1.025 1 2.65508e-223 281.352 1.46198e-220 1.95725 1.023 0.000299994 0.959618 0.613401 0.719637 0.387832 1.95766 124.305 81.2322 18.5625 59.5614 0.00413927 0 -40 10
0.124 3.59673e-09 2.5388e-06 0.035981 0.0359413 0.0120484 1.63488e-06 0.001154 0.0449763 0.000651069 0.0456227 0.846257 101.895 0.24735 0.700233 4.10539 0.05265 0.03873 0.96127 0.0198964 0.00422365 0.0191584 0.00406829 0.00510357 0.00584155 0.204143 0.233662 57.9474 -87.893 125.281 15.9959 145.003 0.000151911 0.267079 192.93 0.310721 0.06739 0.00409474 0.000561552 0.00138242 0.986993 0.991735 -2.97113e-06 -85.6686 0.0929776 31196.8 300.023 0.983523 0.319147 0.788039 0.788034 9.99958 2.98035e-06 1.19213e-05 0.130444 0.967572 0.924411 -0.0132934 4.89051e-06 0.500053 -1.83575e-20 6.75355e-24 -1.83507e-20 0.00139504 0.997818 8.59234e-05 0.152542 2.85165 0.00139504 0.998786 0.629374 0.00103904 0.00187955 0.000859234 0.455666 0.00187955 0.43147 0.000126274 1.02 0.887282 0.534792 0.285501 1.71612e-07 3.05386e-09 2397.8 3352.01 -0.0722495 0.482115 0.277748 0.267978 -0.590659 -0.169467 0.447026 -0.26883 -0.178182 1.026 1 1.61039e-223 281.413 8.87054e-221 1.95753 1.024 0.000299994 0.959217 0.613489 0.71855 0.38788 1.95794 124.319 81.2419 18.5631 59.5661 0.00413885 0 -40 10
0.125 3.62573e-09 2.5388e-06 0.0361032 0.0360639 0.0120484 1.64806e-06 0.001154 0.045129 0.000651109 0.0457756 0.846272 101.895 0.247349 0.700246 4.10539 0.052651 0.0387301 0.96127 0.0198964 0.00422366 0.0191584 0.00406829 0.00510358 0.00584156 0.204143 0.233663 57.9474 -87.893 125.284 15.9959 145.003 0.000151871 0.267079 192.93 0.310721 0.06739 0.00409473 0.000561551 0.00138242 0.986993 0.991735 -2.97112e-06 -85.6686 0.0929775 31196.8 300.024 0.983523 0.319147 0.787833 0.787828 9.99958 2.98034e-06 1.19213e-05 0.130444 0.967622 0.924438 -0.0132934 4.89049e-06 0.500054 -1.83588e-20 6.75401e-24 -1.83521e-20 0.00139504 0.997818 8.59233e-05 0.152542 2.85165 0.00139504 0.99878 0.629503 0.00103904 0.00187955 0.000859233 0.455666 0.00187955 0.431482 0.000126277 1.02 0.887281 0.534792 0.2855 1.71612e-07 3.05384e-09 2397.78 3351.13 -0.0721844 0.482115 0.277748 0.267924 -0.590668 -0.169467 0.44722 -0.26883 -0.178375 1.027 1 9.7675e-224 281.473 5.38217e-221 1.95781 1.025 0.000299994 0.958818 0.613576 0.717466 0.387928 1.95822 124.334 81.2516 18.5637 59.5709 0.00413843 0 -40 10
0.126 3.65473e-09 2.5388e-06 0.0362254 0.0361864 0.0120483 1.66124e-06 0.001154 0.0452817 0.000651148 0.0459283 0.846287 101.895 0.247348 0.70026 4.1054 0.0526521 0.0387302 0.96127 0.0198964 0.00422367 0.0191584 0.0040683 0.00510359 0.00584158 0.204143 0.233663 57.9475 -87.893 125.288 15.9958 145.003 0.000151832 0.267079 192.93 0.310722 0.0673901 0.00409473 0.00056155 0.00138241 0.986993 0.991735 -2.9711e-06 -85.6686 0.0929773 31196.9 300.024 0.983523 0.319147 0.787628 0.787623 9.99958 2.98033e-06 1.19212e-05 0.130444 0.967672 0.924466 -0.0132934 4.89046e-06 0.500054 -1.83601e-20 6.75446e-24 -1.83534e-20 0.00139504 0.997818 8.59231e-05 0.152542 2.85165 0.00139504 0.998773 0.629632 0.00103904 0.00187955 0.000859231 0.455666 0.00187955 0.431493 0.00012628 1.02 0.88728 0.534793 0.285499 1.71611e-07 3.05382e-09 2397.76 3350.26 -0.0721196 0.482115 0.277747 0.267871 -0.590678 -0.169467 0.447414 -0.268831 -0.178568 1.028 1 5.92429e-224 281.533 3.26561e-221 1.95809 1.026 0.000299994 0.95842 0.613663 0.716385 0.387975 1.9585 124.349 81.2613 18.5642 59.5756 0.004138 0 -40 10
0.127 3.68373e-09 2.5388e-06 0.0363474 0.0363088 0.0120483 1.67442e-06 0.001154 0.0454342 0.000651187 0.0460808 0.846302 101.895 0.247347 0.700273 4.10541 0.0526532 0.0387303 0.96127 0.0198964 0.00422368 0.0191584 0.00406831 0.0051036 0.00584159 0.204144 0.233663 57.9475 -87.893 125.291 15.9958 145.003 0.000151792 0.267079 192.931 0.310723 0.0673902 0.00409472 0.000561549 0.00138241 0.986993 0.991735 -2.97108e-06 -85.6687 0.0929772 31196.9 300.024 0.983523 0.319147 0.787423 0.787418 9.99958 2.98033e-06 1.19212e-05 0.130444 0.967722 0.924493 -0.0132934 4.89044e-06 0.500054 -1.83615e-20 6.75492e-24 -1.83547e-20 0.00139504 0.997818 8.5923e-05 0.152542 2.85165 0.00139504 0.998767 0.629762 0.00103905 0.00187955 0.00085923 0.455667 0.00187955 0.431505 0.000126282 1.02 0.887279 0.534793 0.285497 1.71611e-07 3.0538e-09 2397.75 3349.39 -0.0720549 0.482115 0.277747 0.267817 -0.590688 -0.169467 0.447606 -0.268831 -0.178761 1.029 1 3.59326e-224 281.593 1.9814e-221 1.95837 1.027 0.000299994 0.958024 0.613749 0.715308 0.388023 1.95877 124.364 81.271 18.5648 59.5803 0.00413758 0 -40 10
0.128 3.71273e-09 2.5388e-06 0.0364693 0.036431 0.0120483 1.6876e-06 0.001154 0.0455867 0.000651225 0.0462333 0.846317 101.895 0.247346 0.700287 4.10542 0.0526543 0.0387303 0.96127 0.0198964 0.00422368 0.0191584 0.00406832 0.00510361 0.0058416 0.204144 0.233664 57.9476 -87.893 125.295 15.9958 145.003 0.000151753 0.267078 192.931 0.310723 0.0673903 0.00409472 0.000561548 0.00138241 0.986993 0.991735 -2.97106e-06 -85.6687 0.0929771 31196.9 300.024 0.983523 0.319147 0.787219 0.787214 9.99958 2.98032e-06 1.19212e-05 0.130444 0.967771 0.92452 -0.0132934 4.89042e-06 0.500055 -1.83628e-20 6.75537e-24 -1.8356e-20 0.00139504 0.997818 8.59229e-05 0.152541 2.85165 0.00139504 0.998761 0.629891 0.00103905 0.00187954 0.000859229 0.455667 0.00187955 0.431516 0.000126285 1.02 0.887279 0.534793 0.285496 1.7161e-07 3.05378e-09 2397.73 3348.52 -0.0719905 0.482114 0.277747 0.267764 -0.590698 -0.169467 0.447799 -0.268832 -0.178953 1.03 1 2.17942e-224 281.653 1.2022e-221 1.95864 1.028 0.000299994 0.957629 0.613836 0.714234 0.388071 1.95905 124.379 81.2806 18.5654 59.585 0.00413716 0 -40 10
0.129 3.74173e-09 2.5388e-06 0.0365912 0.0365532 0.0120483 1.70079e-06 0.001154 0.045739 0.000651264 0.0463856 0.846333 101.895 0.247345 0.700301 4.10542 0.0526554 0.0387304 0.96127 0.0198964 0.00422369 0.0191584 0.00406832 0.00510362 0.00584161 0.204145 0.233664 57.9476 -87.893 125.298 15.9957 145.003 0.000151714 0.267078 192.931 0.310724 0.0673904 0.00409471 0.000561547 0.0013824 0.986993 0.991735 -2.97104e-06 -85.6687 0.0929769 31197 300.025 0.983523 0.319147 0.787015 0.787011 9.99958 2.98031e-06 1.19211e-05 0.130444 0.96782 0.924547 -0.0132934 4.8904e-06 0.500055 -1.83641e-20 6.75582e-24 -1.83574e-20 0.00139503 0.997818 8.59228e-05 0.152541 2.85165 0.00139503 0.998755 0.63002 0.00103906 0.00187954 0.000859228 0.455667 0.00187954 0.431528 0.000126288 1.02 0.887278 0.534793 0.285495 1.7161e-07 3.05375e-09 2397.72 3347.66 -0.0719263 0.482114 0.277746 0.267711 -0.590707 -0.169467 0.44799 -0.268832 -0.179144 1.031 1 1.32189e-224 281.712 7.29431e-222 1.95892 1.029 0.000299994 0.957235 0.613923 0.713163 0.388119 1.95933 124.394 81.2902 18.566 59.5897 0.00413674 0 -40 10
0.13 3.77073e-09 2.5388e-06 0.0367129 0.0366753 0.0120483 1.71397e-06 0.001154 0.0458911 0.000651301 0.0465378 0.846348 101.895 0.247343 0.700315 4.10543 0.0526565 0.0387305 0.96127 0.0198964 0.0042237 0.0191584 0.00406833 0.00510363 0.00584162 0.204145 0.233665 57.9477 -87.893 125.302 15.9957 145.003 0.000151675 0.267078 192.931 0.310725 0.0673904 0.00409471 0.000561546 0.0013824 0.986993 0.991735 -2.97102e-06 -85.6687 0.0929768 31197 300.025 0.983523 0.319147 0.786813 0.786808 9.99958 2.98031e-06 1.19211e-05 0.130444 0.96787 0.924573 -0.0132934 4.89037e-06 0.500055 -1.83654e-20 6.75628e-24 -1.83587e-20 0.00139503 0.997818 8.59227e-05 0.152541 2.85164 0.00139503 0.998749 0.630149 0.00103906 0.00187954 0.000859227 0.455668 0.00187954 0.431539 0.00012629 1.02 0.887277 0.534794 0.285494 1.7161e-07 3.05373e-09 2397.7 3346.8 -0.0718623 0.482114 0.277746 0.267658 -0.590717 -0.169467 0.448181 -0.268833 -0.179335 1.032 1 8.01765e-225 281.772 4.42578e-222 1.9592 1.03 0.000299994 0.956842 0.614009 0.712095 0.388166 1.9596 124.408 81.2997 18.5665 59.5944 0.00413633 0 -40 10
0.131 3.79973e-09 2.5388e-06 0.0368345 0.0367973 0.0120483 1.72715e-06 0.001154 0.0460432 0.000651339 0.0466899 0.846364 101.895 0.247342 0.70033 4.10544 0.0526577 0.0387306 0.961269 0.0198964 0.00422371 0.0191584 0.00406834 0.00510364 0.00584163 0.204146 0.233665 57.9478 -87.893 125.305 15.9957 145.003 0.000151636 0.267077 192.932 0.310725 0.0673905 0.00409471 0.000561545 0.0013824 0.986993 0.991736 -2.971e-06 -85.6687 0.0929767 31197 300.025 0.983523 0.319147 0.786611 0.786606 9.99958 2.9803e-06 1.19211e-05 0.130444 0.967918 0.9246 -0.0132934 4.89035e-06 0.500056 -1.83667e-20 6.75673e-24 -1.836e-20 0.00139503 0.997818 8.59225e-05 0.152541 2.85164 0.00139503 0.998743 0.630277 0.00103906 0.00187954 0.000859225 0.455668 0.00187954 0.431551 0.000126293 1.02 0.887276 0.534794 0.285493 1.71609e-07 3.05371e-09 2397.68 3345.94 -0.0717985 0.482114 0.277746 0.267605 -0.590727 -0.169467 0.448371 -0.268833 -0.179525 1.033 1 4.86295e-225 281.831 2.68531e-222 1.95947 1.031 0.000299994 0.956451 0.614096 0.711031 0.388214 1.95988 124.423 81.3093 18.5671 59.5991 0.00413591 0 -40 10
0.132 3.82873e-09 2.5388e-06 0.0369561 0.0369191 0.0120483 1.74033e-06 0.001154 0.0461951 0.000651376 0.0468419 0.84638 101.895 0.247341 0.700344 4.10545 0.0526588 0.0387307 0.961269 0.0198963 0.00422372 0.0191584 0.00406835 0.00510366 0.00584164 0.204146 0.233666 57.9478 -87.893 125.309 15.9956 145.003 0.000151597 0.267077 192.932 0.310726 0.0673906 0.0040947 0.000561544 0.00138239 0.986993 0.991736 -2.97098e-06 -85.6687 0.0929766 31197 300.025 0.983523 0.319147 0.786409 0.786405 9.99958 2.98029e-06 1.19211e-05 0.130444 0.967967 0.924627 -0.0132934 4.89033e-06 0.500056 -1.83681e-20 6.75718e-24 -1.83613e-20 0.00139503 0.997818 8.59224e-05 0.15254 2.85164 0.00139503 0.998737 0.630406 0.00103907 0.00187953 0.000859224 0.455668 0.00187954 0.431562 0.000126295 1.02 0.887275 0.534794 0.285492 1.71609e-07 3.05369e-09 2397.67 3345.08 -0.0717349 0.482114 0.277745 0.267553 -0.590736 -0.169468 0.448561 -0.268834 -0.179714 1.034 1 2.94953e-225 281.89 1.62929e-222 1.95975 1.032 0.000299994 0.956061 0.614182 0.70997 0.388261 1.96015 124.438 81.3188 18.5677 59.6037 0.0041355 0 -40 10
0.133 3.85773e-09 2.5388e-06 0.0370775 0.0370409 0.0120482 1.75351e-06 0.001154 0.0463469 0.000651413 0.0469937 0.846396 101.895 0.24734 0.700359 4.10546 0.05266 0.0387307 0.961269 0.0198963 0.00422373 0.0191583 0.00406835 0.00510367 0.00584165 0.204147 0.233666 57.9479 -87.893 125.312 15.9956 145.003 0.000151558 0.267077 192.932 0.310726 0.0673907 0.0040947 0.000561543 0.00138239 0.986993 0.991736 -2.97097e-06 -85.6687 0.0929764 31197.1 300.026 0.983523 0.319147 0.786209 0.786204 9.99958 2.98028e-06 1.1921e-05 0.130444 0.968016 0.924653 -0.0132934 4.89031e-06 0.500057 -1.83694e-20 6.75763e-24 -1.83626e-20 0.00139503 0.997818 8.59223e-05 0.15254 2.85164 0.00139503 0.998731 0.630535 0.00103907 0.00187953 0.000859223 0.455669 0.00187953 0.431574 0.000126298 1.02 0.887275 0.534794 0.285491 1.71609e-07 3.05367e-09 2397.65 3344.23 -0.0716715 0.482114 0.277745 0.2675 -0.590746 -0.169468 0.44875 -0.268834 -0.179903 1.035 1 1.78898e-225 281.949 9.88562e-223 1.96003 1.033 0.000299994 0.955672 0.614268 0.708912 0.388309 1.96043 124.453 81.3282 18.5683 59.6083 0.00413508 0 -40 10
0.134 3.88672e-09 2.5388e-06 0.0371989 0.0371626 0.0120482 1.76669e-06 0.001154 0.0464986 0.000651449 0.0471455 0.846412 101.895 0.247339 0.700374 4.10547 0.0526612 0.0387308 0.961269 0.0198963 0.00422374 0.0191583 0.00406836 0.00510368 0.00584166 0.204147 0.233667 57.9479 -87.893 125.315 15.9956 145.003 0.00015152 0.267077 192.932 0.310727 0.0673907 0.00409469 0.000561543 0.00138239 0.986993 0.991736 -2.97095e-06 -85.6688 0.0929763 31197.1 300.026 0.983523 0.319147 0.786009 0.786004 9.99958 2.98028e-06 1.1921e-05 0.130445 0.968064 0.92468 -0.0132934 4.89029e-06 0.500057 -1.83707e-20 6.75808e-24 -1.83639e-20 0.00139503 0.997818 8.59222e-05 0.15254 2.85164 0.00139503 0.998725 0.630664 0.00103908 0.00187953 0.000859222 0.455669 0.00187953 0.431585 0.000126301 1.02 0.887274 0.534794 0.285489 1.71608e-07 3.05365e-09 2397.64 3343.38 -0.0716084 0.482114 0.277745 0.267448 -0.590755 -0.169468 0.448938 -0.268834 -0.180091 1.036 1 1.08507e-225 282.008 5.99802e-223 1.9603 1.034 0.000299994 0.955285 0.614354 0.707858 0.388356 1.9607 124.467 81.3377 18.5688 59.613 0.00413467 0 -40 10
0.135 3.91572e-09 2.5388e-06 0.0373201 0.0372841 0.0120482 1.77987e-06 0.001154 0.0466502 0.000651485 0.0472971 0.846428 101.895 0.247338 0.700389 4.10548 0.0526623 0.0387309 0.961269 0.0198963 0.00422375 0.0191583 0.00406837 0.00510369 0.00584168 0.204148 0.233667 57.948 -87.893 125.319 15.9955 145.003 0.000151481 0.267076 192.933 0.310728 0.0673908 0.00409469 0.000561542 0.00138239 0.986994 0.991736 -2.97093e-06 -85.6688 0.0929762 31197.1 300.026 0.983523 0.319147 0.785809 0.785805 9.99958 2.98027e-06 1.1921e-05 0.130445 0.968113 0.924706 -0.0132934 4.89027e-06 0.500057 -1.8372e-20 6.75853e-24 -1.83652e-20 0.00139502 0.997818 8.59221e-05 0.15254 2.85164 0.00139503 0.998719 0.630793 0.00103908 0.00187953 0.000859221 0.455669 0.00187953 0.431597 0.000126304 1.02 0.887273 0.534795 0.285488 1.71608e-07 3.05364e-09 2397.62 3342.53 -0.0715454 0.482114 0.277744 0.267396 -0.590765 -0.169468 0.449126 -0.268835 -0.180278 1.037 1 6.58129e-226 282.066 3.63925e-223 1.96058 1.035 0.000299994 0.954899 0.61444 0.706807 0.388403 1.96098 124.482 81.3471 18.5694 59.6176 0.00413426 0 -40 10
0.136 3.94472e-09 2.5388e-06 0.0374413 0.0374056 0.0120482 1.79306e-06 0.001154 0.0468016 0.000651521 0.0474485 0.846444 101.895 0.247336 0.700404 4.10548 0.0526635 0.038731 0.961269 0.0198963 0.00422376 0.0191583 0.00406838 0.0051037 0.00584169 0.204148 0.233668 57.948 -87.8931 125.322 15.9955 145.003 0.000151443 0.267076 192.933 0.310728 0.0673909 0.00409468 0.000561541 0.00138238 0.986994 0.991736 -2.97091e-06 -85.6688 0.0929761 31197.2 300.027 0.983523 0.319147 0.78561 0.785606 9.99958 2.98026e-06 1.19209e-05 0.130445 0.968161 0.924732 -0.0132934 4.89025e-06 0.500058 -1.83733e-20 6.75898e-24 -1.83665e-20 0.00139502 0.997818 8.5922e-05 0.15254 2.85164 0.00139502 0.998713 0.630921 0.00103909 0.00187953 0.00085922 0.45567 0.00187953 0.431608 0.000126306 1.02 0.887272 0.534795 0.285487 1.71607e-07 3.05362e-09 2397.61 3341.69 -0.0714827 0.482114 0.277744 0.267344 -0.590774 -0.169468 0.449313 -0.268835 -0.180465 1.038 1 3.99176e-226 282.124 2.20808e-223 1.96085 1.036 0.000299994 0.954514 0.614526 0.705759 0.388451 1.96125 124.497 81.3565 18.5699 59.6222 0.00413385 0 -40 10
0.137 3.97372e-09 2.5388e-06 0.0375623 0.037527 0.0120482 1.80624e-06 0.001154 0.0469529 0.000651557 0.0475999 0.846461 101.895 0.247335 0.700419 4.10549 0.0526647 0.0387311 0.961269 0.0198963 0.00422377 0.0191583 0.00406839 0.00510372 0.0058417 0.204149 0.233668 57.9481 -87.8931 125.325 15.9954 145.003 0.000151405 0.267076 192.933 0.310729 0.0673909 0.00409468 0.00056154 0.00138238 0.986994 0.991736 -2.9709e-06 -85.6688 0.0929759 31197.2 300.027 0.983523 0.319147 0.785412 0.785408 9.99958 2.98026e-06 1.19209e-05 0.130445 0.968209 0.924758 -0.0132934 4.89023e-06 0.500058 -1.83746e-20 6.75943e-24 -1.83678e-20 0.00139502 0.997818 8.59219e-05 0.152539 2.85163 0.00139502 0.998707 0.63105 0.00103909 0.00187952 0.000859219 0.45567 0.00187953 0.43162 0.000126309 1.02 0.887271 0.534795 0.285486 1.71607e-07 3.0536e-09 2397.59 3340.85 -0.0714201 0.482113 0.277744 0.267292 -0.590784 -0.169468 0.449499 -0.268835 -0.180651 1.039 1 2.42112e-226 282.182 1.33973e-223 1.96112 1.037 0.000299994 0.954131 0.614611 0.704714 0.388498 1.96153 124.511 81.3658 18.5705 59.6267 0.00413345 0 -40 10
0.138 4.00272e-09 2.5388e-06 0.0376833 0.0376482 0.0120482 1.81942e-06 0.001154 0.0471041 0.000651592 0.0477511 0.846477 101.894 0.247334 0.700435 4.1055 0.052666 0.0387312 0.961269 0.0198963 0.00422378 0.0191583 0.00406839 0.00510373 0.00584171 0.204149 0.233669 57.9482 -87.8931 125.329 15.9954 145.003 0.000151367 0.267076 192.933 0.310729 0.067391 0.00409468 0.000561539 0.00138238 0.986994 0.991736 -2.97088e-06 -85.6688 0.0929758 31197.2 300.027 0.983523 0.319147 0.785215 0.78521 9.99958 2.98025e-06 1.19209e-05 0.130445 0.968257 0.924784 -0.0132934 4.89021e-06 0.500059 -1.83759e-20 6.75988e-24 -1.83691e-20 0.00139502 0.997818 8.59218e-05 0.152539 2.85163 0.00139502 0.998701 0.631179 0.0010391 0.00187952 0.000859218 0.45567 0.00187952 0.431631 0.000126312 1.02 0.887271 0.534795 0.285485 1.71607e-07 3.05358e-09 2397.57 3340.01 -0.0713578 0.482113 0.277743 0.267241 -0.590793 -0.169468 0.449685 -0.268836 -0.180837 1.04 1 1.46848e-226 282.24 8.12869e-224 1.9614 1.038 0.000299994 0.953748 0.614697 0.703672 0.388545 1.9618 124.526 81.3752 18.5711 59.6313 0.00413304 0 -40 10
0.139 4.03172e-09 2.5388e-06 0.0378042 0.0377694 0.0120482 1.8326e-06 0.001154 0.0472552 0.000651627 0.0479022 0.846494 101.894 0.247333 0.70045 4.10551 0.0526672 0.0387312 0.961269 0.0198963 0.00422379 0.0191583 0.0040684 0.00510374 0.00584173 0.20415 0.233669 57.9482 -87.8931 125.332 15.9954 145.003 0.000151329 0.267075 192.933 0.31073 0.0673911 0.00409467 0.000561538 0.00138237 0.986994 0.991736 -2.97086e-06 -85.6688 0.0929757 31197.3 300.027 0.983523 0.319147 0.785018 0.785013 9.99958 2.98024e-06 1.19209e-05 0.130445 0.968305 0.92481 -0.0132934 4.89019e-06 0.500059 -1.83772e-20 6.76033e-24 -1.83704e-20 0.00139502 0.997818 8.59217e-05 0.152539 2.85163 0.00139502 0.998695 0.631307 0.0010391 0.00187952 0.000859217 0.45567 0.00187952 0.431642 0.000126314 1.02 0.88727 0.534795 0.285484 1.71606e-07 3.05356e-09 2397.56 3339.17 -0.0712957 0.482113 0.277743 0.267189 -0.590803 -0.169468 0.44987 -0.268836 -0.181022 1.041 1 8.90681e-227 282.298 4.932e-224 1.96167 1.039 0.000299994 0.953368 0.614782 0.702634 0.388592 1.96207 124.54 81.3844 18.5716 59.6358 0.00413264 0 -40 10
0.14 4.06072e-09 2.5388e-06 0.0379249 0.0378905 0.0120482 1.84578e-06 0.001154 0.0474062 0.000651661 0.0480532 0.846511 101.894 0.247332 0.700466 4.10552 0.0526685 0.0387313 0.961269 0.0198962 0.0042238 0.0191583 0.00406841 0.00510375 0.00584174 0.20415 0.23367 57.9483 -87.8931 125.336 15.9953 145.003 0.000151291 0.267075 192.934 0.31073 0.0673912 0.00409467 0.000561537 0.00138237 0.986994 0.991736 -2.97084e-06 -85.6688 0.0929756 31197.3 300.028 0.983523 0.319147 0.784822 0.784817 9.99958 2.98024e-06 1.19208e-05 0.130445 0.968352 0.924836 -0.0132934 4.89017e-06 0.50006 -1.83785e-20 6.76078e-24 -1.83717e-20 0.00139502 0.997818 8.59216e-05 0.152539 2.85163 0.00139502 0.99869 0.631436 0.00103911 0.00187952 0.000859216 0.455671 0.00187952 0.431654 0.000126317 1.02 0.887269 0.534796 0.285483 1.71606e-07 3.05354e-09 2397.54 3338.34 -0.0712338 0.482113 0.277742 0.267138 -0.590812 -0.169468 0.450055 -0.268836 -0.181206 1.042 1 5.40225e-227 282.356 2.99243e-224 1.96194 1.04 0.000299994 0.952988 0.614867 0.701599 0.388639 1.96234 124.555 81.3937 18.5722 59.6404 0.00413223 0 -40 10
0.141 4.08971e-09 2.5388e-06 0.0380456 0.0380114 0.0120481 1.85896e-06 0.001154 0.047557 0.000651696 0.0482041 0.846527 101.894 0.24733 0.700482 4.10553 0.0526697 0.0387314 0.961269 0.0198962 0.00422381 0.0191582 0.00406842 0.00510377 0.00584175 0.204151 0.23367 57.9483 -87.8931 125.339 15.9953 145.003 0.000151253 0.267075 192.934 0.310731 0.0673912 0.00409466 0.000561536 0.00138237 0.986994 0.991736 -2.97083e-06 -85.6688 0.0929755 31197.3 300.028 0.983523 0.319147 0.784627 0.784622 9.99958 2.98023e-06 1.19208e-05 0.130445 0.9684 0.924862 -0.0132934 4.89015e-06 0.50006 -1.83797e-20 6.76122e-24 -1.8373e-20 0.00139502 0.997818 8.59214e-05 0.152539 2.85163 0.00139502 0.998684 0.631564 0.00103911 0.00187952 0.000859214 0.455671 0.00187952 0.431665 0.00012632 1.02 0.887269 0.534796 0.285482 1.71606e-07 3.05353e-09 2397.53 3337.51 -0.0711721 0.482113 0.277742 0.267087 -0.590822 -0.169468 0.450239 -0.268836 -0.18139 1.043 1 3.27663e-227 282.413 1.81562e-224 1.96222 1.041 0.000299994 0.952609 0.614953 0.700566 0.388686 1.96261 124.569 81.403 18.5727 59.6449 0.00413183 0 -40 10
0.142 4.11871e-09 2.5388e-06 0.0381662 0.0381323 0.0120481 1.87214e-06 0.001154 0.0477077 0.00065173 0.0483548 0.846544 101.894 0.247329 0.700498 4.10554 0.052671 0.0387315 0.961268 0.0198962 0.00422382 0.0191582 0.00406843 0.00510378 0.00584176 0.204151 0.233671 57.9484 -87.8931 125.342 15.9953 145.003 0.000151216 0.267075 192.934 0.310732 0.0673913 0.00409466 0.000561535 0.00138236 0.986994 0.991736 -2.97081e-06 -85.6689 0.0929754 31197.4 300.028 0.983523 0.319147 0.784432 0.784427 9.99958 2.98022e-06 1.19208e-05 0.130445 0.968447 0.924888 -0.0132934 4.89014e-06 0.50006 -1.8381e-20 6.76167e-24 -1.83743e-20 0.00139501 0.997818 8.59213e-05 0.152538 2.85163 0.00139501 0.998678 0.631692 0.00103912 0.00187951 0.000859213 0.455671 0.00187952 0.431677 0.000126323 1.02 0.887268 0.534796 0.285481 1.71605e-07 3.05351e-09 2397.51 3336.68 -0.0711106 0.482113 0.277742 0.267036 -0.590831 -0.169468 0.450422 -0.268837 -0.181574 1.044 1 1.98738e-227 282.47 1.10161e-224 1.96249 1.042 0.000299994 0.952232 0.615038 0.699538 0.388732 1.96289 124.584 81.4122 18.5733 59.6494 0.00413143 0 -40 10
0.143 4.14771e-09 2.5388e-06 0.0382866 0.0382531 0.0120481 1.88532e-06 0.001154 0.0478583 0.000651764 0.0485055 0.846561 101.894 0.247328 0.700514 4.10555 0.0526723 0.0387316 0.961268 0.0198962 0.00422383 0.0191582 0.00406844 0.00510379 0.00584178 0.204152 0.233671 57.9484 -87.8931 125.345 15.9952 145.003 0.000151178 0.267074 192.934 0.310732 0.0673914 0.00409466 0.000561535 0.00138236 0.986994 0.991736 -2.9708e-06 -85.6689 0.0929753 31197.4 300.029 0.983523 0.319147 0.784237 0.784233 9.99958 2.98022e-06 1.19208e-05 0.130446 0.968494 0.924913 -0.0132934 4.89012e-06 0.500061 -1.83823e-20 6.76212e-24 -1.83756e-20 0.00139501 0.997818 8.59212e-05 0.152538 2.85163 0.00139501 0.998673 0.631821 0.00103912 0.00187951 0.000859212 0.455672 0.00187951 0.431688 0.000126325 1.02 0.887267 0.534796 0.28548 1.71605e-07 3.05349e-09 2397.49 3335.86 -0.0710493 0.482113 0.277741 0.266985 -0.59084 -0.169468 0.450605 -0.268837 -0.181756 1.045 1 1.20541e-227 282.527 6.68386e-225 1.96276 1.043 0.000299994 0.951856 0.615123 0.698512 0.388779 1.96316 124.598 81.4213 18.5738 59.6539 0.00413103 0 -40 10
0.144 4.17671e-09 2.5388e-06 0.038407 0.0383737 0.0120481 1.8985e-06 0.001154 0.0480088 0.000651797 0.048656 0.846578 101.894 0.247326 0.700531 4.10556 0.0526736 0.0387317 0.961268 0.0198962 0.00422385 0.0191582 0.00406845 0.00510381 0.00584179 0.204152 0.233672 57.9485 -87.8931 125.349 15.9952 145.003 0.000151141 0.267074 192.935 0.310733 0.0673914 0.00409465 0.000561534 0.00138236 0.986994 0.991736 -2.97078e-06 -85.6689 0.0929752 31197.4 300.029 0.983523 0.319147 0.784044 0.784039 9.99958 2.98021e-06 1.19207e-05 0.130446 0.968541 0.924939 -0.0132934 4.8901e-06 0.500061 -1.83836e-20 6.76256e-24 -1.83768e-20 0.00139501 0.997818 8.59211e-05 0.152538 2.85163 0.00139501 0.998667 0.631949 0.00103913 0.00187951 0.000859211 0.455672 0.00187951 0.4317 0.000126328 1.02 0.887267 0.534796 0.28548 1.71605e-07 3.05347e-09 2397.48 3335.03 -0.0709882 0.482113 0.277741 0.266935 -0.590849 -0.169468 0.450787 -0.268837 -0.181938 1.046 1 7.31115e-228 282.584 4.05534e-225 1.96303 1.044 0.000299993 0.951482 0.615208 0.697489 0.388826 1.96343 124.613 81.4305 18.5744 59.6584 0.00413063 0 -40 10
0.145 4.20571e-09 2.5388e-06 0.0385273 0.0384943 0.0120481 1.91169e-06 0.001154 0.0481591 0.00065183 0.0488064 0.846596 101.894 0.247325 0.700547 4.10557 0.0526749 0.0387318 0.961268 0.0198962 0.00422386 0.0191582 0.00406846 0.00510382 0.0058418 0.204153 0.233672 57.9486 -87.8931 125.352 15.9952 145.003 0.000151104 0.267074 192.935 0.310733 0.0673915 0.00409465 0.000561533 0.00138236 0.986994 0.991736 -2.97076e-06 -85.6689 0.0929751 31197.4 300.029 0.983523 0.319147 0.783851 0.783846 9.99958 2.98021e-06 1.19207e-05 0.130446 0.968588 0.924964 -0.0132934 4.89008e-06 0.500062 -1.83849e-20 6.76301e-24 -1.83781e-20 0.00139501 0.997818 8.5921e-05 0.152538 2.85163 0.00139501 0.998662 0.632077 0.00103914 0.00187951 0.00085921 0.455672 0.00187951 0.431711 0.000126331 1.02 0.887266 0.534797 0.285479 1.71604e-07 3.05346e-09 2397.46 3334.21 -0.0709274 0.482113 0.277741 0.266884 -0.590859 -0.169469 0.450968 -0.268837 -0.18212 1.047 1 4.43444e-228 282.641 2.46052e-225 1.9633 1.045 0.000299993 0.951108 0.615292 0.69647 0.388873 1.9637 124.627 81.4396 18.5749 59.6628 0.00413023 0 -40 10
0.146 4.23471e-09 2.5388e-06 0.0386475 0.0386148 0.0120481 1.92487e-06 0.001154 0.0483094 0.000651863 0.0489566 0.846613 101.894 0.247324 0.700564 4.10558 0.0526762 0.0387319 0.961268 0.0198962 0.00422387 0.0191582 0.00406847 0.00510384 0.00584182 0.204153 0.233673 57.9486 -87.8931 125.355 15.9951 145.003 0.000151067 0.267074 192.935 0.310734 0.0673916 0.00409465 0.000561532 0.00138235 0.986994 0.991736 -2.97075e-06 -85.6689 0.0929749 31197.5 300.029 0.983523 0.319147 0.783659 0.783654 9.99958 2.9802e-06 1.19207e-05 0.130446 0.968635 0.924989 -0.0132934 4.89007e-06 0.500062 -1.83861e-20 6.76345e-24 -1.83794e-20 0.00139501 0.997818 8.59209e-05 0.152538 2.85162 0.00139501 0.998656 0.632206 0.00103914 0.00187951 0.000859209 0.455672 0.00187951 0.431722 0.000126334 1.02 0.887265 0.534797 0.285478 1.71604e-07 3.05344e-09 2397.45 3333.4 -0.0708667 0.482113 0.27774 0.266834 -0.590868 -0.169469 0.451149 -0.268837 -0.182301 1.048 1 2.68962e-228 282.698 1.49289e-225 1.96357 1.046 0.000299993 0.950736 0.615377 0.695453 0.388919 1.96397 124.642 81.4487 18.5755 59.6673 0.00412984 0 -40 10
0.147 4.2637e-09 2.5388e-06 0.0387676 0.0387351 0.0120481 1.93805e-06 0.001154 0.0484595 0.000651896 0.0491068 0.84663 101.894 0.247322 0.700581 4.10559 0.0526776 0.038732 0.961268 0.0198962 0.00422388 0.0191582 0.00406848 0.00510385 0.00584183 0.204154 0.233673 57.9487 -87.8931 125.359 15.9951 145.003 0.00015103 0.267073 192.935 0.310734 0.0673916 0.00409464 0.000561531 0.00138235 0.986994 0.991736 -2.97073e-06 -85.6689 0.0929748 31197.5 300.03 0.983523 0.319147 0.783467 0.783462 9.99958 2.98019e-06 1.19207e-05 0.130446 0.968682 0.925014 -0.0132934 4.89005e-06 0.500063 -1.83874e-20 6.7639e-24 -1.83807e-20 0.00139501 0.997818 8.59208e-05 0.152537 2.85162 0.00139501 0.998651 0.632334 0.00103915 0.00187951 0.000859208 0.455673 0.00187951 0.431734 0.000126336 1.02 0.887265 0.534797 0.285477 1.71604e-07 3.05342e-09 2397.43 3332.58 -0.0708062 0.482112 0.27774 0.266784 -0.590877 -0.169469 0.45133 -0.268838 -0.182481 1.049 1 1.63134e-228 282.754 9.05787e-226 1.96384 1.047 0.000299993 0.950365 0.615461 0.69444 0.388966 1.96424 124.656 81.4578 18.576 59.6717 0.00412945 0 -40 10
0.148 4.2927e-09 2.5388e-06 0.0388876 0.0388554 0.012048 1.95123e-06 0.001154 0.0486095 0.000651928 0.0492568 0.846648 101.894 0.247321 0.700598 4.1056 0.0526789 0.0387321 0.961268 0.0198961 0.00422389 0.0191582 0.00406848 0.00510386 0.00584184 0.204155 0.233674 57.9487 -87.8931 125.362 15.9951 145.003 0.000150993 0.267073 192.935 0.310735 0.0673917 0.00409464 0.00056153 0.00138235 0.986994 0.991736 -2.97072e-06 -85.6689 0.0929747 31197.5 300.03 0.983523 0.319147 0.783276 0.783271 9.99958 2.98019e-06 1.19206e-05 0.130446 0.968728 0.925039 -0.0132934 4.89003e-06 0.500063 -1.83887e-20 6.76434e-24 -1.83819e-20 0.00139501 0.997818 8.59208e-05 0.152537 2.85162 0.00139501 0.998645 0.632462 0.00103915 0.0018795 0.000859208 0.455673 0.00187951 0.431745 0.000126339 1.02 0.887264 0.534797 0.285476 1.71603e-07 3.05341e-09 2397.41 3331.77 -0.0707459 0.482112 0.27774 0.266734 -0.590886 -0.169469 0.451509 -0.268838 -0.18266 1.05 1 9.89457e-229 282.81 5.49572e-226 1.96411 1.048 0.000299993 0.949996 0.615546 0.69343 0.389012 1.96451 124.671 81.4668 18.5766 59.6761 0.00412905 0 -40 10
0.149 4.3217e-09 2.5388e-06 0.0390075 0.0389756 0.012048 1.96441e-06 0.001154 0.0487594 0.00065196 0.0494067 0.846666 101.894 0.24732 0.700615 4.10561 0.0526803 0.0387322 0.961268 0.0198961 0.0042239 0.0191581 0.00406849 0.00510388 0.00584186 0.204155 0.233674 57.9488 -87.8931 125.365 15.995 145.003 0.000150956 0.267073 192.936 0.310735 0.0673917 0.00409463 0.00056153 0.00138235 0.986994 0.991736 -2.9707e-06 -85.6689 0.0929746 31197.5 300.03 0.983523 0.319147 0.783085 0.783081 9.99958 2.98018e-06 1.19206e-05 0.130446 0.968774 0.925064 -0.0132934 4.89002e-06 0.500064 -1.839e-20 6.76478e-24 -1.83832e-20 0.001395 0.997818 8.59207e-05 0.152537 2.85162 0.001395 0.99864 0.63259 0.00103916 0.0018795 0.000859207 0.455673 0.0018795 0.431757 0.000126342 1.02 0.887263 0.534797 0.285475 1.71603e-07 3.05339e-09 2397.4 3330.96 -0.0706859 0.482112 0.277739 0.266684 -0.590895 -0.169469 0.451688 -0.268838 -0.18284 1.051 1 6.00136e-229 282.866 3.33444e-226 1.96438 1.049 0.000299993 0.949627 0.61563 0.692422 0.389058 1.96478 124.685 81.4758 18.5771 59.6805 0.00412866 0 -40 10
0.15 4.3507e-09 2.5388e-06 0.0391273 0.0390956 0.012048 1.97759e-06 0.001154 0.0489091 0.000651992 0.0495565 0.846683 101.894 0.247318 0.700633 4.10562 0.0526817 0.0387323 0.961268 0.0198961 0.00422391 0.0191581 0.0040685 0.00510389 0.00584187 0.204156 0.233675 57.9488 -87.8931 125.368 15.995 145.003 0.00015092 0.267073 192.936 0.310736 0.0673918 0.00409463 0.000561529 0.00138234 0.986994 0.991736 -2.97069e-06 -85.6689 0.0929745 31197.6 300.031 0.983523 0.319147 0.782896 0.782891 9.99958 2.98018e-06 1.19206e-05 0.130446 0.96882 0.925089 -0.0132934 4.89e-06 0.500064 -1.83912e-20 6.76523e-24 -1.83845e-20 0.001395 0.997818 8.59206e-05 0.152537 2.85162 0.001395 0.998634 0.632718 0.00103917 0.0018795 0.000859206 0.455674 0.0018795 0.431768 0.000126345 1.02 0.887263 0.534798 0.285474 1.71603e-07 3.05338e-09 2397.38 3330.16 -0.070626 0.482112 0.277739 0.266634 -0.590904 -0.169469 0.451867 -0.268838 -0.183018 1.052 1 3.64001e-229 282.922 2.02312e-226 1.96465 1.05 0.000299993 0.94926 0.615714 0.691418 0.389105 1.96505 124.699 81.4848 18.5776 59.6849 0.00412827 0 -40 10
0.151 4.37969e-09 2.5388e-06 0.039247 0.0392156 0.012048 1.99077e-06 0.001154 0.0490587 0.000652023 0.0497062 0.846701 101.894 0.247317 0.70065 4.10563 0.0526831 0.0387324 0.961268 0.0198961 0.00422393 0.0191581 0.00406851 0.00510391 0.00584189 0.204156 0.233675 57.9489 -87.8931 125.372 15.995 145.003 0.000150883 0.267072 192.936 0.310736 0.0673919 0.00409463 0.000561528 0.00138234 0.986994 0.991736 -2.97067e-06 -85.669 0.0929744 31197.6 300.031 0.983523 0.319147 0.782706 0.782702 9.99958 2.98017e-06 1.19206e-05 0.130446 0.968866 0.925114 -0.0132934 4.88998e-06 0.500065 -1.83925e-20 6.76567e-24 -1.83857e-20 0.001395 0.997818 8.59205e-05 0.152537 2.85162 0.001395 0.998629 0.632846 0.00103917 0.0018795 0.000859205 0.455674 0.0018795 0.431779 0.000126348 1.02 0.887262 0.534798 0.285474 1.71602e-07 3.05336e-09 2397.37 3329.35 -0.0705663 0.482112 0.277739 0.266585 -0.590913 -0.169469 0.452045 -0.268838 -0.183196 1.053 1 2.20778e-229 282.978 1.22749e-226 1.96492 1.051 0.000299993 0.948894 0.615798 0.690417 0.389151 1.96531 124.714 81.4938 18.5782 59.6893 0.00412788 0 -40 10
0.152 4.40869e-09 2.5388e-06 0.0393666 0.0393355 0.012048 2.00395e-06 0.001154 0.0492083 0.000652055 0.0498557 0.846719 101.894 0.247316 0.700668 4.10564 0.0526845 0.0387325 0.961268 0.0198961 0.00422394 0.0191581 0.00406852 0.00510392 0.0058419 0.204157 0.233676 57.949 -87.8931 125.375 15.9949 145.003 0.000150847 0.267072 192.936 0.310737 0.0673919 0.00409462 0.000561527 0.00138234 0.986994 0.991736 -2.97066e-06 -85.669 0.0929743 31197.6 300.031 0.983523 0.319147 0.782518 0.782513 9.99958 2.98016e-06 1.19206e-05 0.130447 0.968912 0.925139 -0.0132934 4.88997e-06 0.500065 -1.83937e-20 6.76611e-24 -1.8387e-20 0.001395 0.997819 8.59204e-05 0.152537 2.85162 0.001395 0.998624 0.632974 0.00103918 0.0018795 0.000859204 0.455674 0.0018795 0.431791 0.000126351 1.02 0.887262 0.534798 0.285473 1.71602e-07 3.05335e-09 2397.35 3328.55 -0.0705068 0.482112 0.277738 0.266536 -0.590923 -0.169469 0.452222 -0.268838 -0.183373 1.054 1 1.33908e-229 283.033 7.4476e-227 1.96519 1.052 0.000299993 0.948529 0.615882 0.689419 0.389197 1.96558 124.728 81.5027 18.5787 59.6936 0.00412749 0 -40 10
0.153 4.43769e-09 2.5388e-06 0.0394861 0.0394552 0.012048 2.01713e-06 0.001154 0.0493576 0.000652086 0.0500051 0.846737 101.894 0.247314 0.700686 4.10565 0.0526859 0.0387326 0.961267 0.0198961 0.00422395 0.0191581 0.00406853 0.00510394 0.00584192 0.204157 0.233677 57.949 -87.8931 125.378 15.9949 145.003 0.000150811 0.267072 192.936 0.310737 0.067392 0.00409462 0.000561527 0.00138234 0.986994 0.991736 -2.97065e-06 -85.669 0.0929742 31197.6 300.032 0.983523 0.319147 0.78233 0.782325 9.99958 2.98016e-06 1.19205e-05 0.130447 0.968958 0.925163 -0.0132934 4.88995e-06 0.500066 -1.8395e-20 6.76655e-24 -1.83882e-20 0.001395 0.997819 8.59203e-05 0.152536 2.85162 0.001395 0.998619 0.633102 0.00103919 0.00187949 0.000859203 0.455674 0.0018795 0.431802 0.000126353 1.02 0.887261 0.534798 0.285472 1.71602e-07 3.05333e-09 2397.34 3327.75 -0.0704476 0.482112 0.277738 0.266486 -0.590932 -0.169469 0.452399 -0.268838 -0.18355 1.055 1 8.12196e-230 283.088 4.5187e-227 1.96546 1.053 0.000299993 0.948165 0.615966 0.688424 0.389243 1.96585 124.743 81.5116 18.5792 59.698 0.00412711 0 -40 10
0.154 4.46669e-09 2.5388e-06 0.0396055 0.0395749 0.012048 2.03031e-06 0.001154 0.0495069 0.000652116 0.0501544 0.846755 101.894 0.247313 0.700704 4.10566 0.0526873 0.0387327 0.961267 0.019896 0.00422396 0.0191581 0.00406854 0.00510395 0.00584193 0.204158 0.233677 57.9491 -87.8931 125.381 15.9949 145.003 0.000150774 0.267072 192.936 0.310738 0.067392 0.00409462 0.000561526 0.00138233 0.986994 0.991736 -2.97063e-06 -85.669 0.0929741 31197.7 300.032 0.983523 0.319147 0.782143 0.782138 9.99958 2.98015e-06 1.19205e-05 0.130447 0.969003 0.925188 -0.0132934 4.88994e-06 0.500066 -1.83963e-20 6.76699e-24 -1.83895e-20 0.001395 0.997819 8.59202e-05 0.152536 2.85162 0.001395 0.998613 0.63323 0.00103919 0.00187949 0.000859202 0.455675 0.00187949 0.431813 0.000126356 1.02 0.887261 0.534798 0.285471 1.71601e-07 3.05332e-09 2397.32 3326.96 -0.0703885 0.482112 0.277738 0.266437 -0.590941 -0.169469 0.452575 -0.268838 -0.183726 1.056 1 4.92622e-230 283.144 2.74164e-227 1.96572 1.054 0.000299993 0.947803 0.61605 0.687433 0.389289 1.96612 124.757 81.5205 18.5798 59.7023 0.00412672 0 -40 10
0.155 4.49568e-09 2.53881e-06 0.0397249 0.0396945 0.012048 2.04349e-06 0.001154 0.0496561 0.000652147 0.0503036 0.846774 101.894 0.247311 0.700722 4.10568 0.0526888 0.0387328 0.961267 0.019896 0.00422398 0.0191581 0.00406855 0.00510397 0.00584195 0.204159 0.233678 57.9491 -87.8931 125.384 15.9948 145.003 0.000150738 0.267072 192.937 0.310738 0.0673921 0.00409461 0.000561525 0.00138233 0.986994 0.991736 -2.97062e-06 -85.669 0.092974 31197.7 300.032 0.983523 0.319147 0.781956 0.781951 9.99958 2.98015e-06 1.19205e-05 0.130447 0.969049 0.925212 -0.0132934 4.88992e-06 0.500067 -1.83975e-20 6.76743e-24 -1.83907e-20 0.001395 0.997819 8.59201e-05 0.152536 2.85161 0.001395 0.998608 0.633358 0.0010392 0.00187949 0.000859201 0.455675 0.00187949 0.431825 0.000126359 1.02 0.88726 0.534798 0.28547 1.71601e-07 3.0533e-09 2397.3 3326.16 -0.0703296 0.482112 0.277737 0.266388 -0.590949 -0.169469 0.45275 -0.268838 -0.183902 1.057 1 2.9879e-230 283.199 1.66344e-227 1.96599 1.055 0.000299993 0.947442 0.616134 0.686444 0.389335 1.96638 124.771 81.5293 18.5803 59.7066 0.00412634 0 -40 10
0.156 4.52468e-09 2.53881e-06 0.0398441 0.0398139 0.0120479 2.05667e-06 0.001154 0.0498051 0.000652177 0.0504527 0.846792 101.894 0.24731 0.700741 4.10569 0.0526902 0.0387329 0.961267 0.019896 0.00422399 0.019158 0.00406856 0.00510398 0.00584196 0.204159 0.233678 57.9492 -87.8931 125.388 15.9948 145.003 0.000150703 0.267071 192.937 0.310739 0.0673922 0.00409461 0.000561524 0.00138233 0.986994 0.991736 -2.9706e-06 -85.669 0.0929739 31197.7 300.033 0.983523 0.319147 0.78177 0.781765 9.99958 2.98014e-06 1.19205e-05 0.130447 0.969094 0.925237 -0.0132934 4.88991e-06 0.500067 -1.83988e-20 6.76787e-24 -1.8392e-20 0.001395 0.997819 8.592e-05 0.152536 2.85161 0.001395 0.998603 0.633486 0.00103921 0.00187949 0.0008592 0.455675 0.00187949 0.431836 0.000126362 1.02 0.887259 0.534798 0.28547 1.71601e-07 3.05329e-09 2397.29 3325.37 -0.0702709 0.482112 0.277737 0.26634 -0.590958 -0.169469 0.452925 -0.268838 -0.184077 1.058 1 1.81225e-230 283.253 1.00926e-227 1.96626 1.056 0.000299993 0.947082 0.616217 0.685458 0.389381 1.96665 124.785 81.5381 18.5808 59.711 0.00412596 0 -40 10
0.157 4.55368e-09 2.53881e-06 0.0399632 0.0399333 0.0120479 2.06985e-06 0.001154 0.049954 0.000652207 0.0506016 0.846811 101.894 0.247308 0.700759 4.1057 0.0526917 0.038733 0.961267 0.019896 0.004224 0.019158 0.00406857 0.005104 0.00584198 0.20416 0.233679 57.9492 -87.8931 125.391 15.9948 145.003 0.000150667 0.267071 192.937 0.310739 0.0673922 0.00409461 0.000561524 0.00138233 0.986994 0.991736 -2.97059e-06 -85.669 0.0929738 31197.7 300.033 0.983523 0.319147 0.781584 0.78158 9.99958 2.98014e-06 1.19204e-05 0.130447 0.969139 0.925261 -0.0132934 4.8899e-06 0.500068 -1.84e-20 6.76831e-24 -1.83932e-20 0.00139499 0.997819 8.59199e-05 0.152536 2.85161 0.00139499 0.998598 0.633613 0.00103921 0.00187949 0.000859199 0.455675 0.00187949 0.431848 0.000126365 1.02 0.887259 0.534799 0.285469 1.71601e-07 3.05328e-09 2397.27 3324.58 -0.0702124 0.482112 0.277737 0.266291 -0.590967 -0.16947 0.4531 -0.268839 -0.184251 1.059 1 1.09919e-230 283.308 6.12346e-228 1.96653 1.057 0.000299993 0.946723 0.6163 0.684475 0.389427 1.96692 124.8 81.5469 18.5813 59.7152 0.00412558 0 -40 10
0.158 4.58267e-09 2.53881e-06 0.0400823 0.0400526 0.0120479 2.08303e-06 0.001154 0.0501028 0.000652237 0.0507505 0.846829 101.894 0.247307 0.700778 4.10571 0.0526932 0.0387331 0.961267 0.019896 0.00422401 0.019158 0.00406858 0.00510401 0.00584199 0.204161 0.23368 57.9493 -87.8931 125.394 15.9947 145.003 0.000150631 0.267071 192.937 0.31074 0.0673923 0.0040946 0.000561523 0.00138232 0.986994 0.991736 -2.97058e-06 -85.669 0.0929738 31197.8 300.033 0.983523 0.319147 0.781399 0.781395 9.99958 2.98013e-06 1.19204e-05 0.130447 0.969184 0.925285 -0.0132934 4.88988e-06 0.500068 -1.84013e-20 6.76875e-24 -1.83945e-20 0.00139499 0.997819 8.59199e-05 0.152536 2.85161 0.00139499 0.998593 0.633741 0.00103922 0.00187949 0.000859199 0.455676 0.00187949 0.431859 0.000126368 1.02 0.887258 0.534799 0.285468 1.716e-07 3.05326e-09 2397.26 3323.8 -0.0701542 0.482112 0.277736 0.266243 -0.590976 -0.16947 0.453274 -0.268839 -0.184425 1.06 1 6.66691e-231 283.363 3.71529e-228 1.96679 1.058 0.000299993 0.946366 0.616384 0.683495 0.389473 1.96718 124.814 81.5557 18.5819 59.7195 0.0041252 0 -40 10
0.159 4.61167e-09 2.53881e-06 0.0402012 0.0401718 0.0120479 2.09621e-06 0.001154 0.0502515 0.000652266 0.0508992 0.846848 101.894 0.247305 0.700797 4.10572 0.0526947 0.0387332 0.961267 0.019896 0.00422403 0.019158 0.0040686 0.00510403 0.00584201 0.204161 0.23368 57.9494 -87.8931 125.397 15.9947 145.003 0.000150596 0.267071 192.937 0.31074 0.0673923 0.0040946 0.000561522 0.00138232 0.986994 0.991736 -2.97057e-06 -85.669 0.0929737 31197.8 300.034 0.983523 0.319147 0.781215 0.78121 9.99958 2.98013e-06 1.19204e-05 0.130447 0.969229 0.925309 -0.0132934 4.88987e-06 0.500069 -1.84025e-20 6.76919e-24 -1.83957e-20 0.00139499 0.997819 8.59198e-05 0.152535 2.85161 0.00139499 0.998588 0.633869 0.00103923 0.00187949 0.000859198 0.455676 0.00187949 0.43187 0.00012637 1.02 0.887258 0.534799 0.285468 1.716e-07 3.05325e-09 2397.24 3323.01 -0.0700961 0.482111 0.277736 0.266195 -0.590985 -0.16947 0.453447 -0.268839 -0.184598 1.061 1 4.04369e-231 283.417 2.25417e-228 1.96706 1.059 0.000299993 0.946009 0.616467 0.682518 0.389518 1.96745 124.828 81.5644 18.5824 59.7238 0.00412482 0 -40 10
0.16 4.64067e-09 2.53881e-06 0.04032 0.0402909 0.0120479 2.10939e-06 0.001154 0.0504001 0.000652296 0.0510477 0.846867 101.894 0.247304 0.700816 4.10573 0.0526962 0.0387333 0.961267 0.019896 0.00422404 0.019158 0.00406861 0.00510405 0.00584202 0.204162 0.233681 57.9494 -87.8931 125.4 15.9947 145.003 0.00015056 0.267071 192.938 0.31074 0.0673924 0.0040946 0.000561522 0.00138232 0.986994 0.991736 -2.97055e-06 -85.669 0.0929736 31197.8 300.034 0.983523 0.319147 0.781031 0.781027 9.99958 2.98012e-06 1.19204e-05 0.130448 0.969274 0.925333 -0.0132934 4.88986e-06 0.500069 -1.84037e-20 6.76962e-24 -1.8397e-20 0.00139499 0.997819 8.59197e-05 0.152535 2.85161 0.00139499 0.998583 0.633996 0.00103924 0.00187948 0.000859197 0.455676 0.00187949 0.431882 0.000126373 1.02 0.887257 0.534799 0.285467 1.716e-07 3.05324e-09 2397.22 3322.23 -0.0700382 0.482111 0.277736 0.266146 -0.590994 -0.16947 0.453619 -0.268839 -0.184771 1.062 1 2.45262e-231 283.471 1.36767e-228 1.96732 1.06 0.000299993 0.945654 0.61655 0.681544 0.389564 1.96771 124.842 81.5731 18.5829 59.728 0.00412444 0 -40 10
0.161 4.66966e-09 2.53881e-06 0.0404388 0.0404098 0.0120479 2.12257e-06 0.001154 0.0505485 0.000652325 0.0511962 0.846886 101.894 0.247302 0.700835 4.10575 0.0526977 0.0387335 0.961267 0.0198959 0.00422405 0.019158 0.00406862 0.00510406 0.00584204 0.204163 0.233682 57.9495 -87.8931 125.403 15.9946 145.003 0.000150525 0.26707 192.938 0.310741 0.0673924 0.00409459 0.000561521 0.00138232 0.986994 0.991736 -2.97054e-06 -85.6691 0.0929735 31197.8 300.034 0.983524 0.319147 0.780848 0.780844 9.99958 2.98012e-06 1.19204e-05 0.130448 0.969318 0.925357 -0.0132934 4.88984e-06 0.50007 -1.8405e-20 6.77006e-24 -1.83982e-20 0.00139499 0.997819 8.59196e-05 0.152535 2.85161 0.00139499 0.998578 0.634124 0.00103924 0.00187948 0.000859196 0.455676 0.00187948 0.431893 0.000126376 1.02 0.887257 0.534799 0.285466 1.71599e-07 3.05322e-09 2397.21 3321.46 -0.0699804 0.482111 0.277735 0.266098 -0.591003 -0.16947 0.453791 -0.268839 -0.184943 1.063 1 1.48759e-231 283.525 8.29804e-229 1.96759 1.061 0.000299993 0.9453 0.616633 0.680573 0.38961 1.96798 124.856 81.5818 18.5834 59.7323 0.00412406 0 -40 10
0.162 4.69866e-09 2.53881e-06 0.0405574 0.0405287 0.0120479 2.13575e-06 0.001154 0.0506968 0.000652354 0.0513446 0.846905 101.894 0.247301 0.700855 4.10576 0.0526992 0.0387336 0.961266 0.0198959 0.00422407 0.0191579 0.00406863 0.00510408 0.00584205 0.204163 0.233682 57.9495 -87.8932 125.406 15.9946 145.003 0.00015049 0.26707 192.938 0.310741 0.0673925 0.00409459 0.00056152 0.00138232 0.986994 0.991736 -2.97053e-06 -85.6691 0.0929734 31197.9 300.035 0.983524 0.319147 0.780666 0.780661 9.99958 2.98011e-06 1.19203e-05 0.130448 0.969363 0.925381 -0.0132934 4.88983e-06 0.50007 -1.84062e-20 6.7705e-24 -1.83994e-20 0.00139499 0.997819 8.59195e-05 0.152535 2.85161 0.00139499 0.998573 0.634251 0.00103925 0.00187948 0.000859195 0.455676 0.00187948 0.431904 0.000126379 1.02 0.887256 0.534799 0.285466 1.71599e-07 3.05321e-09 2397.19 3320.68 -0.0699229 0.482111 0.277735 0.266051 -0.591011 -0.16947 0.453963 -0.268838 -0.185115 1.064 1 9.02268e-232 283.579 5.03465e-229 1.96785 1.062 0.000299993 0.944947 0.616716 0.679605 0.389655 1.96824 124.87 81.5905 18.5839 59.7365 0.00412369 0 -40 10
0.163 4.72765e-09 2.53881e-06 0.040676 0.0406475 0.0120478 2.14893e-06 0.001154 0.050845 0.000652382 0.0514928 0.846924 101.894 0.247299 0.700874 4.10577 0.0527008 0.0387337 0.961266 0.0198959 0.00422408 0.0191579 0.00406864 0.0051041 0.00584207 0.204164 0.233683 57.9496 -87.8932 125.41 15.9946 145.003 0.000150455 0.26707 192.938 0.310742 0.0673925 0.00409459 0.00056152 0.00138231 0.986994 0.991736 -2.97051e-06 -85.6691 0.0929733 31197.9 300.035 0.983524 0.319147 0.780484 0.780479 9.99958 2.98011e-06 1.19203e-05 0.130448 0.969407 0.925404 -0.0132935 4.88982e-06 0.500071 -1.84074e-20 6.77093e-24 -1.84007e-20 0.00139499 0.997819 8.59194e-05 0.152535 2.85161 0.00139499 0.998568 0.634379 0.00103926 0.00187948 0.000859194 0.455677 0.00187948 0.431916 0.000126382 1.02 0.887256 0.534799 0.285465 1.71599e-07 3.0532e-09 2397.18 3319.91 -0.0698656 0.482111 0.277734 0.266003 -0.59102 -0.16947 0.454134 -0.268838 -0.185286 1.065 1 5.47253e-232 283.632 3.05466e-229 1.96812 1.063 0.000299993 0.944596 0.616799 0.67864 0.389701 1.96851 124.885 81.5991 18.5845 59.7407 0.00412331 0 -40 10
0.164 4.75665e-09 2.53881e-06 0.0407945 0.0407662 0.0120478 2.16211e-06 0.001154 0.0509931 0.000652411 0.0516409 0.846943 101.894 0.247298 0.700894 4.10578 0.0527023 0.0387338 0.961266 0.0198959 0.00422409 0.0191579 0.00406865 0.00510411 0.00584209 0.204165 0.233684 57.9497 -87.8932 125.413 15.9945 145.003 0.00015042 0.26707 192.938 0.310742 0.0673926 0.00409459 0.000561519 0.00138231 0.986994 0.991736 -2.9705e-06 -85.6691 0.0929732 31197.9 300.036 0.983524 0.319147 0.780303 0.780298 9.99958 2.9801e-06 1.19203e-05 0.130448 0.969451 0.925428 -0.0132935 4.88981e-06 0.500071 -1.84087e-20 6.77137e-24 -1.84019e-20 0.00139499 0.997819 8.59194e-05 0.152535 2.85161 0.00139499 0.998563 0.634506 0.00103927 0.00187948 0.000859194 0.455677 0.00187948 0.431927 0.000126385 1.02 0.887256 0.5348 0.285464 1.71599e-07 3.05319e-09 2397.16 3319.14 -0.0698085 0.482111 0.277734 0.265956 -0.591029 -0.16947 0.454304 -0.268838 -0.185456 1.066 1 3.31926e-232 283.686 1.85334e-229 1.96838 1.064 0.000299993 0.944245 0.616881 0.677677 0.389746 1.96877 124.899 81.6077 18.585 59.7449 0.00412294 0 -40 10
0.165 4.78565e-09 2.53881e-06 0.0409128 0.0408848 0.0120478 2.17529e-06 0.001154 0.0511411 0.000652439 0.0517889 0.846963 101.894 0.247296 0.700914 4.1058 0.0527039 0.0387339 0.961266 0.0198959 0.00422411 0.0191579 0.00406866 0.00510413 0.0058421 0.204165 0.233684 57.9497 -87.8932 125.416 15.9945 145.003 0.000150385 0.26707 192.938 0.310743 0.0673926 0.00409458 0.000561518 0.00138231 0.986995 0.991737 -2.97049e-06 -85.6691 0.0929731 31197.9 300.036 0.983524 0.319147 0.780122 0.780117 9.99958 2.9801e-06 1.19203e-05 0.130448 0.969495 0.925452 -0.0132935 4.8898e-06 0.500072 -1.84099e-20 6.7718e-24 -1.84031e-20 0.00139499 0.997819 8.59193e-05 0.152534 2.85161 0.00139499 0.998558 0.634634 0.00103927 0.00187948 0.000859193 0.455677 0.00187948 0.431938 0.000126388 1.02 0.887255 0.5348 0.285464 1.71598e-07 3.05317e-09 2397.14 3318.37 -0.0697515 0.482111 0.277734 0.265908 -0.591038 -0.16947 0.454474 -0.268838 -0.185626 1.067 1 2.01323e-232 283.739 1.12447e-229 1.96865 1.065 0.000299993 0.943896 0.616964 0.676718 0.389791 1.96903 124.913 81.6163 18.5855 59.7491 0.00412257 0 -40 10
0.166 4.81464e-09 2.53881e-06 0.0410311 0.0410033 0.0120478 2.18847e-06 0.001154 0.0512889 0.000652467 0.0519368 0.846982 101.894 0.247295 0.700934 4.10581 0.0527055 0.038734 0.961266 0.0198959 0.00422412 0.0191579 0.00406867 0.00510415 0.00584212 0.204166 0.233685 57.9498 -87.8932 125.419 15.9944 145.003 0.00015035 0.267069 192.938 0.310743 0.0673927 0.00409458 0.000561518 0.00138231 0.986995 0.991737 -2.97048e-06 -85.6691 0.0929731 31198 300.036 0.983524 0.319147 0.779942 0.779937 9.99958 2.98009e-06 1.19203e-05 0.130448 0.969539 0.925475 -0.0132935 4.88978e-06 0.500073 -1.84111e-20 6.77224e-24 -1.84044e-20 0.00139498 0.997819 8.59192e-05 0.152534 2.8516 0.00139498 0.998553 0.634761 0.00103928 0.00187947 0.000859192 0.455677 0.00187948 0.431949 0.000126391 1.02 0.887255 0.5348 0.285463 1.71598e-07 3.05316e-09 2397.13 3317.6 -0.0696948 0.482111 0.277733 0.265861 -0.591046 -0.16947 0.454643 -0.268838 -0.185796 1.068 1 1.22109e-232 283.792 6.82245e-230 1.96891 1.066 0.000299993 0.943548 0.617046 0.675762 0.389837 1.9693 124.927 81.6248 18.586 59.7533 0.0041222 0 -40 10
0.167 4.84364e-09 2.53881e-06 0.0411493 0.0411217 0.0120478 2.20165e-06 0.001154 0.0514366 0.000652495 0.0520845 0.847002 101.894 0.247293 0.700954 4.10582 0.0527071 0.0387342 0.961266 0.0198958 0.00422414 0.0191579 0.00406869 0.00510417 0.00584214 0.204167 0.233686 57.9498 -87.8932 125.422 15.9944 145.003 0.000150316 0.267069 192.939 0.310743 0.0673927 0.00409458 0.000561517 0.00138231 0.986995 0.991737 -2.97047e-06 -85.6691 0.092973 31198 300.037 0.983524 0.319147 0.779762 0.779758 9.99958 2.98009e-06 1.19202e-05 0.130449 0.969583 0.925498 -0.0132935 4.88977e-06 0.500073 -1.84124e-20 6.77267e-24 -1.84056e-20 0.00139498 0.997819 8.59191e-05 0.152534 2.8516 0.00139498 0.998548 0.634888 0.00103929 0.00187947 0.000859191 0.455678 0.00187947 0.431961 0.000126394 1.02 0.887254 0.5348 0.285462 1.71598e-07 3.05315e-09 2397.11 3316.84 -0.0696382 0.482111 0.277733 0.265814 -0.591055 -0.16947 0.454811 -0.268838 -0.185964 1.069 1 7.40627e-233 283.845 4.13935e-230 1.96917 1.067 0.000299993 0.943201 0.617128 0.674808 0.389882 1.96956 124.941 81.6333 18.5865 59.7574 0.00412183 0 -40 10
0.168 4.87263e-09 2.53881e-06 0.0412674 0.04124 0.0120478 2.21483e-06 0.001154 0.0515842 0.000652522 0.0522322 0.847021 101.894 0.247291 0.700974 4.10583 0.0527087 0.0387343 0.961266 0.0198958 0.00422415 0.0191578 0.0040687 0.00510418 0.00584216 0.204167 0.233686 57.9499 -87.8932 125.425 15.9944 145.003 0.000150281 0.267069 192.939 0.310744 0.0673928 0.00409457 0.000561516 0.0013823 0.986995 0.991737 -2.97046e-06 -85.6691 0.0929729 31198 300.037 0.983524 0.319147 0.779583 0.779579 9.99958 2.98008e-06 1.19202e-05 0.130449 0.969627 0.925522 -0.0132935 4.88976e-06 0.500074 -1.84136e-20 6.7731e-24 -1.84068e-20 0.00139498 0.997819 8.59191e-05 0.152534 2.8516 0.00139498 0.998544 0.635015 0.0010393 0.00187947 0.000859191 0.455678 0.00187947 0.431972 0.000126397 1.02 0.887254 0.5348 0.285462 1.71598e-07 3.05314e-09 2397.1 3316.08 -0.0695819 0.482111 0.277733 0.265767 -0.591063 -0.16947 0.454979 -0.268838 -0.186133 1.07 1 4.49213e-233 283.898 2.51145e-230 1.96944 1.068 0.000299993 0.942855 0.617211 0.673858 0.389927 1.96982 124.955 81.6418 18.587 59.7616 0.00412146 0 -40 10
0.169 4.90163e-09 2.53881e-06 0.0413854 0.0413582 0.0120478 2.22801e-06 0.001154 0.0517317 0.000652549 0.0523797 0.847041 101.894 0.24729 0.700995 4.10585 0.0527103 0.0387344 0.961266 0.0198958 0.00422417 0.0191578 0.00406871 0.0051042 0.00584217 0.204168 0.233687 57.9499 -87.8932 125.428 15.9943 145.003 0.000150247 0.267069 192.939 0.310744 0.0673928 0.00409457 0.000561516 0.0013823 0.986995 0.991737 -2.97044e-06 -85.6691 0.0929728 31198 300.037 0.983524 0.319147 0.779405 0.7794 9.99958 2.98008e-06 1.19202e-05 0.130449 0.96967 0.925545 -0.0132935 4.88975e-06 0.500074 -1.84148e-20 6.77354e-24 -1.8408e-20 0.00139498 0.997819 8.5919e-05 0.152534 2.8516 0.00139498 0.998539 0.635143 0.00103931 0.00187947 0.00085919 0.455678 0.00187947 0.431983 0.000126399 1.02 0.887253 0.5348 0.285461 1.71597e-07 3.05313e-09 2397.08 3315.32 -0.0695257 0.482111 0.277732 0.26572 -0.591072 -0.169471 0.455147 -0.268838 -0.1863 1.071 1 2.72461e-233 283.951 1.52375e-230 1.9697 1.069 0.000299993 0.94251 0.617293 0.67291 0.389972 1.97008 124.969 81.6503 18.5875 59.7657 0.0041211 0 -40 10
0.17 4.93063e-09 2.53881e-06 0.0415033 0.0414763 0.0120478 2.24119e-06 0.001154 0.0518791 0.000652576 0.0525271 0.847061 101.894 0.247288 0.701016 4.10586 0.052712 0.0387345 0.961265 0.0198958 0.00422418 0.0191578 0.00406872 0.00510422 0.00584219 0.204169 0.233688 57.95 -87.8932 125.431 15.9943 145.003 0.000150213 0.267069 192.939 0.310745 0.0673929 0.00409457 0.000561515 0.0013823 0.986995 0.991737 -2.97043e-06 -85.6691 0.0929727 31198 300.038 0.983524 0.319147 0.779227 0.779223 9.99958 2.98007e-06 1.19202e-05 0.130449 0.969713 0.925568 -0.0132935 4.88974e-06 0.500075 -1.8416e-20 6.77397e-24 -1.84092e-20 0.00139498 0.997819 8.59189e-05 0.152534 2.8516 0.00139498 0.998534 0.63527 0.00103931 0.00187947 0.000859189 0.455678 0.00187947 0.431995 0.000126402 1.02 0.887253 0.5348 0.285461 1.71597e-07 3.05312e-09 2397.07 3314.57 -0.0694697 0.482111 0.277732 0.265674 -0.591081 -0.169471 0.455314 -0.268838 -0.186467 1.072 1 1.65256e-233 284.003 9.24498e-231 1.96996 1.07 0.000299993 0.942167 0.617375 0.671965 0.390017 1.97035 124.983 81.6587 18.588 59.7698 0.00412073 0 -40 10
0.171 4.95962e-09 2.53881e-06 0.0416211 0.0415943 0.0120477 2.25437e-06 0.001154 0.0520263 0.000652603 0.0526744 0.847081 101.894 0.247286 0.701036 4.10587 0.0527136 0.0387347 0.961265 0.0198958 0.0042242 0.0191578 0.00406873 0.00510424 0.00584221 0.204169 0.233688 57.9501 -87.8932 125.434 15.9943 145.004 0.000150178 0.267069 192.939 0.310745 0.0673929 0.00409457 0.000561515 0.0013823 0.986995 0.991737 -2.97042e-06 -85.6691 0.0929727 31198.1 300.038 0.983524 0.319147 0.77905 0.779046 9.99958 2.98007e-06 1.19202e-05 0.130449 0.969757 0.925591 -0.0132935 4.88973e-06 0.500076 -1.84172e-20 6.7744e-24 -1.84104e-20 0.00139498 0.997819 8.59188e-05 0.152534 2.8516 0.00139498 0.998529 0.635397 0.00103932 0.00187947 0.000859188 0.455678 0.00187947 0.432006 0.000126405 1.02 0.887253 0.5348 0.28546 1.71597e-07 3.05311e-09 2397.05 3313.82 -0.0694139 0.482111 0.277732 0.265627 -0.591089 -0.169471 0.45548 -0.268838 -0.186634 1.073 1 1.00233e-233 284.056 5.60914e-231 1.97022 1.071 0.000299993 0.941824 0.617457 0.671023 0.390062 1.97061 124.997 81.6671 18.5885 59.7739 0.00412037 0 -40 10
0.172 4.98862e-09 2.53881e-06 0.0417388 0.0417122 0.0120477 2.26755e-06 0.001154 0.0521735 0.00065263 0.0528215 0.847101 101.894 0.247285 0.701057 4.10589 0.0527153 0.0387348 0.961265 0.0198957 0.00422421 0.0191578 0.00406875 0.00510426 0.00584223 0.20417 0.233689 57.9501 -87.8932 125.437 15.9942 145.004 0.000150144 0.267068 192.939 0.310745 0.067393 0.00409456 0.000561514 0.0013823 0.986995 0.991737 -2.97041e-06 -85.6692 0.0929726 31198.1 300.039 0.983524 0.319147 0.778874 0.778869 9.99958 2.98007e-06 1.19202e-05 0.130449 0.9698 0.925614 -0.0132935 4.88972e-06 0.500076 -1.84184e-20 6.77483e-24 -1.84117e-20 0.00139498 0.997819 8.59188e-05 0.152533 2.8516 0.00139498 0.998525 0.635524 0.00103933 0.00187947 0.000859188 0.455679 0.00187947 0.432017 0.000126408 1.02 0.887252 0.5348 0.28546 1.71597e-07 3.0531e-09 2397.03 3313.06 -0.0693583 0.482111 0.277731 0.265581 -0.591098 -0.169471 0.455646 -0.268837 -0.1868 1.074 1 6.07943e-234 284.108 3.40319e-231 1.97049 1.072 0.000299993 0.941483 0.617538 0.670084 0.390107 1.97087 125.011 81.6755 18.589 59.778 0.00412001 0 -40 10
0.173 5.01761e-09 2.53881e-06 0.0418564 0.04183 0.0120477 2.28073e-06 0.001154 0.0523205 0.000652656 0.0529686 0.847121 101.894 0.247283 0.701079 4.1059 0.052717 0.0387349 0.961265 0.0198957 0.00422423 0.0191578 0.00406876 0.00510427 0.00584224 0.204171 0.23369 57.9502 -87.8932 125.44 15.9942 145.004 0.00015011 0.267068 192.94 0.310746 0.067393 0.00409456 0.000561513 0.00138229 0.986995 0.991737 -2.9704e-06 -85.6692 0.0929725 31198.1 300.039 0.983524 0.319147 0.778698 0.778693 9.99958 2.98006e-06 1.19201e-05 0.13045 0.969843 0.925637 -0.0132935 4.88971e-06 0.500077 -1.84196e-20 6.77526e-24 -1.84129e-20 0.00139498 0.997819 8.59187e-05 0.152533 2.8516 0.00139498 0.99852 0.635651 0.00103934 0.00187947 0.000859187 0.455679 0.00187947 0.432028 0.000126411 1.02 0.887252 0.534801 0.285459 1.71596e-07 3.05309e-09 2397.02 3312.32 -0.0693028 0.48211 0.277731 0.265535 -0.591106 -0.169471 0.455811 -0.268837 -0.186966 1.075 1 3.68736e-234 284.16 2.06479e-231 1.97075 1.073 0.000299993 0.941143 0.61762 0.669147 0.390152 1.97113 125.025 81.6839 18.5895 59.7821 0.00411964 0 -40 10
0.174 5.04661e-09 2.53881e-06 0.0419739 0.0419477 0.0120477 2.29391e-06 0.001154 0.0524674 0.000652683 0.0531155 0.847141 101.894 0.247281 0.7011 4.10591 0.0527186 0.038735 0.961265 0.0198957 0.00422424 0.0191577 0.00406877 0.00510429 0.00584226 0.204172 0.23369 57.9502 -87.8932 125.443 15.9942 145.004 0.000150077 0.267068 192.94 0.310746 0.0673931 0.00409456 0.000561513 0.00138229 0.986995 0.991737 -2.97039e-06 -85.6692 0.0929724 31198.1 300.04 0.983524 0.319147 0.778522 0.778518 9.99958 2.98006e-06 1.19201e-05 0.13045 0.969885 0.92566 -0.0132935 4.8897e-06 0.500077 -1.84209e-20 6.77569e-24 -1.84141e-20 0.00139498 0.997819 8.59186e-05 0.152533 2.8516 0.00139498 0.998516 0.635778 0.00103935 0.00187946 0.000859186 0.455679 0.00187947 0.43204 0.000126414 1.02 0.887252 0.534801 0.285459 1.71596e-07 3.05308e-09 2397 3311.57 -0.0692476 0.48211 0.277731 0.265489 -0.591115 -0.169471 0.455976 -0.268837 -0.187131 1.076 1 2.2365e-234 284.212 1.25275e-231 1.97101 1.074 0.000299993 0.940804 0.617702 0.668214 0.390197 1.97139 125.039 81.6922 18.59 59.7862 0.00411928 0 -40 10
0.175 5.0756e-09 2.53881e-06 0.0420913 0.0420654 0.0120477 2.30709e-06 0.001154 0.0526142 0.000652709 0.0532623 0.847162 101.894 0.24728 0.701122 4.10593 0.0527204 0.0387352 0.961265 0.0198957 0.00422426 0.0191577 0.00406878 0.00510431 0.00584228 0.204172 0.233691 57.9503 -87.8932 125.446 15.9941 145.004 0.000150043 0.267068 192.94 0.310746 0.0673931 0.00409456 0.000561512 0.00138229 0.986995 0.991737 -2.97038e-06 -85.6692 0.0929724 31198.1 300.04 0.983524 0.319147 0.778347 0.778343 9.99958 2.98005e-06 1.19201e-05 0.13045 0.969928 0.925682 -0.0132935 4.88969e-06 0.500078 -1.84221e-20 6.77612e-24 -1.84153e-20 0.00139497 0.997819 8.59186e-05 0.152533 2.8516 0.00139497 0.998511 0.635905 0.00103936 0.00187946 0.000859186 0.455679 0.00187946 0.432051 0.000126417 1.02 0.887251 0.534801 0.285458 1.71596e-07 3.05307e-09 2396.99 3310.83 -0.0691925 0.48211 0.27773 0.265443 -0.591123 -0.169471 0.45614 -0.268837 -0.187295 1.077 1 1.35651e-234 284.263 7.60072e-232 1.97127 1.075 0.000299993 0.940466 0.617783 0.667283 0.390242 1.97165 125.053 81.7005 18.5905 59.7902 0.00411892 0 -40 10
0.176 5.1046e-09 2.53881e-06 0.0422087 0.0421829 0.0120477 2.32027e-06 0.001154 0.0527608 0.000652735 0.053409 0.847182 101.894 0.247278 0.701143 4.10594 0.0527221 0.0387353 0.961265 0.0198957 0.00422427 0.0191577 0.0040688 0.00510433 0.0058423 0.204173 0.233692 57.9504 -87.8932 125.449 15.9941 145.004 0.000150009 0.267068 192.94 0.310747 0.0673932 0.00409455 0.000561512 0.00138229 0.986995 0.991737 -2.97037e-06 -85.6692 0.0929723 31198.2 300.04 0.983524 0.319147 0.778173 0.778169 9.99958 2.98005e-06 1.19201e-05 0.13045 0.969971 0.925705 -0.0132935 4.88968e-06 0.500079 -1.84233e-20 6.77655e-24 -1.84165e-20 0.00139497 0.997819 8.59185e-05 0.152533 2.8516 0.00139497 0.998507 0.636032 0.00103937 0.00187946 0.000859185 0.455679 0.00187946 0.432062 0.00012642 1.02 0.887251 0.534801 0.285458 1.71596e-07 3.05306e-09 2396.97 3310.09 -0.0691376 0.48211 0.27773 0.265397 -0.591131 -0.169471 0.456303 -0.268837 -0.187459 1.078 1 8.22762e-235 284.315 4.61152e-232 1.97153 1.076 0.000299993 0.940129 0.617865 0.666355 0.390286 1.97191 125.067 81.7088 18.591 59.7943 0.00411857 0 -40 10
0.177 5.13359e-09 2.53881e-06 0.0423259 0.0423003 0.0120477 2.33345e-06 0.001154 0.0529074 0.00065276 0.0535556 0.847203 101.894 0.247276 0.701165 4.10596 0.0527238 0.0387354 0.961265 0.0198957 0.00422429 0.0191577 0.00406881 0.00510435 0.00584232 0.204174 0.233693 57.9504 -87.8932 125.452 15.9941 145.004 0.000149976 0.267068 192.94 0.310747 0.0673932 0.00409455 0.000561511 0.00138229 0.986995 0.991737 -2.97036e-06 -85.6692 0.0929722 31198.2 300.041 0.983524 0.319147 0.777999 0.777995 9.99958 2.98004e-06 1.19201e-05 0.13045 0.970013 0.925727 -0.0132935 4.88967e-06 0.500079 -1.84245e-20 6.77698e-24 -1.84177e-20 0.00139497 0.997819 8.59184e-05 0.152533 2.8516 0.00139497 0.998502 0.636159 0.00103937 0.00187946 0.000859184 0.45568 0.00187946 0.432073 0.000126423 1.02 0.887251 0.534801 0.285457 1.71595e-07 3.05305e-09 2396.95 3309.35 -0.0690829 0.48211 0.27773 0.265352 -0.59114 -0.169471 0.456466 -0.268836 -0.187622 1.079 1 4.9903e-235 284.366 2.7979e-232 1.97179 1.077 0.000299993 0.939794 0.617946 0.66543 0.390331 1.97217 125.081 81.7171 18.5915 59.7983 0.00411821 0 -40 10
0.178 5.16259e-09 2.53881e-06 0.0424431 0.0424177 0.0120477 2.34663e-06 0.001154 0.0530538 0.000652786 0.053702 0.847223 101.894 0.247274 0.701187 4.10597 0.0527255 0.0387356 0.961264 0.0198956 0.0042243 0.0191577 0.00406882 0.00510437 0.00584234 0.204175 0.233693 57.9505 -87.8932 125.455 15.994 145.004 0.000149942 0.267067 192.94 0.310747 0.0673932 0.00409455 0.000561511 0.00138228 0.986995 0.991737 -2.97035e-06 -85.6692 0.0929721 31198.2 300.041 0.983524 0.319147 0.777826 0.777822 9.99958 2.98004e-06 1.19201e-05 0.13045 0.970055 0.92575 -0.0132935 4.88967e-06 0.50008 -1.84257e-20 6.77741e-24 -1.84189e-20 0.00139497 0.997819 8.59184e-05 0.152533 2.85159 0.00139497 0.998498 0.636286 0.00103938 0.00187946 0.000859184 0.45568 0.00187946 0.432085 0.000126426 1.02 0.88725 0.534801 0.285457 1.71595e-07 3.05304e-09 2396.94 3308.61 -0.0690284 0.48211 0.277729 0.265306 -0.591148 -0.169471 0.456629 -0.268836 -0.187785 1.08 1 3.02677e-235 284.417 1.69754e-232 1.97205 1.078 0.000299993 0.939459 0.618027 0.664508 0.390376 1.97243 125.094 81.7253 18.592 59.8023 0.00411785 0 -40 10
0.179 5.19158e-09 2.53881e-06 0.0425601 0.0425349 0.0120476 2.35981e-06 0.001154 0.0532001 0.000652811 0.0538483 0.847244 101.894 0.247273 0.701209 4.10599 0.0527273 0.0387357 0.961264 0.0198956 0.00422432 0.0191576 0.00406883 0.00510439 0.00584236 0.204176 0.233694 57.9505 -87.8932 125.458 15.994 145.004 0.000149909 0.267067 192.94 0.310748 0.0673933 0.00409455 0.00056151 0.00138228 0.986995 0.991737 -2.97034e-06 -85.6692 0.0929721 31198.2 300.042 0.983524 0.319147 0.777654 0.777649 9.99958 2.98004e-06 1.192e-05 0.13045 0.970098 0.925772 -0.0132935 4.88966e-06 0.500081 -1.84269e-20 6.77784e-24 -1.84201e-20 0.00139497 0.997819 8.59183e-05 0.152533 2.85159 0.00139497 0.998493 0.636412 0.00103939 0.00187946 0.000859183 0.45568 0.00187946 0.432096 0.000126429 1.02 0.88725 0.534801 0.285456 1.71595e-07 3.05303e-09 2396.92 3307.88 -0.0689741 0.48211 0.277729 0.265261 -0.591156 -0.169471 0.456791 -0.268836 -0.187947 1.081 1 1.83583e-235 284.468 1.02993e-232 1.97231 1.079 0.000299993 0.939126 0.618108 0.663588 0.39042 1.97269 125.108 81.7335 18.5925 59.8063 0.0041175 0 -40 10
0.18 5.22058e-09 2.53881e-06 0.0426771 0.042652 0.0120476 2.37299e-06 0.001154 0.0533463 0.000652836 0.0539946 0.847265 101.894 0.247271 0.701232 4.106 0.0527291 0.0387359 0.961264 0.0198956 0.00422434 0.0191576 0.00406885 0.00510441 0.00584238 0.204176 0.233695 57.9506 -87.8932 125.461 15.994 145.004 0.000149876 0.267067 192.94 0.310748 0.0673933 0.00409454 0.000561509 0.00138228 0.986995 0.991737 -2.97033e-06 -85.6692 0.092972 31198.2 300.042 0.983524 0.319147 0.777482 0.777477 9.99958 2.98003e-06 1.192e-05 0.130451 0.97014 0.925794 -0.0132935 4.88965e-06 0.500081 -1.8428e-20 6.77827e-24 -1.84213e-20 0.00139497 0.997819 8.59182e-05 0.152532 2.85159 0.00139497 0.998489 0.636539 0.0010394 0.00187946 0.000859182 0.45568 0.00187946 0.432107 0.000126432 1.02 0.88725 0.534801 0.285456 1.71595e-07 3.05302e-09 2396.91 3307.15 -0.06892 0.48211 0.277729 0.265216 -0.591165 -0.169471 0.456952 -0.268836 -0.188109 1.082 1 1.11349e-235 284.519 6.24878e-233 1.97257 1.08 0.000299993 0.938794 0.618189 0.662671 0.390465 1.97294 125.122 81.7417 18.593 59.8103 0.00411715 0 -40 10
0.181 5.24957e-09 2.53881e-06 0.0427939 0.0427691 0.0120476 2.38617e-06 0.001154 0.0534924 0.000652861 0.0541407 0.847286 101.894 0.247269 0.701254 4.10602 0.0527308 0.038736 0.961264 0.0198956 0.00422435 0.0191576 0.00406886 0.00510443 0.0058424 0.204177 0.233696 57.9506 -87.8932 125.464 15.9939 145.004 0.000149843 0.267067 192.941 0.310749 0.0673934 0.00409454 0.000561509 0.00138228 0.986995 0.991737 -2.97032e-06 -85.6692 0.0929719 31198.2 300.043 0.983524 0.319147 0.77731 0.777306 9.99958 2.98003e-06 1.192e-05 0.130451 0.970181 0.925817 -0.0132935 4.88964e-06 0.500082 -1.84292e-20 6.77869e-24 -1.84225e-20 0.00139497 0.997819 8.59182e-05 0.152532 2.85159 0.00139497 0.998484 0.636666 0.00103941 0.00187946 0.000859182 0.45568 0.00187946 0.432118 0.000126435 1.02 0.887249 0.534801 0.285456 1.71595e-07 3.05301e-09 2396.89 3306.42 -0.068866 0.48211 0.277728 0.265171 -0.591173 -0.169471 0.457113 -0.268835 -0.18827 1.083 1 6.75364e-236 284.57 3.79125e-233 1.97282 1.081 0.000299993 0.938463 0.61827 0.661757 0.390509 1.9732 125.136 81.7498 18.5934 59.8143 0.0041168 0 -40 10
0.182 5.27857e-09 2.53881e-06 0.0429107 0.042886 0.0120476 2.39935e-06 0.001154 0.0536384 0.000652886 0.0542867 0.847307 101.894 0.247267 0.701277 4.10603 0.0527326 0.0387361 0.961264 0.0198956 0.00422437 0.0191576 0.00406887 0.00510445 0.00584241 0.204178 0.233697 57.9507 -87.8932 125.467 15.9939 145.004 0.00014981 0.267067 192.941 0.310749 0.0673934 0.00409454 0.000561508 0.00138228 0.986995 0.991737 -2.97031e-06 -85.6692 0.0929719 31198.3 300.043 0.983524 0.319147 0.77714 0.777135 9.99958 2.98002e-06 1.192e-05 0.130451 0.970223 0.925839 -0.0132935 4.88963e-06 0.500083 -1.84304e-20 6.77912e-24 -1.84236e-20 0.00139497 0.997819 8.59181e-05 0.152532 2.85159 0.00139497 0.99848 0.636792 0.00103942 0.00187945 0.000859181 0.45568 0.00187946 0.43213 0.000126438 1.02 0.887249 0.534801 0.285455 1.71594e-07 3.053e-09 2396.87 3305.69 -0.0688122 0.48211 0.277728 0.265126 -0.591181 -0.169472 0.457273 -0.268835 -0.188431 1.084 1 4.09629e-236 284.621 2.30022e-233 1.97308 1.082 0.000299993 0.938133 0.618351 0.660846 0.390553 1.97346 125.15 81.758 18.5939 59.8183 0.00411644 0 -40 10
0.183 5.30756e-09 2.53881e-06 0.0430274 0.0430029 0.0120476 2.41253e-06 0.001154 0.0537842 0.000652911 0.0544325 0.847328 101.894 0.247266 0.7013 4.10605 0.0527344 0.0387363 0.961264 0.0198955 0.00422438 0.0191576 0.00406889 0.00510447 0.00584243 0.204179 0.233697 57.9508 -87.8932 125.47 15.9939 145.004 0.000149777 0.267067 192.941 0.310749 0.0673935 0.00409454 0.000561508 0.00138228 0.986995 0.991737 -2.9703e-06 -85.6692 0.0929718 31198.3 300.043 0.983524 0.319147 0.776969 0.776965 9.99958 2.98002e-06 1.192e-05 0.130451 0.970265 0.925861 -0.0132935 4.88963e-06 0.500083 -1.84316e-20 6.77954e-24 -1.84248e-20 0.00139497 0.997819 8.5918e-05 0.152532 2.85159 0.00139497 0.998476 0.636919 0.00103943 0.00187945 0.00085918 0.455681 0.00187945 0.432141 0.000126441 1.02 0.887249 0.534801 0.285455 1.71594e-07 3.05299e-09 2396.86 3304.97 -0.0687586 0.48211 0.277728 0.265081 -0.591189 -0.169472 0.457433 -0.268835 -0.188591 1.085 1 2.48453e-236 284.671 1.39558e-233 1.97334 1.083 0.000299993 0.937804 0.618431 0.659937 0.390598 1.97372 125.163 81.7661 18.5944 59.8222 0.00411609 0 -40 10
0.184 5.33655e-09 2.53881e-06 0.043144 0.0431196 0.0120476 2.42571e-06 0.001154 0.0539299 0.000652935 0.0545783 0.84735 101.894 0.247264 0.701323 4.10606 0.0527363 0.0387364 0.961264 0.0198955 0.0042244 0.0191575 0.0040689 0.00510449 0.00584245 0.20418 0.233698 57.9508 -87.8932 125.473 15.9938 145.004 0.000149744 0.267067 192.941 0.310749 0.0673935 0.00409453 0.000561507 0.00138227 0.986995 0.991737 -2.97029e-06 -85.6692 0.0929717 31198.3 300.044 0.983524 0.319147 0.776799 0.776795 9.99958 2.98002e-06 1.192e-05 0.130451 0.970306 0.925883 -0.0132935 4.88962e-06 0.500084 -1.84328e-20 6.77997e-24 -1.8426e-20 0.00139497 0.997819 8.5918e-05 0.152532 2.85159 0.00139497 0.998471 0.637045 0.00103944 0.00187945 0.00085918 0.455681 0.00187945 0.432152 0.000126444 1.02 0.887248 0.534802 0.285454 1.71594e-07 3.05299e-09 2396.84 3304.25 -0.0687052 0.48211 0.277727 0.265037 -0.591198 -0.169472 0.457592 -0.268835 -0.188751 1.086 1 1.50694e-236 284.721 8.46724e-234 1.9736 1.084 0.000299993 0.937476 0.618512 0.659031 0.390642 1.97397 125.177 81.7741 18.5949 59.8261 0.00411575 0 -40 10
0.185 5.36555e-09 2.53881e-06 0.0432604 0.0432363 0.0120476 2.43889e-06 0.001154 0.0540756 0.000652959 0.0547239 0.847371 101.894 0.247262 0.701346 4.10608 0.0527381 0.0387366 0.961263 0.0198955 0.00422442 0.0191575 0.00406892 0.00510451 0.00584248 0.20418 0.233699 57.9509 -87.8932 125.476 15.9938 145.004 0.000149712 0.267066 192.941 0.31075 0.0673935 0.00409453 0.000561507 0.00138227 0.986995 0.991737 -2.97028e-06 -85.6693 0.0929717 31198.3 300.044 0.983524 0.319147 0.77663 0.776626 9.99958 2.98001e-06 1.19199e-05 0.130451 0.970348 0.925905 -0.0132935 4.88961e-06 0.500085 -1.8434e-20 6.78039e-24 -1.84272e-20 0.00139497 0.997819 8.59179e-05 0.152532 2.85159 0.00139497 0.998467 0.637172 0.00103945 0.00187945 0.000859179 0.455681 0.00187945 0.432163 0.000126447 1.02 0.887248 0.534802 0.285454 1.71594e-07 3.05298e-09 2396.83 3303.53 -0.0686519 0.48211 0.277727 0.264992 -0.591206 -0.169472 0.457751 -0.268834 -0.18891 1.087 1 9.14006e-237 284.771 5.13721e-234 1.97386 1.085 0.000299992 0.937149 0.618592 0.658128 0.390686 1.97423 125.191 81.7822 18.5954 59.8301 0.0041154 0 -40 10
0.186 5.39454e-09 2.53881e-06 0.0433768 0.0433529 0.0120475 2.45206e-06 0.001154 0.054221 0.000652983 0.0548694 0.847393 101.894 0.24726 0.701369 4.10609 0.0527399 0.0387367 0.961263 0.0198955 0.00422444 0.0191575 0.00406893 0.00510453 0.0058425 0.204181 0.2337 57.9509 -87.8932 125.479 15.9937 145.004 0.000149679 0.267066 192.941 0.31075 0.0673936 0.00409453 0.000561506 0.00138227 0.986995 0.991737 -2.97028e-06 -85.6693 0.0929716 31198.3 300.045 0.983524 0.319147 0.776462 0.776457 9.99958 2.98001e-06 1.19199e-05 0.130452 0.970389 0.925926 -0.0132935 4.88961e-06 0.500085 -1.84352e-20 6.78082e-24 -1.84284e-20 0.00139496 0.997819 8.59179e-05 0.152532 2.85159 0.00139496 0.998463 0.637298 0.00103946 0.00187945 0.000859179 0.455681 0.00187945 0.432174 0.00012645 1.02 0.887248 0.534802 0.285454 1.71594e-07 3.05297e-09 2396.81 3302.81 -0.0685989 0.48211 0.277727 0.264948 -0.591214 -0.169472 0.457909 -0.268834 -0.189068 1.088 1 5.54373e-237 284.821 3.11683e-234 1.97411 1.086 0.000299992 0.936823 0.618673 0.657228 0.39073 1.97449 125.205 81.7902 18.5958 59.834 0.00411505 0 -40 10
0.187 5.42354e-09 2.53881e-06 0.0434931 0.0434693 0.0120475 2.46524e-06 0.001154 0.0543664 0.000653007 0.0550148 0.847414 101.894 0.247258 0.701393 4.10611 0.0527418 0.0387369 0.961263 0.0198954 0.00422445 0.0191575 0.00406894 0.00510455 0.00584252 0.204182 0.233701 57.951 -87.8932 125.481 15.9937 145.004 0.000149647 0.267066 192.941 0.31075 0.0673936 0.00409453 0.000561506 0.00138227 0.986995 0.991737 -2.97027e-06 -85.6693 0.0929715 31198.3 300.045 0.983524 0.319147 0.776294 0.776289 9.99958 2.98001e-06 1.19199e-05 0.130452 0.97043 0.925948 -0.0132935 4.8896e-06 0.500086 -1.84363e-20 6.78124e-24 -1.84296e-20 0.00139496 0.997819 8.59178e-05 0.152532 2.85159 0.00139496 0.998459 0.637425 0.00103947 0.00187945 0.000859178 0.455681 0.00187945 0.432186 0.000126453 1.02 0.887248 0.534802 0.285453 1.71593e-07 3.05296e-09 2396.79 3302.1 -0.068546 0.48211 0.277726 0.264904 -0.591222 -0.169472 0.458066 -0.268834 -0.189226 1.089 1 3.36244e-237 284.871 1.89103e-234 1.97437 1.087 0.000299992 0.936499 0.618753 0.65633 0.390774 1.97474 125.218 81.7982 18.5963 59.8379 0.00411471 0 -40 10
0.188 5.45253e-09 2.53881e-06 0.0436093 0.0435857 0.0120475 2.47842e-06 0.001154 0.0545117 0.000653031 0.0551601 0.847436 101.894 0.247256 0.701416 4.10612 0.0527437 0.038737 0.961263 0.0198954 0.00422447 0.0191575 0.00406896 0.00510458 0.00584254 0.204183 0.233701 57.9511 -87.8932 125.484 15.9937 145.004 0.000149615 0.267066 192.941 0.310751 0.0673936 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97026e-06 -85.6693 0.0929715 31198.4 300.046 0.983524 0.319147 0.776126 0.776121 9.99958 2.98e-06 1.19199e-05 0.130452 0.970471 0.92597 -0.0132935 4.88959e-06 0.500087 -1.84375e-20 6.78167e-24 -1.84307e-20 0.00139496 0.997819 8.59177e-05 0.152531 2.85159 0.00139496 0.998454 0.637551 0.00103948 0.00187945 0.000859177 0.455681 0.00187945 0.432197 0.000126456 1.02 0.887247 0.534802 0.285453 1.71593e-07 3.05296e-09 2396.78 3301.39 -0.0684933 0.48211 0.277726 0.26486 -0.59123 -0.169472 0.458223 -0.268833 -0.189384 1.09 1 2.03942e-237 284.921 1.14732e-234 1.97463 1.088 0.000299992 0.936175 0.618833 0.655435 0.390818 1.975 125.232 81.8062 18.5968 59.8418 0.00411436 0 -40 10
0.189 5.48152e-09 2.53881e-06 0.0437255 0.043702 0.0120475 2.4916e-06 0.001154 0.0546568 0.000653054 0.0553053 0.847458 101.894 0.247254 0.70144 4.10614 0.0527456 0.0387372 0.961263 0.0198954 0.00422449 0.0191574 0.00406897 0.0051046 0.00584256 0.204184 0.233702 57.9511 -87.8933 125.487 15.9936 145.004 0.000149582 0.267066 192.942 0.310751 0.0673937 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97025e-06 -85.6693 0.0929714 31198.4 300.046 0.983524 0.319147 0.775959 0.775954 9.99958 2.98e-06 1.19199e-05 0.130452 0.970512 0.925991 -0.0132935 4.88959e-06 0.500088 -1.84387e-20 6.78209e-24 -1.84319e-20 0.00139496 0.997819 8.59177e-05 0.152531 2.85159 0.00139496 0.99845 0.637677 0.00103949 0.00187945 0.000859177 0.455682 0.00187945 0.432208 0.000126459 1.02 0.887247 0.534802 0.285453 1.71593e-07 3.05295e-09 2396.76 3300.68 -0.0684407 0.48211 0.277726 0.264816 -0.591238 -0.169472 0.45838 -0.268833 -0.189541 1.091 1 1.23697e-237 284.97 6.96093e-235 1.97488 1.089 0.000299992 0.935853 0.618913 0.654543 0.390862 1.97525 125.246 81.8141 18.5973 59.8457 0.00411402 0 -40 10
0.19 5.51052e-09 2.53881e-06 0.0438415 0.0438182 0.0120475 2.50478e-06 0.001154 0.0548019 0.000653078 0.0554503 0.84748 101.894 0.247253 0.701464 4.10616 0.0527475 0.0387373 0.961263 0.0198954 0.00422451 0.0191574 0.00406899 0.00510462 0.00584258 0.204185 0.233703 57.9512 -87.8933 125.49 15.9936 145.004 0.00014955 0.267066 192.942 0.310751 0.0673937 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97024e-06 -85.6693 0.0929714 31198.4 300.047 0.983524 0.319147 0.775793 0.775788 9.99958 2.98e-06 1.19199e-05 0.130452 0.970552 0.926013 -0.0132935 4.88958e-06 0.500088 -1.84399e-20 6.78251e-24 -1.84331e-20 0.00139496 0.997819 8.59176e-05 0.152531 2.85159 0.00139496 0.998446 0.637804 0.0010395 0.00187945 0.000859176 0.455682 0.00187945 0.432219 0.000126462 1.02 0.887247 0.534802 0.285452 1.71593e-07 3.05294e-09 2396.75 3299.97 -0.0683884 0.482109 0.277725 0.264772 -0.591246 -0.169472 0.458536 -0.268832 -0.189697 1.092 1 7.50262e-238 285.019 4.2233e-235 1.97514 1.09 0.000299992 0.935532 0.618993 0.653653 0.390906 1.97551 125.259 81.8221 18.5977 59.8495 0.00411368 0 -40 10
0.191 5.53951e-09 2.53881e-06 0.0439574 0.0439343 0.0120475 2.51796e-06 0.001154 0.0549468 0.000653101 0.0555953 0.847502 101.894 0.247251 0.701488 4.10617 0.0527494 0.0387375 0.961263 0.0198954 0.00422452 0.0191574 0.004069 0.00510464 0.0058426 0.204186 0.233704 57.9512 -87.8933 125.493 15.9936 145.004 0.000149518 0.267066 192.942 0.310752 0.0673938 0.00409452 0.000561504 0.00138226 0.986995 0.991737 -2.97023e-06 -85.6693 0.0929713 31198.4 300.047 0.983524 0.319147 0.775627 0.775622 9.99958 2.97999e-06 1.19199e-05 0.130453 0.970593 0.926034 -0.0132935 4.88958e-06 0.500089 -1.8441e-20 6.78293e-24 -1.84342e-20 0.00139496 0.997819 8.59176e-05 0.152531 2.85159 0.00139496 0.998442 0.63793 0.00103951 0.00187944 0.000859176 0.455682 0.00187945 0.43223 0.000126465 1.02 0.887247 0.534802 0.285452 1.71593e-07 3.05294e-09 2396.73 3299.26 -0.0683362 0.482109 0.277725 0.264729 -0.591254 -0.169472 0.458691 -0.268832 -0.189853 1.093 1 4.55057e-238 285.069 2.56233e-235 1.97539 1.091 0.000299992 0.935211 0.619073 0.652766 0.39095 1.97576 125.273 81.83 18.5982 59.8534 0.00411334 0 -40 10
0.192 5.56851e-09 2.53881e-06 0.0440733 0.0440503 0.0120475 2.53114e-06 0.001154 0.0550916 0.000653124 0.0557401 0.847524 101.894 0.247249 0.701513 4.10619 0.0527513 0.0387376 0.961262 0.0198953 0.00422454 0.0191574 0.00406902 0.00510466 0.00584262 0.204187 0.233705 57.9513 -87.8933 125.496 15.9935 145.004 0.000149487 0.267065 192.942 0.310752 0.0673938 0.00409452 0.000561504 0.00138226 0.986995 0.991737 -2.97023e-06 -85.6693 0.0929712 31198.4 300.048 0.983524 0.319147 0.775461 0.775457 9.99958 2.97999e-06 1.19199e-05 0.130453 0.970633 0.926056 -0.0132935 4.88957e-06 0.50009 -1.84422e-20 6.78336e-24 -1.84354e-20 0.00139496 0.997819 8.59175e-05 0.152531 2.85159 0.00139496 0.998438 0.638056 0.00103952 0.00187944 0.000859175 0.455682 0.00187944 0.432241 0.000126469 1.02 0.887247 0.534802 0.285452 1.71593e-07 3.05293e-09 2396.71 3298.56 -0.0682842 0.482109 0.277725 0.264685 -0.591262 -0.169472 0.458846 -0.268832 -0.190009 1.094 1 2.76006e-238 285.118 1.5546e-235 1.97565 1.092 0.000299992 0.934892 0.619153 0.651882 0.390993 1.97602 125.287 81.8378 18.5987 59.8572 0.004113 0 -40 10
0.193 5.5975e-09 2.53881e-06 0.044189 0.0441662 0.0120475 2.54432e-06 0.001154 0.0552362 0.000653147 0.0558848 0.847546 101.894 0.247247 0.701537 4.10621 0.0527532 0.0387378 0.961262 0.0198953 0.00422456 0.0191574 0.00406903 0.00510469 0.00584264 0.204187 0.233706 57.9513 -87.8933 125.499 15.9935 145.004 0.000149455 0.267065 192.942 0.310752 0.0673938 0.00409451 0.000561503 0.00138226 0.986995 0.991737 -2.97022e-06 -85.6693 0.0929712 31198.4 300.048 0.983524 0.319147 0.775297 0.775292 9.99958 2.97999e-06 1.19198e-05 0.130453 0.970674 0.926077 -0.0132935 4.88957e-06 0.500091 -1.84434e-20 6.78378e-24 -1.84366e-20 0.00139496 0.997819 8.59175e-05 0.152531 2.85158 0.00139496 0.998434 0.638182 0.00103953 0.00187944 0.000859175 0.455682 0.00187944 0.432253 0.000126472 1.02 0.887246 0.534802 0.285452 1.71592e-07 3.05292e-09 2396.7 3297.86 -0.0682324 0.482109 0.277724 0.264642 -0.59127 -0.169472 0.459001 -0.268831 -0.190163 1.095 1 1.67406e-238 285.166 9.43196e-236 1.9759 1.093 0.000299992 0.934574 0.619232 0.651 0.391037 1.97627 125.3 81.8457 18.5992 59.861 0.00411266 0 -40 10
0.194 5.62649e-09 2.53881e-06 0.0443046 0.044282 0.0120474 2.5575e-06 0.001154 0.0553808 0.00065317 0.0560294 0.847568 101.894 0.247245 0.701562 4.10622 0.0527552 0.0387379 0.961262 0.0198953 0.00422458 0.0191573 0.00406905 0.00510471 0.00584267 0.204188 0.233707 57.9514 -87.8933 125.501 15.9935 145.004 0.000149423 0.267065 192.942 0.310752 0.0673939 0.00409451 0.000561503 0.00138226 0.986995 0.991737 -2.97021e-06 -85.6693 0.0929711 31198.4 300.049 0.983524 0.319147 0.775132 0.775128 9.99958 2.97998e-06 1.19198e-05 0.130453 0.970714 0.926098 -0.0132935 4.88956e-06 0.500091 -1.84445e-20 6.7842e-24 -1.84377e-20 0.00139496 0.997819 8.59174e-05 0.152531 2.85158 0.00139496 0.99843 0.638308 0.00103954 0.00187944 0.000859174 0.455682 0.00187944 0.432264 0.000126475 1.02 0.887246 0.534802 0.285451 1.71592e-07 3.05292e-09 2396.68 3297.16 -0.0681807 0.482109 0.277724 0.264599 -0.591278 -0.169472 0.459155 -0.268831 -0.190318 1.096 1 1.01537e-238 285.215 5.72249e-236 1.97616 1.094 0.000299992 0.934257 0.619312 0.650121 0.391081 1.97653 125.314 81.8535 18.5996 59.8649 0.00411232 0 -40 10
0.195 5.65549e-09 2.53881e-06 0.0444202 0.0443977 0.0120474 2.57068e-06 0.001154 0.0555253 0.000653192 0.0561739 0.847591 101.894 0.247243 0.701586 4.10624 0.0527572 0.0387381 0.961262 0.0198953 0.0042246 0.0191573 0.00406906 0.00510473 0.00584269 0.204189 0.233708 57.9515 -87.8933 125.504 15.9934 145.004 0.000149392 0.267065 192.942 0.310753 0.0673939 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.9702e-06 -85.6693 0.0929711 31198.5 300.049 0.983524 0.319147 0.774969 0.774964 9.99958 2.97998e-06 1.19198e-05 0.130453 0.970754 0.926119 -0.0132935 4.88956e-06 0.500092 -1.84457e-20 6.78462e-24 -1.84389e-20 0.00139496 0.997819 8.59174e-05 0.152531 2.85158 0.00139496 0.998426 0.638434 0.00103955 0.00187944 0.000859174 0.455682 0.00187944 0.432275 0.000126478 1.02 0.887246 0.534802 0.285451 1.71592e-07 3.05291e-09 2396.67 3296.47 -0.0681292 0.482109 0.277724 0.264556 -0.591286 -0.169473 0.459308 -0.26883 -0.190472 1.097 1 6.15852e-239 285.264 3.4719e-236 1.97641 1.095 0.000299992 0.933941 0.619391 0.649245 0.391124 1.97678 125.327 81.8613 18.6001 59.8687 0.00411199 0 -40 10
0.196 5.68448e-09 2.53881e-06 0.0445357 0.0445133 0.0120474 2.58385e-06 0.001154 0.0556696 0.000653215 0.0563182 0.847613 101.894 0.247241 0.701611 4.10626 0.0527591 0.0387383 0.961262 0.0198952 0.00422462 0.0191573 0.00406908 0.00510475 0.00584271 0.20419 0.233708 57.9515 -87.8933 125.507 15.9934 145.004 0.00014936 0.267065 192.942 0.310753 0.0673939 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.9702e-06 -85.6693 0.092971 31198.5 300.05 0.983524 0.319147 0.774806 0.774801 9.99958 2.97998e-06 1.19198e-05 0.130453 0.970794 0.92614 -0.0132935 4.88955e-06 0.500093 -1.84468e-20 6.78504e-24 -1.84401e-20 0.00139496 0.997819 8.59173e-05 0.152531 2.85158 0.00139496 0.998422 0.63856 0.00103956 0.00187944 0.000859173 0.455683 0.00187944 0.432286 0.000126481 1.02 0.887246 0.534802 0.285451 1.71592e-07 3.05291e-09 2396.65 3295.77 -0.0680779 0.482109 0.277723 0.264513 -0.591294 -0.169473 0.459461 -0.26883 -0.190625 1.098 1 3.73533e-239 285.312 2.10644e-236 1.97666 1.096 0.000299992 0.933626 0.619471 0.648371 0.391168 1.97703 125.341 81.8691 18.6005 59.8725 0.00411165 0 -40 10
0.197 5.71347e-09 2.53881e-06 0.044651 0.0446289 0.0120474 2.59703e-06 0.001154 0.0558138 0.000653237 0.0564624 0.847636 101.894 0.247239 0.701637 4.10627 0.0527611 0.0387384 0.961262 0.0198952 0.00422463 0.0191573 0.00406909 0.00510478 0.00584273 0.204191 0.233709 57.9516 -87.8933 125.51 15.9934 145.004 0.000149329 0.267065 192.942 0.310753 0.067394 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.97019e-06 -85.6693 0.092971 31198.5 300.05 0.983524 0.319147 0.774643 0.774638 9.99958 2.97997e-06 1.19198e-05 0.130454 0.970834 0.926161 -0.0132935 4.88955e-06 0.500094 -1.8448e-20 6.78546e-24 -1.84412e-20 0.00139496 0.997819 8.59173e-05 0.152531 2.85158 0.00139496 0.998418 0.638686 0.00103957 0.00187944 0.000859173 0.455683 0.00187944 0.432297 0.000126484 1.02 0.887246 0.534802 0.285451 1.71592e-07 3.0529e-09 2396.63 3295.08 -0.0680268 0.482109 0.277723 0.26447 -0.591302 -0.169473 0.459613 -0.26883 -0.190778 1.099 1 2.26559e-239 285.36 1.278e-236 1.97692 1.097 0.000299992 0.933312 0.61955 0.6475 0.391211 1.97729 125.354 81.8769 18.601 59.8762 0.00411132 0 -40 10
0.198 5.74246e-09 2.53881e-06 0.0447663 0.0447443 0.0120474 2.61021e-06 0.001154 0.0559579 0.000653259 0.0566066 0.847659 101.894 0.247237 0.701662 4.10629 0.0527631 0.0387386 0.961261 0.0198952 0.00422465 0.0191572 0.00406911 0.0051048 0.00584276 0.204192 0.23371 57.9516 -87.8933 125.513 15.9933 145.004 0.000149298 0.267065 192.943 0.310753 0.067394 0.00409451 0.000561501 0.00138225 0.986995 0.991737 -2.97018e-06 -85.6693 0.0929709 31198.5 300.051 0.983524 0.319147 0.774481 0.774476 9.99958 2.97997e-06 1.19198e-05 0.130454 0.970874 0.926182 -0.0132935 4.88954e-06 0.500094 -1.84492e-20 6.78588e-24 -1.84424e-20 0.00139496 0.997819 8.59172e-05 0.15253 2.85158 0.00139496 0.998414 0.638812 0.00103958 0.00187944 0.000859172 0.455683 0.00187944 0.432308 0.000126487 1.02 0.887246 0.534802 0.28545 1.71591e-07 3.05289e-09 2396.62 3294.39 -0.0679758 0.482109 0.277723 0.264428 -0.59131 -0.169473 0.459765 -0.268829 -0.19093 1.1 1 1.37415e-239 285.408 7.75377e-237 1.97717 1.098 0.000299992 0.932999 0.619629 0.646631 0.391255 1.97754 125.368 81.8846 18.6015 59.88 0.00411099 0 -40 10
0.199 5.77146e-09 2.53881e-06 0.0448815 0.0448596 0.0120474 2.62339e-06 0.001154 0.0561019 0.000653281 0.0567506 0.847681 101.894 0.247235 0.701687 4.10631 0.0527651 0.0387388 0.961261 0.0198952 0.00422467 0.0191572 0.00406912 0.00510482 0.00584278 0.204193 0.233711 57.9517 -87.8933 125.515 15.9933 145.004 0.000149266 0.267065 192.943 0.310754 0.067394 0.0040945 0.000561501 0.00138225 0.986995 0.991737 -2.97018e-06 -85.6693 0.0929709 31198.5 300.051 0.983524 0.319147 0.774319 0.774315 9.99958 2.97997e-06 1.19198e-05 0.130454 0.970913 0.926203 -0.0132935 4.88954e-06 0.500095 -1.84503e-20 6.78629e-24 -1.84435e-20 0.00139496 0.997819 8.59172e-05 0.15253 2.85158 0.00139496 0.99841 0.638938 0.00103959 0.00187944 0.000859172 0.455683 0.00187944 0.432319 0.00012649 1.02 0.887245 0.534802 0.28545 1.71591e-07 3.05289e-09 2396.6 3293.71 -0.067925 0.482109 0.277722 0.264385 -0.591317 -0.169473 0.459916 -0.268829 -0.191082 1.101 1 8.33466e-240 285.456 4.70429e-237 1.97742 1.099 0.000299992 0.932688 0.619708 0.645765 0.391298 1.97779 125.381 81.8923 18.6019 59.8838 0.00411065 0 -40 10
0.2 5.80045e-09 2.53881e-06 0.0449966 0.0449749 0.0120474 2.63657e-06 0.001154 0.0562458 0.000653303 0.0568945 0.847704 101.894 0.247233 0.701713 4.10633 0.0527672 0.0387389 0.961261 0.0198952 0.00422469 0.0191572 0.00406914 0.00510485 0.0058428 0.204194 0.233712 57.9518 -87.8933 125.518 15.9933 145.004 0.000149235 0.267065 192.943 0.310754 0.067394 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97017e-06 -85.6693 0.0929708 31198.5 300.052 0.983524 0.319147 0.774158 0.774154 9.99958 2.97997e-06 1.19198e-05 0.130454 0.970953 0.926224 -0.0132935 4.88954e-06 0.500096 -1.84515e-20 6.78671e-24 -1.84447e-20 0.00139495 0.997819 8.59171e-05 0.15253 2.85158 0.00139495 0.998406 0.639064 0.0010396 0.00187944 0.000859171 0.455683 0.00187944 0.432331 0.000126493 1.02 0.887245 0.534802 0.28545 1.71591e-07 3.05288e-09 2396.59 3293.02 -0.0678744 0.482109 0.277722 0.264343 -0.591325 -0.169473 0.460067 -0.268828 -0.191234 1.102 1 5.05522e-240 285.504 2.85414e-237 1.97768 1.1 0.000299992 0.932377 0.619787 0.644902 0.391341 1.97804 125.395 81.9 18.6024 59.8875 0.00411032 0 -40 10
0.201 5.82944e-09 2.53881e-06 0.0451116 0.04509 0.0120473 2.64975e-06 0.001154 0.0563895 0.000653324 0.0570382 0.847727 101.894 0.247231 0.701739 4.10634 0.0527692 0.0387391 0.961261 0.0198951 0.00422471 0.0191572 0.00406916 0.00510487 0.00584283 0.204195 0.233713 57.9518 -87.8933 125.521 15.9932 145.004 0.000149204 0.267064 192.943 0.310754 0.0673941 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97016e-06 -85.6693 0.0929708 31198.5 300.052 0.983524 0.319147 0.773998 0.773993 9.99958 2.97996e-06 1.19197e-05 0.130454 0.970992 0.926244 -0.0132935 4.88953e-06 0.500097 -1.84526e-20 6.78713e-24 -1.84458e-20 0.00139495 0.997819 8.59171e-05 0.15253 2.85158 0.00139495 0.998403 0.63919 0.00103961 0.00187944 0.000859171 0.455683 0.00187944 0.432342 0.000126496 1.02 0.887245 0.534802 0.28545 1.71591e-07 3.05288e-09 2396.57 3292.34 -0.067824 0.482109 0.277722 0.264301 -0.591333 -0.169473 0.460217 -0.268828 -0.191385 1.103 1 3.06615e-240 285.552 1.73163e-237 1.97793 1.101 0.000299992 0.932067 0.619866 0.644041 0.391385 1.9783 125.408 81.9076 18.6028 59.8912 0.00410999 0 -40 10
0.202 5.85844e-09 2.53881e-06 0.0452265 0.0452051 0.0120473 2.66293e-06 0.001154 0.0565332 0.000653346 0.0571819 0.84775 101.894 0.247229 0.701765 4.10636 0.0527713 0.0387393 0.961261 0.0198951 0.00422473 0.0191571 0.00406917 0.0051049 0.00584285 0.204196 0.233714 57.9519 -87.8933 125.524 15.9932 145.004 0.000149174 0.267064 192.943 0.310754 0.0673941 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97016e-06 -85.6694 0.0929707 31198.6 300.053 0.983524 0.319147 0.773838 0.773833 9.99958 2.97996e-06 1.19197e-05 0.130455 0.971031 0.926265 -0.0132935 4.88953e-06 0.500098 -1.84538e-20 6.78755e-24 -1.8447e-20 0.00139495 0.997819 8.5917e-05 0.15253 2.85158 0.00139495 0.998399 0.639316 0.00103962 0.00187943 0.00085917 0.455683 0.00187944 0.432353 0.000126499 1.02 0.887245 0.534803 0.28545 1.71591e-07 3.05287e-09 2396.56 3291.66 -0.0677737 0.482109 0.277721 0.264258 -0.591341 -0.169473 0.460367 -0.268827 -0.191535 1.104 1 1.85971e-240 285.599 1.0506e-237 1.97818 1.102 0.000299992 0.931758 0.619945 0.643182 0.391428 1.97855 125.422 81.9153 18.6033 59.8949 0.00410967 0 -40 10
0.203 5.88743e-09 2.53881e-06 0.0453414 0.04532 0.0120473 2.6761e-06 0.001154 0.0566767 0.000653367 0.0573255 0.847774 101.894 0.247227 0.701791 4.10638 0.0527733 0.0387394 0.961261 0.0198951 0.00422475 0.0191571 0.00406919 0.00510492 0.00584287 0.204197 0.233715 57.9519 -87.8933 125.527 15.9932 145.004 0.000149143 0.267064 192.943 0.310755 0.0673941 0.0040945 0.000561499 0.00138225 0.986995 0.991737 -2.97015e-06 -85.6694 0.0929707 31198.6 300.053 0.983524 0.319147 0.773678 0.773674 9.99958 2.97996e-06 1.19197e-05 0.130455 0.97107 0.926285 -0.0132935 4.88953e-06 0.500098 -1.84549e-20 6.78796e-24 -1.84481e-20 0.00139495 0.997819 8.5917e-05 0.15253 2.85158 0.00139495 0.998395 0.639441 0.00103963 0.00187943 0.00085917 0.455684 0.00187943 0.432364 0.000126503 1.02 0.887245 0.534803 0.285449 1.71591e-07 3.05287e-09 2396.54 3290.98 -0.0677236 0.482109 0.277721 0.264217 -0.591348 -0.169473 0.460517 -0.268827 -0.191685 1.105 1 1.12797e-240 285.647 6.37406e-238 1.97843 1.103 0.000299992 0.931451 0.620024 0.642327 0.391471 1.9788 125.435 81.9229 18.6037 59.8987 0.00410934 0 -40 10
0.204 5.91642e-09 2.53881e-06 0.0454561 0.0454349 0.0120473 2.68928e-06 0.001154 0.0568201 0.000653389 0.0574689 0.847797 101.894 0.247225 0.701817 4.1064 0.0527754 0.0387396 0.96126 0.0198951 0.00422477 0.0191571 0.0040692 0.00510495 0.0058429 0.204198 0.233716 57.952 -87.8933 125.529 15.9931 145.004 0.000149112 0.267064 192.943 0.310755 0.0673942 0.00409449 0.000561499 0.00138225 0.986995 0.991737 -2.97014e-06 -85.6694 0.0929706 31198.6 300.054 0.983524 0.319147 0.77352 0.773515 9.99958 2.97995e-06 1.19197e-05 0.130455 0.971109 0.926306 -0.0132935 4.88953e-06 0.500099 -1.8456e-20 6.78838e-24 -1.84493e-20 0.00139495 0.997819 8.5917e-05 0.15253 2.85158 0.00139495 0.998391 0.639567 0.00103964 0.00187943 0.00085917 0.455684 0.00187943 0.432375 0.000126506 1.02 0.887245 0.534803 0.285449 1.71591e-07 3.05287e-09 2396.52 3290.31 -0.0676736 0.482109 0.277721 0.264175 -0.591356 -0.169473 0.460665 -0.268826 -0.191834 1.106 1 6.8415e-241 285.694 3.86719e-238 1.97868 1.104 0.000299992 0.931144 0.620102 0.641474 0.391514 1.97905 125.449 81.9304 18.6042 59.9023 0.00410901 0 -40 10
0.205 5.94541e-09 2.53881e-06 0.0455707 0.0455497 0.0120473 2.70246e-06 0.001154 0.0569634 0.00065341 0.0576122 0.84782 101.894 0.247223 0.701843 4.10642 0.0527775 0.0387398 0.96126 0.019895 0.00422479 0.0191571 0.00406922 0.00510497 0.00584292 0.204199 0.233717 57.952 -87.8933 125.532 15.9931 145.004 0.000149082 0.267064 192.943 0.310755 0.0673942 0.00409449 0.000561499 0.00138225 0.986995 0.991737 -2.97014e-06 -85.6694 0.0929706 31198.6 300.054 0.983524 0.319147 0.773361 0.773357 9.99958 2.97995e-06 1.19197e-05 0.130455 0.971148 0.926326 -0.0132935 4.88952e-06 0.5001 -1.84572e-20 6.78879e-24 -1.84504e-20 0.00139495 0.997819 8.59169e-05 0.15253 2.85158 0.00139495 0.998387 0.639693 0.00103965 0.00187943 0.000859169 0.455684 0.00187943 0.432386 0.000126509 1.02 0.887245 0.534803 0.285449 1.7159e-07 3.05286e-09 2396.51 3289.63 -0.0676238 0.482109 0.27772 0.264133 -0.591364 -0.169473 0.460814 -0.268826 -0.191983 1.107 1 4.14958e-241 285.741 2.34626e-238 1.97893 1.105 0.000299992 0.930839 0.620181 0.640623 0.391557 1.9793 125.462 81.938 18.6046 59.906 0.00410869 0 -40 10
0.206 5.9744e-09 2.53881e-06 0.0456853 0.0456644 0.0120473 2.71564e-06 0.001154 0.0571066 0.000653431 0.0577554 0.847844 101.894 0.24722 0.70187 4.10644 0.0527796 0.03874 0.96126 0.019895 0.00422481 0.0191571 0.00406924 0.005105 0.00584295 0.2042 0.233718 57.9521 -87.8933 125.535 15.993 145.004 0.000149051 0.267064 192.943 0.310755 0.0673942 0.00409449 0.000561498 0.00138224 0.986995 0.991737 -2.97013e-06 -85.6694 0.0929705 31198.6 300.055 0.983524 0.319147 0.773203 0.773199 9.99958 2.97995e-06 1.19197e-05 0.130455 0.971187 0.926346 -0.0132935 4.88952e-06 0.500101 -1.84583e-20 6.78921e-24 -1.84515e-20 0.00139495 0.997819 8.59169e-05 0.15253 2.85158 0.00139495 0.998384 0.639818 0.00103966 0.00187943 0.000859169 0.455684 0.00187943 0.432397 0.000126512 1.02 0.887245 0.534803 0.285449 1.7159e-07 3.05286e-09 2396.49 3288.96 -0.0675742 0.482109 0.27772 0.264092 -0.591371 -0.169473 0.460961 -0.268825 -0.192132 1.108 1 2.51685e-241 285.788 1.42349e-238 1.97919 1.106 0.000299992 0.930534 0.620259 0.639775 0.3916 1.97955 125.476 81.9455 18.6051 59.9097 0.00410836 0 -40 10
0.207 6.0034e-09 2.53881e-06 0.0457997 0.045779 0.0120473 2.72882e-06 0.001154 0.0572496 0.000653451 0.0578985 0.847867 101.894 0.247218 0.701897 4.10646 0.0527817 0.0387401 0.96126 0.019895 0.00422483 0.019157 0.00406925 0.00510502 0.00584297 0.204201 0.233719 57.9522 -87.8933 125.537 15.993 145.004 0.000149021 0.267064 192.943 0.310756 0.0673942 0.00409449 0.000561498 0.00138224 0.986995 0.991737 -2.97013e-06 -85.6694 0.0929705 31198.6 300.056 0.983524 0.319147 0.773046 0.773041 9.99958 2.97995e-06 1.19197e-05 0.130456 0.971225 0.926367 -0.0132935 4.88952e-06 0.500102 -1.84595e-20 6.78962e-24 -1.84527e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.99838 0.639944 0.00103967 0.00187943 0.000859168 0.455684 0.00187943 0.432408 0.000126515 1.02 0.887245 0.534803 0.285449 1.7159e-07 3.05285e-09 2396.48 3288.29 -0.0675248 0.482109 0.27772 0.26405 -0.591379 -0.169473 0.461109 -0.268824 -0.192279 1.109 1 1.52655e-241 285.834 8.63641e-239 1.97944 1.107 0.000299992 0.93023 0.620337 0.638929 0.391643 1.9798 125.489 81.953 18.6055 59.9134 0.00410804 0 -40 10
0.208 6.03239e-09 2.53881e-06 0.0459141 0.0458935 0.0120473 2.74199e-06 0.001154 0.0573926 0.000653472 0.0580415 0.847891 101.894 0.247216 0.701924 4.10647 0.0527839 0.0387403 0.96126 0.019895 0.00422485 0.019157 0.00406927 0.00510505 0.005843 0.204202 0.23372 57.9522 -87.8933 125.54 15.993 145.004 0.000148991 0.267064 192.943 0.310756 0.0673943 0.00409449 0.000561498 0.00138224 0.986995 0.991737 -2.97012e-06 -85.6694 0.0929704 31198.6 300.056 0.983524 0.319147 0.772889 0.772884 9.99958 2.97994e-06 1.19197e-05 0.130456 0.971264 0.926387 -0.0132935 4.88952e-06 0.500103 -1.84606e-20 6.79004e-24 -1.84538e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.998376 0.640069 0.00103969 0.00187943 0.000859168 0.455684 0.00187943 0.432419 0.000126518 1.02 0.887244 0.534803 0.285449 1.7159e-07 3.05285e-09 2396.46 3287.63 -0.0674755 0.482109 0.277719 0.264009 -0.591387 -0.169473 0.461255 -0.268824 -0.192427 1.11 1 9.25897e-242 285.881 5.23976e-239 1.97969 1.108 0.000299992 0.929928 0.620416 0.638086 0.391686 1.98005 125.502 81.9605 18.606 59.917 0.00410772 0 -40 10
0.209 6.06138e-09 2.53881e-06 0.0460283 0.0460079 0.0120472 2.75517e-06 0.001154 0.0575354 0.000653493 0.0581843 0.847915 101.894 0.247214 0.701951 4.10649 0.052786 0.0387405 0.961259 0.0198949 0.00422488 0.019157 0.00406929 0.00510507 0.00584302 0.204203 0.233721 57.9523 -87.8933 125.543 15.9929 145.004 0.000148961 0.267064 192.944 0.310756 0.0673943 0.00409449 0.000561497 0.00138224 0.986995 0.991737 -2.97012e-06 -85.6694 0.0929704 31198.6 300.057 0.983524 0.319147 0.772733 0.772728 9.99958 2.97994e-06 1.19197e-05 0.130456 0.971302 0.926407 -0.0132935 4.88952e-06 0.500103 -1.84617e-20 6.79045e-24 -1.84549e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.998373 0.640195 0.0010397 0.00187943 0.000859168 0.455684 0.00187943 0.43243 0.000126521 1.02 0.887244 0.534803 0.285449 1.7159e-07 3.05285e-09 2396.44 3286.96 -0.0674264 0.482109 0.277719 0.263968 -0.591394 -0.169474 0.461402 -0.268823 -0.192574 1.111 1 5.61585e-242 285.928 3.17899e-239 1.97994 1.109 0.000299992 0.929626 0.620494 0.637246 0.391729 1.9803 125.516 81.968 18.6064 59.9206 0.0041074 0 -40 10
0.21 6.09037e-09 2.53881e-06 0.0461425 0.0461222 0.0120472 2.76835e-06 0.001154 0.0576782 0.000653513 0.0583271 0.847939 101.893 0.247212 0.701978 4.10651 0.0527882 0.0387407 0.961259 0.0198949 0.0042249 0.019157 0.00406931 0.0051051 0.00584305 0.204204 0.233722 57.9523 -87.8933 125.546 15.9929 145.004 0.000148931 0.267064 192.944 0.310756 0.0673943 0.00409449 0.000561497 0.00138224 0.986995 0.991737 -2.97011e-06 -85.6694 0.0929704 31198.6 300.057 0.983524 0.319147 0.772577 0.772572 9.99958 2.97994e-06 1.19197e-05 0.130456 0.97134 0.926427 -0.0132935 4.88951e-06 0.500104 -1.84628e-20 6.79086e-24 -1.84561e-20 0.00139495 0.997819 8.59167e-05 0.15253 2.85158 0.00139495 0.998369 0.64032 0.00103971 0.00187943 0.000859167 0.455684 0.00187943 0.432442 0.000126524 1.02 0.887244 0.534803 0.285449 1.7159e-07 3.05284e-09 2396.43 3286.3 -0.0673775 0.482109 0.277719 0.263927 -0.591402 -0.169474 0.461547 -0.268823 -0.19272 1.112 1 3.40618e-242 285.974 1.92871e-239 1.98019 1.11 0.000299992 0.929326 0.620572 0.636408 0.391772 1.98055 125.529 81.9754 18.6069 59.9243 0.00410708 0 -40 10
0.211 6.11936e-09 2.53881e-06 0.0462566 0.0462364 0.0120472 2.78153e-06 0.001154 0.0578208 0.000653533 0.0584697 0.847963 101.893 0.24721 0.702005 4.10653 0.0527903 0.0387409 0.961259 0.0198949 0.00422492 0.0191569 0.00406932 0.00510512 0.00584307 0.204205 0.233723 57.9524 -87.8933 125.548 15.9929 145.004 0.000148901 0.267063 192.944 0.310756 0.0673943 0.00409448 0.000561497 0.00138224 0.986995 0.991737 -2.9701e-06 -85.6694 0.0929703 31198.7 300.058 0.983524 0.319147 0.772422 0.772417 9.99958 2.97994e-06 1.19196e-05 0.130457 0.971378 0.926447 -0.0132935 4.88951e-06 0.500105 -1.8464e-20 6.79128e-24 -1.84572e-20 0.00139495 0.997819 8.59167e-05 0.152529 2.85158 0.00139495 0.998365 0.640445 0.00103972 0.00187943 0.000859167 0.455684 0.00187943 0.432453 0.000126528 1.02 0.887244 0.534803 0.285449 1.7159e-07 3.05284e-09 2396.41 3285.64 -0.0673287 0.482109 0.277719 0.263886 -0.591409 -0.169474 0.461693 -0.268822 -0.192866 1.113 1 2.06595e-242 286.02 1.17016e-239 1.98043 1.111 0.000299992 0.929026 0.62065 0.635572 0.391814 1.9808 125.542 81.9829 18.6073 59.9279 0.00410676 0 -40 10
0.212 6.14836e-09 2.53881e-06 0.0463706 0.0463505 0.0120472 2.79471e-06 0.001154 0.0579633 0.000653554 0.0586122 0.847987 101.893 0.247207 0.702033 4.10655 0.0527925 0.0387411 0.961259 0.0198948 0.00422494 0.0191569 0.00406934 0.00510515 0.0058431 0.204206 0.233724 57.9525 -87.8933 125.551 15.9928 145.004 0.000148871 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986995 0.991737 -2.9701e-06 -85.6694 0.0929703 31198.7 300.058 0.983524 0.319147 0.772267 0.772262 9.99958 2.97993e-06 1.19196e-05 0.130457 0.971416 0.926467 -0.0132935 4.88951e-06 0.500106 -1.84651e-20 6.79169e-24 -1.84583e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.998362 0.640571 0.00103973 0.00187943 0.000859166 0.455685 0.00187943 0.432464 0.000126531 1.02 0.887244 0.534803 0.285449 1.7159e-07 3.05284e-09 2396.4 3284.98 -0.0672801 0.482109 0.277718 0.263845 -0.591417 -0.169474 0.461838 -0.268822 -0.193012 1.114 1 1.25306e-242 286.066 7.09941e-240 1.98068 1.112 0.000299992 0.928728 0.620727 0.634739 0.391857 1.98104 125.556 81.9902 18.6077 59.9315 0.00410644 0 -40 10
0.213 6.17735e-09 2.53881e-06 0.0464845 0.0464646 0.0120472 2.80788e-06 0.001154 0.0581056 0.000653574 0.0587546 0.848011 101.893 0.247205 0.702061 4.10657 0.0527947 0.0387412 0.961259 0.0198948 0.00422496 0.0191569 0.00406936 0.00510518 0.00584312 0.204207 0.233725 57.9525 -87.8933 125.554 15.9928 145.004 0.000148841 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986995 0.991737 -2.97009e-06 -85.6694 0.0929702 31198.7 300.059 0.983524 0.319147 0.772113 0.772108 9.99958 2.97993e-06 1.19196e-05 0.130457 0.971454 0.926486 -0.0132935 4.88951e-06 0.500107 -1.84662e-20 6.7921e-24 -1.84594e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.998358 0.640696 0.00103974 0.00187943 0.000859166 0.455685 0.00187943 0.432475 0.000126534 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05283e-09 2396.38 3284.33 -0.0672316 0.482109 0.277718 0.263804 -0.591424 -0.169474 0.461982 -0.268821 -0.193157 1.115 1 7.60022e-243 286.112 4.30724e-240 1.98093 1.113 0.000299992 0.92843 0.620805 0.633908 0.3919 1.98129 125.569 81.9976 18.6082 59.9351 0.00410613 0 -40 10
0.214 6.20634e-09 2.53881e-06 0.0465983 0.0465785 0.0120472 2.82106e-06 0.001154 0.0582479 0.000653593 0.0588969 0.848035 101.893 0.247203 0.702089 4.10659 0.0527969 0.0387414 0.961259 0.0198948 0.00422498 0.0191568 0.00406938 0.0051052 0.00584315 0.204208 0.233726 57.9526 -87.8933 125.556 15.9928 145.004 0.000148811 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986995 0.991737 -2.97009e-06 -85.6694 0.0929702 31198.7 300.06 0.983524 0.319147 0.771959 0.771954 9.99958 2.97993e-06 1.19196e-05 0.130457 0.971492 0.926506 -0.0132935 4.88951e-06 0.500108 -1.84673e-20 6.79251e-24 -1.84606e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.998355 0.640821 0.00103975 0.00187943 0.000859166 0.455685 0.00187943 0.432486 0.000126537 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05283e-09 2396.36 3283.67 -0.0671834 0.482108 0.277718 0.263764 -0.591432 -0.169474 0.462126 -0.26882 -0.193301 1.116 1 4.60977e-243 286.158 2.61322e-240 1.98118 1.114 0.000299991 0.928134 0.620883 0.63308 0.391942 1.98154 125.582 82.005 18.6086 59.9387 0.00410581 0 -40 10
0.215 6.23533e-09 2.53881e-06 0.046712 0.0466923 0.0120472 2.83424e-06 0.001154 0.05839 0.000653613 0.0590391 0.84806 101.893 0.247201 0.702117 4.10661 0.0527991 0.0387416 0.961258 0.0198948 0.004225 0.0191568 0.0040694 0.00510523 0.00584318 0.204209 0.233727 57.9526 -87.8934 125.559 15.9927 145.004 0.000148782 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561495 0.00138224 0.986995 0.991737 -2.97009e-06 -85.6694 0.0929702 31198.7 300.06 0.983524 0.319147 0.771806 0.771801 9.99958 2.97993e-06 1.19196e-05 0.130457 0.97153 0.926526 -0.0132935 4.88951e-06 0.500109 -1.84685e-20 6.79292e-24 -1.84617e-20 0.00139495 0.997819 8.59165e-05 0.152529 2.85157 0.00139495 0.998351 0.640946 0.00103977 0.00187943 0.000859165 0.455685 0.00187943 0.432497 0.00012654 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05283e-09 2396.35 3283.02 -0.0671352 0.482108 0.277717 0.263724 -0.591439 -0.169474 0.462269 -0.26882 -0.193445 1.117 1 2.79597e-243 286.203 1.58545e-240 1.98143 1.115 0.000299991 0.927838 0.62096 0.632254 0.391985 1.98179 125.595 82.0123 18.6091 59.9422 0.0041055 0 -40 10
0.216 6.26432e-09 2.53881e-06 0.0468257 0.0468061 0.0120471 2.84742e-06 0.001154 0.0585321 0.000653633 0.0591811 0.848084 101.893 0.247199 0.702145 4.10663 0.0528014 0.0387418 0.961258 0.0198947 0.00422503 0.0191568 0.00406941 0.00510526 0.0058432 0.20421 0.233728 57.9527 -87.8934 125.562 15.9927 145.004 0.000148752 0.267063 192.944 0.310757 0.0673945 0.00409448 0.000561495 0.00138223 0.986996 0.991737 -2.97008e-06 -85.6694 0.0929701 31198.7 300.061 0.983524 0.319147 0.771653 0.771648 9.99958 2.97993e-06 1.19196e-05 0.130458 0.971567 0.926545 -0.0132935 4.88951e-06 0.50011 -1.84696e-20 6.79333e-24 -1.84628e-20 0.00139495 0.997819 8.59165e-05 0.152529 2.85157 0.00139495 0.998348 0.641071 0.00103978 0.00187942 0.000859165 0.455685 0.00187943 0.432508 0.000126543 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05283e-09 2396.33 3282.37 -0.0670873 0.482108 0.277717 0.263683 -0.591447 -0.169474 0.462412 -0.268819 -0.193589 1.118 1 1.69584e-243 286.249 9.61896e-241 1.98168 1.116 0.000299991 0.927544 0.621038 0.631431 0.392027 1.98204 125.609 82.0196 18.6095 59.9458 0.00410518 0 -40 10
0.217 6.29331e-09 2.53881e-06 0.0469392 0.0469198 0.0120471 2.8606e-06 0.001154 0.058674 0.000653652 0.0593231 0.848109 101.893 0.247196 0.702173 4.10665 0.0528036 0.038742 0.961258 0.0198947 0.00422505 0.0191568 0.00406943 0.00510529 0.00584323 0.204211 0.233729 57.9528 -87.8934 125.564 15.9927 145.004 0.000148723 0.267063 192.944 0.310758 0.0673945 0.00409448 0.000561495 0.00138223 0.986996 0.991737 -2.97008e-06 -85.6694 0.0929701 31198.7 300.061 0.983524 0.319147 0.771501 0.771496 9.99958 2.97992e-06 1.19196e-05 0.130458 0.971605 0.926565 -0.0132935 4.88951e-06 0.500111 -1.84707e-20 6.79374e-24 -1.84639e-20 0.00139494 0.997819 8.59165e-05 0.152529 2.85157 0.00139494 0.998344 0.641196 0.00103979 0.00187942 0.000859165 0.455685 0.00187942 0.432519 0.000126547 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05282e-09 2396.32 3281.72 -0.0670395 0.482108 0.277717 0.263643 -0.591454 -0.169474 0.462554 -0.268818 -0.193732 1.119 1 1.02858e-243 286.294 5.83584e-241 1.98192 1.117 0.000299991 0.92725 0.621115 0.63061 0.392069 1.98228 125.622 82.0269 18.6099 59.9493 0.00410487 0 -40 10
0.218 6.3223e-09 2.53881e-06 0.0470527 0.0470333 0.0120471 2.87377e-06 0.001154 0.0588158 0.000653672 0.0594649 0.848134 101.893 0.247194 0.702202 4.10667 0.0528059 0.0387422 0.961258 0.0198947 0.00422507 0.0191567 0.00406945 0.00510531 0.00584326 0.204213 0.23373 57.9528 -87.8934 125.567 15.9926 145.004 0.000148694 0.267063 192.944 0.310758 0.0673945 0.00409447 0.000561495 0.00138223 0.986996 0.991737 -2.97007e-06 -85.6694 0.09297 31198.7 300.062 0.983524 0.319147 0.771349 0.771344 9.99958 2.97992e-06 1.19196e-05 0.130458 0.971642 0.926584 -0.0132935 4.88951e-06 0.500112 -1.84718e-20 6.79415e-24 -1.8465e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998341 0.641321 0.0010398 0.00187942 0.000859164 0.455685 0.00187942 0.43253 0.00012655 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05282e-09 2396.3 3281.08 -0.0669918 0.482108 0.277716 0.263603 -0.591461 -0.169474 0.462696 -0.268818 -0.193874 1.12 1 6.23864e-244 286.339 3.54062e-241 1.98217 1.118 0.000299991 0.926958 0.621192 0.629792 0.392112 1.98253 125.635 82.0341 18.6103 59.9529 0.00410456 0 -40 10
0.219 6.35129e-09 2.53881e-06 0.047166 0.0471468 0.0120471 2.88695e-06 0.001154 0.0589575 0.000653691 0.0596066 0.848158 101.893 0.247192 0.702231 4.1067 0.0528081 0.0387424 0.961258 0.0198947 0.00422509 0.0191567 0.00406947 0.00510534 0.00584328 0.204214 0.233731 57.9529 -87.8934 125.569 15.9926 145.004 0.000148665 0.267063 192.944 0.310758 0.0673945 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.97007e-06 -85.6694 0.09297 31198.7 300.063 0.983524 0.319147 0.771198 0.771193 9.99958 2.97992e-06 1.19196e-05 0.130458 0.971679 0.926604 -0.0132935 4.88951e-06 0.500112 -1.84729e-20 6.79456e-24 -1.84661e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998338 0.641446 0.00103981 0.00187942 0.000859164 0.455685 0.00187942 0.432541 0.000126553 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05282e-09 2396.28 3280.44 -0.0669444 0.482108 0.277716 0.263564 -0.591469 -0.169474 0.462837 -0.268817 -0.194017 1.121 1 3.78393e-244 286.384 2.1481e-241 1.98242 1.119 0.000299991 0.926666 0.62127 0.628976 0.392154 1.98278 125.648 82.0414 18.6108 59.9564 0.00410425 0 -40 10
0.22 6.38028e-09 2.53881e-06 0.0472793 0.0472602 0.0120471 2.90013e-06 0.001154 0.0590991 0.00065371 0.0597482 0.848183 101.893 0.24719 0.702259 4.10672 0.0528104 0.0387426 0.961257 0.0198946 0.00422512 0.0191567 0.00406949 0.00510537 0.00584331 0.204215 0.233732 57.9529 -87.8934 125.572 15.9926 145.005 0.000148636 0.267063 192.944 0.310758 0.0673945 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.97006e-06 -85.6694 0.09297 31198.7 300.063 0.983524 0.319147 0.771047 0.771042 9.99958 2.97992e-06 1.19196e-05 0.130459 0.971716 0.926623 -0.0132935 4.88951e-06 0.500113 -1.8474e-20 6.79497e-24 -1.84672e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998334 0.641571 0.00103982 0.00187942 0.000859164 0.455685 0.00187942 0.432552 0.000126556 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05282e-09 2396.27 3279.8 -0.0668971 0.482108 0.277716 0.263524 -0.591476 -0.169474 0.462978 -0.268816 -0.194158 1.122 1 2.29507e-244 286.429 1.30325e-241 1.98266 1.12 0.000299991 0.926375 0.621347 0.628163 0.392196 1.98302 125.661 82.0486 18.6112 59.9599 0.00410394 0 -40 10
0.221 6.40928e-09 2.53881e-06 0.0473925 0.0473735 0.0120471 2.91331e-06 0.001154 0.0592406 0.000653729 0.0598897 0.848208 101.893 0.247187 0.702288 4.10674 0.0528127 0.0387428 0.961257 0.0198946 0.00422514 0.0191567 0.00406951 0.0051054 0.00584334 0.204216 0.233734 57.953 -87.8934 125.575 15.9925 145.005 0.000148607 0.267063 192.944 0.310758 0.0673946 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.97006e-06 -85.6694 0.0929699 31198.8 300.064 0.983524 0.319147 0.770897 0.770892 9.99958 2.97992e-06 1.19196e-05 0.130459 0.971753 0.926642 -0.0132935 4.88951e-06 0.500114 -1.84751e-20 6.79538e-24 -1.84684e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998331 0.641696 0.00103984 0.00187942 0.000859163 0.455685 0.00187942 0.432563 0.000126559 1.02 0.887244 0.534803 0.285448 1.71589e-07 3.05282e-09 2396.25 3279.16 -0.0668499 0.482108 0.277715 0.263484 -0.591483 -0.169474 0.463119 -0.268816 -0.194299 1.123 1 1.39203e-244 286.474 7.90685e-242 1.98291 1.121 0.000299991 0.926086 0.621424 0.627351 0.392238 1.98327 125.674 82.0557 18.6116 59.9634 0.00410363 0 -40 10
0.222 6.43827e-09 2.53881e-06 0.0475055 0.0474867 0.0120471 2.92648e-06 0.001154 0.0593819 0.000653748 0.0600311 0.848233 101.893 0.247185 0.702318 4.10676 0.052815 0.038743 0.961257 0.0198946 0.00422516 0.0191566 0.00406953 0.00510543 0.00584337 0.204217 0.233735 57.9531 -87.8934 125.577 15.9925 145.005 0.000148578 0.267063 192.944 0.310758 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97006e-06 -85.6694 0.0929699 31198.8 300.065 0.983524 0.319147 0.770747 0.770742 9.99958 2.97991e-06 1.19196e-05 0.130459 0.97179 0.926661 -0.0132935 4.88951e-06 0.500115 -1.84763e-20 6.79579e-24 -1.84695e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998327 0.641821 0.00103985 0.00187942 0.000859163 0.455685 0.00187942 0.432574 0.000126563 1.02 0.887244 0.534803 0.285448 1.71588e-07 3.05282e-09 2396.23 3278.52 -0.0668029 0.482108 0.277715 0.263445 -0.591491 -0.169475 0.463259 -0.268815 -0.19444 1.124 1 8.44309e-245 286.518 4.79709e-242 1.98316 1.122 0.000299991 0.925797 0.621501 0.626543 0.392281 1.98351 125.688 82.0629 18.6121 59.9669 0.00410333 0 -40 10
0.223 6.46726e-09 2.53881e-06 0.0476185 0.0475998 0.0120471 2.93966e-06 0.001154 0.0595232 0.000653767 0.0601723 0.848258 101.893 0.247183 0.702347 4.10678 0.0528174 0.0387432 0.961257 0.0198945 0.00422519 0.0191566 0.00406954 0.00510546 0.0058434 0.204218 0.233736 57.9531 -87.8934 125.58 15.9924 145.005 0.000148549 0.267063 192.944 0.310759 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97005e-06 -85.6694 0.0929699 31198.8 300.065 0.983524 0.319147 0.770598 0.770593 9.99958 2.97991e-06 1.19195e-05 0.130459 0.971827 0.926681 -0.0132935 4.88951e-06 0.500116 -1.84774e-20 6.79619e-24 -1.84706e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998324 0.641946 0.00103986 0.00187942 0.000859163 0.455686 0.00187942 0.432585 0.000126566 1.02 0.887244 0.534803 0.285448 1.71588e-07 3.05281e-09 2396.22 3277.89 -0.0667561 0.482108 0.277715 0.263405 -0.591498 -0.169475 0.463398 -0.268814 -0.19458 1.125 1 5.12099e-245 286.563 2.91039e-242 1.9834 1.123 0.000299991 0.925509 0.621577 0.625736 0.392323 1.98376 125.701 82.07 18.6125 59.9704 0.00410302 0 -40 10
0.224 6.49625e-09 2.53881e-06 0.0477314 0.0477128 0.012047 2.95284e-06 0.001154 0.0596643 0.000653786 0.0603135 0.848284 101.893 0.24718 0.702377 4.1068 0.0528197 0.0387434 0.961257 0.0198945 0.00422521 0.0191566 0.00406956 0.00510549 0.00584342 0.204219 0.233737 57.9532 -87.8934 125.582 15.9924 145.005 0.00014852 0.267062 192.945 0.310759 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97005e-06 -85.6694 0.0929698 31198.8 300.066 0.983524 0.319147 0.770449 0.770444 9.99958 2.97991e-06 1.19195e-05 0.13046 0.971863 0.9267 -0.0132935 4.88951e-06 0.500117 -1.84785e-20 6.7966e-24 -1.84717e-20 0.00139494 0.997819 8.59162e-05 0.152529 2.85157 0.00139494 0.998321 0.642071 0.00103987 0.00187942 0.000859162 0.455686 0.00187942 0.432596 0.000126569 1.02 0.887244 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.2 3277.25 -0.0667094 0.482108 0.277714 0.263366 -0.591505 -0.169475 0.463537 -0.268814 -0.19472 1.126 1 3.10604e-245 286.607 1.76573e-242 1.98365 1.124 0.000299991 0.925223 0.621654 0.624932 0.392365 1.984 125.714 82.0772 18.6129 59.9738 0.00410271 0 -40 10
0.225 6.52524e-09 2.53881e-06 0.0478443 0.0478257 0.012047 2.96602e-06 0.001154 0.0598053 0.000653804 0.0604545 0.848309 101.893 0.247178 0.702406 4.10683 0.0528221 0.0387436 0.961256 0.0198945 0.00422524 0.0191565 0.00406958 0.00510551 0.00584345 0.204221 0.233738 57.9532 -87.8934 125.585 15.9924 145.005 0.000148492 0.267062 192.945 0.310759 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97005e-06 -85.6694 0.0929698 31198.8 300.066 0.983524 0.319147 0.770301 0.770296 9.99958 2.97991e-06 1.19195e-05 0.13046 0.9719 0.926719 -0.0132935 4.88951e-06 0.500118 -1.84796e-20 6.79701e-24 -1.84728e-20 0.00139494 0.997819 8.59162e-05 0.152529 2.85157 0.00139494 0.998318 0.642196 0.00103989 0.00187942 0.000859162 0.455686 0.00187942 0.432607 0.000126572 1.02 0.887244 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.19 3276.62 -0.0666629 0.482108 0.277714 0.263327 -0.591512 -0.169475 0.463676 -0.268813 -0.194859 1.127 1 1.88391e-245 286.651 1.07127e-242 1.98389 1.125 0.000299991 0.924937 0.621731 0.624131 0.392407 1.98425 125.727 82.0843 18.6133 59.9773 0.00410241 0 -40 10
0.226 6.55423e-09 2.53881e-06 0.047957 0.0479386 0.012047 2.97919e-06 0.001154 0.0599462 0.000653823 0.0605954 0.848334 101.893 0.247176 0.702436 4.10685 0.0528244 0.0387438 0.961256 0.0198945 0.00422526 0.0191565 0.0040696 0.00510554 0.00584348 0.204222 0.233739 57.9533 -87.8934 125.588 15.9923 145.005 0.000148463 0.267062 192.945 0.310759 0.0673947 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97004e-06 -85.6695 0.0929698 31198.8 300.067 0.983524 0.319147 0.770153 0.770148 9.99958 2.97991e-06 1.19195e-05 0.13046 0.971936 0.926737 -0.0132935 4.88952e-06 0.500119 -1.84807e-20 6.79741e-24 -1.84739e-20 0.00139494 0.997819 8.59162e-05 0.152529 2.85157 0.00139494 0.998314 0.64232 0.0010399 0.00187942 0.000859162 0.455686 0.00187942 0.432618 0.000126575 1.02 0.887244 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.17 3275.99 -0.0666165 0.482108 0.277714 0.263288 -0.59152 -0.169475 0.463814 -0.268812 -0.194998 1.128 1 1.14265e-245 286.695 6.49937e-243 1.98414 1.126 0.000299991 0.924652 0.621807 0.623332 0.392449 1.98449 125.74 82.0913 18.6137 59.9807 0.00410211 0 -40 10
0.227 6.58322e-09 2.53881e-06 0.0480696 0.0480513 0.012047 2.99237e-06 0.001154 0.060087 0.000653841 0.0607362 0.84836 101.893 0.247173 0.702466 4.10687 0.0528268 0.0387441 0.961256 0.0198944 0.00422528 0.0191565 0.00406962 0.00510557 0.00584351 0.204223 0.23374 57.9533 -87.8934 125.59 15.9923 145.005 0.000148435 0.267062 192.945 0.310759 0.0673947 0.00409446 0.000561492 0.00138223 0.986996 0.991737 -2.97004e-06 -85.6695 0.0929698 31198.8 300.068 0.983524 0.319147 0.770006 0.770001 9.99958 2.97991e-06 1.19195e-05 0.13046 0.971972 0.926756 -0.0132935 4.88952e-06 0.50012 -1.84818e-20 6.79782e-24 -1.8475e-20 0.00139494 0.997819 8.59162e-05 0.152528 2.85157 0.00139494 0.998311 0.642445 0.00103991 0.00187942 0.000859162 0.455686 0.00187942 0.432629 0.000126579 1.02 0.887244 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.15 3275.37 -0.0665703 0.482108 0.277713 0.263249 -0.591527 -0.169475 0.463951 -0.268812 -0.195137 1.129 1 6.93051e-246 286.739 3.94316e-243 1.98438 1.127 0.000299991 0.924368 0.621884 0.622535 0.39249 1.98474 125.753 82.0984 18.6142 59.9841 0.00410181 0 -40 10
0.228 6.61221e-09 2.53881e-06 0.0481821 0.048164 0.012047 3.00555e-06 0.001154 0.0602277 0.000653859 0.0608769 0.848386 101.893 0.247171 0.702496 4.10689 0.0528292 0.0387443 0.961256 0.0198944 0.00422531 0.0191565 0.00406964 0.0051056 0.00584354 0.204224 0.233742 57.9534 -87.8934 125.593 15.9923 145.005 0.000148407 0.267062 192.945 0.310759 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97004e-06 -85.6695 0.0929697 31198.8 300.068 0.983524 0.319147 0.769859 0.769854 9.99958 2.9799e-06 1.19195e-05 0.130461 0.972009 0.926775 -0.0132935 4.88952e-06 0.500121 -1.84829e-20 6.79822e-24 -1.84761e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998308 0.642569 0.00103992 0.00187942 0.000859161 0.455686 0.00187942 0.43264 0.000126582 1.02 0.887244 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.14 3274.74 -0.0665243 0.482108 0.277713 0.263211 -0.591534 -0.169475 0.464088 -0.268811 -0.195275 1.13 1 4.20356e-246 286.783 2.39231e-243 1.98463 1.128 0.000299991 0.924085 0.62196 0.62174 0.392532 1.98498 125.766 82.1054 18.6146 59.9876 0.0041015 0 -40 10
0.229 6.6412e-09 2.53881e-06 0.0482946 0.0482765 0.012047 3.01873e-06 0.001154 0.0603683 0.000653877 0.0610175 0.848411 101.893 0.247168 0.702526 4.10691 0.0528316 0.0387445 0.961256 0.0198944 0.00422533 0.0191564 0.00406966 0.00510563 0.00584357 0.204225 0.233743 57.9535 -87.8934 125.595 15.9922 145.005 0.000148378 0.267062 192.945 0.310759 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97003e-06 -85.6695 0.0929697 31198.8 300.069 0.983524 0.319147 0.769713 0.769708 9.99958 2.9799e-06 1.19195e-05 0.130461 0.972045 0.926794 -0.0132935 4.88952e-06 0.500122 -1.84839e-20 6.79863e-24 -1.84771e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998305 0.642694 0.00103993 0.00187942 0.000859161 0.455686 0.00187942 0.432651 0.000126585 1.02 0.887244 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.12 3274.12 -0.0664784 0.482108 0.277713 0.263172 -0.591541 -0.169475 0.464225 -0.26881 -0.195412 1.131 1 2.54959e-246 286.826 1.45141e-243 1.98487 1.129 0.000299991 0.923803 0.622037 0.620948 0.392574 1.98522 125.779 82.1124 18.615 59.991 0.0041012 0 -40 10
0.23 6.67019e-09 2.53881e-06 0.048407 0.048389 0.012047 3.0319e-06 0.001154 0.0605087 0.000653895 0.061158 0.848437 101.893 0.247166 0.702557 4.10694 0.052834 0.0387447 0.961255 0.0198943 0.00422536 0.0191564 0.00406968 0.00510567 0.0058436 0.204227 0.233744 57.9535 -87.8934 125.598 15.9922 145.005 0.00014835 0.267062 192.945 0.31076 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97003e-06 -85.6695 0.0929697 31198.8 300.07 0.983524 0.319147 0.769567 0.769562 9.99958 2.9799e-06 1.19195e-05 0.130461 0.97208 0.926812 -0.0132935 4.88952e-06 0.500123 -1.8485e-20 6.79903e-24 -1.84782e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998301 0.642819 0.00103995 0.00187942 0.000859161 0.455686 0.00187942 0.432662 0.000126588 1.02 0.887245 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.11 3273.5 -0.0664326 0.482108 0.277712 0.263134 -0.591548 -0.169475 0.464361 -0.268809 -0.195549 1.132 1 1.5464e-246 286.87 8.80564e-244 1.98511 1.13 0.000299991 0.923522 0.622113 0.620158 0.392616 1.98547 125.792 82.1194 18.6154 59.9944 0.00410091 0 -40 10
0.231 6.69918e-09 2.53881e-06 0.0485192 0.0485014 0.012047 3.04508e-06 0.001154 0.060649 0.000653913 0.0612984 0.848463 101.893 0.247164 0.702588 4.10696 0.0528364 0.0387449 0.961255 0.0198943 0.00422538 0.0191564 0.0040697 0.0051057 0.00584363 0.204228 0.233745 57.9536 -87.8934 125.6 15.9922 145.005 0.000148322 0.267062 192.945 0.31076 0.0673947 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97003e-06 -85.6695 0.0929697 31198.8 300.07 0.983524 0.319147 0.769421 0.769417 9.99958 2.9799e-06 1.19195e-05 0.130461 0.972116 0.926831 -0.0132935 4.88953e-06 0.500124 -1.84861e-20 6.79944e-24 -1.84793e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998298 0.642943 0.00103996 0.00187942 0.000859161 0.455686 0.00187942 0.432673 0.000126592 1.02 0.887245 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.09 3272.88 -0.0663871 0.482108 0.277712 0.263095 -0.591555 -0.169475 0.464497 -0.268808 -0.195686 1.133 1 9.37942e-247 286.913 5.34235e-244 1.98536 1.131 0.000299991 0.923242 0.622189 0.619371 0.392657 1.98571 125.805 82.1264 18.6158 59.9978 0.00410061 0 -40 10
0.232 6.72817e-09 2.53881e-06 0.0486314 0.0486137 0.0120469 3.05826e-06 0.001154 0.0607893 0.000653931 0.0614386 0.848489 101.893 0.247161 0.702618 4.10698 0.0528389 0.0387451 0.961255 0.0198943 0.00422541 0.0191563 0.00406972 0.00510573 0.00584366 0.204229 0.233746 57.9536 -87.8934 125.603 15.9921 145.005 0.000148294 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97002e-06 -85.6695 0.0929696 31198.8 300.071 0.983524 0.319147 0.769277 0.769272 9.99958 2.9799e-06 1.19195e-05 0.130462 0.972152 0.926849 -0.0132935 4.88953e-06 0.500125 -1.84872e-20 6.79984e-24 -1.84804e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998295 0.643067 0.00103997 0.00187942 0.00085916 0.455686 0.00187942 0.432684 0.000126595 1.02 0.887245 0.534803 0.285449 1.71588e-07 3.05281e-09 2396.07 3272.27 -0.0663416 0.482108 0.277712 0.263057 -0.591562 -0.169475 0.464632 -0.268808 -0.195822 1.134 1 5.68891e-247 286.956 3.24118e-244 1.9856 1.132 0.000299991 0.922963 0.622265 0.618586 0.392699 1.98595 125.818 82.1333 18.6162 60.0011 0.00410031 0 -40 10
0.233 6.75716e-09 2.53881e-06 0.0487435 0.0487259 0.0120469 3.07143e-06 0.001154 0.0609294 0.000653949 0.0615787 0.848515 101.893 0.247159 0.702649 4.10701 0.0528413 0.0387454 0.961255 0.0198942 0.00422543 0.0191563 0.00406975 0.00510576 0.00584369 0.20423 0.233748 57.9537 -87.8934 125.605 15.9921 145.005 0.000148266 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97002e-06 -85.6695 0.0929696 31198.8 300.072 0.983524 0.319147 0.769132 0.769128 9.99958 2.9799e-06 1.19195e-05 0.130462 0.972188 0.926868 -0.0132935 4.88953e-06 0.500126 -1.84883e-20 6.80024e-24 -1.84815e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998292 0.643192 0.00103999 0.00187942 0.00085916 0.455686 0.00187942 0.432695 0.000126598 1.02 0.887245 0.534803 0.285449 1.71587e-07 3.05281e-09 2396.06 3271.65 -0.0662964 0.482108 0.277711 0.263019 -0.591569 -0.169475 0.464767 -0.268807 -0.195957 1.135 1 3.4505e-247 286.999 1.96641e-244 1.98584 1.133 0.000299991 0.922685 0.622341 0.617803 0.392741 1.98619 125.831 82.1402 18.6166 60.0045 0.00410001 0 -40 10
0.234 6.78615e-09 2.53881e-06 0.0488555 0.048838 0.0120469 3.08461e-06 0.001154 0.0610694 0.000653966 0.0617188 0.848542 101.893 0.247156 0.70268 4.10703 0.0528438 0.0387456 0.961254 0.0198942 0.00422546 0.0191563 0.00406977 0.00510579 0.00584372 0.204232 0.233749 57.9538 -87.8934 125.608 15.9921 145.005 0.000148239 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97002e-06 -85.6695 0.0929696 31198.8 300.073 0.983524 0.319147 0.768988 0.768984 9.99958 2.9799e-06 1.19195e-05 0.130462 0.972223 0.926886 -0.0132935 4.88953e-06 0.500127 -1.84894e-20 6.80065e-24 -1.84826e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998289 0.643316 0.00104 0.00187942 0.00085916 0.455686 0.00187942 0.432706 0.000126601 1.02 0.887245 0.534803 0.28545 1.71587e-07 3.05281e-09 2396.04 3271.04 -0.0662512 0.482108 0.277711 0.262981 -0.591576 -0.169475 0.464901 -0.268806 -0.196093 1.136 1 2.09283e-247 287.042 1.19301e-244 1.98608 1.134 0.000299991 0.922408 0.622417 0.617022 0.392782 1.98644 125.844 82.1471 18.617 60.0079 0.00409972 0 -40 10
0.235 6.81514e-09 2.53881e-06 0.0489674 0.04895 0.0120469 3.09779e-06 0.001154 0.0612093 0.000653984 0.0618587 0.848568 101.893 0.247154 0.702712 4.10706 0.0528462 0.0387458 0.961254 0.0198942 0.00422548 0.0191562 0.00406979 0.00510582 0.00584375 0.204233 0.23375 57.9538 -87.8934 125.61 15.992 145.005 0.000148211 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97002e-06 -85.6695 0.0929696 31198.9 300.073 0.983524 0.319147 0.768845 0.76884 9.99958 2.97989e-06 1.19195e-05 0.130462 0.972258 0.926905 -0.0132935 4.88954e-06 0.500128 -1.84905e-20 6.80105e-24 -1.84837e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998286 0.64344 0.00104001 0.00187942 0.00085916 0.455686 0.00187942 0.432717 0.000126605 1.02 0.887245 0.534802 0.28545 1.71587e-07 3.05281e-09 2396.03 3270.43 -0.0662063 0.482108 0.277711 0.262943 -0.591583 -0.169475 0.465035 -0.268805 -0.196227 1.137 1 1.26937e-247 287.085 7.23795e-245 1.98633 1.135 0.000299991 0.922131 0.622492 0.616244 0.392824 1.98668 125.857 82.154 18.6175 60.0112 0.00409943 0 -40 10
0.236 6.84412e-09 2.53881e-06 0.0490792 0.0490619 0.0120469 3.11097e-06 0.001154 0.0613491 0.000654001 0.0619985 0.848594 101.893 0.247151 0.702743 4.10708 0.0528487 0.038746 0.961254 0.0198941 0.00422551 0.0191562 0.00406981 0.00510585 0.00584378 0.204234 0.233751 57.9539 -87.8934 125.613 15.992 145.005 0.000148184 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97001e-06 -85.6695 0.0929695 31198.9 300.074 0.983524 0.319147 0.768702 0.768697 9.99958 2.97989e-06 1.19195e-05 0.130463 0.972294 0.926923 -0.0132935 4.88954e-06 0.50013 -1.84915e-20 6.80145e-24 -1.84847e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998283 0.643565 0.00104002 0.00187941 0.00085916 0.455686 0.00187942 0.432728 0.000126608 1.02 0.887245 0.534802 0.28545 1.71587e-07 3.05281e-09 2396.01 3269.82 -0.0661615 0.482108 0.27771 0.262906 -0.59159 -0.169476 0.465169 -0.268805 -0.196362 1.138 1 7.6991e-248 287.128 4.39123e-245 1.98657 1.136 0.000299991 0.921856 0.622568 0.615468 0.392865 1.98692 125.87 82.1608 18.6179 60.0145 0.00409913 0 -40 10
0.237 6.87311e-09 2.53881e-06 0.049191 0.0491738 0.0120469 3.12414e-06 0.001154 0.0614887 0.000654018 0.0621381 0.848621 101.893 0.247149 0.702775 4.1071 0.0528512 0.0387463 0.961254 0.0198941 0.00422554 0.0191562 0.00406983 0.00510588 0.00584381 0.204235 0.233753 57.9539 -87.8934 125.615 15.9919 145.005 0.000148156 0.267062 192.945 0.31076 0.0673948 0.00409446 0.00056149 0.00138222 0.986996 0.991737 -2.97001e-06 -85.6695 0.0929695 31198.9 300.075 0.983524 0.319147 0.768559 0.768555 9.99958 2.97989e-06 1.19195e-05 0.130463 0.972329 0.926941 -0.0132935 4.88954e-06 0.500131 -1.84926e-20 6.80185e-24 -1.84858e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.99828 0.643689 0.00104004 0.00187941 0.000859159 0.455687 0.00187941 0.432738 0.000126611 1.02 0.887245 0.534802 0.28545 1.71587e-07 3.05281e-09 2395.99 3269.22 -0.0661168 0.482108 0.27771 0.262868 -0.591597 -0.169476 0.465302 -0.268804 -0.196496 1.139 1 4.66974e-248 287.17 2.66413e-245 1.98681 1.137 0.000299991 0.921582 0.622644 0.614694 0.392906 1.98716 125.883 82.1677 18.6183 60.0179 0.00409884 0 -40 10
0.238 6.9021e-09 2.53881e-06 0.0493026 0.0492855 0.0120469 3.13732e-06 0.001154 0.0616283 0.000654035 0.0622777 0.848647 101.893 0.247146 0.702807 4.10713 0.0528537 0.0387465 0.961254 0.0198941 0.00422556 0.0191562 0.00406985 0.00510592 0.00584385 0.204237 0.233754 57.954 -87.8934 125.618 15.9919 145.005 0.000148129 0.267062 192.945 0.31076 0.0673948 0.00409446 0.00056149 0.00138222 0.986996 0.991737 -2.97001e-06 -85.6695 0.0929695 31198.9 300.075 0.983524 0.319147 0.768417 0.768413 9.99958 2.97989e-06 1.19195e-05 0.130463 0.972364 0.926959 -0.0132935 4.88955e-06 0.500132 -1.84937e-20 6.80225e-24 -1.84869e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998277 0.643813 0.00104005 0.00187941 0.000859159 0.455687 0.00187941 0.432749 0.000126614 1.02 0.887245 0.534802 0.28545 1.71587e-07 3.05281e-09 2395.98 3268.61 -0.0660723 0.482108 0.27771 0.26283 -0.591604 -0.169476 0.465434 -0.268803 -0.196629 1.14 1 2.83234e-248 287.213 1.61631e-245 1.98705 1.138 0.00029999 0.921308 0.622719 0.613923 0.392948 1.9874 125.896 82.1745 18.6187 60.0212 0.00409855 0 -40 10
0.239 6.93109e-09 2.53881e-06 0.0494142 0.0493972 0.0120468 3.1505e-06 0.001154 0.0617677 0.000654052 0.0624172 0.848674 101.893 0.247144 0.702838 4.10715 0.0528563 0.0387467 0.961253 0.0198941 0.00422559 0.0191561 0.00406987 0.00510595 0.00584388 0.204238 0.233755 57.9541 -87.8934 125.62 15.9919 145.005 0.000148101 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991737 -2.97001e-06 -85.6695 0.0929695 31198.9 300.076 0.983524 0.319147 0.768276 0.768271 9.99958 2.97989e-06 1.19195e-05 0.130463 0.972399 0.926977 -0.0132935 4.88955e-06 0.500133 -1.84948e-20 6.80265e-24 -1.8488e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998274 0.643937 0.00104006 0.00187941 0.000859159 0.455687 0.00187941 0.43276 0.000126618 1.02 0.887246 0.534802 0.28545 1.71587e-07 3.05282e-09 2395.96 3268.01 -0.0660279 0.482108 0.27771 0.262793 -0.591611 -0.169476 0.465566 -0.268802 -0.196762 1.141 1 1.7179e-248 287.255 9.80607e-246 1.98729 1.139 0.00029999 0.921035 0.622795 0.613154 0.392989 1.98764 125.909 82.1812 18.6191 60.0245 0.00409826 0 -40 10
0.24 6.96008e-09 2.53881e-06 0.0495256 0.0495087 0.0120468 3.16367e-06 0.001154 0.0619071 0.000654069 0.0625565 0.848701 101.893 0.247141 0.70287 4.10718 0.0528588 0.038747 0.961253 0.019894 0.00422562 0.0191561 0.0040699 0.00510598 0.00584391 0.204239 0.233756 57.9541 -87.8934 125.623 15.9918 145.005 0.000148074 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991737 -2.97001e-06 -85.6695 0.0929695 31198.9 300.077 0.983524 0.319147 0.768135 0.76813 9.99958 2.97989e-06 1.19194e-05 0.130464 0.972433 0.926995 -0.0132935 4.88956e-06 0.500134 -1.84958e-20 6.80305e-24 -1.8489e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998271 0.644061 0.00104008 0.00187941 0.000859159 0.455687 0.00187941 0.432771 0.000126621 1.02 0.887246 0.534802 0.285451 1.71587e-07 3.05282e-09 2395.95 3267.41 -0.0659837 0.482108 0.277709 0.262756 -0.591618 -0.169476 0.465698 -0.268801 -0.196894 1.142 1 1.04196e-248 287.297 5.94927e-246 1.98753 1.14 0.00029999 0.920764 0.62287 0.612387 0.39303 1.98788 125.921 82.188 18.6195 60.0278 0.00409797 0 -40 10
0.241 6.98907e-09 2.53881e-06 0.049637 0.0496202 0.0120468 3.17685e-06 0.001154 0.0620463 0.000654086 0.0626958 0.848728 101.893 0.247139 0.702903 4.1072 0.0528614 0.0387472 0.961253 0.019894 0.00422564 0.0191561 0.00406992 0.00510602 0.00584394 0.204241 0.233758 57.9542 -87.8934 125.625 15.9918 145.005 0.000148047 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991737 -2.97e-06 -85.6695 0.0929694 31198.9 300.078 0.983524 0.319147 0.767994 0.76799 9.99958 2.97989e-06 1.19194e-05 0.130464 0.972468 0.927013 -0.0132935 4.88956e-06 0.500135 -1.84969e-20 6.80345e-24 -1.84901e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998268 0.644185 0.00104009 0.00187941 0.000859159 0.455687 0.00187941 0.432782 0.000126624 1.02 0.887246 0.534802 0.285451 1.71587e-07 3.05282e-09 2395.93 3266.81 -0.0659397 0.482108 0.277709 0.262719 -0.591625 -0.169476 0.465829 -0.2688 -0.197026 1.143 1 6.3198e-249 287.339 3.60938e-246 1.98777 1.141 0.00029999 0.920493 0.622945 0.611622 0.393071 1.98812 125.934 82.1948 18.6199 60.031 0.00409768 0 -40 10
0.242 7.01806e-09 2.53881e-06 0.0497483 0.0497316 0.0120468 3.19003e-06 0.001154 0.0621854 0.000654103 0.0628349 0.848755 101.893 0.247136 0.702935 4.10723 0.0528639 0.0387474 0.961253 0.019894 0.00422567 0.019156 0.00406994 0.00510605 0.00584397 0.204242 0.233759 57.9542 -87.8935 125.627 15.9918 145.005 0.00014802 0.267061 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991737 -2.97e-06 -85.6695 0.0929694 31198.9 300.078 0.983524 0.319147 0.767854 0.76785 9.99958 2.97989e-06 1.19194e-05 0.130464 0.972503 0.927031 -0.0132935 4.88956e-06 0.500136 -1.8498e-20 6.80385e-24 -1.84912e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998265 0.644309 0.0010401 0.00187941 0.000859158 0.455687 0.00187941 0.432793 0.000126627 1.02 0.887246 0.534802 0.285451 1.71587e-07 3.05282e-09 2395.91 3266.22 -0.0658958 0.482108 0.277709 0.262682 -0.591631 -0.169476 0.46596 -0.268799 -0.197158 1.144 1 3.83315e-249 287.381 2.18978e-246 1.98801 1.142 0.00029999 0.920223 0.62302 0.61086 0.393113 1.98836 125.947 82.2015 18.6203 60.0343 0.00409739 0 -40 10
0.243 7.04705e-09 2.53881e-06 0.0498595 0.0498429 0.0120468 3.2032e-06 0.001154 0.0623244 0.00065412 0.0629739 0.848782 101.893 0.247133 0.702968 4.10725 0.0528665 0.0387477 0.961252 0.0198939 0.0042257 0.019156 0.00406996 0.00510608 0.00584401 0.204243 0.23376 57.9543 -87.8935 125.63 15.9917 145.005 0.000147993 0.267061 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991737 -2.97e-06 -85.6695 0.0929694 31198.9 300.079 0.983524 0.319147 0.767714 0.76771 9.99958 2.97989e-06 1.19194e-05 0.130465 0.972537 0.927049 -0.0132935 4.88957e-06 0.500137 -1.84991e-20 6.80425e-24 -1.84923e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998262 0.644433 0.00104012 0.00187941 0.000859158 0.455687 0.00187941 0.432804 0.000126631 1.02 0.887246 0.534802 0.285451 1.71587e-07 3.05282e-09 2395.9 3265.62 -0.065852 0.482108 0.277708 0.262645 -0.591638 -0.169476 0.46609 -0.268799 -0.197289 1.145 1 2.32493e-249 287.422 1.32852e-246 1.98825 1.143 0.00029999 0.919954 0.623095 0.6101 0.393154 1.9886 125.96 82.2082 18.6207 60.0376 0.00409711 0 -40 10
0.244 7.07604e-09 2.53881e-06 0.0499706 0.0499541 0.0120468 3.21638e-06 0.001154 0.0624633 0.000654136 0.0631128 0.848809 101.893 0.247131 0.703 4.10728 0.0528691 0.0387479 0.961252 0.0198939 0.00422572 0.019156 0.00406998 0.00510612 0.00584404 0.204245 0.233762 57.9544 -87.8935 125.632 15.9917 145.005 0.000147966 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991737 -2.97e-06 -85.6695 0.0929694 31198.9 300.08 0.983524 0.319147 0.767575 0.767571 9.99958 2.97988e-06 1.19194e-05 0.130465 0.972572 0.927067 -0.0132935 4.88957e-06 0.500138 -1.85001e-20 6.80465e-24 -1.84933e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998259 0.644557 0.00104013 0.00187941 0.000859158 0.455687 0.00187941 0.432815 0.000126634 1.02 0.887246 0.534802 0.285451 1.71587e-07 3.05282e-09 2395.88 3265.03 -0.0658084 0.482108 0.277708 0.262608 -0.591645 -0.169476 0.46622 -0.268798 -0.19742 1.146 1 1.41014e-249 287.464 8.06004e-247 1.98849 1.144 0.00029999 0.919686 0.62317 0.609342 0.393195 1.98884 125.973 82.2148 18.6211 60.0408 0.00409682 0 -40 10
0.245 7.10502e-09 2.53881e-06 0.0500816 0.0500652 0.0120468 3.22956e-06 0.001154 0.062602 0.000654153 0.0632516 0.848836 101.893 0.247128 0.703033 4.1073 0.0528717 0.0387482 0.961252 0.0198938 0.00422575 0.0191559 0.00407001 0.00510615 0.00584407 0.204246 0.233763 57.9544 -87.8935 125.635 15.9917 145.005 0.00014794 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991737 -2.97e-06 -85.6695 0.0929694 31198.9 300.08 0.983524 0.319147 0.767437 0.767432 9.99958 2.97988e-06 1.19194e-05 0.130465 0.972606 0.927084 -0.0132935 4.88958e-06 0.500139 -1.85012e-20 6.80505e-24 -1.84944e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998256 0.644681 0.00104014 0.00187941 0.000859158 0.455687 0.00187941 0.432826 0.000126637 1.02 0.887246 0.534802 0.285452 1.71587e-07 3.05282e-09 2395.87 3264.44 -0.0657649 0.482108 0.277708 0.262572 -0.591652 -0.169476 0.466349 -0.268797 -0.19755 1.147 1 8.55292e-250 287.505 4.88995e-247 1.98873 1.145 0.00029999 0.919419 0.623245 0.608586 0.393236 1.98908 125.985 82.2215 18.6215 60.0441 0.00409654 0 -40 10
0.246 7.13401e-09 2.53881e-06 0.0501926 0.0501762 0.0120468 3.24273e-06 0.001154 0.0627407 0.000654169 0.0633903 0.848863 101.893 0.247126 0.703066 4.10733 0.0528743 0.0387484 0.961252 0.0198938 0.00422578 0.0191559 0.00407003 0.00510618 0.00584411 0.204247 0.233764 57.9545 -87.8935 125.637 15.9916 145.005 0.000147913 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991737 -2.97e-06 -85.6695 0.0929693 31198.9 300.081 0.983524 0.319147 0.767298 0.767294 9.99958 2.97988e-06 1.19194e-05 0.130465 0.97264 0.927102 -0.0132935 4.88958e-06 0.500141 -1.85022e-20 6.80544e-24 -1.84954e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998253 0.644805 0.00104016 0.00187941 0.000859158 0.455687 0.00187941 0.432837 0.00012664 1.02 0.887247 0.534802 0.285452 1.71587e-07 3.05283e-09 2395.85 3263.85 -0.0657216 0.482108 0.277707 0.262535 -0.591659 -0.169476 0.466478 -0.268796 -0.19768 1.148 1 5.18761e-250 287.547 2.96669e-247 1.98897 1.146 0.00029999 0.919153 0.62332 0.607833 0.393277 1.98932 125.998 82.2281 18.6218 60.0473 0.00409626 0 -40 10
0.247 7.163e-09 2.53881e-06 0.0503034 0.0502872 0.0120467 3.25591e-06 0.001154 0.0628793 0.000654185 0.0635288 0.848891 101.893 0.247123 0.703099 4.10736 0.0528769 0.0387486 0.961251 0.0198938 0.00422581 0.0191559 0.00407005 0.00510622 0.00584414 0.204249 0.233766 57.9545 -87.8935 125.64 15.9916 145.005 0.000147886 0.267061 192.946 0.310761 0.0673949 0.00409445 0.000561489 0.00138221 0.986996 0.991737 -2.97e-06 -85.6695 0.0929693 31198.9 300.082 0.983524 0.319147 0.76716 0.767156 9.99958 2.97988e-06 1.19194e-05 0.130466 0.972674 0.927119 -0.0132935 4.88959e-06 0.500142 -1.85033e-20 6.80584e-24 -1.84965e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998251 0.644929 0.00104017 0.00187941 0.000859158 0.455687 0.00187941 0.432847 0.000126644 1.02 0.887247 0.534802 0.285452 1.71587e-07 3.05283e-09 2395.83 3263.27 -0.0656785 0.482108 0.277707 0.262499 -0.591665 -0.169476 0.466606 -0.268795 -0.19781 1.149 1 3.14645e-250 287.588 1.79986e-247 1.98921 1.147 0.00029999 0.918887 0.623395 0.607081 0.393317 1.98956 126.011 82.2348 18.6222 60.0505 0.00409597 0 -40 10
0.248 7.19199e-09 2.53881e-06 0.0504142 0.050398 0.0120467 3.26909e-06 0.001154 0.0630177 0.000654202 0.0636673 0.848918 101.893 0.24712 0.703133 4.10738 0.0528796 0.0387489 0.961251 0.0198937 0.00422584 0.0191558 0.00407008 0.00510625 0.00584417 0.20425 0.233767 57.9546 -87.8935 125.642 15.9916 145.005 0.00014786 0.267061 192.946 0.310761 0.0673949 0.00409445 0.000561489 0.00138221 0.986996 0.991737 -2.97e-06 -85.6695 0.0929693 31198.9 300.083 0.983524 0.319147 0.767023 0.767018 9.99958 2.97988e-06 1.19194e-05 0.130466 0.972708 0.927137 -0.0132935 4.88959e-06 0.500143 -1.85044e-20 6.80624e-24 -1.84976e-20 0.00139493 0.997819 8.59158e-05 0.152528 2.85156 0.00139493 0.998248 0.645052 0.00104018 0.00187941 0.000859158 0.455687 0.00187941 0.432858 0.000126647 1.02 0.887247 0.534802 0.285452 1.71587e-07 3.05283e-09 2395.82 3262.68 -0.0656354 0.482108 0.277707 0.262462 -0.591672 -0.169476 0.466734 -0.268794 -0.197939 1.15 1 1.90842e-250 287.629 1.09196e-247 1.98945 1.148 0.00029999 0.918623 0.623469 0.606332 0.393358 1.9898 126.024 82.2413 18.6226 60.0537 0.00409569 0 -40 10
0.249 7.22098e-09 2.53881e-06 0.0505248 0.0505088 0.0120467 3.28226e-06 0.001154 0.063156 0.000654218 0.0638056 0.848946 101.893 0.247118 0.703166 4.10741 0.0528822 0.0387491 0.961251 0.0198937 0.00422586 0.0191558 0.0040701 0.00510629 0.00584421 0.204252 0.233768 57.9547 -87.8935 125.644 15.9915 145.005 0.000147833 0.267061 192.946 0.310761 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929693 31198.9 300.084 0.983524 0.319147 0.766886 0.766882 9.99958 2.97988e-06 1.19194e-05 0.130466 0.972742 0.927154 -0.0132935 4.8896e-06 0.500144 -1.85054e-20 6.80663e-24 -1.84986e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998245 0.645176 0.0010402 0.00187941 0.000859157 0.455687 0.00187941 0.432869 0.00012665 1.02 0.887247 0.534802 0.285453 1.71587e-07 3.05283e-09 2395.8 3262.1 -0.0655926 0.482108 0.277706 0.262426 -0.591679 -0.169477 0.466862 -0.268793 -0.198067 1.151 1 1.15751e-250 287.67 6.6248e-248 1.98969 1.149 0.00029999 0.918359 0.623544 0.605586 0.393399 1.99003 126.036 82.2479 18.623 60.0569 0.00409541 0 -40 10
0.25 7.24997e-09 2.53881e-06 0.0506354 0.0506194 0.0120467 3.29544e-06 0.001154 0.0632942 0.000654234 0.0639439 0.848974 101.893 0.247115 0.7032 4.10744 0.0528849 0.0387494 0.961251 0.0198937 0.00422589 0.0191558 0.00407012 0.00510632 0.00584424 0.204253 0.23377 57.9547 -87.8935 125.647 15.9915 145.005 0.000147807 0.267061 192.946 0.310761 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929693 31198.9 300.084 0.983524 0.319147 0.76675 0.766745 9.99958 2.97988e-06 1.19194e-05 0.130467 0.972776 0.927172 -0.0132935 4.8896e-06 0.500145 -1.85065e-20 6.80703e-24 -1.84997e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998242 0.6453 0.00104021 0.00187941 0.000859157 0.455687 0.00187941 0.43288 0.000126654 1.02 0.887247 0.534802 0.285453 1.71586e-07 3.05284e-09 2395.79 3261.52 -0.0655498 0.482108 0.277706 0.26239 -0.591685 -0.169477 0.466989 -0.268792 -0.198195 1.152 1 7.02067e-251 287.71 4.01919e-248 1.98993 1.15 0.00029999 0.918096 0.623618 0.604841 0.39344 1.99027 126.049 82.2545 18.6234 60.0601 0.00409513 0 -40 10
0.251 7.27895e-09 2.53881e-06 0.0507459 0.05073 0.0120467 3.30861e-06 0.001154 0.0634324 0.00065425 0.064082 0.849002 101.893 0.247112 0.703234 4.10746 0.0528876 0.0387496 0.96125 0.0198936 0.00422592 0.0191557 0.00407015 0.00510636 0.00584428 0.204254 0.233771 57.9548 -87.8935 125.649 15.9915 145.005 0.000147781 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929693 31198.9 300.085 0.983524 0.319147 0.766614 0.766609 9.99958 2.97988e-06 1.19194e-05 0.130467 0.972809 0.927189 -0.0132935 4.88961e-06 0.500146 -1.85075e-20 6.80743e-24 -1.85007e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998239 0.645423 0.00104022 0.00187941 0.000859157 0.455687 0.00187941 0.432891 0.000126657 1.02 0.887248 0.534802 0.285453 1.71586e-07 3.05284e-09 2395.77 3260.94 -0.0655073 0.482108 0.277706 0.262354 -0.591692 -0.169477 0.467116 -0.268791 -0.198323 1.153 1 4.25825e-251 287.751 2.4384e-248 1.99016 1.151 0.00029999 0.917835 0.623693 0.604098 0.39348 1.99051 126.062 82.261 18.6238 60.0633 0.00409485 0 -40 10
0.252 7.30794e-09 2.53881e-06 0.0508563 0.0508405 0.0120467 3.32179e-06 0.00115401 0.0635704 0.000654265 0.06422 0.849029 101.893 0.24711 0.703268 4.10749 0.0528903 0.0387499 0.96125 0.0198936 0.00422595 0.0191557 0.00407017 0.0051064 0.00584431 0.204256 0.233772 57.9548 -87.8935 125.651 15.9914 145.005 0.000147755 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929693 31198.9 300.086 0.983524 0.319147 0.766478 0.766474 9.99958 2.97988e-06 1.19194e-05 0.130467 0.972843 0.927206 -0.0132935 4.88962e-06 0.500148 -1.85086e-20 6.80782e-24 -1.85018e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998237 0.645547 0.00104024 0.00187941 0.000859157 0.455687 0.00187941 0.432902 0.00012666 1.02 0.887248 0.534802 0.285454 1.71586e-07 3.05284e-09 2395.75 3260.37 -0.0654648 0.482108 0.277705 0.262318 -0.591699 -0.169477 0.467242 -0.26879 -0.19845 1.154 1 2.58276e-251 287.792 1.47935e-248 1.9904 1.152 0.00029999 0.917574 0.623767 0.603358 0.393521 1.99075 126.075 82.2675 18.6242 60.0664 0.00409457 0 -40 10
0.253 7.33693e-09 2.53881e-06 0.0509666 0.0509509 0.0120467 3.33497e-06 0.00115401 0.0637082 0.000654281 0.0643579 0.849057 101.892 0.247107 0.703302 4.10752 0.052893 0.0387502 0.96125 0.0198936 0.00422598 0.0191557 0.00407019 0.00510643 0.00584435 0.204257 0.233774 57.9549 -87.8935 125.654 15.9914 145.005 0.000147729 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929693 31198.9 300.087 0.983524 0.319147 0.766343 0.766338 9.99958 2.97988e-06 1.19194e-05 0.130467 0.972876 0.927224 -0.0132935 4.88962e-06 0.500149 -1.85096e-20 6.80822e-24 -1.85028e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998234 0.64567 0.00104025 0.00187941 0.000859157 0.455687 0.00187941 0.432913 0.000126664 1.02 0.887248 0.534802 0.285454 1.71586e-07 3.05284e-09 2395.74 3259.79 -0.0654225 0.482108 0.277705 0.262283 -0.591705 -0.169477 0.467368 -0.26879 -0.198577 1.155 1 1.56652e-251 287.832 8.97504e-249 1.99064 1.153 0.00029999 0.917314 0.623841 0.60262 0.393562 1.99098 126.087 82.274 18.6246 60.0696 0.0040943 0 -40 10
0.254 7.36592e-09 2.53881e-06 0.0510768 0.0510612 0.0120466 3.34814e-06 0.00115401 0.063846 0.000654297 0.0644957 0.849085 101.892 0.247104 0.703336 4.10754 0.0528957 0.0387504 0.96125 0.0198935 0.00422601 0.0191556 0.00407022 0.00510647 0.00584438 0.204259 0.233775 57.955 -87.8935 125.656 15.9913 145.005 0.000147703 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.087 0.983525 0.319147 0.766208 0.766204 9.99958 2.97988e-06 1.19194e-05 0.130468 0.972909 0.927241 -0.0132935 4.88963e-06 0.50015 -1.85107e-20 6.80861e-24 -1.85039e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998231 0.645794 0.00104026 0.00187941 0.000859157 0.455687 0.00187941 0.432923 0.000126667 1.02 0.887248 0.534802 0.285454 1.71586e-07 3.05285e-09 2395.72 3259.22 -0.0653804 0.482108 0.277705 0.262247 -0.591712 -0.169477 0.467493 -0.268789 -0.198704 1.156 1 9.50144e-252 287.872 5.44504e-249 1.99088 1.154 0.00029999 0.917054 0.623915 0.601884 0.393602 1.99122 126.1 82.2805 18.6249 60.0727 0.00409402 0 -40 10
0.255 7.3949e-09 2.53881e-06 0.0511869 0.0511714 0.0120466 3.36132e-06 0.00115401 0.0639837 0.000654312 0.0646334 0.849114 101.892 0.247102 0.70337 4.10757 0.0528984 0.0387507 0.961249 0.0198935 0.00422604 0.0191556 0.00407024 0.0051065 0.00584442 0.20426 0.233777 57.955 -87.8935 125.658 15.9913 145.005 0.000147677 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.088 0.983525 0.319147 0.766074 0.76607 9.99958 2.97988e-06 1.19194e-05 0.130468 0.972943 0.927258 -0.0132935 4.88963e-06 0.500151 -1.85117e-20 6.809e-24 -1.85049e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998228 0.645917 0.00104028 0.00187941 0.000859157 0.455687 0.00187941 0.432934 0.00012667 1.02 0.887248 0.534802 0.285454 1.71586e-07 3.05285e-09 2395.7 3258.65 -0.0653384 0.482108 0.277705 0.262212 -0.591718 -0.169477 0.467618 -0.268788 -0.19883 1.157 1 5.76292e-252 287.912 3.30344e-249 1.99111 1.155 0.00029999 0.916796 0.623989 0.60115 0.393643 1.99146 126.113 82.2869 18.6253 60.0759 0.00409375 0 -40 10
0.256 7.42389e-09 2.53881e-06 0.051297 0.0512816 0.0120466 3.3745e-06 0.00115401 0.0641212 0.000654328 0.064771 0.849142 101.892 0.247099 0.703405 4.1076 0.0529011 0.0387509 0.961249 0.0198935 0.00422607 0.0191555 0.00407027 0.00510654 0.00584445 0.204262 0.233778 57.9551 -87.8935 125.661 15.9913 145.005 0.000147651 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.089 0.983525 0.319147 0.76594 0.765936 9.99958 2.97988e-06 1.19194e-05 0.130468 0.972976 0.927275 -0.0132935 4.88964e-06 0.500153 -1.85128e-20 6.8094e-24 -1.8506e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998226 0.646041 0.00104029 0.00187941 0.000859157 0.455687 0.00187941 0.432945 0.000126674 1.02 0.887249 0.534801 0.285455 1.71586e-07 3.05285e-09 2395.69 3258.08 -0.0652965 0.482108 0.277704 0.262176 -0.591725 -0.169477 0.467743 -0.268787 -0.198955 1.158 1 3.49538e-252 287.952 2.00415e-249 1.99135 1.156 0.00029999 0.916539 0.624063 0.600418 0.393683 1.99169 126.125 82.2933 18.6257 60.079 0.00409347 0 -40 10
0.257 7.45288e-09 2.53881e-06 0.051407 0.0513916 0.0120466 3.38767e-06 0.00115401 0.0642587 0.000654343 0.0649084 0.84917 101.892 0.247096 0.70344 4.10763 0.0529039 0.0387512 0.961249 0.0198934 0.0042261 0.0191555 0.00407029 0.00510658 0.00584449 0.204263 0.23378 57.9551 -87.8935 125.663 15.9912 145.005 0.000147625 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.09 0.983525 0.319147 0.765807 0.765802 9.99958 2.97987e-06 1.19194e-05 0.130469 0.973009 0.927292 -0.0132935 4.88965e-06 0.500154 -1.85138e-20 6.80979e-24 -1.8507e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998223 0.646164 0.00104031 0.00187941 0.000859157 0.455687 0.00187941 0.432956 0.000126677 1.02 0.887249 0.534801 0.285455 1.71586e-07 3.05286e-09 2395.67 3257.51 -0.0652548 0.482108 0.277704 0.262141 -0.591731 -0.169477 0.467867 -0.268786 -0.199081 1.159 1 2.12006e-252 287.992 1.21589e-249 1.99159 1.157 0.000299989 0.916282 0.624137 0.599688 0.393724 1.99193 126.138 82.2997 18.6261 60.0821 0.0040932 0 -40 10
0.258 7.48187e-09 2.53881e-06 0.0515168 0.0515016 0.0120466 3.40085e-06 0.00115401 0.064396 0.000654359 0.0650458 0.849199 101.892 0.247093 0.703475 4.10766 0.0529067 0.0387515 0.961249 0.0198934 0.00422613 0.0191555 0.00407032 0.00510661 0.00584453 0.204265 0.233781 57.9552 -87.8935 125.665 15.9912 145.005 0.0001476 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.091 0.983525 0.319147 0.765674 0.76567 9.99958 2.97987e-06 1.19194e-05 0.130469 0.973042 0.927309 -0.0132935 4.88965e-06 0.500155 -1.85149e-20 6.81018e-24 -1.85081e-20 0.00139493 0.997819 8.59157e-05 0.152527 2.85156 0.00139493 0.99822 0.646287 0.00104032 0.00187941 0.000859157 0.455687 0.00187941 0.432967 0.00012668 1.02 0.887249 0.534801 0.285455 1.71586e-07 3.05286e-09 2395.66 3256.95 -0.0652133 0.482108 0.277704 0.262106 -0.591738 -0.169477 0.467991 -0.268785 -0.199205 1.16 1 1.28588e-252 288.032 7.37666e-250 1.99182 1.158 0.000299989 0.916026 0.624211 0.598961 0.393764 1.99216 126.15 82.3061 18.6265 60.0852 0.00409293 0 -40 10
0.259 7.51085e-09 2.53881e-06 0.0516266 0.0516114 0.0120466 3.41402e-06 0.00115401 0.0645332 0.000654374 0.065183 0.849227 101.892 0.247091 0.70351 4.10768 0.0529094 0.0387517 0.961248 0.0198933 0.00422616 0.0191554 0.00407034 0.00510665 0.00584456 0.204266 0.233782 57.9553 -87.8935 125.668 15.9912 145.005 0.000147574 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.092 0.983525 0.319147 0.765542 0.765537 9.99958 2.97987e-06 1.19194e-05 0.130469 0.973074 0.927325 -0.0132935 4.88966e-06 0.500156 -1.85159e-20 6.81057e-24 -1.85091e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998218 0.646411 0.00104033 0.00187941 0.000859156 0.455687 0.00187941 0.432978 0.000126683 1.02 0.887249 0.534801 0.285456 1.71586e-07 3.05286e-09 2395.64 3256.38 -0.0651718 0.482108 0.277703 0.262071 -0.591744 -0.169477 0.468114 -0.268784 -0.19933 1.161 1 7.79926e-253 288.072 4.47531e-250 1.99206 1.159 0.000299989 0.915771 0.624285 0.598236 0.393804 1.9924 126.163 82.3125 18.6268 60.0883 0.00409266 0 -40 10
0.26 7.53984e-09 2.53881e-06 0.0517363 0.0517212 0.0120466 3.4272e-06 0.00115401 0.0646704 0.000654389 0.0653202 0.849256 101.892 0.247088 0.703545 4.10771 0.0529122 0.038752 0.961248 0.0198933 0.00422619 0.0191554 0.00407037 0.00510669 0.0058446 0.204268 0.233784 57.9553 -87.8935 125.67 15.9911 145.005 0.000147549 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.092 0.983525 0.319147 0.76541 0.765405 9.99958 2.97987e-06 1.19194e-05 0.13047 0.973107 0.927342 -0.0132935 4.88967e-06 0.500158 -1.85169e-20 6.81097e-24 -1.85101e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998215 0.646534 0.00104035 0.00187941 0.000859156 0.455687 0.00187941 0.432988 0.000126687 1.02 0.88725 0.534801 0.285456 1.71586e-07 3.05287e-09 2395.62 3255.82 -0.0651305 0.482108 0.277703 0.262036 -0.591751 -0.169477 0.468237 -0.268783 -0.199454 1.162 1 4.73049e-253 288.111 2.71511e-250 1.99229 1.16 0.000299989 0.915517 0.624359 0.597512 0.393845 1.99263 126.176 82.3188 18.6272 60.0914 0.00409239 0 -40 10
0.261 7.56883e-09 2.53881e-06 0.0518459 0.0518309 0.0120466 3.44038e-06 0.00115401 0.0648074 0.000654404 0.0654572 0.849285 101.892 0.247085 0.70358 4.10774 0.052915 0.0387523 0.961248 0.0198933 0.00422622 0.0191554 0.00407039 0.00510673 0.00584464 0.204269 0.233785 57.9554 -87.8935 125.672 15.9911 145.005 0.000147524 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991737 -2.96999e-06 -85.6695 0.0929692 31198.9 300.093 0.983525 0.319147 0.765278 0.765274 9.99958 2.97987e-06 1.19194e-05 0.13047 0.97314 0.927359 -0.0132935 4.88968e-06 0.500159 -1.8518e-20 6.81136e-24 -1.85112e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998213 0.646657 0.00104036 0.00187941 0.000859156 0.455687 0.00187941 0.432999 0.00012669 1.02 0.88725 0.534801 0.285457 1.71586e-07 3.05287e-09 2395.61 3255.26 -0.0650894 0.482108 0.277703 0.262001 -0.591757 -0.169477 0.468359 -0.268782 -0.199577 1.163 1 2.86919e-253 288.15 1.64722e-250 1.99253 1.161 0.000299989 0.915264 0.624432 0.596791 0.393885 1.99287 126.188 82.3252 18.6276 60.0945 0.00409212 0 -40 10
0.262 7.59781e-09 2.53881e-06 0.0519554 0.0519405 0.0120465 3.45355e-06 0.00115401 0.0649443 0.000654419 0.0655941 0.849313 101.892 0.247082 0.703616 4.10777 0.0529178 0.0387526 0.961247 0.0198932 0.00422625 0.0191553 0.00407042 0.00510677 0.00584467 0.204271 0.233787 57.9554 -87.8935 125.675 15.9911 145.005 0.000147498 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.96999e-06 -85.6695 0.0929692 31199 300.094 0.983525 0.319147 0.765147 0.765142 9.99958 2.97987e-06 1.19194e-05 0.13047 0.973172 0.927376 -0.0132935 4.88968e-06 0.50016 -1.8519e-20 6.81175e-24 -1.85122e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.99821 0.64678 0.00104038 0.00187941 0.000859156 0.455687 0.00187941 0.43301 0.000126693 1.02 0.88725 0.534801 0.285457 1.71586e-07 3.05288e-09 2395.59 3254.71 -0.0650484 0.482108 0.277702 0.261967 -0.591764 -0.169477 0.468481 -0.268781 -0.1997 1.164 1 1.74025e-253 288.19 9.9934e-251 1.99276 1.162 0.000299989 0.915012 0.624506 0.596072 0.393925 1.9931 126.201 82.3315 18.628 60.0975 0.00409185 0 -40 10
0.263 7.6268e-09 2.53881e-06 0.0520648 0.05205 0.0120465 3.46673e-06 0.00115401 0.0650811 0.000654434 0.0657309 0.849342 101.892 0.247079 0.703652 4.1078 0.0529207 0.0387528 0.961247 0.0198932 0.00422628 0.0191553 0.00407044 0.0051068 0.00584471 0.204272 0.233788 57.9555 -87.8935 125.677 15.991 145.005 0.000147473 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.96999e-06 -85.6695 0.0929692 31199 300.095 0.983525 0.319147 0.765016 0.765012 9.99958 2.97987e-06 1.19194e-05 0.130471 0.973205 0.927392 -0.0132935 4.88969e-06 0.500161 -1.85201e-20 6.81214e-24 -1.85132e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998208 0.646903 0.00104039 0.00187941 0.000859156 0.455687 0.00187941 0.433021 0.000126697 1.02 0.887251 0.534801 0.285457 1.71586e-07 3.05288e-09 2395.58 3254.15 -0.0650075 0.482108 0.277702 0.261932 -0.59177 -0.169478 0.468603 -0.26878 -0.199823 1.165 1 1.05551e-253 288.229 6.06284e-251 1.993 1.163 0.000299989 0.914761 0.624579 0.595355 0.393965 1.99334 126.213 82.3377 18.6283 60.1006 0.00409158 0 -40 10
0.264 7.65579e-09 2.53881e-06 0.0521742 0.0521594 0.0120465 3.4799e-06 0.00115401 0.0652177 0.000654449 0.0658676 0.849371 101.892 0.247076 0.703687 4.10783 0.0529235 0.0387531 0.961247 0.0198932 0.00422632 0.0191553 0.00407047 0.00510684 0.00584475 0.204274 0.23379 57.9556 -87.8935 125.679 15.991 145.005 0.000147448 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.96999e-06 -85.6695 0.0929692 31199 300.096 0.983525 0.319147 0.764886 0.764882 9.99958 2.97987e-06 1.19194e-05 0.130471 0.973237 0.927409 -0.0132935 4.8897e-06 0.500163 -1.85211e-20 6.81253e-24 -1.85143e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998205 0.647026 0.00104041 0.00187941 0.000859156 0.455687 0.00187941 0.433032 0.0001267 1.02 0.887251 0.534801 0.285458 1.71586e-07 3.05289e-09 2395.56 3253.6 -0.0649668 0.482108 0.277702 0.261898 -0.591776 -0.169478 0.468724 -0.268779 -0.199945 1.166 1 6.40202e-254 288.268 3.67823e-251 1.99323 1.164 0.000299989 0.91451 0.624652 0.59464 0.394005 1.99357 126.226 82.344 18.6287 60.1036 0.00409131 0 -40 10
0.265 7.68477e-09 2.53881e-06 0.0522834 0.0522687 0.0120465 3.49308e-06 0.00115401 0.0653543 0.000654463 0.0660042 0.8494 101.892 0.247074 0.703723 4.10786 0.0529264 0.0387534 0.961247 0.0198931 0.00422635 0.0191552 0.00407049 0.00510688 0.00584479 0.204275 0.233791 57.9556 -87.8935 125.681 15.991 145.005 0.000147423 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.96999e-06 -85.6695 0.0929692 31199 300.097 0.983525 0.319147 0.764756 0.764752 9.99958 2.97987e-06 1.19194e-05 0.130471 0.973269 0.927425 -0.0132935 4.88971e-06 0.500164 -1.85221e-20 6.81292e-24 -1.85153e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998202 0.647149 0.00104042 0.00187941 0.000859156 0.455687 0.00187941 0.433042 0.000126704 1.02 0.887251 0.534801 0.285458 1.71586e-07 3.05289e-09 2395.54 3253.04 -0.0649262 0.482108 0.277701 0.261863 -0.591783 -0.169478 0.468845 -0.268778 -0.200067 1.167 1 3.88302e-254 288.307 2.23152e-251 1.99347 1.165 0.000299989 0.91426 0.624726 0.593928 0.394045 1.99381 126.238 82.3502 18.6291 60.1067 0.00409105 0 -40 10
0.266 7.71376e-09 2.53881e-06 0.0523926 0.052378 0.0120465 3.50625e-06 0.00115401 0.0654908 0.000654478 0.0661406 0.84943 101.892 0.247071 0.70376 4.10789 0.0529292 0.0387537 0.961246 0.0198931 0.00422638 0.0191552 0.00407052 0.00510692 0.00584483 0.204277 0.233793 57.9557 -87.8935 125.684 15.9909 145.005 0.000147398 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.96999e-06 -85.6695 0.0929692 31199 300.097 0.983525 0.319147 0.764627 0.764622 9.99958 2.97987e-06 1.19194e-05 0.130471 0.973301 0.927442 -0.0132935 4.88971e-06 0.500165 -1.85231e-20 6.81331e-24 -1.85163e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.9982 0.647272 0.00104043 0.00187941 0.000859156 0.455687 0.00187941 0.433053 0.000126707 1.02 0.887251 0.534801 0.285458 1.71586e-07 3.05289e-09 2395.53 3252.49 -0.0648858 0.482108 0.277701 0.261829 -0.591789 -0.169478 0.468965 -0.268777 -0.200188 1.168 1 2.35517e-254 288.345 1.35383e-251 1.9937 1.166 0.000299989 0.914011 0.624799 0.593217 0.394085 1.99404 126.251 82.3565 18.6294 60.1097 0.00409078 0 -40 10
0.267 7.74275e-09 2.53881e-06 0.0525017 0.0524871 0.0120465 3.51943e-06 0.00115401 0.0656271 0.000654493 0.066277 0.849459 101.892 0.247068 0.703796 4.10792 0.0529321 0.038754 0.961246 0.019893 0.00422641 0.0191551 0.00407055 0.00510696 0.00584486 0.204278 0.233795 57.9557 -87.8935 125.686 15.9909 145.005 0.000147373 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.96999e-06 -85.6695 0.0929692 31199 300.098 0.983525 0.319147 0.764498 0.764493 9.99958 2.97987e-06 1.19194e-05 0.130472 0.973333 0.927458 -0.0132935 4.88972e-06 0.500167 -1.85242e-20 6.8137e-24 -1.85174e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998197 0.647395 0.00104045 0.00187941 0.000859156 0.455687 0.00187941 0.433064 0.00012671 1.02 0.887252 0.534801 0.285459 1.71586e-07 3.0529e-09 2395.51 3251.94 -0.0648454 0.482108 0.277701 0.261795 -0.591795 -0.169478 0.469085 -0.268776 -0.200309 1.169 1 1.42848e-254 288.384 8.21344e-252 1.99393 1.167 0.000299989 0.913763 0.624872 0.592508 0.394125 1.99427 126.263 82.3627 18.6298 60.1127 0.00409052 0 -40 10
0.268 7.77173e-09 2.53881e-06 0.0526107 0.0525962 0.0120465 3.53261e-06 0.00115401 0.0657633 0.000654507 0.0664133 0.849488 101.892 0.247065 0.703832 4.10795 0.052935 0.0387542 0.961246 0.019893 0.00422644 0.0191551 0.00407057 0.005107 0.0058449 0.20428 0.233796 57.9558 -87.8936 125.688 15.9908 145.006 0.000147348 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.099 0.983525 0.319147 0.764369 0.764365 9.99958 2.97987e-06 1.19194e-05 0.130472 0.973365 0.927474 -0.0132935 4.88973e-06 0.500168 -1.85252e-20 6.81409e-24 -1.85184e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998195 0.647518 0.00104046 0.00187941 0.000859156 0.455687 0.00187941 0.433075 0.000126714 1.02 0.887252 0.534801 0.285459 1.71586e-07 3.0529e-09 2395.5 3251.4 -0.0648053 0.482108 0.2777 0.261761 -0.591802 -0.169478 0.469205 -0.268774 -0.20043 1.17 1 8.66419e-255 288.422 4.98295e-252 1.99417 1.168 0.000299989 0.913516 0.624945 0.591802 0.394165 1.9945 126.276 82.3689 18.6302 60.1157 0.00409025 0 -40 10
0.269 7.80072e-09 2.53881e-06 0.0527196 0.0527052 0.0120464 3.54578e-06 0.00115401 0.0658995 0.000654522 0.0665494 0.849518 101.892 0.247062 0.703869 4.10798 0.0529379 0.0387545 0.961245 0.019893 0.00422648 0.0191551 0.0040706 0.00510704 0.00584494 0.204282 0.233798 57.9558 -87.8936 125.69 15.9908 145.006 0.000147324 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.1 0.983525 0.319147 0.764241 0.764237 9.99958 2.97987e-06 1.19194e-05 0.130472 0.973397 0.927491 -0.0132935 4.88974e-06 0.500169 -1.85262e-20 6.81448e-24 -1.85194e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998193 0.647641 0.00104048 0.00187941 0.000859156 0.455687 0.00187941 0.433086 0.000126717 1.02 0.887252 0.5348 0.28546 1.71586e-07 3.05291e-09 2395.48 3250.85 -0.0647652 0.482108 0.2777 0.261727 -0.591808 -0.169478 0.469324 -0.268773 -0.20055 1.171 1 5.2551e-255 288.461 3.02307e-252 1.9944 1.169 0.000299989 0.91327 0.625018 0.591097 0.394205 1.99474 126.288 82.375 18.6305 60.1187 0.00408999 0 -40 10
0.27 7.8297e-09 2.53881e-06 0.0528284 0.0528141 0.0120464 3.55896e-06 0.00115401 0.0660355 0.000654536 0.0666854 0.849547 101.892 0.247059 0.703906 4.10801 0.0529408 0.0387548 0.961245 0.0198929 0.00422651 0.019155 0.00407063 0.00510708 0.00584498 0.204283 0.233799 57.9559 -87.8936 125.693 15.9908 145.006 0.000147299 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.101 0.983525 0.319147 0.764114 0.764109 9.99958 2.97987e-06 1.19194e-05 0.130473 0.973429 0.927507 -0.0132935 4.88975e-06 0.500171 -1.85272e-20 6.81486e-24 -1.85204e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.99819 0.647764 0.00104049 0.00187941 0.000859156 0.455687 0.00187941 0.433096 0.00012672 1.02 0.887253 0.5348 0.28546 1.71586e-07 3.05291e-09 2395.46 3250.31 -0.0647253 0.482108 0.2777 0.261693 -0.591814 -0.169478 0.469443 -0.268772 -0.20067 1.172 1 3.18738e-255 288.499 1.83404e-252 1.99463 1.17 0.000299989 0.913024 0.625091 0.590395 0.394245 1.99497 126.301 82.3812 18.6309 60.1217 0.00408973 0 -40 10
0.271 7.85869e-09 2.53881e-06 0.0529371 0.0529229 0.0120464 3.57213e-06 0.00115401 0.0661714 0.00065455 0.0668214 0.849577 101.892 0.247056 0.703943 4.10804 0.0529437 0.0387551 0.961245 0.0198929 0.00422654 0.019155 0.00407065 0.00510712 0.00584502 0.204285 0.233801 57.956 -87.8936 125.695 15.9907 145.006 0.000147274 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.102 0.983525 0.319147 0.763986 0.763982 9.99958 2.97987e-06 1.19194e-05 0.130473 0.97346 0.927523 -0.0132935 4.88975e-06 0.500172 -1.85283e-20 6.81525e-24 -1.85215e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998188 0.647886 0.00104051 0.00187941 0.000859156 0.455687 0.00187941 0.433107 0.000126724 1.02 0.887253 0.5348 0.285461 1.71586e-07 3.05292e-09 2395.45 3249.77 -0.0646856 0.482108 0.2777 0.26166 -0.59182 -0.169478 0.469561 -0.268771 -0.200789 1.173 1 1.93324e-255 288.537 1.11268e-252 1.99487 1.171 0.000299989 0.91278 0.625163 0.589694 0.394284 1.9952 126.313 82.3873 18.6313 60.1247 0.00408947 0 -40 10
0.272 7.88768e-09 2.53881e-06 0.0530458 0.0530316 0.0120464 3.58531e-06 0.00115401 0.0663072 0.000654564 0.0669572 0.849607 101.892 0.247053 0.70398 4.10807 0.0529466 0.0387554 0.961245 0.0198928 0.00422658 0.0191549 0.00407068 0.00510716 0.00584506 0.204286 0.233802 57.956 -87.8936 125.697 15.9907 145.006 0.00014725 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.103 0.983525 0.319147 0.76386 0.763855 9.99958 2.97987e-06 1.19194e-05 0.130473 0.973492 0.927539 -0.0132935 4.88976e-06 0.500173 -1.85293e-20 6.81564e-24 -1.85225e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998185 0.648009 0.00104052 0.00187941 0.000859156 0.455687 0.00187941 0.433118 0.000126727 1.02 0.887253 0.5348 0.285461 1.71586e-07 3.05292e-09 2395.43 3249.23 -0.064646 0.482108 0.277699 0.261626 -0.591827 -0.169478 0.469679 -0.26877 -0.200908 1.174 1 1.17257e-255 288.575 6.75041e-253 1.9951 1.172 0.000299989 0.912536 0.625236 0.588996 0.394324 1.99543 126.325 82.3934 18.6316 60.1276 0.00408921 0 -40 10
0.273 7.91666e-09 2.53881e-06 0.0531543 0.0531402 0.0120464 3.59848e-06 0.00115401 0.0664429 0.000654578 0.0670929 0.849636 101.892 0.24705 0.704017 4.1081 0.0529496 0.0387557 0.961244 0.0198928 0.00422661 0.0191549 0.00407071 0.0051072 0.0058451 0.204288 0.233804 57.9561 -87.8936 125.699 15.9907 145.006 0.000147226 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.104 0.983525 0.319147 0.763733 0.763729 9.99958 2.97987e-06 1.19194e-05 0.130474 0.973523 0.927555 -0.0132935 4.88977e-06 0.500175 -1.85303e-20 6.81603e-24 -1.85235e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998183 0.648132 0.00104054 0.00187941 0.000859156 0.455687 0.00187941 0.433129 0.00012673 1.02 0.887254 0.5348 0.285461 1.71586e-07 3.05293e-09 2395.41 3248.69 -0.0646065 0.482108 0.277699 0.261593 -0.591833 -0.169478 0.469796 -0.268769 -0.201027 1.175 1 7.112e-256 288.613 4.09534e-253 1.99533 1.173 0.000299989 0.912293 0.625309 0.588299 0.394364 1.99567 126.338 82.3995 18.632 60.1306 0.00408895 0 -40 10
0.274 7.94565e-09 2.53881e-06 0.0532628 0.0532488 0.0120464 3.61166e-06 0.00115401 0.0665785 0.000654593 0.0672285 0.849666 101.892 0.247047 0.704054 4.10814 0.0529526 0.038756 0.961244 0.0198928 0.00422664 0.0191549 0.00407074 0.00510724 0.00584514 0.20429 0.233806 57.9561 -87.8936 125.702 15.9906 145.006 0.000147201 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.105 0.983525 0.319147 0.763607 0.763603 9.99958 2.97987e-06 1.19194e-05 0.130474 0.973554 0.927571 -0.0132935 4.88978e-06 0.500176 -1.85313e-20 6.81641e-24 -1.85245e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.99818 0.648254 0.00104055 0.00187941 0.000859156 0.455687 0.00187941 0.433139 0.000126734 1.02 0.887254 0.5348 0.285462 1.71586e-07 3.05293e-09 2395.4 3248.16 -0.0645671 0.482108 0.277699 0.261559 -0.591839 -0.169478 0.469913 -0.268768 -0.201145 1.176 1 4.31365e-256 288.65 2.48456e-253 1.99556 1.174 0.000299989 0.91205 0.625381 0.587605 0.394403 1.9959 126.35 82.4055 18.6323 60.1335 0.00408869 0 -40 10
0.275 7.97463e-09 2.53881e-06 0.0533712 0.0533572 0.0120464 3.62483e-06 0.00115401 0.066714 0.000654607 0.067364 0.849696 101.892 0.247044 0.704092 4.10817 0.0529555 0.0387563 0.961244 0.0198927 0.00422668 0.0191548 0.00407076 0.00510729 0.00584518 0.204291 0.233807 57.9562 -87.8936 125.704 15.9906 145.006 0.000147177 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97e-06 -85.6695 0.0929692 31199 300.106 0.983525 0.319147 0.763482 0.763477 9.99958 2.97987e-06 1.19194e-05 0.130475 0.973585 0.927587 -0.0132935 4.88979e-06 0.500177 -1.85323e-20 6.8168e-24 -1.85255e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998178 0.648377 0.00104057 0.00187941 0.000859156 0.455687 0.00187941 0.43315 0.000126737 1.02 0.887254 0.5348 0.285462 1.71586e-07 3.05294e-09 2395.38 3247.62 -0.0645279 0.482108 0.277698 0.261526 -0.591845 -0.169478 0.47003 -0.268767 -0.201263 1.177 1 2.61636e-256 288.688 1.50734e-253 1.99579 1.175 0.000299988 0.911809 0.625454 0.586913 0.394443 1.99613 126.363 82.4116 18.6327 60.1365 0.00408844 0 -40 10
0.276 8.00362e-09 2.53881e-06 0.0534795 0.0534656 0.0120464 3.63801e-06 0.00115401 0.0668493 0.00065462 0.0674994 0.849726 101.892 0.247041 0.70413 4.1082 0.0529585 0.0387566 0.961243 0.0198927 0.00422671 0.0191548 0.00407079 0.00510733 0.00584522 0.204293 0.233809 57.9563 -87.8936 125.706 15.9906 145.006 0.000147153 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97001e-06 -85.6695 0.0929692 31199 300.106 0.983525 0.319147 0.763357 0.763352 9.99958 2.97987e-06 1.19194e-05 0.130475 0.973617 0.927603 -0.0132935 4.8898e-06 0.500179 -1.85333e-20 6.81718e-24 -1.85265e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998176 0.648499 0.00104058 0.00187941 0.000859156 0.455687 0.00187941 0.433161 0.00012674 1.02 0.887254 0.5348 0.285463 1.71586e-07 3.05295e-09 2395.37 3247.09 -0.0644888 0.482108 0.277698 0.261493 -0.591851 -0.169478 0.470146 -0.268766 -0.201381 1.178 1 1.5869e-256 288.726 9.1447e-254 1.99603 1.176 0.000299988 0.911568 0.625526 0.586222 0.394482 1.99636 126.375 82.4176 18.633 60.1394 0.00408818 0 -40 10
0.277 8.0326e-09 2.53881e-06 0.0535877 0.0535739 0.0120463 3.65118e-06 0.00115401 0.0669846 0.000654634 0.0676346 0.849757 101.892 0.247038 0.704167 4.10823 0.0529615 0.0387569 0.961243 0.0198926 0.00422674 0.0191547 0.00407082 0.00510737 0.00584526 0.204295 0.233811 57.9563 -87.8936 125.708 15.9905 145.006 0.000147129 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97001e-06 -85.6695 0.0929692 31199 300.107 0.983525 0.319147 0.763232 0.763227 9.99958 2.97987e-06 1.19194e-05 0.130475 0.973648 0.927619 -0.0132935 4.88981e-06 0.50018 -1.85344e-20 6.81757e-24 -1.85275e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998173 0.648622 0.0010406 0.00187941 0.000859156 0.455687 0.00187941 0.433171 0.000126744 1.02 0.887255 0.5348 0.285463 1.71586e-07 3.05295e-09 2395.35 3246.56 -0.0644499 0.482108 0.277698 0.26146 -0.591857 -0.169479 0.470262 -0.268765 -0.201498 1.179 1 9.62505e-257 288.763 5.5479e-254 1.99626 1.177 0.000299988 0.911329 0.625598 0.585534 0.394522 1.99659 126.387 82.4236 18.6334 60.1423 0.00408792 0 -40 10
0.278 8.06159e-09 2.53881e-06 0.0536958 0.0536821 0.0120463 3.66436e-06 0.00115401 0.0671198 0.000654648 0.0677698 0.849787 101.892 0.247035 0.704205 4.10826 0.0529645 0.0387572 0.961243 0.0198926 0.00422678 0.0191547 0.00407085 0.00510741 0.0058453 0.204296 0.233812 57.9564 -87.8936 125.71 15.9905 145.006 0.000147105 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97001e-06 -85.6695 0.0929692 31199 300.108 0.983525 0.319147 0.763108 0.763103 9.99958 2.97987e-06 1.19194e-05 0.130476 0.973678 0.927635 -0.0132935 4.88982e-06 0.500182 -1.85354e-20 6.81795e-24 -1.85286e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998171 0.648744 0.00104061 0.00187941 0.000859156 0.455687 0.00187941 0.433182 0.000126747 1.02 0.887255 0.5348 0.285464 1.71586e-07 3.05296e-09 2395.33 3246.03 -0.0644111 0.482108 0.277697 0.261427 -0.591863 -0.169479 0.470377 -0.268764 -0.201614 1.18 1 5.83789e-257 288.8 3.3658e-254 1.99649 1.178 0.000299988 0.91109 0.625671 0.584848 0.394561 1.99682 126.4 82.4296 18.6338 60.1452 0.00408767 0 -40 10
0.279 8.09057e-09 2.53881e-06 0.0538038 0.0537902 0.0120463 3.67753e-06 0.00115401 0.0672548 0.000654662 0.0679049 0.849817 101.892 0.247032 0.704244 4.1083 0.0529675 0.0387575 0.961242 0.0198925 0.00422681 0.0191547 0.00407088 0.00510745 0.00584535 0.204298 0.233814 57.9564 -87.8936 125.712 15.9904 145.006 0.000147081 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97001e-06 -85.6695 0.0929692 31199 300.109 0.983525 0.319147 0.762984 0.762979 9.99958 2.97987e-06 1.19194e-05 0.130476 0.973709 0.92765 -0.0132935 4.88983e-06 0.500183 -1.85364e-20 6.81834e-24 -1.85296e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998169 0.648867 0.00104062 0.00187941 0.000859156 0.455687 0.00187941 0.433193 0.000126751 1.02 0.887256 0.5348 0.285464 1.71586e-07 3.05296e-09 2395.32 3245.5 -0.0643724 0.482108 0.277697 0.261394 -0.591869 -0.169479 0.470492 -0.268763 -0.20173 1.181 1 3.54086e-257 288.837 2.04196e-254 1.99672 1.179 0.000299988 0.910851 0.625743 0.584163 0.394601 1.99705 126.412 82.4356 18.6341 60.1481 0.00408742 0 -40 10
0.28 8.11956e-09 2.53881e-06 0.0539118 0.0538982 0.0120463 3.69071e-06 0.00115401 0.0673897 0.000654675 0.0680398 0.849848 101.892 0.247029 0.704282 4.10833 0.0529706 0.0387578 0.961242 0.0198925 0.00422685 0.0191546 0.00407091 0.0051075 0.00584539 0.2043 0.233816 57.9565 -87.8936 125.715 15.9904 145.006 0.000147057 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97001e-06 -85.6695 0.0929692 31199 300.11 0.983525 0.319147 0.76286 0.762856 9.99958 2.97987e-06 1.19194e-05 0.130476 0.97374 0.927666 -0.0132935 4.88984e-06 0.500185 -1.85374e-20 6.81872e-24 -1.85306e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998167 0.648989 0.00104064 0.00187941 0.000859156 0.455687 0.00187941 0.433204 0.000126754 1.02 0.887256 0.534799 0.285465 1.71586e-07 3.05297e-09 2395.3 3244.98 -0.0643338 0.482108 0.277697 0.261362 -0.591876 -0.169479 0.470607 -0.268761 -0.201846 1.182 1 2.14764e-257 288.874 1.23881e-254 1.99695 1.18 0.000299988 0.910614 0.625815 0.583481 0.39464 1.99728 126.424 82.4415 18.6345 60.151 0.00408716 0 -40 10
0.281 8.14854e-09 2.53881e-06 0.0540196 0.0540061 0.0120463 3.70388e-06 0.00115401 0.0675246 0.000654689 0.0681746 0.849878 101.892 0.247026 0.70432 4.10836 0.0529736 0.0387581 0.961242 0.0198925 0.00422688 0.0191546 0.00407093 0.00510754 0.00584543 0.204302 0.233817 57.9566 -87.8936 125.717 15.9904 145.006 0.000147034 0.267061 192.946 0.310762 0.067395 0.00409444 0.000561488 0.00138221 0.986996 0.991738 -2.97002e-06 -85.6695 0.0929692 31198.9 300.111 0.983525 0.319147 0.762737 0.762733 9.99958 2.97987e-06 1.19194e-05 0.130477 0.973771 0.927682 -0.0132935 4.88985e-06 0.500186 -1.85384e-20 6.81911e-24 -1.85316e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998164 0.649111 0.00104065 0.00187941 0.000859156 0.455687 0.00187941 0.433214 0.000126757 1.02 0.887256 0.534799 0.285465 1.71586e-07 3.05298e-09 2395.29 3244.45 -0.0642954 0.482108 0.277696 0.261329 -0.591882 -0.169479 0.470721 -0.26876 -0.201962 1.183 1 1.30261e-257 288.911 7.51559e-255 1.99718 1.181 0.000299988 0.910378 0.625887 0.5828 0.394679 1.99751 126.437 82.4474 18.6348 60.1539 0.00408691 0 -40 10
0.282 8.17753e-09 2.53881e-06 0.0541274 0.054114 0.0120463 3.71706e-06 0.00115401 0.0676593 0.000654702 0.0683094 0.849909 101.892 0.247023 0.704359 4.1084 0.0529767 0.0387584 0.961242 0.0198924 0.00422692 0.0191545 0.00407096 0.00510758 0.00584547 0.204303 0.233819 57.9566 -87.8936 125.719 15.9903 145.006 0.00014701 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97002e-06 -85.6695 0.0929692 31198.9 300.112 0.983525 0.319147 0.762615 0.76261 9.99958 2.97987e-06 1.19194e-05 0.130477 0.973801 0.927697 -0.0132935 4.88986e-06 0.500187 -1.85394e-20 6.81949e-24 -1.85326e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.998162 0.649234 0.00104067 0.00187941 0.000859156 0.455687 0.00187941 0.433225 0.000126761 1.02 0.887257 0.534799 0.285466 1.71586e-07 3.05298e-09 2395.27 3243.93 -0.0642571 0.482108 0.277696 0.261297 -0.591888 -0.169479 0.470835 -0.268759 -0.202077 1.184 1 7.90072e-258 288.948 4.55954e-255 1.99741 1.182 0.000299988 0.910142 0.625959 0.582122 0.394719 1.99774 126.449 82.4533 18.6352 60.1568 0.00408666 0 -40 10
0.283 8.20651e-09 2.53881e-06 0.0542351 0.0542217 0.0120463 3.73023e-06 0.00115401 0.0677939 0.000654716 0.068444 0.849939 101.892 0.24702 0.704398 4.10843 0.0529797 0.0387588 0.961241 0.0198924 0.00422695 0.0191545 0.00407099 0.00510763 0.00584551 0.204305 0.233821 57.9567 -87.8936 125.721 15.9903 145.006 0.000146986 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97002e-06 -85.6695 0.0929692 31198.9 300.113 0.983525 0.319147 0.762492 0.762488 9.99958 2.97987e-06 1.19194e-05 0.130477 0.973832 0.927713 -0.0132935 4.88987e-06 0.500189 -1.85404e-20 6.81987e-24 -1.85336e-20 0.00139493 0.997819 8.59156e-05 0.152527 2.85156 0.00139493 0.99816 0.649356 0.00104069 0.00187941 0.000859156 0.455687 0.00187941 0.433236 0.000126764 1.02 0.887257 0.534799 0.285466 1.71586e-07 3.05299e-09 2395.25 3243.41 -0.064219 0.482108 0.277696 0.261264 -0.591894 -0.169479 0.470949 -0.268758 -0.202191 1.185 1 4.79203e-258 288.985 2.76617e-255 1.99764 1.183 0.000299988 0.909907 0.62603 0.581446 0.394758 1.99797 126.461 82.4592 18.6355 60.1596 0.00408641 0 -40 10
0.284 8.2355e-09 2.53881e-06 0.0543427 0.0543294 0.0120463 3.74341e-06 0.00115401 0.0679284 0.000654729 0.0685785 0.84997 101.892 0.247017 0.704437 4.10846 0.0529828 0.0387591 0.961241 0.0198923 0.00422699 0.0191544 0.00407102 0.00510767 0.00584556 0.204307 0.233822 57.9568 -87.8936 125.723 15.9903 145.006 0.000146963 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97002e-06 -85.6695 0.0929692 31198.9 300.114 0.983525 0.319147 0.76237 0.762366 9.99958 2.97987e-06 1.19194e-05 0.130478 0.973862 0.927728 -0.0132935 4.88988e-06 0.50019 -1.85414e-20 6.82026e-24 -1.85346e-20 0.00139493 0.997819 8.59157e-05 0.152527 2.85156 0.00139493 0.998158 0.649478 0.0010407 0.00187941 0.000859157 0.455687 0.00187941 0.433246 0.000126768 1.02 0.887257 0.534799 0.285467 1.71586e-07 3.05299e-09 2395.24 3242.89 -0.064181 0.482108 0.277696 0.261232 -0.5919 -0.169479 0.471062 -0.268757 -0.202306 1.186 1 2.90651e-258 289.021 1.67817e-255 1.99787 1.184 0.000299988 0.909673 0.626102 0.580771 0.394797 1.9982 126.473 82.4651 18.6358 60.1625 0.00408616 0 -40 10
0.285 8.26448e-09 2.53881e-06 0.0544502 0.054437 0.0120462 3.75658e-06 0.00115401 0.0680628 0.000654742 0.0687129 0.850001 101.892 0.247014 0.704476 4.1085 0.0529859 0.0387594 0.961241 0.0198923 0.00422703 0.0191544 0.00407105 0.00510772 0.0058456 0.204309 0.233824 57.9568 -87.8936 125.725 15.9902 145.006 0.00014694 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97002e-06 -85.6695 0.0929692 31198.9 300.115 0.983525 0.319147 0.762249 0.762244 9.99958 2.97987e-06 1.19194e-05 0.130478 0.973892 0.927744 -0.0132935 4.88989e-06 0.500192 -1.85424e-20 6.82064e-24 -1.85356e-20 0.00139493 0.997819 8.59157e-05 0.152527 2.85156 0.00139493 0.998155 0.6496 0.00104072 0.00187941 0.000859157 0.455687 0.00187941 0.433257 0.000126771 1.02 0.887258 0.534799 0.285467 1.71586e-07 3.053e-09 2395.22 3242.38 -0.0641431 0.482108 0.277695 0.2612 -0.591905 -0.169479 0.471174 -0.268756 -0.202419 1.187 1 1.76289e-258 289.057 1.01811e-255 1.9981 1.185 0.000299988 0.909439 0.626174 0.580098 0.394836 1.99843 126.486 82.4709 18.6362 60.1653 0.00408591 0 -40 10
0.286 8.29347e-09 2.53881e-06 0.0545577 0.0545445 0.0120462 3.76976e-06 0.00115401 0.0681971 0.000654755 0.0688472 0.850032 101.891 0.247011 0.704515 4.10853 0.052989 0.0387597 0.96124 0.0198922 0.00422706 0.0191544 0.00407108 0.00510776 0.00584564 0.20431 0.233826 57.9569 -87.8936 125.727 15.9902 145.006 0.000146916 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97003e-06 -85.6695 0.0929692 31198.9 300.116 0.983525 0.319147 0.762128 0.762123 9.99958 2.97987e-06 1.19194e-05 0.130478 0.973922 0.927759 -0.0132935 4.8899e-06 0.500193 -1.85434e-20 6.82102e-24 -1.85366e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998153 0.649722 0.00104073 0.00187941 0.000859157 0.455687 0.00187941 0.433268 0.000126774 1.02 0.887258 0.534799 0.285468 1.71586e-07 3.05301e-09 2395.2 3241.86 -0.0641053 0.482108 0.277695 0.261168 -0.591911 -0.169479 0.471287 -0.268754 -0.202533 1.188 1 1.06925e-258 289.094 6.17662e-256 1.99833 1.186 0.000299988 0.909207 0.626246 0.579428 0.394875 1.99866 126.498 82.4768 18.6365 60.1681 0.00408566 0 -40 10
0.287 8.32245e-09 2.53881e-06 0.054665 0.0546519 0.0120462 3.78293e-06 0.00115401 0.0683313 0.000654769 0.0689814 0.850063 101.891 0.247008 0.704554 4.10856 0.0529921 0.03876 0.96124 0.0198922 0.0042271 0.0191543 0.00407111 0.00510781 0.00584569 0.204312 0.233828 57.9569 -87.8936 125.73 15.9902 145.006 0.000146893 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97003e-06 -85.6695 0.0929692 31198.9 300.117 0.983525 0.319147 0.762007 0.762003 9.99958 2.97988e-06 1.19194e-05 0.130479 0.973952 0.927774 -0.0132935 4.88991e-06 0.500195 -1.85444e-20 6.8214e-24 -1.85376e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998151 0.649844 0.00104075 0.00187941 0.000859157 0.455687 0.00187941 0.433278 0.000126778 1.02 0.887259 0.534799 0.285468 1.71586e-07 3.05302e-09 2395.19 3241.35 -0.0640677 0.482108 0.277695 0.261136 -0.591917 -0.169479 0.471399 -0.268753 -0.202646 1.189 1 6.48531e-259 289.13 3.74721e-256 1.99855 1.187 0.000299988 0.908975 0.626317 0.578759 0.394914 1.99888 126.51 82.4826 18.6369 60.171 0.00408542 0 -40 10
0.288 8.35144e-09 2.53881e-06 0.0547723 0.0547592 0.0120462 3.79611e-06 0.00115401 0.0684653 0.000654782 0.0691155 0.850094 101.891 0.247005 0.704594 4.1086 0.0529953 0.0387604 0.96124 0.0198921 0.00422714 0.0191543 0.00407114 0.00510785 0.00584573 0.204314 0.233829 57.957 -87.8936 125.732 15.9901 145.006 0.00014687 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97003e-06 -85.6695 0.0929692 31198.9 300.118 0.983525 0.319147 0.761887 0.761883 9.99958 2.97988e-06 1.19194e-05 0.130479 0.973982 0.927789 -0.0132935 4.88992e-06 0.500196 -1.85454e-20 6.82178e-24 -1.85386e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998149 0.649966 0.00104076 0.00187941 0.000859157 0.455687 0.00187941 0.433289 0.000126781 1.02 0.887259 0.534799 0.285469 1.71586e-07 3.05302e-09 2395.17 3240.84 -0.0640302 0.482108 0.277694 0.261104 -0.591923 -0.169479 0.47151 -0.268752 -0.202759 1.19 1 3.93354e-259 289.166 2.27334e-256 1.99878 1.188 0.000299988 0.908744 0.626389 0.578092 0.394953 1.99911 126.522 82.4884 18.6372 60.1738 0.00408517 0 -40 10
0.289 8.38042e-09 2.53881e-06 0.0548794 0.0548665 0.0120462 3.80928e-06 0.00115401 0.0685993 0.000654795 0.0692495 0.850126 101.891 0.247002 0.704633 4.10863 0.0529984 0.0387607 0.961239 0.0198921 0.00422717 0.0191542 0.00407117 0.0051079 0.00584578 0.204316 0.233831 57.9571 -87.8936 125.734 15.9901 145.006 0.000146847 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97003e-06 -85.6695 0.0929692 31198.9 300.119 0.983525 0.319147 0.761767 0.761763 9.99958 2.97988e-06 1.19194e-05 0.13048 0.974012 0.927805 -0.0132935 4.88993e-06 0.500198 -1.85464e-20 6.82216e-24 -1.85396e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998147 0.650088 0.00104078 0.00187941 0.000859157 0.455687 0.00187941 0.4333 0.000126785 1.02 0.887259 0.534798 0.285469 1.71586e-07 3.05303e-09 2395.16 3240.33 -0.0639928 0.482108 0.277694 0.261072 -0.591929 -0.169479 0.471621 -0.268751 -0.202871 1.191 1 2.38581e-259 289.202 1.37918e-256 1.99901 1.189 0.000299988 0.908514 0.62646 0.577427 0.394992 1.99934 126.535 82.4942 18.6376 60.1766 0.00408493 0 -40 10
0.29 8.40941e-09 2.53881e-06 0.0549865 0.0549736 0.0120462 3.82246e-06 0.00115401 0.0687332 0.000654808 0.0693834 0.850157 101.891 0.246998 0.704673 4.10867 0.0530016 0.038761 0.961239 0.0198921 0.00422721 0.0191542 0.0040712 0.00510794 0.00584582 0.204318 0.233833 57.9571 -87.8936 125.736 15.9901 145.006 0.000146824 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561488 0.00138221 0.986996 0.991738 -2.97004e-06 -85.6695 0.0929693 31198.9 300.12 0.983524 0.319147 0.761648 0.761643 9.99958 2.97988e-06 1.19194e-05 0.13048 0.974042 0.92782 -0.0132935 4.88994e-06 0.500199 -1.85474e-20 6.82255e-24 -1.85406e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998144 0.65021 0.00104079 0.00187941 0.000859157 0.455687 0.00187941 0.43331 0.000126788 1.02 0.88726 0.534798 0.28547 1.71586e-07 3.05304e-09 2395.14 3239.82 -0.0639556 0.482108 0.277694 0.261041 -0.591935 -0.169479 0.471732 -0.26875 -0.202983 1.192 1 1.44707e-259 289.238 8.36713e-257 1.99924 1.19 0.000299987 0.908284 0.626531 0.576764 0.395031 1.99957 126.547 82.4999 18.6379 60.1794 0.00408468 0 -40 10
0.291 8.43839e-09 2.53881e-06 0.0550935 0.0550807 0.0120462 3.83563e-06 0.00115401 0.0688669 0.00065482 0.0695171 0.850188 101.891 0.246995 0.704713 4.1087 0.0530047 0.0387614 0.961239 0.019892 0.00422725 0.0191541 0.00407123 0.00510799 0.00584587 0.204319 0.233835 57.9572 -87.8936 125.738 15.99 145.006 0.000146801 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991738 -2.97004e-06 -85.6695 0.0929693 31198.9 300.121 0.983524 0.319147 0.761529 0.761524 9.99958 2.97988e-06 1.19194e-05 0.13048 0.974071 0.927835 -0.0132935 4.88995e-06 0.500201 -1.85484e-20 6.82293e-24 -1.85416e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998142 0.650332 0.00104081 0.00187941 0.000859157 0.455687 0.00187941 0.433321 0.000126791 1.02 0.88726 0.534798 0.285471 1.71586e-07 3.05304e-09 2395.12 3239.31 -0.0639185 0.482108 0.277693 0.261009 -0.591941 -0.169479 0.471842 -0.268749 -0.203095 1.193 1 8.77691e-260 289.273 5.07613e-257 1.99947 1.191 0.000299987 0.908056 0.626602 0.576103 0.39507 1.9998 126.559 82.5057 18.6382 60.1822 0.00408444 0 -40 10
0.292 8.46737e-09 2.53881e-06 0.0552004 0.0551877 0.0120461 3.84881e-06 0.00115401 0.0690005 0.000654833 0.0696508 0.85022 101.891 0.246992 0.704753 4.10874 0.0530079 0.0387617 0.961238 0.019892 0.00422728 0.0191541 0.00407126 0.00510803 0.00584591 0.204321 0.233836 57.9572 -87.8936 125.74 15.99 145.006 0.000146778 0.267061 192.946 0.310762 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991738 -2.97004e-06 -85.6695 0.0929693 31198.9 300.122 0.983524 0.319147 0.76141 0.761406 9.99958 2.97988e-06 1.19194e-05 0.130481 0.974101 0.92785 -0.0132935 4.88996e-06 0.500202 -1.85494e-20 6.82331e-24 -1.85425e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.99814 0.650454 0.00104082 0.00187941 0.000859157 0.455687 0.00187941 0.433332 0.000126795 1.02 0.887261 0.534798 0.285471 1.71586e-07 3.05305e-09 2395.11 3238.81 -0.0638815 0.482108 0.277693 0.260978 -0.591947 -0.16948 0.471952 -0.268747 -0.203206 1.194 1 5.32346e-260 289.309 3.07955e-257 1.99969 1.192 0.000299987 0.907828 0.626674 0.575444 0.395109 2.00002 126.571 82.5114 18.6386 60.1849 0.0040842 0 -40 10
0.293 8.49636e-09 2.53881e-06 0.0553073 0.0552946 0.0120461 3.86198e-06 0.00115401 0.0691341 0.000654846 0.0697843 0.850251 101.891 0.246989 0.704794 4.10878 0.0530111 0.038762 0.961238 0.0198919 0.00422732 0.019154 0.00407129 0.00510808 0.00584596 0.204323 0.233838 57.9573 -87.8936 125.742 15.9899 145.006 0.000146755 0.267061 192.946 0.310761 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991738 -2.97005e-06 -85.6695 0.0929693 31198.9 300.123 0.983524 0.319147 0.761292 0.761288 9.99958 2.97988e-06 1.19194e-05 0.130481 0.974131 0.927865 -0.0132935 4.88998e-06 0.500204 -1.85504e-20 6.82368e-24 -1.85435e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998138 0.650576 0.00104084 0.00187941 0.000859157 0.455687 0.00187941 0.433342 0.000126798 1.02 0.887261 0.534798 0.285472 1.71586e-07 3.05306e-09 2395.09 3238.31 -0.0638447 0.482108 0.277693 0.260946 -0.591952 -0.16948 0.472062 -0.268746 -0.203317 1.195 1 3.22884e-260 289.344 1.86829e-257 1.99992 1.193 0.000299987 0.907601 0.626745 0.574787 0.395148 2.00025 126.583 82.5171 18.6389 60.1877 0.00408395 0 -40 10
0.294 8.52534e-09 2.53881e-06 0.055414 0.0554014 0.0120461 3.87515e-06 0.00115401 0.0692675 0.000654859 0.0699178 0.850283 101.891 0.246986 0.704834 4.10881 0.0530143 0.0387624 0.961238 0.0198919 0.00422736 0.019154 0.00407132 0.00510813 0.005846 0.204325 0.23384 57.9574 -87.8936 125.744 15.9899 145.006 0.000146732 0.267061 192.946 0.310761 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991738 -2.97005e-06 -85.6695 0.0929693 31198.9 300.124 0.983524 0.319147 0.761174 0.76117 9.99958 2.97988e-06 1.19194e-05 0.130482 0.97416 0.92788 -0.0132935 4.88999e-06 0.500206 -1.85513e-20 6.82406e-24 -1.85445e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998136 0.650697 0.00104085 0.00187941 0.000859157 0.455687 0.00187941 0.433353 0.000126802 1.02 0.887261 0.534798 0.285472 1.71587e-07 3.05307e-09 2395.08 3237.81 -0.0638079 0.482108 0.277692 0.260915 -0.591958 -0.16948 0.472171 -0.268745 -0.203427 1.196 1 1.95839e-260 289.38 1.13344e-257 2.00015 1.194 0.000299987 0.907375 0.626816 0.574132 0.395187 2.00048 126.595 82.5228 18.6393 60.1905 0.00408371 0 -40 10
0.295 8.55432e-09 2.53881e-06 0.0555207 0.0555081 0.0120461 3.88833e-06 0.00115401 0.0694008 0.000654871 0.0700511 0.850315 101.891 0.246982 0.704875 4.10885 0.0530175 0.0387627 0.961237 0.0198918 0.0042274 0.019154 0.00407136 0.00510817 0.00584605 0.204327 0.233842 57.9574 -87.8937 125.746 15.9899 145.006 0.00014671 0.267061 192.946 0.310761 0.067395 0.00409445 0.000561489 0.00138221 0.986996 0.991738 -2.97005e-06 -85.6695 0.0929693 31198.9 300.125 0.983524 0.319147 0.761057 0.761052 9.99958 2.97988e-06 1.19194e-05 0.130482 0.974189 0.927895 -0.0132935 4.89e-06 0.500207 -1.85523e-20 6.82444e-24 -1.85455e-20 0.00139493 0.997819 8.59157e-05 0.152528 2.85156 0.00139493 0.998134 0.650819 0.00104087 0.00187941 0.000859157 0.455687 0.00187941 0.433364 0.000126805 1.02 0.887262 0.534798 0.285473 1.71587e-07 3.05307e-09 2395.06 3237.31 -0.0637713 0.482108 0.277692 0.260884 -0.591964 -0.16948 0.47228 -0.268744 -0.203537 1.197 1 1.18783e-260 289.415 6.87627e-258 2.00038 1.195 0.000299987 0.907149 0.626887 0.573478 0.395225 2.0007 126.607 82.5284 18.6396 60.1932 0.00408347 0 -40 10
0.296 8.58331e-09 2.53881e-06 0.0556272 0.0556147 0.0120461 3.9015e-06 0.00115401 0.0695341 0.000654884 0.0701843 0.850347 101.891 0.246979 0.704915 4.10888 0.0530207 0.038763 0.961237 0.0198918 0.00422744 0.0191539 0.00407139 0.00510822 0.00584609 0.204329 0.233844 57.9575 -87.8937 125.748 15.9898 145.006 0.000146687 0.267061 192.946 0.310761 0.0673949 0.00409445 0.000561489 0.00138221 0.986996 0.991738 -2.97006e-06 -85.6695 0.0929693 31198.9 300.126 0.983524 0.319147 0.76094 0.760935 9.99958 2.97988e-06 1.19194e-05 0.130482 0.974218 0.927909 -0.0132935 4.89001e-06 0.500209 -1.85533e-20 6.82482e-24 -1.85465e-20 0.00139493 0.997819 8.59158e-05 0.152528 2.85156 0.00139493 0.998132 0.650941 0.00104089 0.00187941 0.000859158 0.455687 0.00187941 0.433374 0.000126808 1.02 0.887262 0.534798 0.285474 1.71587e-07 3.05308e-09 2395.04 3236.81 -0.0637349 0.482108 0.277692 0.260853 -0.59197 -0.16948 0.472388 -0.268742 -0.203647 1.198 1 7.20452e-261 289.45 4.17165e-258 2.0006 1.196 0.000299987 0.906924 0.626958 0.572826 0.395264 2.00093 126.62 82.5341 18.6399 60.196 0.00408323 0 -40 10
0.297 8.61229e-09 2.53882e-06 0.0557337 0.0557213 0.0120461 3.91468e-06 0.00115401 0.0696672 0.000654896 0.0703175 0.850379 101.891 0.246976 0.704956 4.10892 0.053024 0.0387634 0.961237 0.0198917 0.00422748 0.0191539 0.00407142 0.00510827 0.00584614 0.204331 0.233846 57.9575 -87.8937 125.75 15.9898 145.006 0.000146665 0.267061 192.946 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991738 -2.97006e-06 -85.6695 0.0929693 31198.9 300.127 0.983524 0.319147 0.760823 0.760819 9.99958 2.97988e-06 1.19194e-05 0.130483 0.974248 0.927924 -0.0132935 4.89002e-06 0.50021 -1.85543e-20 6.8252e-24 -1.85475e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.99813 0.651062 0.0010409 0.00187941 0.000859158 0.455687 0.00187941 0.433385 0.000126812 1.02 0.887263 0.534798 0.285474 1.71587e-07 3.05309e-09 2395.03 3236.31 -0.0636985 0.482108 0.277692 0.260822 -0.591975 -0.16948 0.472496 -0.268741 -0.203756 1.199 1 4.36977e-261 289.485 2.53083e-258 2.00083 1.197 0.000299987 0.9067 0.627028 0.572177 0.395303 2.00115 126.632 82.5397 18.6402 60.1987 0.00408299 0 -40 10
0.298 8.64127e-09 2.53882e-06 0.0558401 0.0558277 0.0120461 3.92785e-06 0.00115401 0.0698002 0.000654909 0.0704505 0.850411 101.891 0.246973 0.704997 4.10896 0.0530272 0.0387637 0.961236 0.0198917 0.00422751 0.0191538 0.00407145 0.00510832 0.00584619 0.204333 0.233847 57.9576 -87.8937 125.752 15.9898 145.006 0.000146642 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991738 -2.97006e-06 -85.6695 0.0929693 31198.9 300.128 0.983524 0.319147 0.760707 0.760703 9.99958 2.97988e-06 1.19194e-05 0.130483 0.974277 0.927939 -0.0132935 4.89003e-06 0.500212 -1.85553e-20 6.82558e-24 -1.85484e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998128 0.651184 0.00104092 0.00187941 0.000859158 0.455687 0.00187941 0.433395 0.000126815 1.02 0.887263 0.534797 0.285475 1.71587e-07 3.0531e-09 2395.01 3235.82 -0.0636623 0.482108 0.277691 0.260791 -0.591981 -0.16948 0.472604 -0.26874 -0.203865 1.2 1 2.6504e-261 289.52 1.53538e-258 2.00105 1.198 0.000299987 0.906477 0.627099 0.571529 0.395341 2.00138 126.644 82.5453 18.6406 60.2014 0.00408276 0 -40 10
0.299 8.67026e-09 2.53882e-06 0.0559464 0.0559341 0.0120461 3.94103e-06 0.00115401 0.0699331 0.000654921 0.0705834 0.850443 101.891 0.24697 0.705038 4.10899 0.0530305 0.0387641 0.961236 0.0198916 0.00422755 0.0191538 0.00407148 0.00510836 0.00584623 0.204335 0.233849 57.9577 -87.8937 125.754 15.9897 145.006 0.00014662 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991738 -2.97007e-06 -85.6695 0.0929694 31198.9 300.129 0.983524 0.319147 0.760591 0.760587 9.99958 2.97988e-06 1.19194e-05 0.130483 0.974305 0.927954 -0.0132935 4.89005e-06 0.500213 -1.85563e-20 6.82595e-24 -1.85494e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998126 0.651305 0.00104093 0.00187941 0.000859158 0.455687 0.00187941 0.433406 0.000126819 1.02 0.887264 0.534797 0.285475 1.71587e-07 3.05311e-09 2394.99 3235.32 -0.0636262 0.482108 0.277691 0.260761 -0.591987 -0.16948 0.472711 -0.268739 -0.203974 1.201 1 1.60755e-261 289.555 9.31473e-259 2.00128 1.199 0.000299987 0.906254 0.62717 0.570883 0.39538 2.00161 126.656 82.5509 18.6409 60.2041 0.00408252 0 -40 10
0.3 8.69924e-09 2.53882e-06 0.0560527 0.0560404 0.012046 3.9542e-06 0.00115401 0.0700658 0.000654933 0.0707162 0.850475 101.891 0.246966 0.70508 4.10903 0.0530338 0.0387644 0.961236 0.0198916 0.00422759 0.0191537 0.00407152 0.00510841 0.00584628 0.204336 0.233851 57.9577 -87.8937 125.756 15.9897 145.006 0.000146598 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991738 -2.97007e-06 -85.6695 0.0929694 31198.9 300.13 0.983524 0.319147 0.760476 0.760471 9.99958 2.97988e-06 1.19194e-05 0.130484 0.974334 0.927968 -0.0132935 4.89006e-06 0.500215 -1.85572e-20 6.82633e-24 -1.85504e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998124 0.651427 0.00104095 0.00187941 0.000859158 0.455687 0.00187941 0.433417 0.000126822 1.02 0.887264 0.534797 0.285476 1.71587e-07 3.05311e-09 2394.98 3234.83 -0.0635902 0.482108 0.277691 0.26073 -0.591993 -0.16948 0.472818 -0.268738 -0.204082 1.202 1 9.75026e-262 289.589 5.65098e-259 2.00151 1.2 0.000299987 0.906033 0.62724 0.570239 0.395418 2.00183 126.668 82.5565 18.6412 60.2068 0.00408228 0 -40 10
0.301 8.72822e-09 2.53882e-06 0.0561588 0.0561466 0.012046 3.96737e-06 0.00115401 0.0701985 0.000654946 0.0708489 0.850507 101.891 0.246963 0.705121 4.10907 0.053037 0.0387648 0.961235 0.0198915 0.00422763 0.0191537 0.00407155 0.00510846 0.00584633 0.204338 0.233853 57.9578 -87.8937 125.758 15.9897 145.006 0.000146576 0.267061 192.945 0.310761 0.0673949 0.00409445 0.000561489 0.00138222 0.986996 0.991738 -2.97007e-06 -85.6695 0.0929694 31198.9 300.131 0.983524 0.319147 0.760361 0.760356 9.99958 2.97988e-06 1.19194e-05 0.130484 0.974363 0.927983 -0.0132935 4.89007e-06 0.500217 -1.85582e-20 6.82671e-24 -1.85514e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.998122 0.651548 0.00104096 0.00187941 0.000859158 0.455687 0.00187941 0.433427 0.000126825 1.02 0.887264 0.534797 0.285477 1.71587e-07 3.05312e-09 2394.96 3234.34 -0.0635544 0.482108 0.27769 0.260699 -0.591998 -0.16948 0.472925 -0.268736 -0.20419 1.203 1 5.91383e-262 289.624 3.42829e-259 2.00173 1.201 0.000299987 0.905812 0.627311 0.569596 0.395457 2.00206 126.68 82.562 18.6416 60.2095 0.00408205 0 -40 10
0.302 8.75721e-09 2.53882e-06 0.0562649 0.0562527 0.012046 3.98055e-06 0.00115401 0.0703311 0.000654958 0.0709815 0.85054 101.891 0.24696 0.705163 4.10911 0.0530403 0.0387651 0.961235 0.0198915 0.00422767 0.0191536 0.00407158 0.00510851 0.00584638 0.20434 0.233855 57.9578 -87.8937 125.76 15.9896 145.006 0.000146553 0.267061 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991738 -2.97008e-06 -85.6695 0.0929694 31198.9 300.132 0.983524 0.319147 0.760246 0.760241 9.99958 2.97989e-06 1.19194e-05 0.130485 0.974392 0.927997 -0.0132935 4.89008e-06 0.500218 -1.85592e-20 6.82709e-24 -1.85524e-20 0.00139494 0.997819 8.59158e-05 0.152528 2.85157 0.00139494 0.99812 0.65167 0.00104098 0.00187941 0.000859158 0.455687 0.00187941 0.433438 0.000126829 1.02 0.887265 0.534797 0.285477 1.71587e-07 3.05313e-09 2394.95 3233.86 -0.0635187 0.482108 0.27769 0.260669 -0.592004 -0.16948 0.473031 -0.268735 -0.204297 1.204 1 3.58692e-262 289.658 2.07984e-259 2.00196 1.202 0.000299987 0.905592 0.627381 0.568956 0.395495 2.00228 126.692 82.5676 18.6419 60.2122 0.00408181 0 -40 10
0.303 8.78619e-09 2.53882e-06 0.0563709 0.0563588 0.012046 3.99372e-06 0.00115401 0.0704636 0.00065497 0.0711139 0.850572 101.891 0.246956 0.705204 4.10914 0.0530436 0.0387655 0.961234 0.0198914 0.00422771 0.0191536 0.00407161 0.00510856 0.00584642 0.204342 0.233857 57.9579 -87.8937 125.762 15.9896 145.006 0.000146531 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991738 -2.97008e-06 -85.6695 0.0929694 31198.9 300.134 0.983524 0.319147 0.760132 0.760127 9.99958 2.97989e-06 1.19194e-05 0.130485 0.97442 0.928012 -0.0132935 4.8901e-06 0.50022 -1.85602e-20 6.82746e-24 -1.85533e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998118 0.651791 0.001041 0.00187941 0.000859159 0.455687 0.00187941 0.433448 0.000126832 1.02 0.887265 0.534797 0.285478 1.71587e-07 3.05314e-09 2394.93 3233.37 -0.0634831 0.482108 0.27769 0.260639 -0.592009 -0.16948 0.473137 -0.268734 -0.204405 1.205 1 2.17558e-262 289.693 1.26178e-259 2.00218 1.203 0.000299987 0.905372 0.627452 0.568317 0.395534 2.0025 126.704 82.5731 18.6422 60.2149 0.00408158 0 -40 10
0.304 8.81517e-09 2.53882e-06 0.0564768 0.0564647 0.012046 4.0069e-06 0.00115401 0.0705959 0.000654982 0.0712463 0.850605 101.891 0.246953 0.705246 4.10918 0.053047 0.0387659 0.961234 0.0198914 0.00422775 0.0191535 0.00407165 0.00510861 0.00584647 0.204344 0.233859 57.958 -87.8937 125.764 15.9895 145.006 0.000146509 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991738 -2.97008e-06 -85.6695 0.0929694 31198.9 300.135 0.983524 0.319147 0.760018 0.760013 9.99958 2.97989e-06 1.19194e-05 0.130486 0.974449 0.928026 -0.0132935 4.89011e-06 0.500222 -1.85611e-20 6.82784e-24 -1.85543e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998116 0.651913 0.00104101 0.00187941 0.000859159 0.455687 0.00187941 0.433459 0.000126836 1.02 0.887266 0.534797 0.285478 1.71587e-07 3.05315e-09 2394.91 3232.88 -0.0634476 0.482108 0.277689 0.260609 -0.592015 -0.16948 0.473242 -0.268733 -0.204511 1.206 1 1.31955e-262 289.727 7.65485e-260 2.00241 1.204 0.000299986 0.905153 0.627522 0.567681 0.395572 2.00273 126.716 82.5786 18.6425 60.2176 0.00408134 0 -40 10
0.305 8.84416e-09 2.53882e-06 0.0565826 0.0565706 0.012046 4.02007e-06 0.00115401 0.0707282 0.000654994 0.0713786 0.850637 101.891 0.24695 0.705288 4.10922 0.0530503 0.0387662 0.961234 0.0198913 0.00422779 0.0191535 0.00407168 0.00510866 0.00584652 0.204346 0.233861 57.958 -87.8937 125.766 15.9895 145.006 0.000146488 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991738 -2.97009e-06 -85.6695 0.0929695 31198.9 300.136 0.983524 0.319147 0.759904 0.7599 9.99958 2.97989e-06 1.19194e-05 0.130486 0.974477 0.928041 -0.0132935 4.89012e-06 0.500223 -1.85621e-20 6.82821e-24 -1.85553e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998114 0.652034 0.00104103 0.00187941 0.000859159 0.455687 0.00187941 0.43347 0.000126839 1.02 0.887266 0.534797 0.285479 1.71587e-07 3.05316e-09 2394.9 3232.4 -0.0634123 0.482108 0.277689 0.260578 -0.592021 -0.16948 0.473347 -0.268731 -0.204618 1.207 1 8.0035e-263 289.761 4.64397e-260 2.00263 1.205 0.000299986 0.904935 0.627592 0.567046 0.39561 2.00295 126.728 82.5841 18.6429 60.2202 0.00408111 0 -40 10
0.306 8.87314e-09 2.53882e-06 0.0566883 0.0566764 0.012046 4.03324e-06 0.00115401 0.0708604 0.000655006 0.0715108 0.85067 101.891 0.246946 0.705331 4.10926 0.0530536 0.0387666 0.961233 0.0198913 0.00422783 0.0191534 0.00407171 0.00510871 0.00584657 0.204348 0.233863 57.9581 -87.8937 125.768 15.9895 145.006 0.000146466 0.267062 192.945 0.310761 0.0673949 0.00409445 0.00056149 0.00138222 0.986996 0.991738 -2.97009e-06 -85.6695 0.0929695 31198.9 300.137 0.983524 0.319147 0.759791 0.759787 9.99958 2.97989e-06 1.19195e-05 0.130486 0.974505 0.928055 -0.0132935 4.89013e-06 0.500225 -1.85631e-20 6.82859e-24 -1.85562e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998112 0.652155 0.00104104 0.00187941 0.000859159 0.455687 0.00187941 0.43348 0.000126843 1.02 0.887267 0.534796 0.28548 1.71587e-07 3.05316e-09 2394.88 3231.92 -0.063377 0.482108 0.277689 0.260548 -0.592026 -0.169481 0.473452 -0.26873 -0.204724 1.208 1 4.85437e-263 289.795 2.81735e-260 2.00285 1.206 0.000299986 0.904718 0.627662 0.566412 0.395648 2.00318 126.74 82.5895 18.6432 60.2229 0.00408088 0 -40 10
0.307 8.90212e-09 2.53882e-06 0.0567939 0.0567821 0.0120459 4.04642e-06 0.00115401 0.0709924 0.000655018 0.0716428 0.850703 101.891 0.246943 0.705373 4.1093 0.053057 0.0387669 0.961233 0.0198912 0.00422787 0.0191534 0.00407175 0.00510876 0.00584662 0.20435 0.233865 57.9581 -87.8937 125.77 15.9894 145.006 0.000146444 0.267062 192.945 0.31076 0.0673948 0.00409446 0.00056149 0.00138222 0.986996 0.991738 -2.9701e-06 -85.6695 0.0929695 31198.9 300.138 0.983524 0.319147 0.759678 0.759674 9.99958 2.97989e-06 1.19195e-05 0.130487 0.974534 0.928069 -0.0132935 4.89015e-06 0.500227 -1.8564e-20 6.82896e-24 -1.85572e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.99811 0.652276 0.00104106 0.00187941 0.000859159 0.455687 0.00187941 0.433491 0.000126846 1.02 0.887267 0.534796 0.28548 1.71587e-07 3.05317e-09 2394.87 3231.44 -0.0633419 0.482108 0.277689 0.260518 -0.592032 -0.169481 0.473556 -0.268729 -0.204829 1.209 1 2.94432e-263 289.829 1.7092e-260 2.00308 1.207 0.000299986 0.904502 0.627732 0.565781 0.395687 2.0034 126.752 82.595 18.6435 60.2255 0.00408065 0 -40 10
0.308 8.9311e-09 2.53882e-06 0.0568995 0.0568877 0.0120459 4.05959e-06 0.00115401 0.0711243 0.00065503 0.0717748 0.850736 101.891 0.24694 0.705416 4.10934 0.0530604 0.0387673 0.961233 0.0198912 0.00422791 0.0191533 0.00407178 0.00510881 0.00584667 0.204352 0.233867 57.9582 -87.8937 125.772 15.9894 145.006 0.000146422 0.267062 192.945 0.31076 0.0673948 0.00409446 0.00056149 0.00138222 0.986996 0.991738 -2.9701e-06 -85.6695 0.0929695 31198.9 300.139 0.983524 0.319147 0.759566 0.759561 9.99958 2.97989e-06 1.19195e-05 0.130487 0.974562 0.928083 -0.0132935 4.89016e-06 0.500228 -1.8565e-20 6.82934e-24 -1.85582e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998108 0.652397 0.00104108 0.00187941 0.000859159 0.455687 0.00187941 0.433501 0.00012685 1.02 0.887268 0.534796 0.285481 1.71587e-07 3.05318e-09 2394.85 3230.96 -0.063307 0.482108 0.277688 0.260489 -0.592037 -0.169481 0.47366 -0.268727 -0.204935 1.21 1 1.78582e-263 289.863 1.03692e-260 2.0033 1.208 0.000299986 0.904286 0.627802 0.565152 0.395725 2.00362 126.764 82.6004 18.6438 60.2282 0.00408042 0 -40 10
0.309 8.96009e-09 2.53882e-06 0.0570049 0.0569932 0.0120459 4.07277e-06 0.00115401 0.0712562 0.000655041 0.0719066 0.850769 101.891 0.246936 0.705458 4.10937 0.0530637 0.0387677 0.961232 0.0198911 0.00422796 0.0191533 0.00407181 0.00510886 0.00584672 0.204354 0.233869 57.9583 -87.8937 125.774 15.9894 145.006 0.000146401 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991738 -2.9701e-06 -85.6695 0.0929695 31198.9 300.14 0.983524 0.319147 0.759454 0.759449 9.99958 2.97989e-06 1.19195e-05 0.130488 0.97459 0.928098 -0.0132935 4.89017e-06 0.50023 -1.8566e-20 6.82971e-24 -1.85592e-20 0.00139494 0.997819 8.59159e-05 0.152528 2.85157 0.00139494 0.998106 0.652519 0.00104109 0.00187941 0.000859159 0.455686 0.00187941 0.433512 0.000126853 1.02 0.887268 0.534796 0.285482 1.71587e-07 3.05319e-09 2394.83 3230.49 -0.0632721 0.482108 0.277688 0.260459 -0.592043 -0.169481 0.473764 -0.268726 -0.20504 1.211 1 1.08316e-263 289.896 6.29067e-261 2.00353 1.209 0.000299986 0.904071 0.627872 0.564524 0.395763 2.00385 126.776 82.6058 18.6441 60.2308 0.00408019 0 -40 10
0.31 8.98907e-09 2.53882e-06 0.0571103 0.0570986 0.0120459 4.08594e-06 0.00115401 0.0713879 0.000655053 0.0720384 0.850802 101.891 0.246933 0.705501 4.10941 0.0530671 0.0387681 0.961232 0.0198911 0.004228 0.0191532 0.00407185 0.00510891 0.00584677 0.204356 0.233871 57.9583 -87.8937 125.776 15.9893 145.006 0.000146379 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991738 -2.97011e-06 -85.6695 0.0929695 31198.9 300.141 0.983524 0.319147 0.759342 0.759338 9.99958 2.97989e-06 1.19195e-05 0.130488 0.974618 0.928112 -0.0132935 4.89019e-06 0.500232 -1.85669e-20 6.83008e-24 -1.85601e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998104 0.65264 0.00104111 0.00187941 0.00085916 0.455686 0.00187941 0.433522 0.000126856 1.02 0.887269 0.534796 0.285482 1.71587e-07 3.0532e-09 2394.82 3230.01 -0.0632374 0.482108 0.277688 0.260429 -0.592048 -0.169481 0.473867 -0.268725 -0.205144 1.212 1 6.56968e-264 289.93 3.81635e-261 2.00375 1.21 0.000299986 0.903857 0.627942 0.563898 0.395801 2.00407 126.788 82.6112 18.6445 60.2334 0.00407996 0 -40 10
0.311 9.01805e-09 2.53882e-06 0.0572156 0.057204 0.0120459 4.09911e-06 0.00115401 0.0715195 0.000655065 0.07217 0.850835 101.891 0.246929 0.705544 4.10945 0.0530705 0.0387684 0.961232 0.019891 0.00422804 0.0191532 0.00407188 0.00510896 0.00584682 0.204358 0.233873 57.9584 -87.8937 125.778 15.9893 145.006 0.000146358 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991738 -2.97011e-06 -85.6695 0.0929696 31198.9 300.142 0.983524 0.319147 0.759231 0.759227 9.99958 2.97989e-06 1.19195e-05 0.130488 0.974646 0.928126 -0.0132935 4.8902e-06 0.500233 -1.85679e-20 6.83046e-24 -1.85611e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998103 0.652761 0.00104112 0.00187942 0.00085916 0.455686 0.00187941 0.433533 0.00012686 1.02 0.887269 0.534796 0.285483 1.71587e-07 3.05321e-09 2394.8 3229.54 -0.0632027 0.482108 0.277687 0.2604 -0.592054 -0.169481 0.47397 -0.268723 -0.205248 1.213 1 3.98471e-264 289.963 2.31526e-261 2.00397 1.211 0.000299986 0.903643 0.628012 0.563274 0.395839 2.00429 126.8 82.6166 18.6448 60.236 0.00407973 0 -40 10
0.312 9.04703e-09 2.53882e-06 0.0573208 0.0573093 0.0120459 4.11229e-06 0.00115401 0.071651 0.000655076 0.0723015 0.850868 101.891 0.246926 0.705587 4.10949 0.0530739 0.0387688 0.961231 0.019891 0.00422808 0.0191531 0.00407192 0.00510901 0.00584687 0.204361 0.233875 57.9584 -87.8937 125.78 15.9893 145.006 0.000146336 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991738 -2.97012e-06 -85.6695 0.0929696 31198.8 300.144 0.983524 0.319147 0.75912 0.759116 9.99958 2.9799e-06 1.19195e-05 0.130489 0.974673 0.92814 -0.0132935 4.89021e-06 0.500235 -1.85689e-20 6.83083e-24 -1.8562e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998101 0.652882 0.00104114 0.00187942 0.00085916 0.455686 0.00187942 0.433544 0.000126863 1.02 0.88727 0.534796 0.285484 1.71587e-07 3.05322e-09 2394.78 3229.07 -0.0631682 0.482108 0.277687 0.26037 -0.592059 -0.169481 0.474072 -0.268722 -0.205352 1.214 1 2.41685e-264 289.996 1.40459e-261 2.00419 1.212 0.000299986 0.90343 0.628082 0.562651 0.395877 2.00452 126.812 82.622 18.6451 60.2386 0.00407951 0 -40 10
0.313 9.07601e-09 2.53882e-06 0.057426 0.0574144 0.0120459 4.12546e-06 0.00115401 0.0717825 0.000655088 0.0724329 0.850901 101.89 0.246923 0.70563 4.10953 0.0530774 0.0387692 0.961231 0.0198909 0.00422812 0.0191531 0.00407195 0.00510906 0.00584692 0.204363 0.233877 57.9585 -87.8937 125.782 15.9892 145.006 0.000146315 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991738 -2.97012e-06 -85.6695 0.0929696 31198.8 300.145 0.983524 0.319147 0.75901 0.759005 9.99958 2.9799e-06 1.19195e-05 0.130489 0.974701 0.928154 -0.0132935 4.89023e-06 0.500237 -1.85698e-20 6.8312e-24 -1.8563e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998099 0.653003 0.00104116 0.00187942 0.00085916 0.455686 0.00187942 0.433554 0.000126867 1.02 0.88727 0.534795 0.285484 1.71587e-07 3.05323e-09 2394.77 3228.6 -0.0631339 0.482108 0.277687 0.260341 -0.592065 -0.169481 0.474174 -0.268721 -0.205456 1.215 1 1.46589e-264 290.03 8.52121e-262 2.00442 1.213 0.000299986 0.903218 0.628151 0.562031 0.395915 2.00474 126.823 82.6273 18.6454 60.2412 0.00407928 0 -40 10
0.314 9.105e-09 2.53882e-06 0.057531 0.0575195 0.0120459 4.13863e-06 0.00115401 0.0719138 0.000655099 0.0725643 0.850935 101.89 0.246919 0.705674 4.10957 0.0530808 0.0387696 0.96123 0.0198909 0.00422817 0.019153 0.00407199 0.00510912 0.00584697 0.204365 0.233879 57.9586 -87.8937 125.784 15.9892 145.006 0.000146294 0.267062 192.945 0.31076 0.0673948 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97013e-06 -85.6695 0.0929696 31198.8 300.146 0.983524 0.319147 0.758899 0.758895 9.99958 2.9799e-06 1.19195e-05 0.13049 0.974729 0.928168 -0.0132935 4.89024e-06 0.500239 -1.85708e-20 6.83158e-24 -1.8564e-20 0.00139494 0.997819 8.5916e-05 0.152528 2.85157 0.00139494 0.998097 0.653123 0.00104117 0.00187942 0.00085916 0.455686 0.00187942 0.433565 0.00012687 1.02 0.887271 0.534795 0.285485 1.71588e-07 3.05324e-09 2394.75 3228.13 -0.0630996 0.482108 0.277686 0.260312 -0.59207 -0.169481 0.474276 -0.26872 -0.205559 1.216 1 8.89109e-265 290.063 5.16954e-262 2.00464 1.214 0.000299986 0.903007 0.628221 0.561412 0.395953 2.00496 126.835 82.6326 18.6457 60.2438 0.00407906 0 -40 10
0.315 9.13398e-09 2.53882e-06 0.057636 0.0576246 0.0120458 4.15181e-06 0.00115401 0.072045 0.000655111 0.0726955 0.850968 101.89 0.246916 0.705717 4.10961 0.0530843 0.03877 0.96123 0.0198908 0.00422821 0.019153 0.00407202 0.00510917 0.00584702 0.204367 0.233881 57.9586 -87.8937 125.786 15.9891 145.006 0.000146273 0.267062 192.945 0.31076 0.0673947 0.00409446 0.000561491 0.00138222 0.986996 0.991737 -2.97013e-06 -85.6695 0.0929696 31198.8 300.147 0.983524 0.319147 0.75879 0.758785 9.99958 2.9799e-06 1.19195e-05 0.13049 0.974756 0.928182 -0.0132935 4.89025e-06 0.50024 -1.85718e-20 6.83195e-24 -1.85649e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998095 0.653244 0.00104119 0.00187942 0.000859161 0.455686 0.00187942 0.433575 0.000126874 1.02 0.887271 0.534795 0.285486 1.71588e-07 3.05325e-09 2394.74 3227.66 -0.0630655 0.482108 0.277686 0.260283 -0.592075 -0.169481 0.474378 -0.268718 -0.205662 1.217 1 5.39272e-265 290.096 3.13619e-262 2.00486 1.215 0.000299986 0.902796 0.62829 0.560795 0.395991 2.00518 126.847 82.6379 18.646 60.2464 0.00407883 0 -40 10
0.316 9.16296e-09 2.53882e-06 0.0577409 0.0577295 0.0120458 4.16498e-06 0.00115401 0.0721761 0.000655122 0.0728266 0.851002 101.89 0.246912 0.705761 4.10966 0.0530877 0.0387703 0.96123 0.0198908 0.00422825 0.0191529 0.00407206 0.00510922 0.00584707 0.204369 0.233883 57.9587 -87.8937 125.788 15.9891 145.006 0.000146252 0.267062 192.945 0.31076 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97014e-06 -85.6695 0.0929697 31198.8 300.148 0.983524 0.319147 0.75868 0.758676 9.99958 2.9799e-06 1.19195e-05 0.130491 0.974784 0.928195 -0.0132935 4.89027e-06 0.500242 -1.85727e-20 6.83232e-24 -1.85659e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998093 0.653365 0.0010412 0.00187942 0.000859161 0.455686 0.00187942 0.433586 0.000126877 1.02 0.887272 0.534795 0.285487 1.71588e-07 3.05326e-09 2394.72 3227.19 -0.0630315 0.482108 0.277686 0.260254 -0.592081 -0.169481 0.474479 -0.268717 -0.205764 1.218 1 3.27085e-265 290.129 1.90262e-262 2.00508 1.216 0.000299986 0.902586 0.62836 0.56018 0.396029 2.0054 126.859 82.6432 18.6463 60.2489 0.00407861 0 -40 10
0.317 9.19194e-09 2.53882e-06 0.0578456 0.0578343 0.0120458 4.17815e-06 0.00115401 0.0723071 0.000655134 0.0729576 0.851035 101.89 0.246909 0.705805 4.1097 0.0530912 0.0387707 0.961229 0.0198907 0.0042283 0.0191529 0.00407209 0.00510928 0.00584712 0.204371 0.233885 57.9587 -87.8937 125.79 15.9891 145.007 0.000146231 0.267062 192.945 0.31076 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97014e-06 -85.6695 0.0929697 31198.8 300.149 0.983524 0.319147 0.758571 0.758567 9.99958 2.9799e-06 1.19195e-05 0.130491 0.974811 0.928209 -0.0132935 4.89028e-06 0.500244 -1.85737e-20 6.83269e-24 -1.85668e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998092 0.653486 0.00104122 0.00187942 0.000859161 0.455686 0.00187942 0.433596 0.000126881 1.02 0.887272 0.534795 0.285487 1.71588e-07 3.05327e-09 2394.7 3226.73 -0.0629976 0.482108 0.277685 0.260225 -0.592086 -0.169481 0.474579 -0.268716 -0.205866 1.219 1 1.98387e-265 290.161 1.15425e-262 2.00531 1.217 0.000299985 0.902377 0.628429 0.559566 0.396067 2.00562 126.871 82.6485 18.6467 60.2515 0.00407838 0 -40 10
0.318 9.22092e-09 2.53882e-06 0.0579504 0.0579391 0.0120458 4.19133e-06 0.00115401 0.0724379 0.000655145 0.0730885 0.851069 101.89 0.246905 0.705849 4.10974 0.0530947 0.0387711 0.961229 0.0198907 0.00422834 0.0191528 0.00407213 0.00510933 0.00584718 0.204373 0.233887 57.9588 -87.8937 125.792 15.989 145.007 0.00014621 0.267062 192.945 0.310759 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97014e-06 -85.6695 0.0929697 31198.8 300.151 0.983524 0.319147 0.758463 0.758458 9.99958 2.9799e-06 1.19195e-05 0.130492 0.974838 0.928223 -0.0132935 4.8903e-06 0.500246 -1.85746e-20 6.83306e-24 -1.85678e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.99809 0.653607 0.00104124 0.00187942 0.000859161 0.455686 0.00187942 0.433607 0.000126884 1.02 0.887273 0.534795 0.285488 1.71588e-07 3.05327e-09 2394.69 3226.27 -0.0629638 0.482108 0.277685 0.260196 -0.592092 -0.169481 0.47468 -0.268714 -0.205968 1.22 1 1.20328e-265 290.194 7.00247e-263 2.00553 1.218 0.000299985 0.902168 0.628498 0.558954 0.396104 2.00585 126.883 82.6537 18.647 60.254 0.00407816 0 -40 10
0.319 9.2499e-09 2.53882e-06 0.058055 0.0580438 0.0120458 4.2045e-06 0.00115401 0.0725687 0.000655156 0.0732193 0.851103 101.89 0.246902 0.705893 4.10978 0.0530982 0.0387715 0.961228 0.0198906 0.00422838 0.0191528 0.00407216 0.00510938 0.00584723 0.204375 0.233889 57.9589 -87.8937 125.794 15.989 145.007 0.000146189 0.267062 192.945 0.310759 0.0673947 0.00409446 0.000561492 0.00138222 0.986996 0.991737 -2.97015e-06 -85.6695 0.0929697 31198.8 300.152 0.983524 0.319147 0.758354 0.75835 9.99958 2.9799e-06 1.19195e-05 0.130492 0.974865 0.928237 -0.0132935 4.89031e-06 0.500248 -1.85756e-20 6.83343e-24 -1.85687e-20 0.00139494 0.997819 8.59161e-05 0.152528 2.85157 0.00139494 0.998088 0.653727 0.00104125 0.00187942 0.000859161 0.455686 0.00187942 0.433617 0.000126887 1.02 0.887273 0.534795 0.285489 1.71588e-07 3.05328e-09 2394.67 3225.81 -0.0629301 0.482108 0.277685 0.260167 -0.592097 -0.169481 0.47478 -0.268713 -0.206069 1.221 1 7.29825e-266 290.226 4.24816e-263 2.00575 1.219 0.000299985 0.901961 0.628568 0.558344 0.396142 2.00607 126.895 82.659 18.6473 60.2566 0.00407794 0 -40 10
0.32 9.27888e-09 2.53882e-06 0.0581595 0.0581484 0.0120458 4.21767e-06 0.00115401 0.0726994 0.000655167 0.07335 0.851137 101.89 0.246898 0.705937 4.10982 0.0531017 0.0387719 0.961228 0.0198906 0.00422843 0.0191527 0.0040722 0.00510944 0.00584728 0.204377 0.233891 57.9589 -87.8937 125.796 15.989 145.007 0.000146168 0.267062 192.945 0.310759 0.0673947 0.00409446 0.000561492 0.00138223 0.986996 0.991737 -2.97015e-06 -85.6695 0.0929698 31198.8 300.153 0.983524 0.319147 0.758246 0.758242 9.99958 2.97991e-06 1.19195e-05 0.130492 0.974893 0.92825 -0.0132935 4.89032e-06 0.500249 -1.85765e-20 6.8338e-24 -1.85697e-20 0.00139494 0.997819 8.59162e-05 0.152528 2.85157 0.00139494 0.998086 0.653848 0.00104127 0.00187942 0.000859162 0.455686 0.00187942 0.433628 0.000126891 1.02 0.887274 0.534794 0.285489 1.71588e-07 3.05329e-09 2394.65 3225.35 -0.0628966 0.482108 0.277685 0.260139 -0.592102 -0.169481 0.47488 -0.268712 -0.206171 1.222 1 4.42661e-266 290.259 2.57721e-263 2.00597 1.22 0.000299985 0.901754 0.628637 0.557736 0.39618 2.00629 126.906 82.6642 18.6476 60.2591 0.00407772 0 -40 10
0.321 9.30787e-09 2.53882e-06 0.058264 0.0582529 0.0120458 4.23085e-06 0.00115401 0.07283 0.000655178 0.0734806 0.851171 101.89 0.246895 0.705981 4.10986 0.0531052 0.0387723 0.961228 0.0198905 0.00422847 0.0191527 0.00407224 0.00510949 0.00584734 0.20438 0.233893 57.959 -87.8938 125.798 15.9889 145.007 0.000146147 0.267062 192.945 0.310759 0.0673947 0.00409447 0.000561492 0.00138223 0.986996 0.991737 -2.97016e-06 -85.6695 0.0929698 31198.8 300.154 0.983524 0.319147 0.758139 0.758134 9.99958 2.97991e-06 1.19195e-05 0.130493 0.97492 0.928264 -0.0132935 4.89034e-06 0.500251 -1.85775e-20 6.83417e-24 -1.85706e-20 0.00139494 0.997819 8.59162e-05 0.152529 2.85157 0.00139494 0.998085 0.653969 0.00104129 0.00187942 0.000859162 0.455686 0.00187942 0.433638 0.000126894 1.02 0.887274 0.534794 0.28549 1.71588e-07 3.0533e-09 2394.64 3224.89 -0.0628631 0.482108 0.277684 0.26011 -0.592108 -0.169482 0.474979 -0.26871 -0.206271 1.223 1 2.68488e-266 290.291 1.5635e-263 2.00619 1.221 0.000299985 0.901547 0.628706 0.557129 0.396217 2.00651 126.918 82.6694 18.6479 60.2616 0.0040775 0 -40 10
0.322 9.33685e-09 2.53882e-06 0.0583684 0.0583573 0.0120457 4.24402e-06 0.00115401 0.0729604 0.00065519 0.073611 0.851205 101.89 0.246891 0.706026 4.10991 0.0531087 0.0387727 0.961227 0.0198905 0.00422851 0.0191526 0.00407227 0.00510955 0.00584739 0.204382 0.233896 57.959 -87.8938 125.799 15.9889 145.007 0.000146127 0.267062 192.945 0.310759 0.0673947 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97016e-06 -85.6695 0.0929698 31198.8 300.155 0.983524 0.319147 0.758032 0.758027 9.99958 2.97991e-06 1.19195e-05 0.130493 0.974946 0.928277 -0.0132935 4.89035e-06 0.500253 -1.85784e-20 6.83454e-24 -1.85716e-20 0.00139494 0.997819 8.59162e-05 0.152529 2.85157 0.00139494 0.998083 0.654089 0.0010413 0.00187942 0.000859162 0.455686 0.00187942 0.433649 0.000126898 1.02 0.887275 0.534794 0.285491 1.71588e-07 3.05331e-09 2394.62 3224.43 -0.0628298 0.482108 0.277684 0.260082 -0.592113 -0.169482 0.475078 -0.268709 -0.206372 1.224 1 1.62846e-266 290.323 9.48522e-264 2.00641 1.222 0.000299985 0.901342 0.628775 0.556524 0.396255 2.00673 126.93 82.6746 18.6482 60.2642 0.00407728 0 -40 10
0.323 9.36583e-09 2.53882e-06 0.0584726 0.0584617 0.0120457 4.25719e-06 0.00115401 0.0730908 0.000655201 0.0737414 0.851239 101.89 0.246888 0.706071 4.10995 0.0531123 0.0387731 0.961227 0.0198904 0.00422856 0.0191526 0.00407231 0.0051096 0.00584744 0.204384 0.233898 57.9591 -87.8938 125.801 15.9889 145.007 0.000146106 0.267062 192.945 0.310759 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97017e-06 -85.6694 0.0929698 31198.8 300.157 0.983524 0.319147 0.757925 0.75792 9.99958 2.97991e-06 1.19195e-05 0.130494 0.974973 0.928291 -0.0132935 4.89037e-06 0.500255 -1.85794e-20 6.83491e-24 -1.85725e-20 0.00139494 0.997819 8.59162e-05 0.152529 2.85157 0.00139494 0.998081 0.65421 0.00104132 0.00187942 0.000859162 0.455686 0.00187942 0.433659 0.000126901 1.02 0.887275 0.534794 0.285492 1.71588e-07 3.05332e-09 2394.61 3223.98 -0.0627966 0.482108 0.277684 0.260053 -0.592118 -0.169482 0.475176 -0.268707 -0.206472 1.225 1 9.87711e-267 290.356 5.75435e-264 2.00663 1.223 0.000299985 0.901137 0.628844 0.555921 0.396293 2.00695 126.942 82.6797 18.6485 60.2667 0.00407706 0 -40 10
0.324 9.39481e-09 2.53882e-06 0.0585769 0.0585659 0.0120457 4.27037e-06 0.00115401 0.0732211 0.000655212 0.0738717 0.851273 101.89 0.246884 0.706115 4.10999 0.0531158 0.0387735 0.961227 0.0198903 0.0042286 0.0191525 0.00407235 0.00510966 0.0058475 0.204386 0.2339 57.9592 -87.8938 125.803 15.9888 145.007 0.000146085 0.267062 192.945 0.310759 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97017e-06 -85.6694 0.0929699 31198.8 300.158 0.983524 0.319147 0.757818 0.757814 9.99958 2.97991e-06 1.19195e-05 0.130494 0.975 0.928304 -0.0132935 4.89038e-06 0.500257 -1.85803e-20 6.83528e-24 -1.85735e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998079 0.65433 0.00104134 0.00187942 0.000859163 0.455686 0.00187942 0.43367 0.000126905 1.02 0.887276 0.534794 0.285492 1.71588e-07 3.05333e-09 2394.59 3223.53 -0.0627636 0.482108 0.277683 0.260025 -0.592123 -0.169482 0.475275 -0.268706 -0.206571 1.226 1 5.99077e-267 290.388 3.49096e-264 2.00685 1.224 0.000299985 0.900932 0.628913 0.55532 0.39633 2.00717 126.954 82.6849 18.6488 60.2692 0.00407684 0 -40 10
0.325 9.42379e-09 2.53882e-06 0.058681 0.0586701 0.0120457 4.28354e-06 0.00115401 0.0733512 0.000655222 0.0740018 0.851308 101.89 0.246881 0.70616 4.11003 0.0531194 0.0387739 0.961226 0.0198903 0.00422865 0.0191524 0.00407238 0.00510971 0.00584755 0.204388 0.233902 57.9592 -87.8938 125.805 15.9888 145.007 0.000146065 0.267063 192.944 0.310759 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97018e-06 -85.6694 0.0929699 31198.8 300.159 0.983524 0.319147 0.757712 0.757708 9.99958 2.97991e-06 1.19195e-05 0.130495 0.975027 0.928318 -0.0132935 4.8904e-06 0.500259 -1.85813e-20 6.83565e-24 -1.85744e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998078 0.654451 0.00104135 0.00187942 0.000859163 0.455686 0.00187942 0.43368 0.000126908 1.02 0.887276 0.534794 0.285493 1.71588e-07 3.05335e-09 2394.57 3223.07 -0.0627306 0.482108 0.277683 0.259997 -0.592129 -0.169482 0.475373 -0.268705 -0.206671 1.227 1 3.63359e-267 290.419 2.11784e-264 2.00707 1.225 0.000299985 0.900729 0.628982 0.55472 0.396368 2.00739 126.965 82.69 18.6491 60.2716 0.00407663 0 -40 10
0.326 9.45277e-09 2.53882e-06 0.058785 0.0587742 0.0120457 4.29671e-06 0.00115401 0.0734813 0.000655233 0.0741319 0.851342 101.89 0.246877 0.706206 4.11008 0.053123 0.0387743 0.961226 0.0198902 0.00422869 0.0191524 0.00407242 0.00510977 0.0058476 0.204391 0.233904 57.9593 -87.8938 125.807 15.9887 145.007 0.000146045 0.267063 192.944 0.310758 0.0673946 0.00409447 0.000561493 0.00138223 0.986996 0.991737 -2.97018e-06 -85.6694 0.0929699 31198.8 300.16 0.983524 0.319147 0.757606 0.757602 9.99958 2.97991e-06 1.19195e-05 0.130495 0.975053 0.928331 -0.0132935 4.89041e-06 0.50026 -1.85822e-20 6.83602e-24 -1.85754e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998076 0.654571 0.00104137 0.00187942 0.000859163 0.455686 0.00187942 0.433691 0.000126912 1.02 0.887277 0.534794 0.285494 1.71588e-07 3.05336e-09 2394.56 3222.62 -0.0626978 0.482108 0.277683 0.259969 -0.592134 -0.169482 0.47547 -0.268703 -0.20677 1.228 1 2.20388e-267 290.451 1.28481e-264 2.00729 1.226 0.000299985 0.900526 0.62905 0.554122 0.396405 2.00761 126.977 82.6952 18.6494 60.2741 0.00407641 0 -40 10
0.327 9.48175e-09 2.53882e-06 0.058889 0.0588782 0.0120457 4.30989e-06 0.00115401 0.0736112 0.000655244 0.0742619 0.851376 101.89 0.246873 0.706251 4.11012 0.0531265 0.0387747 0.961225 0.0198902 0.00422874 0.0191523 0.00407246 0.00510982 0.00584766 0.204393 0.233906 57.9593 -87.8938 125.809 15.9887 145.007 0.000146024 0.267063 192.944 0.310758 0.0673946 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.97019e-06 -85.6694 0.0929699 31198.8 300.161 0.983524 0.319147 0.757501 0.757497 9.99958 2.97992e-06 1.19196e-05 0.130496 0.97508 0.928345 -0.0132935 4.89043e-06 0.500262 -1.85832e-20 6.83639e-24 -1.85763e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998074 0.654691 0.00104139 0.00187942 0.000859163 0.455685 0.00187942 0.433701 0.000126915 1.02 0.887278 0.534793 0.285495 1.71588e-07 3.05337e-09 2394.54 3222.18 -0.062665 0.482108 0.277682 0.259941 -0.592139 -0.169482 0.475567 -0.268702 -0.206868 1.229 1 1.33672e-267 290.483 7.79449e-265 2.00751 1.227 0.000299985 0.900324 0.629119 0.553526 0.396443 2.00783 126.989 82.7003 18.6497 60.2766 0.0040762 0 -40 10
0.328 9.51073e-09 2.53882e-06 0.0589929 0.0589821 0.0120457 4.32306e-06 0.00115401 0.0737411 0.000655255 0.0743917 0.851411 101.89 0.24687 0.706296 4.11016 0.0531301 0.0387751 0.961225 0.0198901 0.00422879 0.0191523 0.00407249 0.00510988 0.00584771 0.204395 0.233909 57.9594 -87.8938 125.811 15.9887 145.007 0.000146004 0.267063 192.944 0.310758 0.0673946 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.9702e-06 -85.6694 0.09297 31198.7 300.163 0.983524 0.319147 0.757396 0.757392 9.99958 2.97992e-06 1.19196e-05 0.130496 0.975106 0.928358 -0.0132935 4.89044e-06 0.500264 -1.85841e-20 6.83676e-24 -1.85773e-20 0.00139494 0.997819 8.59163e-05 0.152529 2.85157 0.00139494 0.998073 0.654812 0.0010414 0.00187942 0.000859163 0.455685 0.00187942 0.433712 0.000126919 1.02 0.887278 0.534793 0.285495 1.71589e-07 3.05338e-09 2394.52 3221.73 -0.0626324 0.482108 0.277682 0.259913 -0.592144 -0.169482 0.475664 -0.268701 -0.206967 1.23 1 8.10762e-268 290.515 4.72863e-265 2.00773 1.228 0.000299985 0.900122 0.629188 0.552931 0.39648 2.00805 127 82.7053 18.65 60.2791 0.00407598 0 -40 10
0.329 9.53971e-09 2.53882e-06 0.0590966 0.0590859 0.0120457 4.33623e-06 0.00115401 0.0738708 0.000655266 0.0745215 0.851446 101.89 0.246866 0.706342 4.11021 0.0531337 0.0387755 0.961224 0.0198901 0.00422883 0.0191522 0.00407253 0.00510993 0.00584777 0.204397 0.233911 57.9595 -87.8938 125.812 15.9886 145.007 0.000145984 0.267063 192.944 0.310758 0.0673945 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.9702e-06 -85.6694 0.09297 31198.7 300.164 0.983524 0.319147 0.757291 0.757287 9.99958 2.97992e-06 1.19196e-05 0.130497 0.975133 0.928371 -0.0132935 4.89046e-06 0.500266 -1.8585e-20 6.83713e-24 -1.85782e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998071 0.654932 0.00104142 0.00187942 0.000859164 0.455685 0.00187942 0.433722 0.000126922 1.02 0.887279 0.534793 0.285496 1.71589e-07 3.05339e-09 2394.51 3221.28 -0.0625999 0.482108 0.277682 0.259885 -0.592149 -0.169482 0.475761 -0.268699 -0.207065 1.231 1 4.91752e-268 290.546 2.86868e-265 2.00795 1.229 0.000299984 0.899922 0.629256 0.552338 0.396517 2.00826 127.012 82.7104 18.6503 60.2815 0.00407577 0 -40 10
0.33 9.56869e-09 2.53882e-06 0.0592003 0.0591897 0.0120456 4.34941e-06 0.00115401 0.0740004 0.000655276 0.0746511 0.85148 101.89 0.246863 0.706388 4.11025 0.0531374 0.038776 0.961224 0.01989 0.00422888 0.0191522 0.00407257 0.00510999 0.00584783 0.2044 0.233913 57.9595 -87.8938 125.814 15.9886 145.007 0.000145964 0.267063 192.944 0.310758 0.0673945 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.97021e-06 -85.6694 0.09297 31198.7 300.165 0.983524 0.319147 0.757187 0.757183 9.99958 2.97992e-06 1.19196e-05 0.130497 0.975159 0.928384 -0.0132935 4.89047e-06 0.500268 -1.8586e-20 6.83749e-24 -1.85791e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998069 0.655052 0.00104144 0.00187942 0.000859164 0.455685 0.00187942 0.433733 0.000126926 1.02 0.887279 0.534793 0.285497 1.71589e-07 3.0534e-09 2394.49 3220.84 -0.0625675 0.482108 0.277682 0.259857 -0.592154 -0.169482 0.475857 -0.268698 -0.207162 1.232 1 2.98263e-268 290.577 1.74032e-265 2.00817 1.23 0.000299984 0.899722 0.629325 0.551747 0.396555 2.00848 127.024 82.7155 18.6506 60.284 0.00407555 0 -40 10
0.331 9.59767e-09 2.53882e-06 0.059304 0.0592934 0.0120456 4.36258e-06 0.00115401 0.07413 0.000655287 0.0747807 0.851515 101.89 0.246859 0.706433 4.1103 0.053141 0.0387764 0.961224 0.01989 0.00422892 0.0191521 0.00407261 0.00511005 0.00584788 0.204402 0.233915 57.9596 -87.8938 125.816 15.9886 145.007 0.000145944 0.267063 192.944 0.310758 0.0673945 0.00409447 0.000561494 0.00138223 0.986996 0.991737 -2.97021e-06 -85.6694 0.09297 31198.7 300.166 0.983524 0.319147 0.757083 0.757079 9.99958 2.97992e-06 1.19196e-05 0.130497 0.975185 0.928397 -0.0132935 4.89049e-06 0.50027 -1.85869e-20 6.83786e-24 -1.85801e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998068 0.655172 0.00104145 0.00187942 0.000859164 0.455685 0.00187942 0.433743 0.000126929 1.02 0.88728 0.534793 0.285498 1.71589e-07 3.05341e-09 2394.48 3220.4 -0.0625353 0.482108 0.277681 0.25983 -0.59216 -0.169482 0.475953 -0.268696 -0.207259 1.233 1 1.80906e-268 290.609 1.05579e-265 2.00839 1.231 0.000299984 0.899522 0.629393 0.551157 0.396592 2.0087 127.036 82.7205 18.6509 60.2864 0.00407534 0 -40 10
0.332 9.62665e-09 2.53882e-06 0.0594075 0.059397 0.0120456 4.37575e-06 0.00115401 0.0742594 0.000655298 0.0749101 0.85155 101.89 0.246855 0.706479 4.11034 0.0531446 0.0387768 0.961223 0.0198899 0.00422897 0.0191521 0.00407265 0.00511011 0.00584794 0.204404 0.233917 57.9597 -87.8938 125.818 15.9885 145.007 0.000145924 0.267063 192.944 0.310758 0.0673945 0.00409448 0.000561495 0.00138223 0.986996 0.991737 -2.97022e-06 -85.6694 0.0929701 31198.7 300.168 0.983524 0.319147 0.756979 0.756975 9.99958 2.97992e-06 1.19196e-05 0.130498 0.975211 0.928411 -0.0132935 4.8905e-06 0.500272 -1.85879e-20 6.83823e-24 -1.8581e-20 0.00139494 0.997819 8.59164e-05 0.152529 2.85157 0.00139494 0.998066 0.655292 0.00104147 0.00187942 0.000859164 0.455685 0.00187942 0.433753 0.000126933 1.02 0.88728 0.534793 0.285499 1.71589e-07 3.05342e-09 2394.46 3219.96 -0.0625031 0.482108 0.277681 0.259802 -0.592165 -0.169482 0.476048 -0.268695 -0.207356 1.234 1 1.09725e-268 290.64 6.40505e-266 2.00861 1.232 0.000299984 0.899324 0.629461 0.55057 0.396629 2.00892 127.047 82.7255 18.6512 60.2889 0.00407513 0 -40 10
0.333 9.65563e-09 2.53882e-06 0.059511 0.0595005 0.0120456 4.38892e-06 0.00115401 0.0743887 0.000655308 0.0750394 0.851585 101.89 0.246852 0.706526 4.11039 0.0531483 0.0387772 0.961223 0.0198898 0.00422902 0.019152 0.00407269 0.00511016 0.00584799 0.204407 0.23392 57.9597 -87.8938 125.82 15.9885 145.007 0.000145904 0.267063 192.944 0.310758 0.0673945 0.00409448 0.000561495 0.00138223 0.986996 0.991737 -2.97022e-06 -85.6694 0.0929701 31198.7 300.169 0.983524 0.319147 0.756876 0.756872 9.99958 2.97992e-06 1.19196e-05 0.130498 0.975237 0.928424 -0.0132935 4.89052e-06 0.500274 -1.85888e-20 6.83859e-24 -1.8582e-20 0.00139495 0.997819 8.59165e-05 0.152529 2.85157 0.00139495 0.998064 0.655413 0.00104149 0.00187942 0.000859165 0.455685 0.00187942 0.433764 0.000126936 1.02 0.887281 0.534792 0.285499 1.71589e-07 3.05343e-09 2394.44 3219.52 -0.062471 0.482108 0.277681 0.259775 -0.59217 -0.169482 0.476144 -0.268694 -0.207453 1.235 1 6.65514e-269 290.671 3.8857e-266 2.00882 1.233 0.000299984 0.899126 0.62953 0.549983 0.396666 2.00914 127.059 82.7305 18.6515 60.2913 0.00407492 0 -40 10
0.334 9.68461e-09 2.53882e-06 0.0596143 0.0596039 0.0120456 4.4021e-06 0.00115401 0.0745179 0.000655319 0.0751687 0.85162 101.89 0.246848 0.706572 4.11043 0.053152 0.0387776 0.961222 0.0198898 0.00422907 0.0191519 0.00407272 0.00511022 0.00584805 0.204409 0.233922 57.9598 -87.8938 125.822 15.9885 145.007 0.000145884 0.267063 192.944 0.310757 0.0673945 0.00409448 0.000561495 0.00138223 0.986996 0.991737 -2.97023e-06 -85.6694 0.0929701 31198.7 300.17 0.983524 0.319147 0.756773 0.756769 9.99958 2.97993e-06 1.19196e-05 0.130499 0.975263 0.928437 -0.0132935 4.89053e-06 0.500276 -1.85897e-20 6.83896e-24 -1.85829e-20 0.00139495 0.997819 8.59165e-05 0.152529 2.85157 0.00139495 0.998063 0.655533 0.0010415 0.00187942 0.000859165 0.455685 0.00187942 0.433774 0.00012694 1.02 0.887281 0.534792 0.2855 1.71589e-07 3.05344e-09 2394.43 3219.08 -0.0624391 0.482108 0.27768 0.259747 -0.592175 -0.169482 0.476238 -0.268692 -0.207549 1.236 1 4.03655e-269 290.702 2.3573e-266 2.00904 1.234 0.000299984 0.898928 0.629598 0.549399 0.396703 2.00935 127.071 82.7355 18.6518 60.2937 0.00407471 0 -40 10
0.335 9.71359e-09 2.53882e-06 0.0597176 0.0597072 0.0120456 4.41527e-06 0.00115401 0.0746471 0.000655329 0.0752978 0.851655 101.89 0.246844 0.706618 4.11048 0.0531556 0.0387781 0.961222 0.0198897 0.00422911 0.0191519 0.00407276 0.00511028 0.00584811 0.204411 0.233924 57.9598 -87.8938 125.823 15.9884 145.007 0.000145864 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561495 0.00138224 0.986996 0.991737 -2.97024e-06 -85.6694 0.0929702 31198.7 300.172 0.983524 0.319147 0.756671 0.756666 9.99958 2.97993e-06 1.19196e-05 0.130499 0.975289 0.92845 -0.0132935 4.89055e-06 0.500278 -1.85907e-20 6.83933e-24 -1.85838e-20 0.00139495 0.997819 8.59165e-05 0.152529 2.85157 0.00139495 0.998061 0.655653 0.00104152 0.00187943 0.000859165 0.455685 0.00187942 0.433785 0.000126943 1.02 0.887282 0.534792 0.285501 1.71589e-07 3.05345e-09 2394.41 3218.64 -0.0624073 0.482108 0.27768 0.25972 -0.59218 -0.169483 0.476333 -0.268691 -0.207645 1.237 1 2.44829e-269 290.733 1.43008e-266 2.00926 1.235 0.000299984 0.898732 0.629666 0.548816 0.396741 2.00957 127.082 82.7405 18.6521 60.2961 0.0040745 0 -40 10
0.336 9.74257e-09 2.53882e-06 0.0598209 0.0598105 0.0120456 4.42844e-06 0.00115401 0.0747761 0.000655339 0.0754268 0.851691 101.889 0.246841 0.706665 4.11052 0.0531593 0.0387785 0.961221 0.0198897 0.00422916 0.0191518 0.0040728 0.00511034 0.00584817 0.204414 0.233927 57.9599 -87.8938 125.825 15.9884 145.007 0.000145845 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986996 0.991737 -2.97024e-06 -85.6694 0.0929702 31198.7 300.173 0.983524 0.319147 0.756568 0.756564 9.99958 2.97993e-06 1.19196e-05 0.1305 0.975315 0.928463 -0.0132935 4.89057e-06 0.50028 -1.85916e-20 6.83969e-24 -1.85848e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.99806 0.655773 0.00104154 0.00187943 0.000859166 0.455685 0.00187943 0.433795 0.000126946 1.02 0.887283 0.534792 0.285502 1.71589e-07 3.05346e-09 2394.39 3218.21 -0.0623756 0.482108 0.27768 0.259693 -0.592185 -0.169483 0.476427 -0.268689 -0.207741 1.238 1 1.48496e-269 290.763 8.67575e-267 2.00948 1.236 0.000299984 0.898536 0.629734 0.548235 0.396778 2.00979 127.094 82.7454 18.6524 60.2985 0.00407429 0 -40 10
0.337 9.77155e-09 2.53882e-06 0.059924 0.0599137 0.0120455 4.44161e-06 0.00115401 0.074905 0.00065535 0.0755557 0.851726 101.889 0.246837 0.706712 4.11057 0.053163 0.0387789 0.961221 0.0198896 0.00422921 0.0191518 0.00407284 0.0051104 0.00584822 0.204416 0.233929 57.96 -87.8938 125.827 15.9883 145.007 0.000145825 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986996 0.991737 -2.97025e-06 -85.6694 0.0929702 31198.7 300.174 0.983524 0.319147 0.756467 0.756462 9.99958 2.97993e-06 1.19196e-05 0.1305 0.97534 0.928475 -0.0132935 4.89058e-06 0.500282 -1.85925e-20 6.84006e-24 -1.85857e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.998058 0.655892 0.00104155 0.00187943 0.000859166 0.455685 0.00187943 0.433806 0.00012695 1.02 0.887283 0.534792 0.285503 1.71589e-07 3.05348e-09 2394.38 3217.77 -0.062344 0.482109 0.277679 0.259666 -0.59219 -0.169483 0.476521 -0.268688 -0.207836 1.239 1 9.00676e-270 290.794 5.26323e-267 2.00969 1.237 0.000299984 0.89834 0.629802 0.547655 0.396815 2.01001 127.105 82.7503 18.6526 60.3009 0.00407408 0 -40 10
0.338 9.80053e-09 2.53882e-06 0.060027 0.0600167 0.0120455 4.45479e-06 0.00115401 0.0750338 0.00065536 0.0756845 0.851761 101.889 0.246833 0.706758 4.11061 0.0531667 0.0387794 0.961221 0.0198895 0.00422926 0.0191517 0.00407288 0.00511046 0.00584828 0.204418 0.233931 57.96 -87.8938 125.829 15.9883 145.007 0.000145805 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986996 0.991737 -2.97025e-06 -85.6694 0.0929702 31198.7 300.175 0.983524 0.319147 0.756365 0.75636 9.99958 2.97993e-06 1.19196e-05 0.130501 0.975366 0.928488 -0.0132935 4.8906e-06 0.500284 -1.85935e-20 6.84042e-24 -1.85866e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.998056 0.656012 0.00104157 0.00187943 0.000859166 0.455685 0.00187943 0.433816 0.000126953 1.02 0.887284 0.534792 0.285503 1.71589e-07 3.05349e-09 2394.36 3217.34 -0.0623125 0.482109 0.277679 0.259639 -0.592195 -0.169483 0.476614 -0.268686 -0.207931 1.24 1 5.46287e-270 290.825 3.19299e-267 2.00991 1.238 0.000299984 0.898146 0.62987 0.547077 0.396852 2.01022 127.117 82.7553 18.6529 60.3033 0.00407387 0 -40 10
0.339 9.82951e-09 2.53882e-06 0.06013 0.0601198 0.0120455 4.46796e-06 0.00115401 0.0751625 0.00065537 0.0758133 0.851797 101.889 0.24683 0.706805 4.11066 0.0531705 0.0387798 0.96122 0.0198895 0.00422931 0.0191517 0.00407292 0.00511052 0.00584834 0.204421 0.233934 57.9601 -87.8938 125.831 15.9883 145.007 0.000145786 0.267063 192.944 0.310757 0.0673944 0.00409448 0.000561496 0.00138224 0.986996 0.991737 -2.97026e-06 -85.6694 0.0929703 31198.7 300.177 0.983524 0.319147 0.756264 0.756259 9.99958 2.97993e-06 1.19196e-05 0.130501 0.975391 0.928501 -0.0132935 4.89061e-06 0.500286 -1.85944e-20 6.84079e-24 -1.85876e-20 0.00139495 0.997819 8.59166e-05 0.152529 2.85157 0.00139495 0.998055 0.656132 0.00104159 0.00187943 0.000859166 0.455685 0.00187943 0.433826 0.000126957 1.02 0.887284 0.534791 0.285504 1.7159e-07 3.0535e-09 2394.35 3216.91 -0.0622811 0.482109 0.277679 0.259612 -0.5922 -0.169483 0.476708 -0.268685 -0.208026 1.241 1 3.3134e-270 290.855 1.93706e-267 2.01013 1.239 0.000299984 0.897952 0.629938 0.546501 0.396889 2.01044 127.129 82.7602 18.6532 60.3057 0.00407366 0 -40 10
0.34 9.85849e-09 2.53882e-06 0.0602329 0.0602227 0.0120455 4.48113e-06 0.00115401 0.0752911 0.00065538 0.0759419 0.851832 101.889 0.246826 0.706852 4.11071 0.0531742 0.0387802 0.96122 0.0198894 0.00422935 0.0191516 0.00407296 0.00511058 0.0058484 0.204423 0.233936 57.9601 -87.8938 125.832 15.9882 145.007 0.000145766 0.267063 192.944 0.310756 0.0673943 0.00409448 0.000561497 0.00138224 0.986996 0.991737 -2.97026e-06 -85.6694 0.0929703 31198.7 300.178 0.983524 0.319147 0.756163 0.756158 9.99958 2.97994e-06 1.19196e-05 0.130502 0.975417 0.928514 -0.0132935 4.89063e-06 0.500288 -1.85953e-20 6.84115e-24 -1.85885e-20 0.00139495 0.997819 8.59167e-05 0.152529 2.85158 0.00139495 0.998053 0.656252 0.0010416 0.00187943 0.000859167 0.455684 0.00187943 0.433837 0.00012696 1.02 0.887285 0.534791 0.285505 1.7159e-07 3.05351e-09 2394.33 3216.48 -0.0622499 0.482109 0.277679 0.259585 -0.592205 -0.169483 0.4768 -0.268684 -0.20812 1.242 1 2.00968e-270 290.885 1.17514e-267 2.01035 1.24 0.000299984 0.897758 0.630006 0.545926 0.396926 2.01066 127.14 82.765 18.6535 60.308 0.00407346 0 -40 10
0.341 9.88747e-09 2.53882e-06 0.0603357 0.0603255 0.0120455 4.4943e-06 0.00115401 0.0754196 0.000655391 0.0760704 0.851868 101.889 0.246822 0.7069 4.11075 0.0531779 0.0387807 0.961219 0.0198894 0.0042294 0.0191515 0.004073 0.00511064 0.00584846 0.204425 0.233938 57.9602 -87.8938 125.834 15.9882 145.007 0.000145747 0.267064 192.944 0.310756 0.0673943 0.00409449 0.000561497 0.00138224 0.986996 0.991737 -2.97027e-06 -85.6694 0.0929703 31198.7 300.179 0.983524 0.319147 0.756062 0.756058 9.99958 2.97994e-06 1.19196e-05 0.130502 0.975442 0.928526 -0.0132935 4.89065e-06 0.50029 -1.85963e-20 6.84152e-24 -1.85894e-20 0.00139495 0.997819 8.59167e-05 0.152529 2.85158 0.00139495 0.998052 0.656372 0.00104162 0.00187943 0.000859167 0.455684 0.00187943 0.433847 0.000126964 1.02 0.887286 0.534791 0.285506 1.7159e-07 3.05352e-09 2394.31 3216.05 -0.0622187 0.482109 0.277678 0.259558 -0.59221 -0.169483 0.476893 -0.268682 -0.208214 1.243 1 1.21893e-270 290.916 7.12906e-268 2.01056 1.241 0.000299983 0.897566 0.630074 0.545353 0.396963 2.01087 127.152 82.7699 18.6538 60.3104 0.00407325 0 -40 10
0.342 9.91645e-09 2.53882e-06 0.0604384 0.0604283 0.0120455 4.50748e-06 0.00115401 0.075548 0.000655401 0.0761988 0.851904 101.889 0.246818 0.706947 4.1108 0.0531817 0.0387811 0.961219 0.0198893 0.00422945 0.0191515 0.00407304 0.0051107 0.00584852 0.204428 0.233941 57.9603 -87.8938 125.836 15.9882 145.007 0.000145728 0.267064 192.944 0.310756 0.0673943 0.00409449 0.000561497 0.00138224 0.986995 0.991737 -2.97028e-06 -85.6694 0.0929704 31198.6 300.181 0.983524 0.319147 0.755962 0.755958 9.99958 2.97994e-06 1.19197e-05 0.130503 0.975468 0.928539 -0.0132935 4.89066e-06 0.500292 -1.85972e-20 6.84188e-24 -1.85903e-20 0.00139495 0.997819 8.59167e-05 0.15253 2.85158 0.00139495 0.99805 0.656491 0.00104164 0.00187943 0.000859167 0.455684 0.00187943 0.433858 0.000126967 1.02 0.887286 0.534791 0.285507 1.7159e-07 3.05353e-09 2394.3 3215.63 -0.0621877 0.482109 0.277678 0.259532 -0.592215 -0.169483 0.476985 -0.268681 -0.208308 1.244 1 7.3932e-271 290.946 4.32491e-268 2.01078 1.242 0.000299983 0.897374 0.630141 0.544781 0.396999 2.01109 127.163 82.7748 18.6541 60.3127 0.00407305 0 -40 10
0.343 9.94543e-09 2.53882e-06 0.060541 0.060531 0.0120455 4.52065e-06 0.00115401 0.0756763 0.000655411 0.0763271 0.85194 101.889 0.246815 0.706995 4.11085 0.0531855 0.0387816 0.961218 0.0198892 0.0042295 0.0191514 0.00407308 0.00511076 0.00584857 0.20443 0.233943 57.9603 -87.8938 125.838 15.9881 145.007 0.000145708 0.267064 192.943 0.310756 0.0673943 0.00409449 0.000561497 0.00138224 0.986995 0.991737 -2.97028e-06 -85.6694 0.0929704 31198.6 300.182 0.983524 0.319147 0.755862 0.755858 9.99958 2.97994e-06 1.19197e-05 0.130503 0.975493 0.928552 -0.0132935 4.89068e-06 0.500294 -1.85981e-20 6.84224e-24 -1.85913e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.998049 0.656611 0.00104166 0.00187943 0.000859168 0.455684 0.00187943 0.433868 0.000126971 1.02 0.887287 0.534791 0.285508 1.7159e-07 3.05354e-09 2394.28 3215.2 -0.0621567 0.482109 0.277678 0.259505 -0.59222 -0.169483 0.477077 -0.268679 -0.208401 1.245 1 4.4842e-271 290.976 2.62374e-268 2.01099 1.243 0.000299983 0.897183 0.630209 0.544211 0.397036 2.01131 127.175 82.7796 18.6544 60.3151 0.00407284 0 -40 10
0.344 9.97441e-09 2.53882e-06 0.0606436 0.0606336 0.0120455 4.53382e-06 0.00115401 0.0758044 0.000655421 0.0764553 0.851976 101.889 0.246811 0.707042 4.11089 0.0531893 0.038782 0.961218 0.0198892 0.00422955 0.0191514 0.00407312 0.00511082 0.00584863 0.204433 0.233945 57.9604 -87.8938 125.839 15.9881 145.007 0.000145689 0.267064 192.943 0.310756 0.0673943 0.00409449 0.000561497 0.00138224 0.986995 0.991737 -2.97029e-06 -85.6694 0.0929704 31198.6 300.183 0.983524 0.319147 0.755763 0.755759 9.99958 2.97994e-06 1.19197e-05 0.130504 0.975518 0.928564 -0.0132935 4.89069e-06 0.500296 -1.8599e-20 6.84261e-24 -1.85922e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.998047 0.656731 0.00104167 0.00187943 0.000859168 0.455684 0.00187943 0.433878 0.000126974 1.02 0.887287 0.534791 0.285508 1.7159e-07 3.05356e-09 2394.26 3214.78 -0.0621259 0.482109 0.277677 0.259479 -0.592225 -0.169483 0.477168 -0.268678 -0.208494 1.246 1 2.71981e-271 291.006 1.59171e-268 2.01121 1.244 0.000299983 0.896992 0.630276 0.543643 0.397073 2.01152 127.186 82.7844 18.6547 60.3174 0.00407264 0 -40 10
0.345 1.00034e-08 2.53882e-06 0.060746 0.0607361 0.0120454 4.54699e-06 0.00115401 0.0759325 0.000655431 0.0765834 0.852012 101.889 0.246807 0.70709 4.11094 0.053193 0.0387825 0.961218 0.0198891 0.0042296 0.0191513 0.00407316 0.00511088 0.00584869 0.204435 0.233948 57.9604 -87.8938 125.841 15.9881 145.007 0.00014567 0.267064 192.943 0.310756 0.0673943 0.00409449 0.000561498 0.00138224 0.986995 0.991737 -2.9703e-06 -85.6694 0.0929705 31198.6 300.185 0.983524 0.319147 0.755664 0.755659 9.99958 2.97995e-06 1.19197e-05 0.130504 0.975543 0.928577 -0.0132935 4.89071e-06 0.500298 -1.86e-20 6.84297e-24 -1.85931e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.998046 0.65685 0.00104169 0.00187943 0.000859168 0.455684 0.00187943 0.433889 0.000126978 1.02 0.887288 0.53479 0.285509 1.7159e-07 3.05357e-09 2394.25 3214.36 -0.0620952 0.482109 0.277677 0.259452 -0.59223 -0.169483 0.47726 -0.268676 -0.208587 1.247 1 1.64965e-271 291.035 9.65626e-269 2.01143 1.245 0.000299983 0.896802 0.630344 0.543076 0.39711 2.01174 127.198 82.7892 18.6549 60.3198 0.00407244 0 -40 10
0.346 1.00324e-08 2.53882e-06 0.0608484 0.0608385 0.0120454 4.56017e-06 0.00115401 0.0760605 0.000655441 0.0767114 0.852048 101.889 0.246803 0.707138 4.11099 0.0531968 0.0387829 0.961217 0.0198891 0.00422965 0.0191512 0.00407321 0.00511094 0.00584875 0.204438 0.23395 57.9605 -87.8938 125.843 15.988 145.007 0.000145651 0.267064 192.943 0.310756 0.0673942 0.00409449 0.000561498 0.00138224 0.986995 0.991737 -2.9703e-06 -85.6694 0.0929705 31198.6 300.186 0.983524 0.319147 0.755565 0.755561 9.99958 2.97995e-06 1.19197e-05 0.130505 0.975568 0.928589 -0.0132935 4.89073e-06 0.5003 -1.86009e-20 6.84333e-24 -1.8594e-20 0.00139495 0.997819 8.59168e-05 0.15253 2.85158 0.00139495 0.998044 0.65697 0.00104171 0.00187943 0.000859168 0.455684 0.00187943 0.433899 0.000126981 1.02 0.887289 0.53479 0.28551 1.7159e-07 3.05358e-09 2394.23 3213.94 -0.0620646 0.482109 0.277677 0.259426 -0.592234 -0.169483 0.47735 -0.268675 -0.208679 1.248 1 1.00056e-271 291.065 5.85805e-269 2.01164 1.246 0.000299983 0.896613 0.630411 0.542511 0.397146 2.01195 127.21 82.794 18.6552 60.3221 0.00407224 0 -40 10
0.347 1.00613e-08 2.53882e-06 0.0609507 0.0609408 0.0120454 4.57334e-06 0.00115401 0.0761884 0.000655451 0.0768392 0.852084 101.889 0.246799 0.707186 4.11104 0.0532007 0.0387834 0.961217 0.019889 0.0042297 0.0191512 0.00407325 0.005111 0.00584882 0.20444 0.233953 57.9606 -87.8939 125.845 15.988 145.007 0.000145632 0.267064 192.943 0.310755 0.0673942 0.00409449 0.000561498 0.00138224 0.986995 0.991737 -2.97031e-06 -85.6694 0.0929705 31198.6 300.187 0.983524 0.319147 0.755467 0.755462 9.99958 2.97995e-06 1.19197e-05 0.130505 0.975593 0.928602 -0.0132935 4.89074e-06 0.500302 -1.86018e-20 6.8437e-24 -1.8595e-20 0.00139495 0.997819 8.59169e-05 0.15253 2.85158 0.00139495 0.998043 0.657089 0.00104172 0.00187943 0.000859169 0.455684 0.00187943 0.43391 0.000126985 1.02 0.887289 0.53479 0.285511 1.7159e-07 3.05359e-09 2394.22 3213.52 -0.0620341 0.482109 0.277676 0.2594 -0.592239 -0.169483 0.477441 -0.268673 -0.208771 1.249 1 6.06871e-272 291.095 3.55383e-269 2.01186 1.247 0.000299983 0.896424 0.630479 0.541948 0.397183 2.01217 127.221 82.7988 18.6555 60.3244 0.00407203 0 -40 10
0.348 1.00903e-08 2.53882e-06 0.0610529 0.0610431 0.0120454 4.58651e-06 0.00115401 0.0763162 0.00065546 0.076967 0.85212 101.889 0.246796 0.707235 4.11109 0.0532045 0.0387838 0.961216 0.0198889 0.00422975 0.0191511 0.00407329 0.00511107 0.00584888 0.204443 0.233955 57.9606 -87.8939 125.846 15.9879 145.007 0.000145613 0.267064 192.943 0.310755 0.0673942 0.00409449 0.000561499 0.00138225 0.986995 0.991737 -2.97032e-06 -85.6694 0.0929706 31198.6 300.189 0.983524 0.319147 0.755368 0.755364 9.99958 2.97995e-06 1.19197e-05 0.130506 0.975618 0.928614 -0.0132935 4.89076e-06 0.500304 -1.86027e-20 6.84406e-24 -1.85959e-20 0.00139495 0.997819 8.59169e-05 0.15253 2.85158 0.00139495 0.998041 0.657209 0.00104174 0.00187943 0.000859169 0.455684 0.00187943 0.43392 0.000126988 1.02 0.88729 0.53479 0.285512 1.7159e-07 3.0536e-09 2394.2 3213.1 -0.0620037 0.482109 0.277676 0.259374 -0.592244 -0.169483 0.477531 -0.268672 -0.208863 1.25 1 3.68086e-272 291.124 2.15595e-269 2.01207 1.248 0.000299983 0.896236 0.630546 0.541386 0.39722 2.01238 127.233 82.8036 18.6558 60.3267 0.00407183 0 -40 10
0.349 1.01193e-08 2.53882e-06 0.0611551 0.0611453 0.0120454 4.59968e-06 0.00115401 0.0764438 0.00065547 0.0770947 0.852156 101.889 0.246792 0.707283 4.11114 0.0532083 0.0387843 0.961216 0.0198889 0.0042298 0.0191511 0.00407333 0.00511113 0.00584894 0.204445 0.233957 57.9607 -87.8939 125.848 15.9879 145.007 0.000145594 0.267064 192.943 0.310755 0.0673942 0.00409449 0.000561499 0.00138225 0.986995 0.991737 -2.97032e-06 -85.6694 0.0929706 31198.6 300.19 0.983524 0.319147 0.755271 0.755266 9.99958 2.97995e-06 1.19197e-05 0.130506 0.975642 0.928627 -0.0132935 4.89078e-06 0.500306 -1.86036e-20 6.84442e-24 -1.85968e-20 0.00139495 0.997819 8.59169e-05 0.15253 2.85158 0.00139495 0.99804 0.657328 0.00104176 0.00187943 0.000859169 0.455684 0.00187943 0.43393 0.000126992 1.02 0.88729 0.53479 0.285513 1.71591e-07 3.05362e-09 2394.18 3212.68 -0.0619734 0.482109 0.277676 0.259348 -0.592249 -0.169483 0.477621 -0.26867 -0.208954 1.251 1 2.23255e-272 291.154 1.30792e-269 2.01229 1.249 0.000299983 0.896049 0.630613 0.540826 0.397256 2.0126 127.244 82.8083 18.6561 60.329 0.00407163 0 -40 10
0.35 1.01483e-08 2.53882e-06 0.0612571 0.0612474 0.0120454 4.61285e-06 0.00115401 0.0765714 0.00065548 0.0772223 0.852193 101.889 0.246788 0.707332 4.11118 0.0532122 0.0387848 0.961215 0.0198888 0.00422985 0.019151 0.00407337 0.00511119 0.005849 0.204448 0.23396 57.9607 -87.8939 125.85 15.9879 145.007 0.000145576 0.267064 192.943 0.310755 0.0673942 0.0040945 0.000561499 0.00138225 0.986995 0.991737 -2.97033e-06 -85.6694 0.0929706 31198.6 300.192 0.983524 0.319147 0.755173 0.755169 9.99958 2.97996e-06 1.19197e-05 0.130507 0.975667 0.928639 -0.0132935 4.8908e-06 0.500308 -1.86046e-20 6.84478e-24 -1.85977e-20 0.00139495 0.997819 8.5917e-05 0.15253 2.85158 0.00139495 0.998038 0.657448 0.00104178 0.00187943 0.00085917 0.455684 0.00187943 0.433941 0.000126995 1.02 0.887291 0.53479 0.285514 1.71591e-07 3.05363e-09 2394.17 3212.27 -0.0619432 0.482109 0.277676 0.259322 -0.592254 -0.169484 0.477711 -0.268669 -0.209045 1.252 1 1.35411e-272 291.183 7.93461e-270 2.0125 1.25 0.000299983 0.895862 0.630681 0.540267 0.397293 2.01281 127.255 82.813 18.6563 60.3313 0.00407143 0 -40 10
0.351 1.01773e-08 2.53882e-06 0.0613591 0.0613494 0.0120454 4.62603e-06 0.00115401 0.0766989 0.00065549 0.0773498 0.852229 101.889 0.246784 0.70738 4.11123 0.053216 0.0387852 0.961215 0.0198887 0.00422991 0.0191509 0.00407341 0.00511125 0.00584906 0.20445 0.233962 57.9608 -87.8939 125.852 15.9878 145.007 0.000145557 0.267064 192.943 0.310755 0.0673941 0.0040945 0.000561499 0.00138225 0.986995 0.991737 -2.97034e-06 -85.6694 0.0929707 31198.6 300.193 0.983524 0.319147 0.755076 0.755072 9.99958 2.97996e-06 1.19197e-05 0.130508 0.975692 0.928651 -0.0132935 4.89081e-06 0.50031 -1.86055e-20 6.84514e-24 -1.85986e-20 0.00139495 0.997819 8.5917e-05 0.15253 2.85158 0.00139495 0.998037 0.657567 0.00104179 0.00187943 0.00085917 0.455684 0.00187943 0.433951 0.000126999 1.02 0.887292 0.534789 0.285514 1.71591e-07 3.05364e-09 2394.15 3211.85 -0.0619131 0.482109 0.277675 0.259296 -0.592259 -0.169484 0.4778 -0.268667 -0.209136 1.253 1 8.2131e-273 291.212 4.81358e-270 2.01272 1.251 0.000299983 0.895676 0.630748 0.53971 0.397329 2.01302 127.267 82.8177 18.6566 60.3336 0.00407124 0 -40 10
0.352 1.02062e-08 2.53882e-06 0.061461 0.0614513 0.0120454 4.6392e-06 0.00115401 0.0768263 0.000655499 0.0774772 0.852266 101.889 0.24678 0.707429 4.11128 0.0532199 0.0387857 0.961214 0.0198887 0.00422996 0.0191509 0.00407346 0.00511132 0.00584912 0.204453 0.233965 57.9609 -87.8939 125.853 15.9878 145.007 0.000145538 0.267064 192.943 0.310755 0.0673941 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97034e-06 -85.6694 0.0929707 31198.6 300.194 0.983524 0.319147 0.754979 0.754975 9.99958 2.97996e-06 1.19197e-05 0.130508 0.975716 0.928663 -0.0132935 4.89083e-06 0.500312 -1.86064e-20 6.8455e-24 -1.85995e-20 0.00139495 0.997819 8.5917e-05 0.15253 2.85158 0.00139495 0.998036 0.657686 0.00104181 0.00187943 0.00085917 0.455683 0.00187943 0.433961 0.000127002 1.02 0.887292 0.534789 0.285515 1.71591e-07 3.05365e-09 2394.13 3211.44 -0.0618832 0.482109 0.277675 0.25927 -0.592263 -0.169484 0.477889 -0.268666 -0.209227 1.254 1 4.9815e-273 291.241 2.92019e-270 2.01293 1.252 0.000299982 0.89549 0.630815 0.539154 0.397366 2.01324 127.278 82.8224 18.6569 60.3358 0.00407104 0 -40 10
0.353 1.02352e-08 2.53882e-06 0.0615628 0.0615532 0.0120453 4.65237e-06 0.00115401 0.0769535 0.000655509 0.0776044 0.852302 101.889 0.246776 0.707478 4.11133 0.0532238 0.0387862 0.961214 0.0198886 0.00423001 0.0191508 0.0040735 0.00511138 0.00584919 0.204455 0.233967 57.9609 -87.8939 125.855 15.9878 145.007 0.00014552 0.267064 192.943 0.310754 0.0673941 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97035e-06 -85.6693 0.0929707 31198.5 300.196 0.983524 0.319147 0.754883 0.754878 9.99958 2.97996e-06 1.19197e-05 0.130509 0.97574 0.928676 -0.0132935 4.89085e-06 0.500315 -1.86073e-20 6.84587e-24 -1.86005e-20 0.00139495 0.997819 8.59171e-05 0.15253 2.85158 0.00139495 0.998034 0.657806 0.00104183 0.00187944 0.000859171 0.455683 0.00187943 0.433972 0.000127006 1.02 0.887293 0.534789 0.285516 1.71591e-07 3.05366e-09 2394.12 3211.03 -0.0618533 0.482109 0.277675 0.259245 -0.592268 -0.169484 0.477977 -0.268664 -0.209317 1.255 1 3.02143e-273 291.27 1.77155e-270 2.01315 1.253 0.000299982 0.895306 0.630882 0.5386 0.397402 2.01345 127.29 82.8271 18.6572 60.3381 0.00407084 0 -40 10
0.354 1.02642e-08 2.53882e-06 0.0616646 0.061655 0.0120453 4.66554e-06 0.00115401 0.0770807 0.000655519 0.0777316 0.852339 101.889 0.246772 0.707527 4.11138 0.0532277 0.0387866 0.961213 0.0198886 0.00423006 0.0191508 0.00407354 0.00511145 0.00584925 0.204458 0.23397 57.961 -87.8939 125.857 15.9877 145.007 0.000145501 0.267064 192.943 0.310754 0.0673941 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97036e-06 -85.6693 0.0929708 31198.5 300.197 0.983524 0.319147 0.754787 0.754782 9.99958 2.97996e-06 1.19197e-05 0.130509 0.975765 0.928688 -0.0132935 4.89086e-06 0.500317 -1.86082e-20 6.84623e-24 -1.86014e-20 0.00139495 0.997819 8.59171e-05 0.15253 2.85158 0.00139495 0.998033 0.657925 0.00104184 0.00187944 0.000859171 0.455683 0.00187944 0.433982 0.000127009 1.02 0.887294 0.534789 0.285517 1.71591e-07 3.05368e-09 2394.1 3210.62 -0.0618236 0.482109 0.277674 0.259219 -0.592273 -0.169484 0.478066 -0.268663 -0.209407 1.256 1 1.83259e-273 291.299 1.07472e-270 2.01336 1.254 0.000299982 0.895122 0.630949 0.538048 0.397439 2.01367 127.301 82.8318 18.6574 60.3404 0.00407064 0 -40 10
0.355 1.02932e-08 2.53882e-06 0.0617662 0.0617567 0.0120453 4.67871e-06 0.00115401 0.0772078 0.000655528 0.0778587 0.852376 101.889 0.246768 0.707576 4.11143 0.0532316 0.0387871 0.961213 0.0198885 0.00423011 0.0191507 0.00407359 0.00511151 0.00584931 0.20446 0.233972 57.9611 -87.8939 125.858 15.9877 145.007 0.000145483 0.267065 192.943 0.310754 0.067394 0.0040945 0.0005615 0.00138225 0.986995 0.991737 -2.97036e-06 -85.6693 0.0929708 31198.5 300.199 0.983524 0.319147 0.754691 0.754686 9.99958 2.97997e-06 1.19198e-05 0.13051 0.975789 0.9287 -0.0132935 4.89088e-06 0.500319 -1.86091e-20 6.84659e-24 -1.86023e-20 0.00139495 0.997819 8.59171e-05 0.15253 2.85158 0.00139495 0.998031 0.658044 0.00104186 0.00187944 0.000859171 0.455683 0.00187944 0.433992 0.000127013 1.02 0.887294 0.534789 0.285518 1.71591e-07 3.05369e-09 2394.09 3210.21 -0.0617939 0.482109 0.277674 0.259194 -0.592278 -0.169484 0.478154 -0.268661 -0.209496 1.257 1 1.11152e-273 291.328 6.51984e-271 2.01357 1.255 0.000299982 0.894938 0.631016 0.537497 0.397475 2.01388 127.313 82.8364 18.6577 60.3426 0.00407045 0 -40 10
0.356 1.03221e-08 2.53882e-06 0.0618678 0.0618583 0.0120453 4.69188e-06 0.00115401 0.0773347 0.000655538 0.0779856 0.852413 101.889 0.246765 0.707626 4.11148 0.0532355 0.0387876 0.961212 0.0198884 0.00423017 0.0191506 0.00407363 0.00511157 0.00584937 0.204463 0.233975 57.9611 -87.8939 125.86 15.9877 145.007 0.000145464 0.267065 192.943 0.310754 0.067394 0.0040945 0.000561501 0.00138225 0.986995 0.991737 -2.97037e-06 -85.6693 0.0929709 31198.5 300.2 0.983524 0.319147 0.754595 0.754591 9.99958 2.97997e-06 1.19198e-05 0.13051 0.975813 0.928712 -0.0132935 4.8909e-06 0.500321 -1.861e-20 6.84695e-24 -1.86032e-20 0.00139495 0.997819 8.59172e-05 0.15253 2.85158 0.00139495 0.99803 0.658163 0.00104188 0.00187944 0.000859172 0.455683 0.00187944 0.434003 0.000127016 1.02 0.887295 0.534789 0.285519 1.71591e-07 3.0537e-09 2394.07 3209.81 -0.0617644 0.482109 0.277674 0.259168 -0.592282 -0.169484 0.478241 -0.26866 -0.209585 1.258 1 6.74172e-274 291.357 3.95529e-271 2.01379 1.256 0.000299982 0.894755 0.631082 0.536948 0.397512 2.01409 127.324 82.8411 18.658 60.3449 0.00407025 0 -40 10
0.357 1.03511e-08 2.53882e-06 0.0619693 0.0619598 0.0120453 4.70506e-06 0.00115401 0.0774616 0.000655547 0.0781125 0.85245 101.888 0.246761 0.707675 4.11153 0.0532394 0.0387881 0.961212 0.0198884 0.00423022 0.0191506 0.00407367 0.00511164 0.00584944 0.204466 0.233978 57.9612 -87.8939 125.862 15.9876 145.007 0.000145446 0.267065 192.943 0.310754 0.067394 0.0040945 0.000561501 0.00138225 0.986995 0.991737 -2.97038e-06 -85.6693 0.0929709 31198.5 300.202 0.983524 0.319147 0.7545 0.754496 9.99958 2.97997e-06 1.19198e-05 0.130511 0.975837 0.928724 -0.0132935 4.89092e-06 0.500323 -1.86109e-20 6.84731e-24 -1.86041e-20 0.00139496 0.997819 8.59172e-05 0.15253 2.85158 0.00139496 0.998029 0.658282 0.0010419 0.00187944 0.000859172 0.455683 0.00187944 0.434013 0.00012702 1.02 0.887296 0.534788 0.28552 1.71591e-07 3.05372e-09 2394.05 3209.4 -0.061735 0.482109 0.277674 0.259143 -0.592287 -0.169484 0.478329 -0.268658 -0.209674 1.259 1 4.08906e-274 291.386 2.39949e-271 2.014 1.257 0.000299982 0.894573 0.631149 0.5364 0.397548 2.01431 127.336 82.8457 18.6582 60.3471 0.00407006 0 -40 10
0.358 1.03801e-08 2.53882e-06 0.0620707 0.0620612 0.0120453 4.71823e-06 0.00115401 0.0775883 0.000655557 0.0782393 0.852487 101.888 0.246757 0.707725 4.11159 0.0532433 0.0387885 0.961211 0.0198883 0.00423027 0.0191505 0.00407372 0.0051117 0.0058495 0.204468 0.23398 57.9612 -87.8939 125.863 15.9876 145.007 0.000145428 0.267065 192.943 0.310753 0.067394 0.00409451 0.000561501 0.00138225 0.986995 0.991737 -2.97038e-06 -85.6693 0.0929709 31198.5 300.203 0.983524 0.319147 0.754405 0.754401 9.99958 2.97997e-06 1.19198e-05 0.130511 0.975861 0.928736 -0.0132935 4.89093e-06 0.500325 -1.86119e-20 6.84767e-24 -1.8605e-20 0.00139496 0.997819 8.59172e-05 0.152531 2.85158 0.00139496 0.998027 0.658401 0.00104191 0.00187944 0.000859172 0.455683 0.00187944 0.434023 0.000127023 1.02 0.887296 0.534788 0.285521 1.71592e-07 3.05373e-09 2394.04 3209 -0.0617056 0.482109 0.277673 0.259118 -0.592292 -0.169484 0.478416 -0.268657 -0.209763 1.26 1 2.48014e-274 291.414 1.45566e-271 2.01421 1.258 0.000299982 0.894391 0.631216 0.535853 0.397584 2.01452 127.347 82.8503 18.6585 60.3493 0.00406986 0 -40 10
0.359 1.04091e-08 2.53882e-06 0.062172 0.0621626 0.0120453 4.7314e-06 0.00115401 0.077715 0.000655566 0.0783659 0.852524 101.888 0.246753 0.707775 4.11164 0.0532473 0.038789 0.961211 0.0198882 0.00423033 0.0191504 0.00407376 0.00511177 0.00584957 0.204471 0.233983 57.9613 -87.8939 125.865 15.9875 145.007 0.000145409 0.267065 192.942 0.310753 0.067394 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.97039e-06 -85.6693 0.092971 31198.5 300.204 0.983524 0.319147 0.754311 0.754306 9.99958 2.97997e-06 1.19198e-05 0.130512 0.975885 0.928748 -0.0132935 4.89095e-06 0.500328 -1.86128e-20 6.84803e-24 -1.86059e-20 0.00139496 0.997819 8.59173e-05 0.152531 2.85158 0.00139496 0.998026 0.65852 0.00104193 0.00187944 0.000859173 0.455683 0.00187944 0.434034 0.000127027 1.02 0.887297 0.534788 0.285522 1.71592e-07 3.05374e-09 2394.02 3208.6 -0.0616764 0.482109 0.277673 0.259093 -0.592296 -0.169484 0.478502 -0.268655 -0.209851 1.261 1 1.50428e-274 291.443 8.83084e-272 2.01443 1.259 0.000299982 0.89421 0.631282 0.535309 0.39762 2.01473 127.358 82.8549 18.6588 60.3516 0.00406967 0 -40 10
0.36 1.04381e-08 2.53882e-06 0.0622732 0.0622639 0.0120452 4.74457e-06 0.00115401 0.0778415 0.000655575 0.0784925 0.852561 101.888 0.246749 0.707825 4.11169 0.0532512 0.0387895 0.96121 0.0198882 0.00423038 0.0191504 0.0040738 0.00511184 0.00584963 0.204473 0.233985 57.9614 -87.8939 125.867 15.9875 145.007 0.000145391 0.267065 192.942 0.310753 0.0673939 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.9704e-06 -85.6693 0.092971 31198.5 300.206 0.983524 0.319147 0.754217 0.754212 9.99958 2.97998e-06 1.19198e-05 0.130512 0.975909 0.92876 -0.0132935 4.89097e-06 0.50033 -1.86137e-20 6.84838e-24 -1.86068e-20 0.00139496 0.997819 8.59173e-05 0.152531 2.85158 0.00139496 0.998025 0.658639 0.00104195 0.00187944 0.000859173 0.455683 0.00187944 0.434044 0.00012703 1.02 0.887298 0.534788 0.285522 1.71592e-07 3.05375e-09 2394 3208.2 -0.0616473 0.482109 0.277673 0.259067 -0.592301 -0.169484 0.478589 -0.268654 -0.209939 1.262 1 9.12393e-275 291.471 5.35726e-272 2.01464 1.26 0.000299982 0.89403 0.631349 0.534765 0.397657 2.01494 127.37 82.8594 18.6591 60.3538 0.00406948 0 -40 10
0.361 1.0467e-08 2.53882e-06 0.0623744 0.0623651 0.0120452 4.75774e-06 0.00115401 0.077968 0.000655585 0.078619 0.852598 101.888 0.246745 0.707875 4.11174 0.0532552 0.03879 0.96121 0.0198881 0.00423043 0.0191503 0.00407385 0.0051119 0.0058497 0.204476 0.233988 57.9614 -87.8939 125.868 15.9875 145.007 0.000145373 0.267065 192.942 0.310753 0.0673939 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.97041e-06 -85.6693 0.092971 31198.5 300.207 0.983524 0.319147 0.754123 0.754118 9.99958 2.97998e-06 1.19198e-05 0.130513 0.975933 0.928772 -0.0132935 4.89099e-06 0.500332 -1.86146e-20 6.84874e-24 -1.86077e-20 0.00139496 0.997819 8.59173e-05 0.152531 2.85158 0.00139496 0.998023 0.658758 0.00104197 0.00187944 0.000859173 0.455683 0.00187944 0.434054 0.000127034 1.02 0.887298 0.534788 0.285523 1.71592e-07 3.05377e-09 2393.99 3207.8 -0.0616183 0.482109 0.277672 0.259042 -0.592306 -0.169484 0.478675 -0.268652 -0.210027 1.263 1 5.53394e-275 291.499 3.25e-272 2.01485 1.261 0.000299982 0.89385 0.631416 0.534224 0.397693 2.01516 127.381 82.864 18.6593 60.356 0.00406929 0 -40 10
0.362 1.0496e-08 2.53882e-06 0.0624755 0.0624662 0.0120452 4.77091e-06 0.00115401 0.0780943 0.000655594 0.0787453 0.852636 101.888 0.246741 0.707925 4.11179 0.0532592 0.0387905 0.96121 0.019888 0.00423049 0.0191502 0.00407389 0.00511197 0.00584976 0.204479 0.23399 57.9615 -87.8939 125.87 15.9874 145.007 0.000145355 0.267065 192.942 0.310753 0.0673939 0.00409451 0.000561502 0.00138226 0.986995 0.991737 -2.97041e-06 -85.6693 0.0929711 31198.5 300.209 0.983524 0.319147 0.754029 0.754025 9.99958 2.97998e-06 1.19198e-05 0.130513 0.975957 0.928784 -0.0132935 4.89101e-06 0.500334 -1.86155e-20 6.8491e-24 -1.86086e-20 0.00139496 0.997819 8.59174e-05 0.152531 2.85158 0.00139496 0.998022 0.658877 0.00104198 0.00187944 0.000859174 0.455682 0.00187944 0.434065 0.000127037 1.02 0.887299 0.534787 0.285524 1.71592e-07 3.05378e-09 2393.97 3207.4 -0.0615894 0.482109 0.277672 0.259018 -0.59231 -0.169484 0.478761 -0.268651 -0.210114 1.264 1 3.35651e-275 291.527 1.97162e-272 2.01506 1.262 0.000299981 0.893671 0.631482 0.533684 0.397729 2.01537 127.392 82.8685 18.6596 60.3582 0.0040691 0 -40 10
0.363 1.0525e-08 2.53882e-06 0.0625765 0.0625673 0.0120452 4.78409e-06 0.00115401 0.0782206 0.000655603 0.0788716 0.852673 101.888 0.246737 0.707975 4.11184 0.0532632 0.038791 0.961209 0.019888 0.00423054 0.0191502 0.00407394 0.00511204 0.00584983 0.204481 0.233993 57.9615 -87.8939 125.872 15.9874 145.007 0.000145337 0.267065 192.942 0.310753 0.0673939 0.00409451 0.000561503 0.00138226 0.986995 0.991737 -2.97042e-06 -85.6693 0.0929711 31198.5 300.21 0.983524 0.319147 0.753936 0.753932 9.99958 2.97998e-06 1.19198e-05 0.130514 0.975981 0.928795 -0.0132935 4.89102e-06 0.500337 -1.86164e-20 6.84946e-24 -1.86095e-20 0.00139496 0.997819 8.59174e-05 0.152531 2.85158 0.00139496 0.998021 0.658996 0.001042 0.00187944 0.000859174 0.455682 0.00187944 0.434075 0.000127041 1.02 0.8873 0.534787 0.285525 1.71592e-07 3.05379e-09 2393.95 3207 -0.0615605 0.482109 0.277672 0.258993 -0.592315 -0.169484 0.478846 -0.268649 -0.210201 1.265 1 2.03582e-275 291.555 1.19609e-272 2.01528 1.263 0.000299981 0.893493 0.631548 0.533145 0.397765 2.01558 127.404 82.8731 18.6599 60.3604 0.00406891 0 -40 10
0.364 1.0554e-08 2.53882e-06 0.0626774 0.0626682 0.0120452 4.79726e-06 0.00115401 0.0783467 0.000655612 0.0789978 0.85271 101.888 0.246733 0.708026 4.1119 0.0532672 0.0387915 0.961209 0.0198879 0.0042306 0.0191501 0.00407398 0.0051121 0.00584989 0.204484 0.233996 57.9616 -87.8939 125.873 15.9874 145.007 0.000145319 0.267065 192.942 0.310752 0.0673938 0.00409451 0.000561503 0.00138226 0.986995 0.991737 -2.97043e-06 -85.6693 0.0929712 31198.4 300.212 0.983524 0.319147 0.753843 0.753839 9.99958 2.97998e-06 1.19198e-05 0.130515 0.976004 0.928807 -0.0132935 4.89104e-06 0.500339 -1.86173e-20 6.84982e-24 -1.86104e-20 0.00139496 0.997819 8.59174e-05 0.152531 2.85158 0.00139496 0.998019 0.659115 0.00104202 0.00187944 0.000859174 0.455682 0.00187944 0.434085 0.000127044 1.02 0.8873 0.534787 0.285526 1.71592e-07 3.05381e-09 2393.94 3206.61 -0.0615318 0.482109 0.277671 0.258968 -0.59232 -0.169484 0.478931 -0.268648 -0.210288 1.266 1 1.23479e-275 291.583 7.25612e-273 2.01549 1.264 0.000299981 0.893315 0.631615 0.532608 0.397801 2.01579 127.415 82.8776 18.6601 60.3626 0.00406872 0 -40 10
0.365 1.05829e-08 2.53882e-06 0.0627782 0.0627691 0.0120452 4.81043e-06 0.00115401 0.0784728 0.000655622 0.0791238 0.852748 101.888 0.246729 0.708076 4.11195 0.0532712 0.038792 0.961208 0.0198878 0.00423065 0.01915 0.00407403 0.00511217 0.00584996 0.204487 0.233998 57.9617 -87.8939 125.875 15.9873 145.007 0.000145301 0.267065 192.942 0.310752 0.0673938 0.00409451 0.000561503 0.00138226 0.986995 0.991737 -2.97043e-06 -85.6693 0.0929712 31198.4 300.213 0.983524 0.319147 0.753751 0.753746 9.99958 2.97999e-06 1.19198e-05 0.130515 0.976028 0.928819 -0.0132935 4.89106e-06 0.500341 -1.86182e-20 6.85018e-24 -1.86113e-20 0.00139496 0.997819 8.59175e-05 0.152531 2.85158 0.00139496 0.998018 0.659233 0.00104204 0.00187944 0.000859175 0.455682 0.00187944 0.434095 0.000127048 1.02 0.887301 0.534787 0.285527 1.71592e-07 3.05382e-09 2393.92 3206.21 -0.0615032 0.482109 0.277671 0.258943 -0.592324 -0.169485 0.479016 -0.268646 -0.210374 1.267 1 7.48938e-276 291.611 4.40194e-273 2.0157 1.265 0.000299981 0.893138 0.631681 0.532072 0.397837 2.016 127.426 82.8821 18.6604 60.3647 0.00406853 0 -40 10
0.366 1.06119e-08 2.53882e-06 0.062879 0.0628699 0.0120452 4.8236e-06 0.00115401 0.0785987 0.000655631 0.0792498 0.852786 101.888 0.246725 0.708127 4.112 0.0532752 0.0387925 0.961208 0.0198878 0.00423071 0.01915 0.00407407 0.00511224 0.00585002 0.20449 0.234001 57.9617 -87.8939 125.877 15.9873 145.008 0.000145284 0.267065 192.942 0.310752 0.0673938 0.00409452 0.000561504 0.00138226 0.986995 0.991737 -2.97044e-06 -85.6693 0.0929712 31198.4 300.215 0.983524 0.319147 0.753658 0.753654 9.99958 2.97999e-06 1.19198e-05 0.130516 0.976051 0.92883 -0.0132935 4.89108e-06 0.500343 -1.86191e-20 6.85053e-24 -1.86122e-20 0.00139496 0.997819 8.59175e-05 0.152531 2.85159 0.00139496 0.998017 0.659352 0.00104205 0.00187944 0.000859175 0.455682 0.00187944 0.434106 0.000127051 1.02 0.887302 0.534787 0.285528 1.71592e-07 3.05383e-09 2393.91 3205.82 -0.0614747 0.482109 0.277671 0.258919 -0.592329 -0.169485 0.479101 -0.268645 -0.21046 1.268 1 4.54254e-276 291.639 2.67045e-273 2.01591 1.266 0.000299981 0.892961 0.631747 0.531538 0.397873 2.01621 127.438 82.8865 18.6606 60.3669 0.00406834 0 -40 10
0.367 1.06409e-08 2.53882e-06 0.0629797 0.0629706 0.0120452 4.83677e-06 0.00115401 0.0787246 0.00065564 0.0793756 0.852823 101.888 0.246721 0.708178 4.11206 0.0532792 0.038793 0.961207 0.0198877 0.00423076 0.0191499 0.00407412 0.00511231 0.00585009 0.204492 0.234004 57.9618 -87.8939 125.878 15.9873 145.008 0.000145266 0.267066 192.942 0.310752 0.0673938 0.00409452 0.000561504 0.00138226 0.986995 0.991737 -2.97045e-06 -85.6693 0.0929713 31198.4 300.216 0.983524 0.319147 0.753566 0.753562 9.99958 2.97999e-06 1.19199e-05 0.130516 0.976075 0.928842 -0.0132935 4.8911e-06 0.500346 -1.862e-20 6.85089e-24 -1.86131e-20 0.00139496 0.997819 8.59176e-05 0.152531 2.85159 0.00139496 0.998015 0.659471 0.00104207 0.00187944 0.000859176 0.455682 0.00187944 0.434116 0.000127055 1.02 0.887302 0.534786 0.285529 1.71593e-07 3.05385e-09 2393.89 3205.43 -0.0614463 0.482109 0.277671 0.258894 -0.592333 -0.169485 0.479185 -0.268643 -0.210546 1.269 1 2.75519e-276 291.667 1.62003e-273 2.01612 1.267 0.000299981 0.892785 0.631813 0.531005 0.397909 2.01643 127.449 82.891 18.6609 60.3691 0.00406815 0 -40 10
0.368 1.06699e-08 2.53882e-06 0.0630803 0.0630712 0.0120451 4.84994e-06 0.00115401 0.0788503 0.000655649 0.0795014 0.852861 101.888 0.246717 0.708229 4.11211 0.0532833 0.0387935 0.961207 0.0198876 0.00423082 0.0191498 0.00407416 0.00511237 0.00585016 0.204495 0.234006 57.9618 -87.8939 125.88 15.9872 145.008 0.000145248 0.267066 192.942 0.310752 0.0673937 0.00409452 0.000561504 0.00138226 0.986995 0.991737 -2.97046e-06 -85.6693 0.0929713 31198.4 300.218 0.983524 0.319147 0.753475 0.75347 9.99958 2.97999e-06 1.19199e-05 0.130517 0.976098 0.928854 -0.0132935 4.89111e-06 0.500348 -1.86209e-20 6.85125e-24 -1.8614e-20 0.00139496 0.997819 8.59176e-05 0.152531 2.85159 0.00139496 0.998014 0.659589 0.00104209 0.00187945 0.000859176 0.455682 0.00187944 0.434126 0.000127058 1.02 0.887303 0.534786 0.28553 1.71593e-07 3.05386e-09 2393.87 3205.04 -0.061418 0.482109 0.27767 0.25887 -0.592338 -0.169485 0.479269 -0.268641 -0.210632 1.27 1 1.67111e-276 291.694 9.82795e-274 2.01633 1.268 0.000299981 0.89261 0.631879 0.530474 0.397945 2.01664 127.46 82.8955 18.6612 60.3712 0.00406796 0 -40 10
0.369 1.06988e-08 2.53882e-06 0.0631808 0.0631718 0.0120451 4.86311e-06 0.00115401 0.078976 0.000655658 0.079627 0.852899 101.888 0.246713 0.70828 4.11216 0.0532873 0.038794 0.961206 0.0198876 0.00423087 0.0191498 0.00407421 0.00511244 0.00585022 0.204498 0.234009 57.9619 -87.8939 125.882 15.9872 145.008 0.000145231 0.267066 192.942 0.310751 0.0673937 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97047e-06 -85.6693 0.0929714 31198.4 300.219 0.983524 0.319147 0.753383 0.753379 9.99958 2.98e-06 1.19199e-05 0.130517 0.976121 0.928865 -0.0132935 4.89113e-06 0.50035 -1.86218e-20 6.8516e-24 -1.86149e-20 0.00139496 0.997819 8.59176e-05 0.152531 2.85159 0.00139496 0.998013 0.659708 0.00104211 0.00187945 0.000859176 0.455682 0.00187945 0.434136 0.000127062 1.02 0.887304 0.534786 0.285531 1.71593e-07 3.05387e-09 2393.86 3204.65 -0.0613898 0.482109 0.27767 0.258846 -0.592342 -0.169485 0.479353 -0.26864 -0.210717 1.271 1 1.01358e-276 291.722 5.96214e-274 2.01654 1.269 0.000299981 0.892435 0.631945 0.529944 0.397981 2.01685 127.472 82.8999 18.6614 60.3734 0.00406778 0 -40 10
0.37 1.07278e-08 2.53882e-06 0.0632812 0.0632723 0.0120451 4.87628e-06 0.00115401 0.0791015 0.000655667 0.0797526 0.852937 101.888 0.246709 0.708332 4.11222 0.0532914 0.0387945 0.961205 0.0198875 0.00423093 0.0191497 0.00407426 0.00511251 0.00585029 0.2045 0.234012 57.962 -87.8939 125.883 15.9871 145.008 0.000145213 0.267066 192.942 0.310751 0.0673937 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97047e-06 -85.6693 0.0929714 31198.4 300.221 0.983524 0.319147 0.753292 0.753288 9.99958 2.98e-06 1.19199e-05 0.130518 0.976144 0.928877 -0.0132935 4.89115e-06 0.500352 -1.86227e-20 6.85196e-24 -1.86158e-20 0.00139496 0.997819 8.59177e-05 0.152531 2.85159 0.00139496 0.998011 0.659827 0.00104213 0.00187945 0.000859177 0.455682 0.00187945 0.434147 0.000127065 1.02 0.887304 0.534786 0.285532 1.71593e-07 3.05389e-09 2393.84 3204.26 -0.0613617 0.48211 0.27767 0.258821 -0.592347 -0.169485 0.479436 -0.268638 -0.210802 1.272 1 6.14766e-277 291.749 3.61694e-274 2.01676 1.27 0.000299981 0.892261 0.632011 0.529416 0.398017 2.01706 127.483 82.9043 18.6617 60.3755 0.00406759 0 -40 10
0.371 1.07568e-08 2.53882e-06 0.0633816 0.0633727 0.0120451 4.88946e-06 0.00115401 0.079227 0.000655676 0.079878 0.852975 101.888 0.246705 0.708383 4.11227 0.0532955 0.038795 0.961205 0.0198874 0.00423099 0.0191496 0.0040743 0.00511258 0.00585036 0.204503 0.234014 57.962 -87.8939 125.885 15.9871 145.008 0.000145196 0.267066 192.942 0.310751 0.0673937 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97048e-06 -85.6693 0.0929714 31198.4 300.222 0.983524 0.319147 0.753202 0.753197 9.99958 2.98e-06 1.19199e-05 0.130519 0.976167 0.928888 -0.0132935 4.89117e-06 0.500355 -1.86236e-20 6.85232e-24 -1.86167e-20 0.00139496 0.997819 8.59177e-05 0.152531 2.85159 0.00139496 0.99801 0.659945 0.00104214 0.00187945 0.000859177 0.455682 0.00187945 0.434157 0.000127069 1.02 0.887305 0.534786 0.285533 1.71593e-07 3.0539e-09 2393.82 3203.87 -0.0613337 0.48211 0.277669 0.258797 -0.592351 -0.169485 0.479519 -0.268637 -0.210887 1.273 1 3.72874e-277 291.776 2.19422e-274 2.01697 1.271 0.00029998 0.892087 0.632077 0.528889 0.398053 2.01727 127.494 82.9087 18.6619 60.3777 0.0040674 0 -40 10
0.372 1.07858e-08 2.53882e-06 0.0634818 0.063473 0.0120451 4.90263e-06 0.00115401 0.0793523 0.000655685 0.0800034 0.853013 101.888 0.2467 0.708435 4.11233 0.0532996 0.0387955 0.961204 0.0198873 0.00423104 0.0191496 0.00407435 0.00511265 0.00585043 0.204506 0.234017 57.9621 -87.8939 125.886 15.9871 145.008 0.000145178 0.267066 192.941 0.310751 0.0673936 0.00409452 0.000561505 0.00138227 0.986995 0.991737 -2.97049e-06 -85.6693 0.0929715 31198.4 300.224 0.983524 0.319147 0.753111 0.753107 9.99958 2.98e-06 1.19199e-05 0.130519 0.97619 0.9289 -0.0132935 4.89119e-06 0.500357 -1.86245e-20 6.85267e-24 -1.86176e-20 0.00139496 0.997819 8.59177e-05 0.152531 2.85159 0.00139496 0.998009 0.660064 0.00104216 0.00187945 0.000859177 0.455681 0.00187945 0.434167 0.000127073 1.02 0.887306 0.534786 0.285534 1.71593e-07 3.05391e-09 2393.81 3203.49 -0.0613058 0.48211 0.277669 0.258773 -0.592356 -0.169485 0.479602 -0.268635 -0.210971 1.274 1 2.2616e-277 291.804 1.33112e-274 2.01718 1.272 0.00029998 0.891914 0.632143 0.528364 0.398088 2.01748 127.505 82.9131 18.6622 60.3798 0.00406722 0 -40 10
0.373 1.08148e-08 2.53882e-06 0.063582 0.0635732 0.0120451 4.9158e-06 0.00115401 0.0794775 0.000655694 0.0801286 0.853052 101.888 0.246696 0.708486 4.11238 0.0533037 0.0387961 0.961204 0.0198873 0.0042311 0.0191495 0.0040744 0.00511272 0.0058505 0.204509 0.23402 57.9622 -87.8939 125.888 15.987 145.008 0.000145161 0.267066 192.941 0.310751 0.0673936 0.00409453 0.000561506 0.00138227 0.986995 0.991737 -2.9705e-06 -85.6693 0.0929715 31198.3 300.225 0.983524 0.319147 0.753021 0.753017 9.99958 2.98001e-06 1.19199e-05 0.13052 0.976213 0.928911 -0.0132935 4.89121e-06 0.500359 -1.86254e-20 6.85303e-24 -1.86185e-20 0.00139496 0.997819 8.59178e-05 0.152532 2.85159 0.00139496 0.998008 0.660182 0.00104218 0.00187945 0.000859178 0.455681 0.00187945 0.434177 0.000127076 1.02 0.887306 0.534785 0.285535 1.71593e-07 3.05393e-09 2393.79 3203.11 -0.0612781 0.48211 0.277669 0.258749 -0.59236 -0.169485 0.479684 -0.268634 -0.211055 1.275 1 1.37173e-277 291.831 8.07527e-275 2.01739 1.273 0.00029998 0.891742 0.632209 0.52784 0.398124 2.01769 127.517 82.9175 18.6625 60.3819 0.00406704 0 -40 10
0.374 1.08437e-08 2.53882e-06 0.0636821 0.0636733 0.0120451 4.92897e-06 0.00115401 0.0796027 0.000655702 0.0802538 0.85309 101.888 0.246692 0.708538 4.11244 0.0533078 0.0387966 0.961203 0.0198872 0.00423116 0.0191494 0.00407444 0.00511279 0.00585057 0.204512 0.234023 57.9622 -87.894 125.89 15.987 145.008 0.000145143 0.267066 192.941 0.31075 0.0673936 0.00409453 0.000561506 0.00138227 0.986995 0.991737 -2.9705e-06 -85.6693 0.0929716 31198.3 300.227 0.983524 0.319147 0.752932 0.752927 9.99958 2.98001e-06 1.19199e-05 0.13052 0.976236 0.928922 -0.0132935 4.89123e-06 0.500362 -1.86263e-20 6.85339e-24 -1.86194e-20 0.00139496 0.997819 8.59178e-05 0.152532 2.85159 0.00139496 0.998006 0.6603 0.0010422 0.00187945 0.000859178 0.455681 0.00187945 0.434188 0.00012708 1.02 0.887307 0.534785 0.285536 1.71593e-07 3.05394e-09 2393.78 3202.72 -0.0612504 0.48211 0.277668 0.258725 -0.592365 -0.169485 0.479766 -0.268632 -0.211139 1.276 1 8.31995e-278 291.858 4.89886e-275 2.0176 1.274 0.00029998 0.89157 0.632275 0.527318 0.39816 2.0179 127.528 82.9218 18.6627 60.384 0.00406685 0 -40 10
0.375 1.08727e-08 2.53882e-06 0.0637822 0.0637734 0.012045 4.94214e-06 0.00115401 0.0797277 0.000655711 0.0803788 0.853128 101.888 0.246688 0.70859 4.11249 0.0533119 0.0387971 0.961203 0.0198871 0.00423121 0.0191494 0.00407449 0.00511286 0.00585064 0.204514 0.234025 57.9623 -87.894 125.891 15.987 145.008 0.000145126 0.267066 192.941 0.31075 0.0673936 0.00409453 0.000561506 0.00138227 0.986995 0.991737 -2.97051e-06 -85.6693 0.0929716 31198.3 300.228 0.983524 0.319147 0.752842 0.752838 9.99958 2.98001e-06 1.19199e-05 0.130521 0.976259 0.928934 -0.0132935 4.89125e-06 0.500364 -1.86272e-20 6.85374e-24 -1.86203e-20 0.00139496 0.997819 8.59179e-05 0.152532 2.85159 0.00139496 0.998005 0.660419 0.00104221 0.00187945 0.000859179 0.455681 0.00187945 0.434198 0.000127083 1.02 0.887308 0.534785 0.285537 1.71594e-07 3.05395e-09 2393.76 3202.34 -0.0612228 0.48211 0.277668 0.258702 -0.592369 -0.169485 0.479848 -0.268631 -0.211222 1.277 1 5.0463e-278 291.885 2.97189e-275 2.01781 1.275 0.00029998 0.891399 0.63234 0.526797 0.398196 2.01811 127.539 82.9262 18.663 60.3861 0.00406667 0 -40 10
0.376 1.09017e-08 2.53882e-06 0.0638821 0.0638734 0.012045 4.95531e-06 0.00115401 0.0798527 0.00065572 0.0805038 0.853167 101.887 0.246684 0.708642 4.11255 0.053316 0.0387976 0.961202 0.0198871 0.00423127 0.0191493 0.00407454 0.00511293 0.0058507 0.204517 0.234028 57.9623 -87.894 125.893 15.9869 145.008 0.000145109 0.267066 192.941 0.31075 0.0673935 0.00409453 0.000561507 0.00138227 0.986995 0.991737 -2.97052e-06 -85.6693 0.0929716 31198.3 300.23 0.983524 0.319147 0.752753 0.752748 9.99958 2.98001e-06 1.19199e-05 0.130521 0.976282 0.928945 -0.0132935 4.89126e-06 0.500367 -1.86281e-20 6.8541e-24 -1.86212e-20 0.00139497 0.997819 8.59179e-05 0.152532 2.85159 0.00139497 0.998004 0.660537 0.00104223 0.00187945 0.000859179 0.455681 0.00187945 0.434208 0.000127087 1.02 0.887308 0.534785 0.285538 1.71594e-07 3.05397e-09 2393.74 3201.96 -0.0611953 0.48211 0.277668 0.258678 -0.592374 -0.169485 0.47993 -0.268629 -0.211305 1.278 1 3.06074e-278 291.912 1.8029e-275 2.01802 1.276 0.00029998 0.891229 0.632406 0.526278 0.398231 2.01832 127.55 82.9305 18.6632 60.3882 0.00406649 0 -40 10
0.377 1.09307e-08 2.53882e-06 0.063982 0.0639733 0.012045 4.96848e-06 0.00115401 0.0799775 0.000655729 0.0806286 0.853205 101.887 0.24668 0.708695 4.1126 0.0533202 0.0387982 0.961202 0.019887 0.00423133 0.0191492 0.00407458 0.005113 0.00585077 0.20452 0.234031 57.9624 -87.894 125.894 15.9869 145.008 0.000145092 0.267066 192.941 0.31075 0.0673935 0.00409453 0.000561507 0.00138227 0.986995 0.991737 -2.97053e-06 -85.6692 0.0929717 31198.3 300.232 0.983524 0.319147 0.752664 0.75266 9.99958 2.98001e-06 1.192e-05 0.130522 0.976304 0.928956 -0.0132935 4.89128e-06 0.500369 -1.8629e-20 6.85445e-24 -1.86221e-20 0.00139497 0.997819 8.59179e-05 0.152532 2.85159 0.00139497 0.998003 0.660655 0.00104225 0.00187945 0.000859179 0.455681 0.00187945 0.434218 0.00012709 1.02 0.887309 0.534785 0.285538 1.71594e-07 3.05398e-09 2393.73 3201.59 -0.0611679 0.48211 0.277668 0.258654 -0.592378 -0.169485 0.480011 -0.268627 -0.211388 1.279 1 1.85643e-278 291.938 1.09373e-275 2.01823 1.277 0.00029998 0.891059 0.632471 0.52576 0.398267 2.01853 127.561 82.9348 18.6635 60.3903 0.00406631 0 -40 10
0.378 1.09596e-08 2.53882e-06 0.0640818 0.0640731 0.012045 4.98165e-06 0.00115401 0.0801022 0.000655737 0.0807534 0.853244 101.887 0.246676 0.708747 4.11266 0.0533243 0.0387987 0.961201 0.0198869 0.00423139 0.0191492 0.00407463 0.00511308 0.00585084 0.204523 0.234034 57.9625 -87.894 125.896 15.9868 145.008 0.000145075 0.267067 192.941 0.310749 0.0673935 0.00409453 0.000561507 0.00138227 0.986995 0.991737 -2.97054e-06 -85.6692 0.0929717 31198.3 300.233 0.983524 0.319147 0.752576 0.752571 9.99958 2.98002e-06 1.192e-05 0.130523 0.976327 0.928967 -0.0132935 4.8913e-06 0.500371 -1.86298e-20 6.85481e-24 -1.8623e-20 0.00139497 0.997819 8.5918e-05 0.152532 2.85159 0.00139497 0.998002 0.660774 0.00104227 0.00187945 0.00085918 0.455681 0.00187945 0.434229 0.000127094 1.02 0.88731 0.534784 0.285539 1.71594e-07 3.054e-09 2393.71 3201.21 -0.0611406 0.48211 0.277667 0.258631 -0.592382 -0.169485 0.480092 -0.268626 -0.211471 1.28 1 1.12598e-278 291.965 6.63508e-276 2.01844 1.278 0.00029998 0.890889 0.632537 0.525243 0.398303 2.01873 127.573 82.9391 18.6637 60.3924 0.00406612 0 -40 10
0.379 1.09886e-08 2.53883e-06 0.0641815 0.0641729 0.012045 4.99482e-06 0.00115401 0.0802269 0.000655746 0.080878 0.853283 101.887 0.246672 0.708799 4.11272 0.0533285 0.0387992 0.961201 0.0198869 0.00423145 0.0191491 0.00407468 0.00511315 0.00585091 0.204526 0.234037 57.9625 -87.894 125.897 15.9868 145.008 0.000145058 0.267067 192.941 0.310749 0.0673935 0.00409454 0.000561508 0.00138228 0.986995 0.991737 -2.97054e-06 -85.6692 0.0929718 31198.3 300.235 0.983524 0.319147 0.752487 0.752483 9.99958 2.98002e-06 1.192e-05 0.130523 0.976349 0.928979 -0.0132935 4.89132e-06 0.500374 -1.86307e-20 6.85516e-24 -1.86239e-20 0.00139497 0.997819 8.5918e-05 0.152532 2.85159 0.00139497 0.998 0.660892 0.00104229 0.00187945 0.00085918 0.455681 0.00187945 0.434239 0.000127097 1.02 0.887311 0.534784 0.28554 1.71594e-07 3.05401e-09 2393.69 3200.83 -0.0611134 0.48211 0.277667 0.258607 -0.592387 -0.169485 0.480172 -0.268624 -0.211553 1.281 1 6.82943e-279 291.992 4.02516e-276 2.01864 1.279 0.00029998 0.890721 0.632602 0.524728 0.398338 2.01894 127.584 82.9434 18.664 60.3945 0.00406594 0 -40 10
0.38 1.10176e-08 2.53883e-06 0.0642811 0.0642726 0.012045 5.00799e-06 0.00115401 0.0803514 0.000655755 0.0810026 0.853321 101.887 0.246667 0.708852 4.11277 0.0533326 0.0387998 0.9612 0.0198868 0.0042315 0.019149 0.00407473 0.00511322 0.00585099 0.204529 0.234039 57.9626 -87.894 125.899 15.9868 145.008 0.000145041 0.267067 192.941 0.310749 0.0673934 0.00409454 0.000561508 0.00138228 0.986995 0.991737 -2.97055e-06 -85.6692 0.0929718 31198.3 300.236 0.983524 0.319147 0.752399 0.752395 9.99958 2.98002e-06 1.192e-05 0.130524 0.976372 0.92899 -0.0132935 4.89134e-06 0.500376 -1.86316e-20 6.85551e-24 -1.86248e-20 0.00139497 0.997819 8.59181e-05 0.152532 2.85159 0.00139497 0.997999 0.66101 0.0010423 0.00187945 0.000859181 0.455681 0.00187945 0.434249 0.000127101 1.02 0.887311 0.534784 0.285541 1.71594e-07 3.05402e-09 2393.68 3200.46 -0.0610863 0.48211 0.277667 0.258584 -0.592391 -0.169486 0.480253 -0.268623 -0.211635 1.282 1 4.14226e-279 292.018 2.44186e-276 2.01885 1.28 0.00029998 0.890552 0.632668 0.524214 0.398374 2.01915 127.595 82.9477 18.6642 60.3965 0.00406576 0 -40 10
0.381 1.10466e-08 2.53883e-06 0.0643807 0.0643721 0.012045 5.02116e-06 0.00115401 0.0804759 0.000655763 0.081127 0.85336 101.887 0.246663 0.708905 4.11283 0.0533368 0.0388003 0.9612 0.0198867 0.00423156 0.0191489 0.00407478 0.00511329 0.00585106 0.204532 0.234042 57.9626 -87.894 125.901 15.9867 145.008 0.000145024 0.267067 192.941 0.310749 0.0673934 0.00409454 0.000561508 0.00138228 0.986995 0.991737 -2.97056e-06 -85.6692 0.0929719 31198.3 300.238 0.983524 0.319147 0.752312 0.752307 9.99958 2.98002e-06 1.192e-05 0.130524 0.976394 0.929001 -0.0132935 4.89136e-06 0.500379 -1.86325e-20 6.85587e-24 -1.86257e-20 0.00139497 0.997819 8.59181e-05 0.152532 2.85159 0.00139497 0.997998 0.661128 0.00104232 0.00187945 0.000859181 0.45568 0.00187945 0.434259 0.000127104 1.02 0.887312 0.534784 0.285542 1.71594e-07 3.05404e-09 2393.66 3200.09 -0.0610593 0.48211 0.277666 0.25856 -0.592395 -0.169486 0.480333 -0.268621 -0.211717 1.283 1 2.51241e-279 292.044 1.48135e-276 2.01906 1.281 0.000299979 0.890385 0.632733 0.523702 0.398409 2.01936 127.606 82.952 18.6645 60.3986 0.00406559 0 -40 10
0.382 1.10755e-08 2.53883e-06 0.0644802 0.0644716 0.012045 5.03433e-06 0.00115401 0.0806002 0.000655772 0.0812514 0.853399 101.887 0.246659 0.708958 4.11289 0.053341 0.0388008 0.961199 0.0198866 0.00423162 0.0191489 0.00407483 0.00511336 0.00585113 0.204535 0.234045 57.9627 -87.894 125.902 15.9867 145.008 0.000145007 0.267067 192.941 0.310749 0.0673934 0.00409454 0.000561509 0.00138228 0.986995 0.991737 -2.97057e-06 -85.6692 0.0929719 31198.2 300.24 0.983524 0.319147 0.752225 0.75222 9.99958 2.98003e-06 1.192e-05 0.130525 0.976417 0.929012 -0.0132935 4.89138e-06 0.500381 -1.86334e-20 6.85622e-24 -1.86265e-20 0.00139497 0.997819 8.59181e-05 0.152532 2.85159 0.00139497 0.997997 0.661246 0.00104234 0.00187946 0.000859181 0.45568 0.00187945 0.434269 0.000127108 1.02 0.887313 0.534784 0.285543 1.71595e-07 3.05405e-09 2393.64 3199.71 -0.0610324 0.48211 0.277666 0.258537 -0.5924 -0.169486 0.480413 -0.268619 -0.211798 1.284 1 1.52385e-279 292.071 8.98657e-277 2.01927 1.282 0.000299979 0.890218 0.632798 0.523191 0.398445 2.01957 127.617 82.9562 18.6647 60.4007 0.00406541 0 -40 10
0.383 1.11045e-08 2.53883e-06 0.0645796 0.0645711 0.0120449 5.04751e-06 0.00115401 0.0807245 0.00065578 0.0813756 0.853438 101.887 0.246655 0.709011 4.11295 0.0533452 0.0388014 0.961199 0.0198866 0.00423168 0.0191488 0.00407488 0.00511344 0.0058512 0.204538 0.234048 57.9628 -87.894 125.904 15.9867 145.008 0.00014499 0.267067 192.941 0.310748 0.0673934 0.00409454 0.000561509 0.00138228 0.986995 0.991737 -2.97058e-06 -85.6692 0.092972 31198.2 300.241 0.983524 0.319147 0.752138 0.752133 9.99958 2.98003e-06 1.192e-05 0.130526 0.976439 0.929023 -0.0132935 4.8914e-06 0.500384 -1.86343e-20 6.85658e-24 -1.86274e-20 0.00139497 0.997819 8.59182e-05 0.152532 2.85159 0.00139497 0.997996 0.661364 0.00104236 0.00187946 0.000859182 0.45568 0.00187946 0.43428 0.000127111 1.02 0.887313 0.534783 0.285544 1.71595e-07 3.05407e-09 2393.63 3199.34 -0.0610055 0.48211 0.277666 0.258514 -0.592404 -0.169486 0.480492 -0.268618 -0.211879 1.285 1 9.24263e-280 292.097 5.45168e-277 2.01948 1.283 0.000299979 0.890052 0.632863 0.522682 0.39848 2.01978 127.628 82.9604 18.665 60.4027 0.00406523 0 -40 10
0.384 1.11335e-08 2.53883e-06 0.0646789 0.0646704 0.0120449 5.06068e-06 0.00115401 0.0808486 0.000655789 0.0814998 0.853477 101.887 0.246651 0.709064 4.113 0.0533494 0.0388019 0.961198 0.0198865 0.00423174 0.0191487 0.00407492 0.00511351 0.00585127 0.20454 0.234051 57.9628 -87.894 125.905 15.9866 145.008 0.000144974 0.267067 192.94 0.310748 0.0673933 0.00409454 0.000561509 0.00138228 0.986995 0.991737 -2.97058e-06 -85.6692 0.092972 31198.2 300.243 0.983524 0.319147 0.752051 0.752046 9.99958 2.98003e-06 1.192e-05 0.130526 0.976461 0.929034 -0.0132935 4.89142e-06 0.500386 -1.86352e-20 6.85693e-24 -1.86283e-20 0.00139497 0.997819 8.59182e-05 0.152532 2.85159 0.00139497 0.997995 0.661482 0.00104237 0.00187946 0.000859182 0.45568 0.00187946 0.43429 0.000127115 1.02 0.887314 0.534783 0.285545 1.71595e-07 3.05408e-09 2393.61 3198.97 -0.0609788 0.48211 0.277666 0.258491 -0.592408 -0.169486 0.480571 -0.268616 -0.21196 1.286 1 5.60594e-280 292.123 3.30725e-277 2.01969 1.284 0.000299979 0.889886 0.632929 0.522174 0.398515 2.01998 127.64 82.9647 18.6652 60.4047 0.00406505 0 -40 10
0.385 1.11625e-08 2.53883e-06 0.0647781 0.0647697 0.0120449 5.07385e-06 0.00115401 0.0809726 0.000655797 0.0816238 0.853516 101.887 0.246646 0.709117 4.11306 0.0533537 0.0388025 0.961198 0.0198864 0.0042318 0.0191487 0.00407497 0.00511358 0.00585134 0.204543 0.234054 57.9629 -87.894 125.907 15.9866 145.008 0.000144957 0.267067 192.94 0.310748 0.0673933 0.00409454 0.00056151 0.00138228 0.986995 0.991737 -2.97059e-06 -85.6692 0.092972 31198.2 300.244 0.983524 0.319147 0.751964 0.75196 9.99958 2.98003e-06 1.192e-05 0.130527 0.976483 0.929045 -0.0132935 4.89144e-06 0.500388 -1.8636e-20 6.85728e-24 -1.86292e-20 0.00139497 0.997819 8.59183e-05 0.152532 2.85159 0.00139497 0.997993 0.6616 0.00104239 0.00187946 0.000859183 0.45568 0.00187946 0.4343 0.000127118 1.02 0.887315 0.534783 0.285546 1.71595e-07 3.05409e-09 2393.6 3198.61 -0.0609522 0.48211 0.277665 0.258468 -0.592413 -0.169486 0.48065 -0.268615 -0.212041 1.287 1 3.40017e-280 292.149 2.00633e-277 2.0199 1.285 0.000299979 0.889721 0.632994 0.521667 0.398551 2.02019 127.651 82.9689 18.6655 60.4068 0.00406488 0 -40 10
0.386 1.11914e-08 2.53883e-06 0.0648773 0.0648689 0.0120449 5.08702e-06 0.00115401 0.0810966 0.000655805 0.0817478 0.853556 101.887 0.246642 0.709171 4.11312 0.0533579 0.038803 0.961197 0.0198863 0.00423186 0.0191486 0.00407502 0.00511366 0.00585142 0.204546 0.234057 57.963 -87.894 125.908 15.9866 145.008 0.00014494 0.267067 192.94 0.310748 0.0673933 0.00409455 0.00056151 0.00138228 0.986995 0.991737 -2.9706e-06 -85.6692 0.0929721 31198.2 300.246 0.983524 0.319147 0.751878 0.751874 9.99958 2.98004e-06 1.192e-05 0.130528 0.976505 0.929056 -0.0132935 4.89146e-06 0.500391 -1.86369e-20 6.85763e-24 -1.86301e-20 0.00139497 0.997819 8.59183e-05 0.152533 2.85159 0.00139497 0.997992 0.661718 0.00104241 0.00187946 0.000859183 0.45568 0.00187946 0.43431 0.000127122 1.02 0.887316 0.534783 0.285547 1.71595e-07 3.05411e-09 2393.58 3198.24 -0.0609257 0.48211 0.277665 0.258445 -0.592417 -0.169486 0.480729 -0.268613 -0.212121 1.288 1 2.06231e-280 292.175 1.21714e-277 2.0201 1.286 0.000299979 0.889556 0.633059 0.521162 0.398586 2.0204 127.662 82.973 18.6657 60.4088 0.0040647 0 -40 10
0.387 1.12204e-08 2.53883e-06 0.0649763 0.064968 0.0120449 5.10019e-06 0.00115401 0.0812204 0.000655814 0.0818716 0.853595 101.887 0.246638 0.709224 4.11318 0.0533622 0.0388036 0.961196 0.0198863 0.00423192 0.0191485 0.00407507 0.00511373 0.00585149 0.204549 0.23406 57.963 -87.894 125.91 15.9865 145.008 0.000144924 0.267067 192.94 0.310747 0.0673932 0.00409455 0.000561511 0.00138228 0.986995 0.991737 -2.97061e-06 -85.6692 0.0929721 31198.2 300.248 0.983524 0.319147 0.751793 0.751788 9.99958 2.98004e-06 1.19201e-05 0.130528 0.976527 0.929067 -0.0132935 4.89148e-06 0.500393 -1.86378e-20 6.85799e-24 -1.8631e-20 0.00139497 0.997819 8.59184e-05 0.152533 2.85159 0.00139497 0.997991 0.661836 0.00104243 0.00187946 0.000859184 0.45568 0.00187946 0.43432 0.000127125 1.02 0.887316 0.534783 0.285548 1.71595e-07 3.05412e-09 2393.56 3197.87 -0.0608993 0.48211 0.277665 0.258422 -0.592421 -0.169486 0.480807 -0.268611 -0.212201 1.289 1 1.25085e-280 292.201 7.38371e-278 2.02031 1.287 0.000299979 0.889392 0.633124 0.520658 0.398621 2.02061 127.673 82.9772 18.666 60.4108 0.00406452 0 -40 10
0.388 1.12494e-08 2.53883e-06 0.0650753 0.065067 0.0120449 5.11336e-06 0.00115401 0.0813442 0.000655822 0.0819954 0.853634 101.887 0.246634 0.709278 4.11324 0.0533664 0.0388041 0.961196 0.0198862 0.00423198 0.0191484 0.00407512 0.00511381 0.00585156 0.204552 0.234063 57.9631 -87.894 125.911 15.9865 145.008 0.000144907 0.267068 192.94 0.310747 0.0673932 0.00409455 0.000561511 0.00138229 0.986995 0.991737 -2.97062e-06 -85.6692 0.0929722 31198.2 300.249 0.983524 0.319147 0.751707 0.751703 9.99958 2.98004e-06 1.19201e-05 0.130529 0.976549 0.929077 -0.0132935 4.8915e-06 0.500396 -1.86387e-20 6.85834e-24 -1.86318e-20 0.00139497 0.997819 8.59184e-05 0.152533 2.8516 0.00139497 0.99799 0.661953 0.00104245 0.00187946 0.000859184 0.45568 0.00187946 0.434331 0.000127129 1.02 0.887317 0.534782 0.285549 1.71595e-07 3.05414e-09 2393.55 3197.51 -0.0608729 0.48211 0.277664 0.258399 -0.592425 -0.169486 0.480885 -0.26861 -0.21228 1.29 1 7.58681e-281 292.226 4.4793e-278 2.02052 1.288 0.000299979 0.889228 0.633189 0.520156 0.398657 2.02081 127.684 82.9814 18.6662 60.4128 0.00406435 0 -40 10
0.389 1.12784e-08 2.53883e-06 0.0651743 0.065166 0.0120449 5.12653e-06 0.00115401 0.0814678 0.00065583 0.082119 0.853674 101.887 0.246629 0.709332 4.1133 0.0533707 0.0388047 0.961195 0.0198861 0.00423204 0.0191484 0.00407517 0.00511388 0.00585164 0.204555 0.234065 57.9631 -87.894 125.913 15.9864 145.008 0.000144891 0.267068 192.94 0.310747 0.0673932 0.00409455 0.000561511 0.00138229 0.986995 0.991737 -2.97063e-06 -85.6692 0.0929722 31198.2 300.251 0.983524 0.319147 0.751622 0.751617 9.99958 2.98005e-06 1.19201e-05 0.130529 0.976571 0.929088 -0.0132935 4.89152e-06 0.500398 -1.86396e-20 6.85869e-24 -1.86327e-20 0.00139497 0.997819 8.59184e-05 0.152533 2.8516 0.00139497 0.997989 0.662071 0.00104246 0.00187946 0.000859184 0.455679 0.00187946 0.434341 0.000127132 1.02 0.887318 0.534782 0.28555 1.71596e-07 3.05415e-09 2393.53 3197.15 -0.0608467 0.48211 0.277664 0.258376 -0.59243 -0.169486 0.480963 -0.268608 -0.21236 1.291 1 4.60163e-281 292.252 2.71735e-278 2.02073 1.289 0.000299979 0.889065 0.633253 0.519655 0.398692 2.02102 127.695 82.9855 18.6664 60.4148 0.00406418 0 -40 10
0.39 1.13073e-08 2.53883e-06 0.0652731 0.0652648 0.0120448 5.1397e-06 0.00115401 0.0815914 0.000655839 0.0822426 0.853713 101.887 0.246625 0.709386 4.11336 0.053375 0.0388052 0.961195 0.019886 0.00423211 0.0191483 0.00407522 0.00511396 0.00585171 0.204558 0.234068 57.9632 -87.894 125.914 15.9864 145.008 0.000144875 0.267068 192.94 0.310747 0.0673932 0.00409455 0.000561512 0.00138229 0.986995 0.991737 -2.97064e-06 -85.6692 0.0929723 31198.2 300.253 0.983524 0.319147 0.751537 0.751532 9.99958 2.98005e-06 1.19201e-05 0.13053 0.976593 0.929099 -0.0132935 4.89154e-06 0.500401 -1.86405e-20 6.85904e-24 -1.86336e-20 0.00139497 0.997819 8.59185e-05 0.152533 2.8516 0.00139497 0.997988 0.662189 0.00104248 0.00187946 0.000859185 0.455679 0.00187946 0.434351 0.000127136 1.02 0.887318 0.534782 0.285551 1.71596e-07 3.05417e-09 2393.51 3196.79 -0.0608206 0.48211 0.277664 0.258354 -0.592434 -0.169486 0.48104 -0.268606 -0.212439 1.292 1 2.79103e-281 292.278 1.64847e-278 2.02093 1.29 0.000299978 0.888903 0.633318 0.519155 0.398727 2.02123 127.706 82.9897 18.6667 60.4168 0.004064 0 -40 10
0.391 1.13363e-08 2.53883e-06 0.0653718 0.0653636 0.0120448 5.15287e-06 0.00115401 0.0817148 0.000655847 0.0823661 0.853753 101.887 0.246621 0.70944 4.11342 0.0533793 0.0388058 0.961194 0.019886 0.00423217 0.0191482 0.00407527 0.00511403 0.00585178 0.204561 0.234071 57.9633 -87.894 125.916 15.9864 145.008 0.000144858 0.267068 192.94 0.310747 0.0673931 0.00409455 0.000561512 0.00138229 0.986995 0.991737 -2.97064e-06 -85.6692 0.0929723 31198.1 300.254 0.983524 0.319147 0.751452 0.751448 9.99958 2.98005e-06 1.19201e-05 0.130531 0.976614 0.92911 -0.0132935 4.89156e-06 0.500404 -1.86413e-20 6.85939e-24 -1.86345e-20 0.00139497 0.997819 8.59185e-05 0.152533 2.8516 0.00139497 0.997987 0.662307 0.0010425 0.00187946 0.000859185 0.455679 0.00187946 0.434361 0.000127139 1.02 0.887319 0.534782 0.285552 1.71596e-07 3.05418e-09 2393.5 3196.43 -0.0607945 0.48211 0.277663 0.258331 -0.592438 -0.169486 0.481118 -0.268605 -0.212518 1.293 1 1.69285e-281 292.303 1.00004e-278 2.02114 1.291 0.000299978 0.888741 0.633383 0.518657 0.398762 2.02143 127.717 82.9938 18.6669 60.4188 0.00406383 0 -40 10
0.392 1.13653e-08 2.53883e-06 0.0654705 0.0654623 0.0120448 5.16604e-06 0.00115401 0.0818382 0.000655855 0.0824894 0.853793 101.887 0.246616 0.709494 4.11348 0.0533836 0.0388064 0.961194 0.0198859 0.00423223 0.0191481 0.00407533 0.00511411 0.00585186 0.204564 0.234074 57.9633 -87.894 125.917 15.9863 145.008 0.000144842 0.267068 192.94 0.310746 0.0673931 0.00409456 0.000561512 0.00138229 0.986995 0.991737 -2.97065e-06 -85.6692 0.0929724 31198.1 300.256 0.983524 0.319147 0.751368 0.751363 9.99958 2.98005e-06 1.19201e-05 0.130531 0.976636 0.92912 -0.0132935 4.89158e-06 0.500406 -1.86422e-20 6.85975e-24 -1.86354e-20 0.00139497 0.997819 8.59186e-05 0.152533 2.8516 0.00139497 0.997986 0.662424 0.00104252 0.00187946 0.000859186 0.455679 0.00187946 0.434371 0.000127143 1.02 0.88732 0.534782 0.285554 1.71596e-07 3.0542e-09 2393.48 3196.07 -0.0607686 0.48211 0.277663 0.258309 -0.592442 -0.169486 0.481195 -0.268603 -0.212596 1.294 1 1.02676e-281 292.329 6.06668e-279 2.02135 1.292 0.000299978 0.88858 0.633448 0.51816 0.398797 2.02164 127.728 82.9979 18.6672 60.4208 0.00406366 0 -40 10
0.393 1.13943e-08 2.53883e-06 0.0655691 0.065561 0.0120448 5.17921e-06 0.00115401 0.0819614 0.000655863 0.0826127 0.853832 101.886 0.246612 0.709549 4.11354 0.0533879 0.0388069 0.961193 0.0198858 0.00423229 0.0191481 0.00407538 0.00511419 0.00585193 0.204567 0.234077 57.9634 -87.894 125.919 15.9863 145.008 0.000144826 0.267068 192.94 0.310746 0.0673931 0.00409456 0.000561513 0.00138229 0.986995 0.991737 -2.97066e-06 -85.6692 0.0929724 31198.1 300.258 0.983524 0.319147 0.751284 0.751279 9.99958 2.98006e-06 1.19201e-05 0.130532 0.976657 0.929131 -0.0132935 4.8916e-06 0.500409 -1.86431e-20 6.8601e-24 -1.86362e-20 0.00139498 0.997819 8.59186e-05 0.152533 2.8516 0.00139498 0.997984 0.662542 0.00104254 0.00187946 0.000859186 0.455679 0.00187946 0.434381 0.000127147 1.02 0.887321 0.534781 0.285555 1.71596e-07 3.05421e-09 2393.46 3195.71 -0.0607427 0.48211 0.277663 0.258286 -0.592446 -0.169486 0.481271 -0.268602 -0.212675 1.295 1 6.22763e-282 292.354 3.68032e-279 2.02155 1.293 0.000299978 0.888419 0.633512 0.517665 0.398833 2.02185 127.739 83.002 18.6674 60.4228 0.00406349 0 -40 10
0.394 1.14232e-08 2.53883e-06 0.0656676 0.0656595 0.0120448 5.19238e-06 0.00115401 0.0820846 0.000655871 0.0827358 0.853872 101.886 0.246608 0.709603 4.1136 0.0533922 0.0388075 0.961192 0.0198857 0.00423235 0.019148 0.00407543 0.00511426 0.00585201 0.204571 0.23408 57.9634 -87.894 125.92 15.9863 145.008 0.00014481 0.267068 192.94 0.310746 0.067393 0.00409456 0.000561513 0.00138229 0.986995 0.991737 -2.97067e-06 -85.6692 0.0929725 31198.1 300.259 0.983524 0.319147 0.7512 0.751196 9.99958 2.98006e-06 1.19201e-05 0.130533 0.976679 0.929142 -0.0132935 4.89162e-06 0.500411 -1.8644e-20 6.86045e-24 -1.86371e-20 0.00139498 0.997819 8.59187e-05 0.152533 2.8516 0.00139498 0.997983 0.662659 0.00104256 0.00187946 0.000859187 0.455679 0.00187946 0.434391 0.00012715 1.02 0.887321 0.534781 0.285556 1.71596e-07 3.05423e-09 2393.45 3195.35 -0.060717 0.48211 0.277663 0.258264 -0.592451 -0.169486 0.481347 -0.2686 -0.212753 1.296 1 3.77725e-282 292.379 2.23265e-279 2.02176 1.294 0.000299978 0.888259 0.633577 0.517171 0.398868 2.02205 127.75 83.006 18.6677 60.4248 0.00406331 0 -40 10
0.395 1.14522e-08 2.53883e-06 0.0657661 0.065758 0.0120448 5.20555e-06 0.00115401 0.0822076 0.00065588 0.0828589 0.853912 101.886 0.246603 0.709658 4.11366 0.0533965 0.0388081 0.961192 0.0198857 0.00423242 0.0191479 0.00407548 0.00511434 0.00585208 0.204574 0.234083 57.9635 -87.894 125.922 15.9862 145.008 0.000144794 0.267068 192.94 0.310746 0.067393 0.00409456 0.000561513 0.00138229 0.986995 0.991737 -2.97068e-06 -85.6692 0.0929725 31198.1 300.261 0.983524 0.319147 0.751117 0.751112 9.99958 2.98006e-06 1.19201e-05 0.130533 0.9767 0.929152 -0.0132935 4.89164e-06 0.500414 -1.86448e-20 6.8608e-24 -1.8638e-20 0.00139498 0.997819 8.59187e-05 0.152533 2.8516 0.00139498 0.997982 0.662777 0.00104257 0.00187947 0.000859187 0.455679 0.00187946 0.434402 0.000127154 1.02 0.887322 0.534781 0.285557 1.71596e-07 3.05424e-09 2393.43 3195 -0.0606913 0.48211 0.277662 0.258242 -0.592455 -0.169487 0.481424 -0.268598 -0.21283 1.297 1 2.29102e-282 292.404 1.35442e-279 2.02197 1.295 0.000299978 0.8881 0.633641 0.516678 0.398903 2.02226 127.761 83.0101 18.6679 60.4267 0.00406314 0 -40 10
0.396 1.14812e-08 2.53883e-06 0.0658645 0.0658564 0.0120448 5.21872e-06 0.00115401 0.0823306 0.000655888 0.0829819 0.853952 101.886 0.246599 0.709713 4.11372 0.0534009 0.0388087 0.961191 0.0198856 0.00423248 0.0191478 0.00407553 0.00511442 0.00585216 0.204577 0.234086 57.9636 -87.894 125.923 15.9862 145.008 0.000144778 0.267068 192.939 0.310745 0.067393 0.00409456 0.000561514 0.00138229 0.986995 0.991737 -2.97069e-06 -85.6692 0.0929726 31198.1 300.263 0.983524 0.319147 0.751033 0.751029 9.99958 2.98006e-06 1.19201e-05 0.130534 0.976722 0.929163 -0.0132935 4.89166e-06 0.500416 -1.86457e-20 6.86115e-24 -1.86389e-20 0.00139498 0.997819 8.59187e-05 0.152533 2.8516 0.00139498 0.997981 0.662894 0.00104259 0.00187947 0.000859187 0.455679 0.00187947 0.434412 0.000127157 1.02 0.887323 0.534781 0.285558 1.71597e-07 3.05426e-09 2393.42 3194.64 -0.0606657 0.482111 0.277662 0.25822 -0.592459 -0.169487 0.481499 -0.268597 -0.212908 1.298 1 1.38957e-282 292.429 8.21654e-280 2.02217 1.296 0.000299978 0.887941 0.633706 0.516187 0.398938 2.02247 127.772 83.0141 18.6681 60.4287 0.00406297 0 -40 10
0.397 1.15102e-08 2.53883e-06 0.0659627 0.0659547 0.0120448 5.23189e-06 0.00115401 0.0824534 0.000655896 0.0831047 0.853992 101.886 0.246595 0.709768 4.11378 0.0534052 0.0388092 0.961191 0.0198855 0.00423254 0.0191478 0.00407558 0.0051145 0.00585224 0.20458 0.234089 57.9636 -87.894 125.925 15.9862 145.008 0.000144762 0.267068 192.939 0.310745 0.067393 0.00409456 0.000561514 0.0013823 0.986995 0.991737 -2.9707e-06 -85.6691 0.0929726 31198.1 300.264 0.983524 0.319147 0.750951 0.750946 9.99958 2.98007e-06 1.19202e-05 0.130534 0.976743 0.929173 -0.0132935 4.89168e-06 0.500419 -1.86466e-20 6.8615e-24 -1.86397e-20 0.00139498 0.997819 8.59188e-05 0.152533 2.8516 0.00139498 0.99798 0.663012 0.00104261 0.00187947 0.000859188 0.455679 0.00187947 0.434422 0.000127161 1.02 0.887324 0.53478 0.285559 1.71597e-07 3.05427e-09 2393.4 3194.29 -0.0606402 0.482111 0.277662 0.258197 -0.592463 -0.169487 0.481575 -0.268595 -0.212985 1.299 1 8.42818e-283 292.454 4.98452e-280 2.02238 1.297 0.000299978 0.887783 0.63377 0.515697 0.398973 2.02267 127.783 83.0182 18.6684 60.4307 0.0040628 0 -40 10
0.398 1.15391e-08 2.53883e-06 0.0660609 0.0660529 0.0120447 5.24506e-06 0.00115401 0.0825762 0.000655904 0.0832275 0.854032 101.886 0.24659 0.709823 4.11384 0.0534096 0.0388098 0.96119 0.0198854 0.00423261 0.0191477 0.00407564 0.00511457 0.00585231 0.204583 0.234093 57.9637 -87.894 125.926 15.9861 145.008 0.000144746 0.267069 192.939 0.310745 0.0673929 0.00409457 0.000561515 0.0013823 0.986995 0.991737 -2.97071e-06 -85.6691 0.0929727 31198.1 300.266 0.983524 0.319147 0.750868 0.750864 9.99958 2.98007e-06 1.19202e-05 0.130535 0.976764 0.929184 -0.0132935 4.8917e-06 0.500422 -1.86475e-20 6.86185e-24 -1.86406e-20 0.00139498 0.997819 8.59188e-05 0.152534 2.8516 0.00139498 0.997979 0.663129 0.00104263 0.00187947 0.000859188 0.455678 0.00187947 0.434432 0.000127164 1.02 0.887324 0.53478 0.28556 1.71597e-07 3.05429e-09 2393.38 3193.94 -0.0606148 0.482111 0.277661 0.258175 -0.592467 -0.169487 0.48165 -0.268593 -0.213062 1.3 1 5.11195e-283 292.479 3.02383e-280 2.02258 1.298 0.000299977 0.887625 0.633835 0.515208 0.399008 2.02288 127.794 83.0222 18.6686 60.4326 0.00406264 0 -40 10
0.399 1.15681e-08 2.53883e-06 0.0661591 0.0661511 0.0120447 5.25823e-06 0.00115401 0.0826988 0.000655912 0.0833501 0.854073 101.886 0.246586 0.709878 4.1139 0.053414 0.0388104 0.96119 0.0198853 0.00423267 0.0191476 0.00407569 0.00511465 0.00585239 0.204586 0.234096 57.9638 -87.894 125.928 15.9861 145.008 0.00014473 0.267069 192.939 0.310745 0.0673929 0.00409457 0.000561515 0.0013823 0.986995 0.991737 -2.97071e-06 -85.6691 0.0929727 31198 300.268 0.983524 0.319147 0.750786 0.750781 9.99958 2.98007e-06 1.19202e-05 0.130536 0.976785 0.929194 -0.0132935 4.89172e-06 0.500424 -1.86483e-20 6.8622e-24 -1.86415e-20 0.00139498 0.997819 8.59189e-05 0.152534 2.8516 0.00139498 0.997978 0.663246 0.00104265 0.00187947 0.000859189 0.455678 0.00187947 0.434442 0.000127168 1.02 0.887325 0.53478 0.285561 1.71597e-07 3.0543e-09 2393.37 3193.59 -0.0605895 0.482111 0.277661 0.258153 -0.592471 -0.169487 0.481725 -0.268592 -0.213139 1.301 1 3.10056e-283 292.504 1.83438e-280 2.02279 1.299 0.000299977 0.887467 0.633899 0.514721 0.399042 2.02308 127.805 83.0262 18.6688 60.4345 0.00406247 0 -40 10
0.4 1.15971e-08 2.53883e-06 0.0662571 0.0662492 0.0120447 5.2714e-06 0.00115401 0.0828214 0.00065592 0.0834727 0.854113 101.886 0.246582 0.709933 4.11397 0.0534183 0.038811 0.961189 0.0198853 0.00423273 0.0191475 0.00407574 0.00511473 0.00585247 0.204589 0.234099 57.9638 -87.8941 125.929 15.986 145.008 0.000144714 0.267069 192.939 0.310744 0.0673929 0.00409457 0.000561515 0.0013823 0.986995 0.991737 -2.97072e-06 -85.6691 0.0929728 31198 300.27 0.983524 0.319147 0.750704 0.750699 9.99958 2.98008e-06 1.19202e-05 0.130536 0.976806 0.929204 -0.0132935 4.89174e-06 0.500427 -1.86492e-20 6.86255e-24 -1.86423e-20 0.00139498 0.997819 8.59189e-05 0.152534 2.8516 0.00139498 0.997977 0.663364 0.00104266 0.00187947 0.000859189 0.455678 0.00187947 0.434452 0.000127171 1.02 0.887326 0.53478 0.285562 1.71597e-07 3.05432e-09 2393.35 3193.24 -0.0605643 0.482111 0.277661 0.258132 -0.592475 -0.169487 0.4818 -0.26859 -0.213215 1.302 1 1.88058e-283 292.529 1.11282e-280 2.02299 1.3 0.000299977 0.887311 0.633963 0.514235 0.399077 2.02329 127.816 83.0302 18.6691 60.4365 0.0040623 0 -40 10
0.401 1.16261e-08 2.53883e-06 0.0663551 0.0663472 0.0120447 5.28457e-06 0.00115401 0.0829439 0.000655928 0.0835952 0.854153 101.886 0.246577 0.709989 4.11403 0.0534227 0.0388116 0.961188 0.0198852 0.0042328 0.0191475 0.00407579 0.00511481 0.00585254 0.204592 0.234102 57.9639 -87.8941 125.931 15.986 145.008 0.000144698 0.267069 192.939 0.310744 0.0673928 0.00409457 0.000561516 0.0013823 0.986995 0.991737 -2.97073e-06 -85.6691 0.0929728 31198 300.271 0.983524 0.319147 0.750622 0.750617 9.99958 2.98008e-06 1.19202e-05 0.130537 0.976827 0.929215 -0.0132935 4.89176e-06 0.50043 -1.86501e-20 6.8629e-24 -1.86432e-20 0.00139498 0.997819 8.5919e-05 0.152534 2.8516 0.00139498 0.997976 0.663481 0.00104268 0.00187947 0.00085919 0.455678 0.00187947 0.434462 0.000127175 1.02 0.887327 0.53478 0.285563 1.71597e-07 3.05433e-09 2393.33 3192.89 -0.0605392 0.482111 0.277661 0.25811 -0.592479 -0.169487 0.481874 -0.268588 -0.213291 1.303 1 1.14063e-283 292.553 6.75083e-281 2.0232 1.301 0.000299977 0.887155 0.634027 0.51375 0.399112 2.02349 127.827 83.0342 18.6693 60.4384 0.00406213 0 -40 10
0.402 1.1655e-08 2.53883e-06 0.066453 0.0664451 0.0120447 5.29774e-06 0.00115401 0.0830662 0.000655935 0.0837176 0.854194 101.886 0.246573 0.710044 4.11409 0.0534271 0.0388122 0.961188 0.0198851 0.00423286 0.0191474 0.00407585 0.00511489 0.00585262 0.204596 0.234105 57.9639 -87.8941 125.932 15.986 145.008 0.000144683 0.267069 192.939 0.310744 0.0673928 0.00409457 0.000561516 0.0013823 0.986995 0.991737 -2.97074e-06 -85.6691 0.0929729 31198 300.273 0.983524 0.319147 0.75054 0.750536 9.99958 2.98008e-06 1.19202e-05 0.130538 0.976848 0.929225 -0.0132935 4.89178e-06 0.500432 -1.86509e-20 6.86325e-24 -1.86441e-20 0.00139498 0.997819 8.5919e-05 0.152534 2.8516 0.00139498 0.997975 0.663598 0.0010427 0.00187947 0.00085919 0.455678 0.00187947 0.434472 0.000127178 1.02 0.887327 0.534779 0.285564 1.71597e-07 3.05435e-09 2393.32 3192.54 -0.0605142 0.482111 0.27766 0.258088 -0.592483 -0.169487 0.481948 -0.268587 -0.213367 1.304 1 6.91827e-284 292.578 4.09534e-281 2.0234 1.302 0.000299977 0.886999 0.634091 0.513267 0.399147 2.0237 127.838 83.0381 18.6695 60.4403 0.00406197 0 -40 10
0.403 1.1684e-08 2.53883e-06 0.0665508 0.066543 0.0120447 5.31091e-06 0.00115401 0.0831885 0.000655943 0.0838398 0.854234 101.886 0.246568 0.7101 4.11415 0.0534316 0.0388128 0.961187 0.019885 0.00423293 0.0191473 0.0040759 0.00511497 0.0058527 0.204599 0.234108 57.964 -87.8941 125.933 15.9859 145.008 0.000144667 0.267069 192.939 0.310744 0.0673928 0.00409457 0.000561516 0.0013823 0.986995 0.991737 -2.97075e-06 -85.6691 0.0929729 31198 300.275 0.983524 0.319147 0.750459 0.750455 9.99958 2.98008e-06 1.19202e-05 0.130538 0.976869 0.929235 -0.0132935 4.8918e-06 0.500435 -1.86518e-20 6.8636e-24 -1.8645e-20 0.00139498 0.997819 8.59191e-05 0.152534 2.8516 0.00139498 0.997974 0.663715 0.00104272 0.00187947 0.000859191 0.455678 0.00187947 0.434482 0.000127182 1.02 0.887328 0.534779 0.285565 1.71598e-07 3.05436e-09 2393.3 3192.2 -0.0604893 0.482111 0.27766 0.258066 -0.592487 -0.169487 0.482022 -0.268585 -0.213442 1.305 1 4.19615e-284 292.602 2.48441e-281 2.02361 1.303 0.000299977 0.886844 0.634156 0.512785 0.399182 2.0239 127.849 83.0421 18.6698 60.4422 0.0040618 0 -40 10
0.404 1.1713e-08 2.53883e-06 0.0666485 0.0666407 0.0120447 5.32408e-06 0.00115401 0.0833107 0.000655951 0.083962 0.854275 101.886 0.246564 0.710156 4.11422 0.053436 0.0388134 0.961187 0.019885 0.00423299 0.0191472 0.00407595 0.00511505 0.00585278 0.204602 0.234111 57.9641 -87.8941 125.935 15.9859 145.008 0.000144651 0.267069 192.939 0.310743 0.0673928 0.00409458 0.000561517 0.0013823 0.986995 0.991737 -2.97076e-06 -85.6691 0.092973 31198 300.277 0.983524 0.319147 0.750378 0.750374 9.99958 2.98009e-06 1.19202e-05 0.130539 0.97689 0.929246 -0.0132935 4.89182e-06 0.500438 -1.86527e-20 6.86395e-24 -1.86458e-20 0.00139498 0.997819 8.59191e-05 0.152534 2.8516 0.00139498 0.997973 0.663833 0.00104274 0.00187947 0.000859191 0.455678 0.00187947 0.434493 0.000127185 1.02 0.887329 0.534779 0.285566 1.71598e-07 3.05438e-09 2393.28 3191.85 -0.0604644 0.482111 0.27766 0.258045 -0.592491 -0.169487 0.482096 -0.268583 -0.213518 1.306 1 2.54509e-284 292.626 1.50715e-281 2.02381 1.304 0.000299977 0.886689 0.63422 0.512304 0.399217 2.02411 127.86 83.046 18.67 60.4441 0.00406164 0 -40 10
0.405 1.17419e-08 2.53883e-06 0.0667462 0.0667384 0.0120446 5.33725e-06 0.00115401 0.0834327 0.000655959 0.0840841 0.854315 101.886 0.24656 0.710212 4.11428 0.0534404 0.038814 0.961186 0.0198849 0.00423306 0.0191471 0.00407601 0.00511513 0.00585286 0.204605 0.234114 57.9641 -87.8941 125.936 15.9859 145.008 0.000144636 0.267069 192.939 0.310743 0.0673927 0.00409458 0.000561517 0.00138231 0.986995 0.991737 -2.97077e-06 -85.6691 0.092973 31198 300.278 0.983524 0.319147 0.750298 0.750293 9.99958 2.98009e-06 1.19203e-05 0.13054 0.976911 0.929256 -0.0132935 4.89184e-06 0.50044 -1.86536e-20 6.8643e-24 -1.86467e-20 0.00139498 0.997819 8.59192e-05 0.152534 2.8516 0.00139498 0.997972 0.66395 0.00104276 0.00187947 0.000859192 0.455677 0.00187947 0.434503 0.000127189 1.02 0.88733 0.534779 0.285567 1.71598e-07 3.05439e-09 2393.27 3191.51 -0.0604397 0.482111 0.277659 0.258023 -0.592495 -0.169487 0.482169 -0.268582 -0.213593 1.307 1 1.54368e-284 292.651 9.143e-282 2.02402 1.305 0.000299977 0.886535 0.634284 0.511825 0.399251 2.02431 127.871 83.05 18.6702 60.446 0.00406147 0 -40 10
0.406 1.17709e-08 2.53883e-06 0.0668438 0.066836 0.0120446 5.35042e-06 0.00115401 0.0835547 0.000655967 0.0842061 0.854356 101.886 0.246555 0.710268 4.11434 0.0534449 0.0388146 0.961185 0.0198848 0.00423312 0.0191471 0.00407606 0.00511521 0.00585294 0.204608 0.234117 57.9642 -87.8941 125.938 15.9858 145.008 0.00014462 0.267069 192.938 0.310743 0.0673927 0.00409458 0.000561518 0.00138231 0.986995 0.991737 -2.97078e-06 -85.6691 0.0929731 31198 300.28 0.983524 0.319147 0.750218 0.750213 9.99958 2.98009e-06 1.19203e-05 0.13054 0.976931 0.929266 -0.0132935 4.89186e-06 0.500443 -1.86544e-20 6.86465e-24 -1.86476e-20 0.00139498 0.997819 8.59192e-05 0.152534 2.8516 0.00139498 0.997971 0.664067 0.00104277 0.00187947 0.000859192 0.455677 0.00187947 0.434513 0.000127192 1.02 0.88733 0.534779 0.285568 1.71598e-07 3.05441e-09 2393.25 3191.17 -0.060415 0.482111 0.277659 0.258002 -0.592499 -0.169487 0.482242 -0.26858 -0.213667 1.308 1 9.36287e-285 292.675 5.54653e-282 2.02422 1.306 0.000299976 0.886382 0.634347 0.511347 0.399286 2.02451 127.882 83.0539 18.6705 60.4479 0.00406131 0 -40 10
0.407 1.17999e-08 2.53883e-06 0.0669413 0.0669335 0.0120446 5.36359e-06 0.00115401 0.0836766 0.000655974 0.0843279 0.854397 101.886 0.246551 0.710324 4.11441 0.0534493 0.0388152 0.961185 0.0198847 0.00423319 0.019147 0.00407612 0.00511529 0.00585302 0.204612 0.234121 57.9642 -87.8941 125.939 15.9858 145.008 0.000144605 0.26707 192.938 0.310743 0.0673927 0.00409458 0.000561518 0.00138231 0.986995 0.991737 -2.97079e-06 -85.6691 0.0929731 31197.9 300.282 0.983524 0.319147 0.750137 0.750133 9.99958 2.9801e-06 1.19203e-05 0.130541 0.976952 0.929276 -0.0132935 4.89188e-06 0.500446 -1.86553e-20 6.86499e-24 -1.86484e-20 0.00139498 0.997819 8.59192e-05 0.152534 2.8516 0.00139498 0.99797 0.664184 0.00104279 0.00187948 0.000859192 0.455677 0.00187947 0.434523 0.000127196 1.02 0.887331 0.534778 0.285569 1.71598e-07 3.05442e-09 2393.24 3190.83 -0.0603905 0.482111 0.277659 0.257981 -0.592503 -0.169487 0.482315 -0.268578 -0.213742 1.309 1 5.67887e-285 292.699 3.36476e-282 2.02443 1.307 0.000299976 0.886229 0.634411 0.510871 0.399321 2.02472 127.893 83.0578 18.6707 60.4498 0.00406114 0 -40 10
0.408 1.18289e-08 2.53883e-06 0.0670387 0.067031 0.0120446 5.37676e-06 0.00115401 0.0837983 0.000655982 0.0844497 0.854438 101.886 0.246546 0.710381 4.11447 0.0534538 0.0388158 0.961184 0.0198846 0.00423325 0.0191469 0.00407617 0.00511537 0.00585309 0.204615 0.234124 57.9643 -87.8941 125.941 15.9857 145.008 0.000144589 0.26707 192.938 0.310742 0.0673926 0.00409458 0.000561518 0.00138231 0.986995 0.991737 -2.9708e-06 -85.6691 0.0929732 31197.9 300.284 0.983524 0.319147 0.750058 0.750053 9.99958 2.9801e-06 1.19203e-05 0.130542 0.976973 0.929286 -0.0132935 4.89191e-06 0.500448 -1.86561e-20 6.86534e-24 -1.86493e-20 0.00139499 0.997819 8.59193e-05 0.152534 2.85161 0.00139499 0.997969 0.664301 0.00104281 0.00187948 0.000859193 0.455677 0.00187948 0.434533 0.0001272 1.02 0.887332 0.534778 0.28557 1.71598e-07 3.05444e-09 2393.22 3190.49 -0.060366 0.482111 0.277658 0.257959 -0.592507 -0.169487 0.482387 -0.268577 -0.213816 1.31 1 3.44441e-285 292.723 2.0412e-282 2.02463 1.308 0.000299976 0.886077 0.634475 0.510395 0.399355 2.02492 127.904 83.0617 18.6709 60.4517 0.00406098 0 -40 10
0.409 1.18578e-08 2.53883e-06 0.067136 0.0671284 0.0120446 5.38992e-06 0.00115401 0.08392 0.00065599 0.0845714 0.854479 101.885 0.246542 0.710437 4.11454 0.0534583 0.0388164 0.961184 0.0198845 0.00423332 0.0191468 0.00407622 0.00511545 0.00585317 0.204618 0.234127 57.9644 -87.8941 125.942 15.9857 145.008 0.000144574 0.26707 192.938 0.310742 0.0673926 0.00409458 0.000561519 0.00138231 0.986995 0.991737 -2.97081e-06 -85.6691 0.0929732 31197.9 300.286 0.983524 0.319147 0.749978 0.749974 9.99958 2.9801e-06 1.19203e-05 0.130542 0.976993 0.929296 -0.0132935 4.89193e-06 0.500451 -1.8657e-20 6.86569e-24 -1.86501e-20 0.00139499 0.997819 8.59193e-05 0.152535 2.85161 0.00139499 0.997968 0.664418 0.00104283 0.00187948 0.000859193 0.455677 0.00187948 0.434543 0.000127203 1.02 0.887333 0.534778 0.285571 1.71599e-07 3.05445e-09 2393.2 3190.15 -0.0603416 0.482111 0.277658 0.257938 -0.592511 -0.169487 0.482459 -0.268575 -0.21389 1.311 1 2.08914e-285 292.747 1.23828e-282 2.02483 1.309 0.000299976 0.885925 0.634539 0.509921 0.39939 2.02512 127.915 83.0655 18.6711 60.4536 0.00406082 0 -40 10
0.41 1.18868e-08 2.53883e-06 0.0672333 0.0672257 0.0120446 5.40309e-06 0.00115401 0.0840416 0.000655997 0.084693 0.85452 101.885 0.246537 0.710494 4.1146 0.0534628 0.038817 0.961183 0.0198845 0.00423339 0.0191467 0.00407628 0.00511553 0.00585326 0.204621 0.23413 57.9644 -87.8941 125.943 15.9857 145.008 0.000144559 0.26707 192.938 0.310742 0.0673926 0.00409459 0.000561519 0.00138231 0.986995 0.991737 -2.97081e-06 -85.6691 0.0929733 31197.9 300.287 0.983524 0.319147 0.749899 0.749895 9.99958 2.9801e-06 1.19203e-05 0.130543 0.977014 0.929306 -0.0132935 4.89195e-06 0.500454 -1.86579e-20 6.86604e-24 -1.8651e-20 0.00139499 0.997819 8.59194e-05 0.152535 2.85161 0.00139499 0.997967 0.664535 0.00104285 0.00187948 0.000859194 0.455677 0.00187948 0.434553 0.000127207 1.02 0.887334 0.534778 0.285572 1.71599e-07 3.05447e-09 2393.19 3189.81 -0.0603173 0.482111 0.277658 0.257917 -0.592515 -0.169488 0.482531 -0.268573 -0.213964 1.312 1 1.26713e-285 292.771 7.5119e-283 2.02504 1.31 0.000299976 0.885774 0.634603 0.509449 0.399424 2.02533 127.926 83.0694 18.6714 60.4554 0.00406066 0 -40 10
0.411 1.19158e-08 2.53883e-06 0.0673305 0.0673229 0.0120446 5.41626e-06 0.00115401 0.0841631 0.000656005 0.0848145 0.854561 101.885 0.246533 0.71055 4.11467 0.0534673 0.0388176 0.961182 0.0198844 0.00423345 0.0191467 0.00407633 0.00511562 0.00585334 0.204625 0.234133 57.9645 -87.8941 125.945 15.9856 145.008 0.000144544 0.26707 192.938 0.310742 0.0673925 0.00409459 0.00056152 0.00138231 0.986995 0.991737 -2.97082e-06 -85.6691 0.0929733 31197.9 300.289 0.983524 0.319147 0.74982 0.749816 9.99958 2.98011e-06 1.19203e-05 0.130544 0.977034 0.929316 -0.0132935 4.89197e-06 0.500457 -1.86587e-20 6.86639e-24 -1.86519e-20 0.00139499 0.997819 8.59194e-05 0.152535 2.85161 0.00139499 0.997966 0.664651 0.00104287 0.00187948 0.000859194 0.455677 0.00187948 0.434563 0.00012721 1.02 0.887334 0.534777 0.285574 1.71599e-07 3.05449e-09 2393.17 3189.47 -0.0602931 0.482111 0.277658 0.257896 -0.592519 -0.169488 0.482603 -0.268572 -0.214037 1.313 1 7.68551e-286 292.795 4.55702e-283 2.02524 1.311 0.000299976 0.885623 0.634666 0.508977 0.399459 2.02553 127.936 83.0732 18.6716 60.4573 0.0040605 0 -40 10
0.412 1.19448e-08 2.53883e-06 0.0674276 0.06742 0.0120446 5.42943e-06 0.00115401 0.0842845 0.000656013 0.0849359 0.854602 101.885 0.246528 0.710607 4.11473 0.0534718 0.0388182 0.961182 0.0198843 0.00423352 0.0191466 0.00407639 0.0051157 0.00585342 0.204628 0.234137 57.9646 -87.8941 125.946 15.9856 145.008 0.000144528 0.26707 192.938 0.310741 0.0673925 0.00409459 0.00056152 0.00138231 0.986995 0.991737 -2.97083e-06 -85.6691 0.0929734 31197.9 300.291 0.983524 0.319147 0.749741 0.749737 9.99958 2.98011e-06 1.19203e-05 0.130544 0.977054 0.929326 -0.0132935 4.89199e-06 0.500459 -1.86596e-20 6.86673e-24 -1.86527e-20 0.00139499 0.997819 8.59195e-05 0.152535 2.85161 0.00139499 0.997965 0.664768 0.00104289 0.00187948 0.000859195 0.455677 0.00187948 0.434573 0.000127214 1.02 0.887335 0.534777 0.285575 1.71599e-07 3.0545e-09 2393.15 3189.14 -0.060269 0.482111 0.277657 0.257875 -0.592523 -0.169488 0.482674 -0.26857 -0.21411 1.314 1 4.6615e-286 292.818 2.76448e-283 2.02544 1.312 0.000299976 0.885473 0.63473 0.508507 0.399494 2.02573 127.947 83.0771 18.6718 60.4592 0.00406033 0 -40 10
0.413 1.19737e-08 2.53883e-06 0.0675246 0.0675171 0.0120445 5.4426e-06 0.00115401 0.0844058 0.00065602 0.0850572 0.854644 101.885 0.246524 0.710664 4.1148 0.0534763 0.0388189 0.961181 0.0198842 0.00423359 0.0191465 0.00407645 0.00511578 0.0058535 0.204631 0.23414 57.9646 -87.8941 125.948 15.9856 145.008 0.000144513 0.26707 192.938 0.310741 0.0673925 0.00409459 0.00056152 0.00138232 0.986995 0.991737 -2.97084e-06 -85.6691 0.0929734 31197.9 300.293 0.983524 0.319147 0.749663 0.749659 9.99958 2.98011e-06 1.19203e-05 0.130545 0.977074 0.929336 -0.0132934 4.89201e-06 0.500462 -1.86605e-20 6.86708e-24 -1.86536e-20 0.00139499 0.997819 8.59195e-05 0.152535 2.85161 0.00139499 0.997964 0.664885 0.0010429 0.00187948 0.000859195 0.455676 0.00187948 0.434583 0.000127217 1.02 0.887336 0.534777 0.285576 1.71599e-07 3.05452e-09 2393.14 3188.81 -0.060245 0.482111 0.277657 0.257854 -0.592527 -0.169488 0.482745 -0.268568 -0.214183 1.315 1 2.82734e-286 292.842 1.67704e-283 2.02565 1.313 0.000299976 0.885323 0.634793 0.508038 0.399528 2.02594 127.958 83.0809 18.672 60.461 0.00406017 0 -40 10
0.414 1.20027e-08 2.53883e-06 0.0676216 0.0676141 0.0120445 5.45577e-06 0.00115401 0.084527 0.000656028 0.0851784 0.854685 101.885 0.246519 0.710721 4.11486 0.0534808 0.0388195 0.961181 0.0198841 0.00423366 0.0191464 0.0040765 0.00511586 0.00585358 0.204635 0.234143 57.9647 -87.8941 125.949 15.9855 145.009 0.000144498 0.26707 192.938 0.310741 0.0673924 0.00409459 0.000561521 0.00138232 0.986995 0.991737 -2.97085e-06 -85.6691 0.0929735 31197.8 300.295 0.983524 0.319147 0.749585 0.749581 9.99958 2.98012e-06 1.19204e-05 0.130546 0.977095 0.929346 -0.0132934 4.89203e-06 0.500465 -1.86613e-20 6.86743e-24 -1.86545e-20 0.00139499 0.997819 8.59196e-05 0.152535 2.85161 0.00139499 0.997963 0.665002 0.00104292 0.00187948 0.000859196 0.455676 0.00187948 0.434593 0.000127221 1.02 0.887337 0.534777 0.285577 1.71599e-07 3.05453e-09 2393.12 3188.47 -0.060221 0.482111 0.277657 0.257833 -0.592531 -0.169488 0.482816 -0.268566 -0.214255 1.316 1 1.71487e-286 292.865 1.01736e-283 2.02585 1.314 0.000299975 0.885174 0.634857 0.507571 0.399562 2.02614 127.969 83.0847 18.6723 60.4629 0.00406002 0 -40 10
0.415 1.20317e-08 2.53883e-06 0.0677184 0.067711 0.0120445 5.46894e-06 0.00115401 0.0846481 0.000656035 0.0852995 0.854726 101.885 0.246515 0.710779 4.11493 0.0534853 0.0388201 0.96118 0.0198841 0.00423372 0.0191463 0.00407656 0.00511595 0.00585366 0.204638 0.234146 57.9647 -87.8941 125.95 15.9855 145.009 0.000144483 0.26707 192.938 0.310741 0.0673924 0.0040946 0.000561521 0.00138232 0.986995 0.991737 -2.97086e-06 -85.6691 0.0929735 31197.8 300.297 0.983524 0.319147 0.749507 0.749503 9.99958 2.98012e-06 1.19204e-05 0.130547 0.977115 0.929356 -0.0132934 4.89205e-06 0.500468 -1.86622e-20 6.86777e-24 -1.86553e-20 0.00139499 0.997819 8.59196e-05 0.152535 2.85161 0.00139499 0.997962 0.665118 0.00104294 0.00187948 0.000859196 0.455676 0.00187948 0.434603 0.000127224 1.02 0.887338 0.534777 0.285578 1.716e-07 3.05455e-09 2393.1 3188.14 -0.0601972 0.482111 0.277656 0.257812 -0.592535 -0.169488 0.482887 -0.268565 -0.214328 1.317 1 1.04012e-286 292.889 6.17172e-284 2.02605 1.315 0.000299975 0.885026 0.63492 0.507104 0.399597 2.02634 127.98 83.0885 18.6725 60.4647 0.00405986 0 -40 10
0.416 1.20606e-08 2.53883e-06 0.0678152 0.0678078 0.0120445 5.48211e-06 0.00115401 0.0847691 0.000656043 0.0854205 0.854768 101.885 0.24651 0.710836 4.115 0.0534899 0.0388207 0.961179 0.019884 0.00423379 0.0191463 0.00407661 0.00511603 0.00585374 0.204641 0.23415 57.9648 -87.8941 125.952 15.9855 145.009 0.000144468 0.267071 192.938 0.31074 0.0673924 0.0040946 0.000561522 0.00138232 0.986995 0.991737 -2.97087e-06 -85.669 0.0929736 31197.8 300.298 0.983523 0.319147 0.74943 0.749425 9.99958 2.98012e-06 1.19204e-05 0.130547 0.977135 0.929366 -0.0132934 4.89208e-06 0.500471 -1.8663e-20 6.86812e-24 -1.86562e-20 0.00139499 0.997819 8.59197e-05 0.152535 2.85161 0.00139499 0.997961 0.665235 0.00104296 0.00187948 0.000859197 0.455676 0.00187948 0.434613 0.000127228 1.02 0.887338 0.534776 0.285579 1.716e-07 3.05456e-09 2393.09 3187.81 -0.0601734 0.482111 0.277656 0.257792 -0.592538 -0.169488 0.482957 -0.268563 -0.2144 1.318 1 6.30865e-287 292.912 3.74401e-284 2.02625 1.316 0.000299975 0.884878 0.634984 0.506639 0.399631 2.02654 127.991 83.0923 18.6727 60.4665 0.0040597 0 -40 10
0.417 1.20896e-08 2.53883e-06 0.067912 0.0679045 0.0120445 5.49528e-06 0.00115401 0.08489 0.00065605 0.0855414 0.854809 101.885 0.246506 0.710894 4.11506 0.0534945 0.0388214 0.961179 0.0198839 0.00423386 0.0191462 0.00407667 0.00511612 0.00585383 0.204645 0.234153 57.9649 -87.8941 125.953 15.9854 145.009 0.000144453 0.267071 192.937 0.31074 0.0673923 0.0040946 0.000561522 0.00138232 0.986995 0.991737 -2.97088e-06 -85.669 0.0929736 31197.8 300.3 0.983523 0.319147 0.749352 0.749348 9.99958 2.98012e-06 1.19204e-05 0.130548 0.977155 0.929376 -0.0132934 4.8921e-06 0.500474 -1.86639e-20 6.86847e-24 -1.8657e-20 0.00139499 0.997819 8.59197e-05 0.152535 2.85161 0.00139499 0.99796 0.665352 0.00104298 0.00187948 0.000859197 0.455676 0.00187948 0.434623 0.000127231 1.02 0.887339 0.534776 0.28558 1.716e-07 3.05458e-09 2393.07 3187.48 -0.0601497 0.482111 0.277656 0.257771 -0.592542 -0.169488 0.483027 -0.268561 -0.214472 1.319 1 3.82639e-287 292.935 2.27126e-284 2.02646 1.317 0.000299975 0.88473 0.635047 0.506176 0.399666 2.02675 128.001 83.096 18.6729 60.4683 0.00405954 0 -40 10
0.418 1.21186e-08 2.53883e-06 0.0680086 0.0680012 0.0120445 5.50845e-06 0.00115401 0.0850108 0.000656058 0.0856622 0.854851 101.885 0.246501 0.710951 4.11513 0.053499 0.038822 0.961178 0.0198838 0.00423393 0.0191461 0.00407673 0.0051162 0.00585391 0.204648 0.234156 57.9649 -87.8941 125.955 15.9854 145.009 0.000144439 0.267071 192.937 0.31074 0.0673923 0.0040946 0.000561522 0.00138232 0.986994 0.991737 -2.97089e-06 -85.669 0.0929737 31197.8 300.302 0.983523 0.319147 0.749275 0.749271 9.99958 2.98013e-06 1.19204e-05 0.130549 0.977175 0.929386 -0.0132934 4.89212e-06 0.500476 -1.86648e-20 6.86881e-24 -1.86579e-20 0.00139499 0.997819 8.59198e-05 0.152535 2.85161 0.00139499 0.997959 0.665468 0.001043 0.00187949 0.000859198 0.455676 0.00187948 0.434633 0.000127235 1.02 0.88734 0.534776 0.285581 1.716e-07 3.0546e-09 2393.05 3187.15 -0.0601261 0.482111 0.277656 0.257751 -0.592546 -0.169488 0.483097 -0.26856 -0.214543 1.32 1 2.32082e-287 292.959 1.37784e-284 2.02666 1.318 0.000299975 0.884583 0.63511 0.505713 0.3997 2.02695 128.012 83.0998 18.6731 60.4702 0.00405938 0 -40 10
0.419 1.21476e-08 2.53883e-06 0.0681052 0.0680978 0.0120445 5.52162e-06 0.00115401 0.0851315 0.000656065 0.0857829 0.854893 101.885 0.246496 0.711009 4.1152 0.0535036 0.0388226 0.961177 0.0198837 0.004234 0.019146 0.00407678 0.00511629 0.00585399 0.204651 0.23416 57.965 -87.8941 125.956 15.9853 145.009 0.000144424 0.267071 192.937 0.31074 0.0673923 0.0040946 0.000561523 0.00138232 0.986994 0.991737 -2.9709e-06 -85.669 0.0929737 31197.8 300.304 0.983523 0.319147 0.749199 0.749194 9.99958 2.98013e-06 1.19204e-05 0.130549 0.977195 0.929395 -0.0132934 4.89214e-06 0.500479 -1.86656e-20 6.86916e-24 -1.86587e-20 0.00139499 0.997819 8.59198e-05 0.152535 2.85161 0.00139499 0.997958 0.665585 0.00104301 0.00187949 0.000859198 0.455676 0.00187949 0.434643 0.000127238 1.02 0.887341 0.534776 0.285582 1.716e-07 3.05461e-09 2393.04 3186.83 -0.0601026 0.482112 0.277655 0.25773 -0.59255 -0.169488 0.483167 -0.268558 -0.214615 1.321 1 1.40765e-287 292.982 8.3585e-285 2.02686 1.319 0.000299975 0.884437 0.635174 0.505252 0.399734 2.02715 128.023 83.1035 18.6734 60.472 0.00405923 0 -40 10
0.42 1.21765e-08 2.53883e-06 0.0682017 0.0681943 0.0120445 5.53479e-06 0.00115401 0.0852521 0.000656072 0.0859036 0.854935 101.885 0.246492 0.711067 4.11527 0.0535082 0.0388233 0.961177 0.0198836 0.00423407 0.0191459 0.00407684 0.00511637 0.00585408 0.204655 0.234163 57.965 -87.8941 125.957 15.9853 145.009 0.000144409 0.267071 192.937 0.310739 0.0673923 0.0040946 0.000561523 0.00138233 0.986994 0.991737 -2.97091e-06 -85.669 0.0929738 31197.8 300.306 0.983523 0.319147 0.749122 0.749118 9.99958 2.98013e-06 1.19204e-05 0.13055 0.977214 0.929405 -0.0132934 4.89216e-06 0.500482 -1.86665e-20 6.86951e-24 -1.86596e-20 0.00139499 0.997819 8.59199e-05 0.152536 2.85161 0.00139499 0.997958 0.665701 0.00104303 0.00187949 0.000859199 0.455675 0.00187949 0.434653 0.000127242 1.02 0.887342 0.534775 0.285583 1.716e-07 3.05463e-09 2393.02 3186.5 -0.0600792 0.482112 0.277655 0.25771 -0.592554 -0.169488 0.483236 -0.268556 -0.214686 1.322 1 8.53783e-288 293.005 5.07059e-285 2.02706 1.32 0.000299975 0.884291 0.635237 0.504792 0.399769 2.02735 128.034 83.1073 18.6736 60.4738 0.00405907 0 -40 10
0.421 1.22055e-08 2.53883e-06 0.0682981 0.0682908 0.0120444 5.54795e-06 0.00115401 0.0853726 0.00065608 0.0860241 0.854977 101.885 0.246487 0.711125 4.11533 0.0535128 0.0388239 0.961176 0.0198835 0.00423414 0.0191458 0.0040769 0.00511646 0.00585416 0.204658 0.234166 57.9651 -87.8941 125.959 15.9853 145.009 0.000144394 0.267071 192.937 0.310739 0.0673922 0.00409461 0.000561524 0.00138233 0.986994 0.991737 -2.97092e-06 -85.669 0.0929738 31197.7 300.308 0.983523 0.319147 0.749046 0.749041 9.99958 2.98014e-06 1.19204e-05 0.130551 0.977234 0.929415 -0.0132934 4.89218e-06 0.500485 -1.86673e-20 6.86985e-24 -1.86605e-20 0.00139499 0.997819 8.59199e-05 0.152536 2.85161 0.00139499 0.997957 0.665818 0.00104305 0.00187949 0.000859199 0.455675 0.00187949 0.434663 0.000127246 1.02 0.887342 0.534775 0.285585 1.71601e-07 3.05465e-09 2393.01 3186.18 -0.0600559 0.482112 0.277655 0.257689 -0.592558 -0.169488 0.483305 -0.268555 -0.214756 1.323 1 5.17846e-288 293.028 3.07601e-285 2.02727 1.321 0.000299975 0.884145 0.6353 0.504333 0.399803 2.02755 128.045 83.111 18.6738 60.4756 0.00405891 0 -40 10
0.422 1.22345e-08 2.53883e-06 0.0683944 0.0683871 0.0120444 5.56112e-06 0.00115401 0.085493 0.000656087 0.0861445 0.855018 101.885 0.246483 0.711183 4.1154 0.0535174 0.0388246 0.961175 0.0198835 0.00423421 0.0191458 0.00407696 0.00511654 0.00585425 0.204662 0.23417 57.9652 -87.8941 125.96 15.9852 145.009 0.00014438 0.267071 192.937 0.310739 0.0673922 0.00409461 0.000561524 0.00138233 0.986994 0.991737 -2.97093e-06 -85.669 0.0929739 31197.7 300.31 0.983523 0.319147 0.74897 0.748966 9.99958 2.98014e-06 1.19205e-05 0.130552 0.977254 0.929424 -0.0132934 4.8922e-06 0.500488 -1.86682e-20 6.8702e-24 -1.86613e-20 0.00139499 0.997819 8.592e-05 0.152536 2.85161 0.00139499 0.997956 0.665934 0.00104307 0.00187949 0.0008592 0.455675 0.00187949 0.434673 0.000127249 1.02 0.887343 0.534775 0.285586 1.71601e-07 3.05466e-09 2392.99 3185.85 -0.0600327 0.482112 0.277654 0.257669 -0.592561 -0.169488 0.483374 -0.268553 -0.214827 1.324 1 3.14089e-288 293.05 1.86603e-285 2.02747 1.322 0.000299974 0.884 0.635363 0.503876 0.399837 2.02775 128.055 83.1147 18.674 60.4774 0.00405876 0 -40 10
0.423 1.22634e-08 2.53883e-06 0.0684907 0.0684834 0.0120444 5.57429e-06 0.00115401 0.0856133 0.000656094 0.0862648 0.855061 101.885 0.246478 0.711241 4.11547 0.053522 0.0388252 0.961175 0.0198834 0.00423428 0.0191457 0.00407701 0.00511663 0.00585433 0.204665 0.234173 57.9652 -87.8941 125.961 15.9852 145.009 0.000144365 0.267071 192.937 0.310739 0.0673922 0.00409461 0.000561524 0.00138233 0.986994 0.991737 -2.97094e-06 -85.669 0.0929739 31197.7 300.312 0.983523 0.319147 0.748894 0.74889 9.99958 2.98014e-06 1.19205e-05 0.130552 0.977273 0.929434 -0.0132934 4.89223e-06 0.500491 -1.8669e-20 6.87054e-24 -1.86622e-20 0.001395 0.997819 8.592e-05 0.152536 2.85161 0.001395 0.997955 0.666051 0.00104309 0.00187949 0.0008592 0.455675 0.00187949 0.434683 0.000127253 1.02 0.887344 0.534775 0.285587 1.71601e-07 3.05468e-09 2392.97 3185.53 -0.0600095 0.482112 0.277654 0.257649 -0.592565 -0.169488 0.483442 -0.268551 -0.214897 1.325 1 1.90505e-288 293.073 1.132e-285 2.02767 1.323 0.000299974 0.883856 0.635426 0.50342 0.399871 2.02795 128.066 83.1184 18.6742 60.4791 0.0040586 0 -40 10
0.424 1.22924e-08 2.53883e-06 0.0685868 0.0685796 0.0120444 5.58746e-06 0.00115401 0.0857336 0.000656101 0.0863851 0.855103 101.884 0.246473 0.7113 4.11554 0.0535267 0.0388259 0.961174 0.0198833 0.00423435 0.0191456 0.00407707 0.00511672 0.00585441 0.204669 0.234177 57.9653 -87.8941 125.963 15.9852 145.009 0.000144351 0.267072 192.937 0.310738 0.0673921 0.00409461 0.000561525 0.00138233 0.986994 0.991737 -2.97095e-06 -85.669 0.092974 31197.7 300.313 0.983523 0.319147 0.748819 0.748814 9.99958 2.98015e-06 1.19205e-05 0.130553 0.977293 0.929443 -0.0132934 4.89225e-06 0.500494 -1.86699e-20 6.87089e-24 -1.8663e-20 0.001395 0.997819 8.59201e-05 0.152536 2.85161 0.001395 0.997954 0.666167 0.00104311 0.00187949 0.000859201 0.455675 0.00187949 0.434693 0.000127256 1.02 0.887345 0.534775 0.285588 1.71601e-07 3.05469e-09 2392.96 3185.21 -0.0599864 0.482112 0.277654 0.257629 -0.592569 -0.169488 0.483511 -0.268549 -0.214967 1.326 1 1.15547e-288 293.096 6.86716e-286 2.02787 1.324 0.000299974 0.883712 0.635489 0.502965 0.399905 2.02816 128.077 83.122 18.6744 60.4809 0.00405845 0 -40 10
0.425 1.23214e-08 2.53883e-06 0.0686829 0.0686757 0.0120444 5.60063e-06 0.00115401 0.0858537 0.000656109 0.0865052 0.855145 101.884 0.246469 0.711358 4.11561 0.0535313 0.0388265 0.961173 0.0198832 0.00423442 0.0191455 0.00407713 0.0051168 0.0058545 0.204672 0.23418 57.9654 -87.8941 125.964 15.9851 145.009 0.000144336 0.267072 192.937 0.310738 0.0673921 0.00409461 0.000561525 0.00138233 0.986994 0.991737 -2.97096e-06 -85.669 0.0929741 31197.7 300.315 0.983523 0.319147 0.748744 0.748739 9.99958 2.98015e-06 1.19205e-05 0.130554 0.977312 0.929453 -0.0132934 4.89227e-06 0.500497 -1.86707e-20 6.87123e-24 -1.86639e-20 0.001395 0.997819 8.59201e-05 0.152536 2.85161 0.001395 0.997953 0.666283 0.00104313 0.00187949 0.000859201 0.455675 0.00187949 0.434703 0.00012726 1.02 0.887346 0.534774 0.285589 1.71601e-07 3.05471e-09 2392.94 3184.89 -0.0599634 0.482112 0.277654 0.257609 -0.592573 -0.169489 0.483579 -0.268548 -0.215037 1.327 1 7.00828e-289 293.119 4.16588e-286 2.02807 1.325 0.000299974 0.883569 0.635552 0.502511 0.399939 2.02836 128.088 83.1257 18.6747 60.4827 0.0040583 0 -40 10
0.426 1.23504e-08 2.53883e-06 0.068779 0.0687718 0.0120444 5.6138e-06 0.00115401 0.0859737 0.000656116 0.0866252 0.855187 101.884 0.246464 0.711417 4.11568 0.053536 0.0388272 0.961173 0.0198831 0.00423449 0.0191454 0.00407719 0.00511689 0.00585459 0.204676 0.234183 57.9654 -87.8941 125.965 15.9851 145.009 0.000144322 0.267072 192.937 0.310738 0.0673921 0.00409462 0.000561526 0.00138233 0.986994 0.991737 -2.97097e-06 -85.669 0.0929741 31197.7 300.317 0.983523 0.319147 0.748669 0.748665 9.99958 2.98015e-06 1.19205e-05 0.130554 0.977332 0.929462 -0.0132934 4.89229e-06 0.5005 -1.86716e-20 6.87158e-24 -1.86647e-20 0.001395 0.997819 8.59202e-05 0.152536 2.85162 0.001395 0.997952 0.666399 0.00104314 0.00187949 0.000859202 0.455675 0.00187949 0.434713 0.000127263 1.02 0.887346 0.534774 0.28559 1.71601e-07 3.05473e-09 2392.92 3184.57 -0.0599405 0.482112 0.277653 0.257589 -0.592576 -0.169489 0.483646 -0.268546 -0.215107 1.328 1 4.25073e-289 293.141 2.52718e-286 2.02827 1.326 0.000299974 0.883426 0.635615 0.502059 0.399974 2.02856 128.098 83.1294 18.6749 60.4845 0.00405814 0 -40 10
0.427 1.23793e-08 2.53883e-06 0.0688749 0.0688678 0.0120444 5.62697e-06 0.00115401 0.0860937 0.000656123 0.0867452 0.855229 101.884 0.246459 0.711476 4.11575 0.0535406 0.0388278 0.961172 0.019883 0.00423456 0.0191453 0.00407725 0.00511698 0.00585467 0.204679 0.234187 57.9655 -87.8942 125.967 15.985 145.009 0.000144307 0.267072 192.936 0.310738 0.067392 0.00409462 0.000561526 0.00138233 0.986994 0.991737 -2.97098e-06 -85.669 0.0929742 31197.7 300.319 0.983523 0.319147 0.748594 0.74859 9.99958 2.98016e-06 1.19205e-05 0.130555 0.977351 0.929472 -0.0132934 4.89231e-06 0.500502 -1.86724e-20 6.87192e-24 -1.86656e-20 0.001395 0.997819 8.59202e-05 0.152536 2.85162 0.001395 0.997951 0.666516 0.00104316 0.00187949 0.000859202 0.455674 0.00187949 0.434723 0.000127267 1.02 0.887347 0.534774 0.285591 1.71602e-07 3.05474e-09 2392.91 3184.25 -0.0599177 0.482112 0.277653 0.257569 -0.59258 -0.169489 0.483714 -0.268544 -0.215176 1.329 1 2.5782e-289 293.163 1.53308e-286 2.02847 1.327 0.000299974 0.883284 0.635677 0.501608 0.400008 2.02876 128.109 83.133 18.6751 60.4862 0.00405799 0 -40 10
0.428 1.24083e-08 2.53883e-06 0.0689708 0.0689637 0.0120443 5.64014e-06 0.00115401 0.0862135 0.00065613 0.086865 0.855272 101.884 0.246455 0.711535 4.11582 0.0535453 0.0388285 0.961172 0.0198829 0.00423463 0.0191452 0.00407731 0.00511707 0.00585476 0.204683 0.23419 57.9655 -87.8942 125.968 15.985 145.009 0.000144293 0.267072 192.936 0.310737 0.067392 0.00409462 0.000561527 0.00138234 0.986994 0.991737 -2.97099e-06 -85.669 0.0929742 31197.6 300.321 0.983523 0.319147 0.74852 0.748516 9.99958 2.98016e-06 1.19205e-05 0.130556 0.977371 0.929481 -0.0132934 4.89234e-06 0.500505 -1.86733e-20 6.87227e-24 -1.86664e-20 0.001395 0.997819 8.59203e-05 0.152536 2.85162 0.001395 0.99795 0.666632 0.00104318 0.00187949 0.000859203 0.455674 0.00187949 0.434733 0.00012727 1.02 0.887348 0.534774 0.285592 1.71602e-07 3.05476e-09 2392.89 3183.94 -0.059895 0.482112 0.277653 0.257549 -0.592584 -0.169489 0.483781 -0.268542 -0.215245 1.33 1 1.56376e-289 293.186 9.30023e-287 2.02867 1.328 0.000299974 0.883142 0.63574 0.501158 0.400042 2.02896 128.12 83.1366 18.6753 60.488 0.00405784 0 -40 10
0.429 1.24373e-08 2.53883e-06 0.0690666 0.0690595 0.0120443 5.6533e-06 0.00115401 0.0863332 0.000656137 0.0869848 0.855314 101.884 0.24645 0.711594 4.11589 0.05355 0.0388291 0.961171 0.0198828 0.00423471 0.0191452 0.00407737 0.00511715 0.00585484 0.204686 0.234194 57.9656 -87.8942 125.969 15.985 145.009 0.000144279 0.267072 192.936 0.310737 0.067392 0.00409462 0.000561527 0.00138234 0.986994 0.991737 -2.971e-06 -85.669 0.0929743 31197.6 300.323 0.983523 0.319147 0.748446 0.748441 9.99958 2.98016e-06 1.19205e-05 0.130557 0.97739 0.929491 -0.0132934 4.89236e-06 0.500508 -1.86741e-20 6.87261e-24 -1.86673e-20 0.001395 0.997819 8.59203e-05 0.152536 2.85162 0.001395 0.99795 0.666748 0.0010432 0.0018795 0.000859203 0.455674 0.00187949 0.434743 0.000127274 1.02 0.887349 0.534773 0.285594 1.71602e-07 3.05478e-09 2392.87 3183.62 -0.0598724 0.482112 0.277652 0.257529 -0.592587 -0.169489 0.483848 -0.268541 -0.215314 1.331 1 9.48467e-290 293.208 5.64186e-287 2.02887 1.329 0.000299973 0.883001 0.635803 0.500709 0.400076 2.02916 128.131 83.1402 18.6755 60.4897 0.00405769 0 -40 10
0.43 1.24662e-08 2.53883e-06 0.0691623 0.0691552 0.0120443 5.66647e-06 0.00115402 0.0864529 0.000656144 0.0871044 0.855357 101.884 0.246445 0.711653 4.11596 0.0535547 0.0388298 0.96117 0.0198828 0.00423478 0.0191451 0.00407742 0.00511724 0.00585493 0.20469 0.234197 57.9657 -87.8942 125.971 15.9849 145.009 0.000144265 0.267072 192.936 0.310737 0.0673919 0.00409462 0.000561527 0.00138234 0.986994 0.991737 -2.97101e-06 -85.669 0.0929743 31197.6 300.325 0.983523 0.319147 0.748372 0.748368 9.99958 2.98016e-06 1.19206e-05 0.130557 0.977409 0.9295 -0.0132934 4.89238e-06 0.500511 -1.8675e-20 6.87296e-24 -1.86681e-20 0.001395 0.997819 8.59204e-05 0.152537 2.85162 0.001395 0.997949 0.666864 0.00104322 0.0018795 0.000859204 0.455674 0.0018795 0.434753 0.000127277 1.02 0.88735 0.534773 0.285595 1.71602e-07 3.05479e-09 2392.86 3183.31 -0.0598498 0.482112 0.277652 0.257509 -0.592591 -0.169489 0.483915 -0.268539 -0.215382 1.332 1 5.75274e-290 293.23 3.42256e-287 2.02907 1.33 0.000299973 0.88286 0.635866 0.500262 0.40011 2.02936 128.141 83.1438 18.6757 60.4915 0.00405754 0 -40 10
0.431 1.24952e-08 2.53883e-06 0.0692579 0.0692509 0.0120443 5.67964e-06 0.00115402 0.0865724 0.000656151 0.087224 0.855399 101.884 0.246441 0.711712 4.11603 0.0535594 0.0388305 0.96117 0.0198827 0.00423485 0.019145 0.00407748 0.00511733 0.00585502 0.204693 0.234201 57.9657 -87.8942 125.972 15.9849 145.009 0.00014425 0.267072 192.936 0.310736 0.0673919 0.00409463 0.000561528 0.00138234 0.986994 0.991737 -2.97102e-06 -85.669 0.0929744 31197.6 300.327 0.983523 0.319147 0.748299 0.748294 9.99958 2.98017e-06 1.19206e-05 0.130558 0.977428 0.92951 -0.0132934 4.8924e-06 0.500514 -1.86758e-20 6.8733e-24 -1.8669e-20 0.001395 0.997818 8.59204e-05 0.152537 2.85162 0.001395 0.997948 0.66698 0.00104324 0.0018795 0.000859204 0.455674 0.0018795 0.434763 0.000127281 1.02 0.88735 0.534773 0.285596 1.71602e-07 3.05481e-09 2392.84 3182.99 -0.0598273 0.482112 0.277652 0.25749 -0.592595 -0.169489 0.483981 -0.268537 -0.21545 1.333 1 3.48922e-290 293.252 2.07625e-287 2.02927 1.331 0.000299973 0.88272 0.635928 0.499815 0.400144 2.02956 128.152 83.1474 18.6759 60.4932 0.00405739 0 -40 10
0.432 1.25242e-08 2.53883e-06 0.0693535 0.0693465 0.0120443 5.69281e-06 0.00115402 0.0866919 0.000656158 0.0873434 0.855442 101.884 0.246436 0.711772 4.1161 0.0535641 0.0388311 0.961169 0.0198826 0.00423492 0.0191449 0.00407754 0.00511742 0.00585511 0.204697 0.234204 57.9658 -87.8942 125.973 15.9849 145.009 0.000144236 0.267073 192.936 0.310736 0.0673919 0.00409463 0.000561528 0.00138234 0.986994 0.991737 -2.97103e-06 -85.669 0.0929744 31197.6 300.329 0.983523 0.319147 0.748225 0.748221 9.99958 2.98017e-06 1.19206e-05 0.130559 0.977447 0.929519 -0.0132934 4.89242e-06 0.500517 -1.86767e-20 6.87365e-24 -1.86698e-20 0.001395 0.997818 8.59205e-05 0.152537 2.85162 0.001395 0.997947 0.667096 0.00104326 0.0018795 0.000859205 0.455674 0.0018795 0.434773 0.000127285 1.02 0.887351 0.534773 0.285597 1.71602e-07 3.05483e-09 2392.83 3182.68 -0.0598049 0.482112 0.277651 0.25747 -0.592598 -0.169489 0.484048 -0.268535 -0.215518 1.334 1 2.11632e-290 293.275 1.25953e-287 2.02947 1.332 0.000299973 0.88258 0.635991 0.49937 0.400177 2.02976 128.163 83.151 18.6761 60.4949 0.00405724 0 -40 10
0.433 1.25532e-08 2.53883e-06 0.069449 0.069442 0.0120443 5.70598e-06 0.00115402 0.0868113 0.000656166 0.0874628 0.855485 101.884 0.246431 0.711831 4.11617 0.0535688 0.0388318 0.961168 0.0198825 0.004235 0.0191448 0.0040776 0.00511751 0.00585519 0.2047 0.234208 57.9658 -87.8942 125.975 15.9848 145.009 0.000144222 0.267073 192.936 0.310736 0.0673918 0.00409463 0.000561529 0.00138234 0.986994 0.991737 -2.97104e-06 -85.6689 0.0929745 31197.6 300.331 0.983523 0.319147 0.748152 0.748148 9.99958 2.98017e-06 1.19206e-05 0.13056 0.977466 0.929528 -0.0132934 4.89245e-06 0.50052 -1.86775e-20 6.87399e-24 -1.86707e-20 0.001395 0.997818 8.59205e-05 0.152537 2.85162 0.001395 0.997946 0.667212 0.00104328 0.0018795 0.000859205 0.455674 0.0018795 0.434783 0.000127288 1.02 0.887352 0.534772 0.285598 1.71603e-07 3.05484e-09 2392.81 3182.37 -0.0597826 0.482112 0.277651 0.257451 -0.592602 -0.169489 0.484114 -0.268534 -0.215586 1.335 1 1.28361e-290 293.297 7.64074e-288 2.02967 1.333 0.000299973 0.88244 0.636053 0.498927 0.400211 2.02996 128.173 83.1546 18.6763 60.4967 0.00405709 0 -40 10
0.434 1.25821e-08 2.53883e-06 0.0695444 0.0695374 0.0120443 5.71915e-06 0.00115402 0.0869305 0.000656172 0.0875821 0.855528 101.884 0.246426 0.711891 4.11625 0.0535735 0.0388325 0.961167 0.0198824 0.00423507 0.0191447 0.00407766 0.0051176 0.00585528 0.204704 0.234211 57.9659 -87.8942 125.976 15.9848 145.009 0.000144208 0.267073 192.936 0.310736 0.0673918 0.00409463 0.000561529 0.00138234 0.986994 0.991737 -2.97105e-06 -85.6689 0.0929746 31197.6 300.333 0.983523 0.319147 0.748079 0.748075 9.99958 2.98018e-06 1.19206e-05 0.13056 0.977485 0.929537 -0.0132934 4.89247e-06 0.500523 -1.86784e-20 6.87433e-24 -1.86715e-20 0.001395 0.997818 8.59206e-05 0.152537 2.85162 0.001395 0.997945 0.667328 0.00104329 0.0018795 0.000859206 0.455673 0.0018795 0.434793 0.000127292 1.02 0.887353 0.534772 0.285599 1.71603e-07 3.05486e-09 2392.79 3182.06 -0.0597604 0.482112 0.277651 0.257431 -0.592606 -0.169489 0.484179 -0.268532 -0.215654 1.336 1 7.78549e-291 293.318 4.63514e-288 2.02987 1.334 0.000299973 0.882302 0.636116 0.498484 0.400245 2.03016 128.184 83.1581 18.6765 60.4984 0.00405694 0 -40 10
0.435 1.26111e-08 2.53883e-06 0.0696397 0.0696328 0.0120443 5.73232e-06 0.00115402 0.0870497 0.000656179 0.0877013 0.85557 101.884 0.246422 0.711951 4.11632 0.0535783 0.0388332 0.961167 0.0198823 0.00423514 0.0191446 0.00407773 0.00511769 0.00585537 0.204708 0.234215 57.966 -87.8942 125.977 15.9847 145.009 0.000144194 0.267073 192.936 0.310735 0.0673917 0.00409463 0.00056153 0.00138235 0.986994 0.991737 -2.97106e-06 -85.6689 0.0929746 31197.5 300.335 0.983523 0.319147 0.748007 0.748003 9.99958 2.98018e-06 1.19206e-05 0.130561 0.977504 0.929547 -0.0132934 4.89249e-06 0.500526 -1.86792e-20 6.87468e-24 -1.86724e-20 0.001395 0.997818 8.59206e-05 0.152537 2.85162 0.001395 0.997945 0.667444 0.00104331 0.0018795 0.000859206 0.455673 0.0018795 0.434803 0.000127295 1.02 0.887354 0.534772 0.2856 1.71603e-07 3.05488e-09 2392.78 3181.75 -0.0597382 0.482112 0.277651 0.257412 -0.592609 -0.169489 0.484245 -0.26853 -0.215721 1.337 1 4.72214e-291 293.34 2.81184e-288 2.03007 1.335 0.000299973 0.882163 0.636178 0.498043 0.400279 2.03036 128.195 83.1617 18.6768 60.5001 0.00405679 0 -40 10
0.436 1.26401e-08 2.53883e-06 0.069735 0.0697281 0.0120442 5.74548e-06 0.00115402 0.0871688 0.000656186 0.0878203 0.855613 101.884 0.246417 0.71201 4.11639 0.053583 0.0388339 0.961166 0.0198822 0.00423522 0.0191445 0.00407779 0.00511778 0.00585546 0.204711 0.234218 57.966 -87.8942 125.979 15.9847 145.009 0.00014418 0.267073 192.935 0.310735 0.0673917 0.00409464 0.00056153 0.00138235 0.986994 0.991737 -2.97107e-06 -85.6689 0.0929747 31197.5 300.337 0.983523 0.319147 0.747935 0.74793 9.99958 2.98018e-06 1.19206e-05 0.130562 0.977523 0.929556 -0.0132934 4.89251e-06 0.500529 -1.86801e-20 6.87502e-24 -1.86732e-20 0.00139501 0.997818 8.59207e-05 0.152537 2.85162 0.00139501 0.997944 0.66756 0.00104333 0.0018795 0.000859207 0.455673 0.0018795 0.434813 0.000127299 1.02 0.887355 0.534772 0.285602 1.71603e-07 3.05489e-09 2392.76 3181.44 -0.0597162 0.482112 0.27765 0.257393 -0.592613 -0.169489 0.48431 -0.268528 -0.215788 1.338 1 2.86412e-291 293.362 1.70576e-288 2.03027 1.336 0.000299973 0.882026 0.636241 0.497602 0.400313 2.03055 128.205 83.1652 18.677 60.5018 0.00405665 0 -40 10
0.437 1.2669e-08 2.53883e-06 0.0698302 0.0698233 0.0120442 5.75865e-06 0.00115402 0.0872877 0.000656193 0.0879393 0.855656 101.884 0.246412 0.71207 4.11646 0.0535878 0.0388345 0.961165 0.0198821 0.00423529 0.0191444 0.00407785 0.00511787 0.00585555 0.204715 0.234222 57.9661 -87.8942 125.98 15.9847 145.009 0.000144166 0.267073 192.935 0.310735 0.0673917 0.00409464 0.00056153 0.00138235 0.986994 0.991737 -2.97108e-06 -85.6689 0.0929747 31197.5 300.339 0.983523 0.319147 0.747863 0.747858 9.99958 2.98019e-06 1.19206e-05 0.130563 0.977542 0.929565 -0.0132934 4.89254e-06 0.500533 -1.86809e-20 6.87536e-24 -1.86741e-20 0.00139501 0.997818 8.59207e-05 0.152537 2.85162 0.00139501 0.997943 0.667675 0.00104335 0.0018795 0.000859207 0.455673 0.0018795 0.434823 0.000127302 1.02 0.887355 0.534772 0.285603 1.71603e-07 3.05491e-09 2392.74 3181.14 -0.0596942 0.482112 0.27765 0.257373 -0.592616 -0.169489 0.484375 -0.268527 -0.215855 1.339 1 1.73718e-291 293.384 1.03478e-288 2.03047 1.337 0.000299972 0.881888 0.636303 0.497163 0.400347 2.03075 128.216 83.1687 18.6772 60.5035 0.0040565 0 -40 10
0.438 1.2698e-08 2.53883e-06 0.0699253 0.0699184 0.0120442 5.77182e-06 0.00115402 0.0874066 0.0006562 0.0880582 0.8557 101.883 0.246407 0.712131 4.11654 0.0535925 0.0388352 0.961165 0.019882 0.00423536 0.0191444 0.00407791 0.00511796 0.00585564 0.204719 0.234226 57.9662 -87.8942 125.981 15.9846 145.009 0.000144152 0.267073 192.935 0.310734 0.0673916 0.00409464 0.000561531 0.00138235 0.986994 0.991737 -2.97109e-06 -85.6689 0.0929748 31197.5 300.341 0.983523 0.319147 0.747791 0.747786 9.99958 2.98019e-06 1.19207e-05 0.130563 0.97756 0.929574 -0.0132934 4.89256e-06 0.500536 -1.86818e-20 6.87571e-24 -1.86749e-20 0.00139501 0.997818 8.59208e-05 0.152537 2.85162 0.00139501 0.997942 0.667791 0.00104337 0.0018795 0.000859208 0.455673 0.0018795 0.434833 0.000127306 1.02 0.887356 0.534771 0.285604 1.71603e-07 3.05493e-09 2392.73 3180.83 -0.0596723 0.482112 0.27765 0.257354 -0.59262 -0.169489 0.48444 -0.268525 -0.215921 1.34 1 1.05365e-291 293.405 6.27731e-289 2.03067 1.338 0.000299972 0.881752 0.636365 0.496725 0.40038 2.03095 128.227 83.1722 18.6774 60.5052 0.00405635 0 -40 10
0.439 1.2727e-08 2.53883e-06 0.0700203 0.0700135 0.0120442 5.78499e-06 0.00115402 0.0875254 0.000656207 0.088177 0.855743 101.883 0.246403 0.712191 4.11661 0.0535973 0.0388359 0.961164 0.0198819 0.00423544 0.0191443 0.00407797 0.00511805 0.00585573 0.204722 0.234229 57.9662 -87.8942 125.982 15.9846 145.009 0.000144139 0.267073 192.935 0.310734 0.0673916 0.00409464 0.000561531 0.00138235 0.986994 0.991737 -2.9711e-06 -85.6689 0.0929748 31197.5 300.343 0.983523 0.319147 0.747719 0.747715 9.99958 2.98019e-06 1.19207e-05 0.130564 0.977579 0.929583 -0.0132934 4.89258e-06 0.500539 -1.86826e-20 6.87605e-24 -1.86757e-20 0.00139501 0.997818 8.59209e-05 0.152537 2.85162 0.00139501 0.997941 0.667907 0.00104339 0.00187951 0.000859209 0.455673 0.0018795 0.434843 0.000127309 1.02 0.887357 0.534771 0.285605 1.71604e-07 3.05494e-09 2392.71 3180.53 -0.0596505 0.482113 0.277649 0.257335 -0.592624 -0.169489 0.484504 -0.268523 -0.215987 1.341 1 6.39072e-292 293.427 3.80803e-289 2.03087 1.339 0.000299972 0.881615 0.636427 0.496289 0.400414 2.03115 128.237 83.1757 18.6776 60.5069 0.00405621 0 -40 10
0.44 1.27559e-08 2.53883e-06 0.0701153 0.0701085 0.0120442 5.79816e-06 0.00115402 0.0876441 0.000656214 0.0882957 0.855786 101.883 0.246398 0.712251 4.11668 0.0536021 0.0388366 0.961163 0.0198819 0.00423551 0.0191442 0.00407803 0.00511815 0.00585582 0.204726 0.234233 57.9663 -87.8942 125.984 15.9846 145.009 0.000144125 0.267074 192.935 0.310734 0.0673916 0.00409464 0.000561532 0.00138235 0.986994 0.991737 -2.97111e-06 -85.6689 0.0929749 31197.5 300.345 0.983523 0.319147 0.747648 0.747644 9.99958 2.9802e-06 1.19207e-05 0.130565 0.977598 0.929592 -0.0132934 4.8926e-06 0.500542 -1.86835e-20 6.87639e-24 -1.86766e-20 0.00139501 0.997818 8.59209e-05 0.152538 2.85162 0.00139501 0.99794 0.668022 0.00104341 0.00187951 0.000859209 0.455673 0.00187951 0.434853 0.000127313 1.02 0.887358 0.534771 0.285606 1.71604e-07 3.05496e-09 2392.69 3180.22 -0.0596288 0.482113 0.277649 0.257316 -0.592627 -0.16949 0.484569 -0.268521 -0.216053 1.342 1 3.87617e-292 293.448 2.31008e-289 2.03107 1.34 0.000299972 0.881479 0.636489 0.495853 0.400448 2.03135 128.248 83.1792 18.6778 60.5086 0.00405606 0 -40 10
0.441 1.27849e-08 2.53884e-06 0.0702102 0.0702034 0.0120442 5.81132e-06 0.00115402 0.0877627 0.000656221 0.0884143 0.855829 101.883 0.246393 0.712312 4.11676 0.0536069 0.0388373 0.961163 0.0198818 0.00423559 0.0191441 0.00407809 0.00511824 0.00585591 0.20473 0.234236 57.9663 -87.8942 125.985 15.9845 145.009 0.000144111 0.267074 192.935 0.310734 0.0673915 0.00409465 0.000561532 0.00138235 0.986994 0.991737 -2.97112e-06 -85.6689 0.092975 31197.5 300.347 0.983523 0.319147 0.747577 0.747573 9.99958 2.9802e-06 1.19207e-05 0.130566 0.977616 0.929601 -0.0132934 4.89263e-06 0.500545 -1.86843e-20 6.87673e-24 -1.86774e-20 0.00139501 0.997818 8.5921e-05 0.152538 2.85162 0.00139501 0.99794 0.668138 0.00104343 0.00187951 0.00085921 0.455672 0.00187951 0.434863 0.000127316 1.02 0.887359 0.534771 0.285607 1.71604e-07 3.05498e-09 2392.68 3179.92 -0.0596071 0.482113 0.277649 0.257297 -0.592631 -0.16949 0.484633 -0.26852 -0.216119 1.343 1 2.35102e-292 293.469 1.40137e-289 2.03127 1.341 0.000299972 0.881344 0.636552 0.495419 0.400481 2.03155 128.259 83.1826 18.678 60.5102 0.00405592 0 -40 10
0.442 1.28139e-08 2.53884e-06 0.070305 0.0702982 0.0120442 5.82449e-06 0.00115402 0.0878812 0.000656227 0.0885328 0.855873 101.883 0.246388 0.712373 4.11683 0.0536117 0.038838 0.961162 0.0198817 0.00423566 0.019144 0.00407816 0.00511833 0.005856 0.204733 0.23424 57.9664 -87.8942 125.986 15.9845 145.009 0.000144098 0.267074 192.935 0.310733 0.0673915 0.00409465 0.000561533 0.00138236 0.986994 0.991737 -2.97113e-06 -85.6689 0.092975 31197.4 300.349 0.983523 0.319147 0.747506 0.747502 9.99958 2.9802e-06 1.19207e-05 0.130566 0.977635 0.92961 -0.0132934 4.89265e-06 0.500548 -1.86851e-20 6.87708e-24 -1.86783e-20 0.00139501 0.997818 8.5921e-05 0.152538 2.85163 0.00139501 0.997939 0.668254 0.00104344 0.00187951 0.00085921 0.455672 0.00187951 0.434872 0.00012732 1.02 0.88736 0.53477 0.285608 1.71604e-07 3.05499e-09 2392.66 3179.62 -0.0595855 0.482113 0.277649 0.257278 -0.592634 -0.16949 0.484696 -0.268518 -0.216185 1.344 1 1.42596e-292 293.491 8.50121e-290 2.03146 1.342 0.000299972 0.881209 0.636614 0.494986 0.400515 2.03175 128.269 83.1861 18.6782 60.5119 0.00405577 0 -40 10
0.443 1.28429e-08 2.53884e-06 0.0703997 0.0703929 0.0120441 5.83766e-06 0.00115402 0.0879996 0.000656234 0.0886512 0.855916 101.883 0.246383 0.712433 4.1169 0.0536165 0.0388387 0.961161 0.0198816 0.00423574 0.0191439 0.00407822 0.00511842 0.00585609 0.204737 0.234244 57.9665 -87.8942 125.987 15.9845 145.009 0.000144084 0.267074 192.935 0.310733 0.0673915 0.00409465 0.000561533 0.00138236 0.986994 0.991737 -2.97114e-06 -85.6689 0.0929751 31197.4 300.351 0.983523 0.319147 0.747436 0.747432 9.99958 2.98021e-06 1.19207e-05 0.130567 0.977653 0.929619 -0.0132934 4.89267e-06 0.500551 -1.8686e-20 6.87742e-24 -1.86791e-20 0.00139501 0.997818 8.59211e-05 0.152538 2.85163 0.00139501 0.997938 0.668369 0.00104346 0.00187951 0.000859211 0.455672 0.00187951 0.434882 0.000127323 1.02 0.88736 0.53477 0.28561 1.71604e-07 3.05501e-09 2392.64 3179.32 -0.059564 0.482113 0.277648 0.257259 -0.592638 -0.16949 0.48476 -0.268516 -0.21625 1.345 1 8.6489e-293 293.512 5.15712e-290 2.03166 1.343 0.000299972 0.881075 0.636676 0.494554 0.400549 2.03194 128.28 83.1895 18.6784 60.5136 0.00405563 0 -40 10
0.444 1.28718e-08 2.53884e-06 0.0704943 0.0704876 0.0120441 5.85083e-06 0.00115402 0.0881179 0.000656241 0.0887696 0.85596 101.883 0.246379 0.712494 4.11698 0.0536214 0.0388394 0.961161 0.0198815 0.00423582 0.0191438 0.00407828 0.00511852 0.00585619 0.204741 0.234247 57.9665 -87.8942 125.989 15.9844 145.009 0.000144071 0.267074 192.935 0.310733 0.0673914 0.00409465 0.000561534 0.00138236 0.986994 0.991737 -2.97115e-06 -85.6689 0.0929751 31197.4 300.353 0.983523 0.319147 0.747366 0.747361 9.99958 2.98021e-06 1.19207e-05 0.130568 0.977671 0.929628 -0.0132934 4.8927e-06 0.500554 -1.86868e-20 6.87776e-24 -1.868e-20 0.00139501 0.997818 8.59211e-05 0.152538 2.85163 0.00139501 0.997937 0.668485 0.00104348 0.00187951 0.000859211 0.455672 0.00187951 0.434892 0.000127327 1.02 0.887361 0.53477 0.285611 1.71605e-07 3.05503e-09 2392.63 3179.02 -0.0595426 0.482113 0.277648 0.257241 -0.592641 -0.16949 0.484823 -0.268514 -0.216315 1.346 1 5.24582e-293 293.533 3.12848e-290 2.03186 1.344 0.000299971 0.880941 0.636738 0.494123 0.400582 2.03214 128.29 83.193 18.6786 60.5152 0.00405548 0 -40 10
0.445 1.29008e-08 2.53884e-06 0.0705889 0.0705822 0.0120441 5.864e-06 0.00115402 0.0882361 0.000656248 0.0888878 0.856003 101.883 0.246374 0.712555 4.11705 0.0536262 0.0388401 0.96116 0.0198814 0.00423589 0.0191437 0.00407834 0.00511861 0.00585628 0.204744 0.234251 57.9666 -87.8942 125.99 15.9844 145.009 0.000144057 0.267074 192.934 0.310732 0.0673914 0.00409465 0.000561534 0.00138236 0.986994 0.991737 -2.97116e-06 -85.6689 0.0929752 31197.4 300.355 0.983523 0.319147 0.747296 0.747291 9.99958 2.98021e-06 1.19207e-05 0.130569 0.97769 0.929637 -0.0132934 4.89272e-06 0.500557 -1.86877e-20 6.8781e-24 -1.86808e-20 0.00139501 0.997818 8.59212e-05 0.152538 2.85163 0.00139501 0.997937 0.6686 0.0010435 0.00187951 0.000859212 0.455672 0.00187951 0.434902 0.000127331 1.02 0.887362 0.53477 0.285612 1.71605e-07 3.05504e-09 2392.61 3178.72 -0.0595213 0.482113 0.277648 0.257222 -0.592645 -0.16949 0.484886 -0.268513 -0.21638 1.347 1 3.18175e-293 293.554 1.89784e-290 2.03206 1.345 0.000299971 0.880808 0.6368 0.493694 0.400616 2.03234 128.301 83.1964 18.6788 60.5169 0.00405534 0 -40 10
0.446 1.29298e-08 2.53884e-06 0.0706834 0.0706767 0.0120441 5.87716e-06 0.00115402 0.0883543 0.000656254 0.0890059 0.856047 101.883 0.246369 0.712616 4.11713 0.0536311 0.0388408 0.961159 0.0198813 0.00423597 0.0191436 0.00407841 0.00511871 0.00585637 0.204748 0.234255 57.9667 -87.8942 125.991 15.9843 145.009 0.000144044 0.267074 192.934 0.310732 0.0673914 0.00409466 0.000561534 0.00138236 0.986994 0.991737 -2.97117e-06 -85.6689 0.0929753 31197.4 300.357 0.983523 0.319147 0.747226 0.747222 9.99958 2.98022e-06 1.19208e-05 0.13057 0.977708 0.929646 -0.0132934 4.89274e-06 0.500561 -1.86885e-20 6.87844e-24 -1.86816e-20 0.00139501 0.997818 8.59212e-05 0.152538 2.85163 0.00139501 0.997936 0.668716 0.00104352 0.00187951 0.000859212 0.455672 0.00187951 0.434912 0.000127334 1.02 0.887363 0.534769 0.285613 1.71605e-07 3.05506e-09 2392.59 3178.42 -0.0595001 0.482113 0.277647 0.257203 -0.592648 -0.16949 0.484949 -0.268511 -0.216445 1.348 1 1.92983e-293 293.575 1.15129e-290 2.03226 1.346 0.000299971 0.880675 0.636861 0.493265 0.400649 2.03254 128.312 83.1998 18.679 60.5185 0.0040552 0 -40 10
0.447 1.29587e-08 2.53884e-06 0.0707778 0.0707712 0.0120441 5.89033e-06 0.00115402 0.0884723 0.000656261 0.0891239 0.856091 101.883 0.246364 0.712678 4.1172 0.0536359 0.0388416 0.961158 0.0198812 0.00423605 0.0191435 0.00407847 0.0051188 0.00585646 0.204752 0.234258 57.9667 -87.8942 125.992 15.9843 145.009 0.00014403 0.267074 192.934 0.310732 0.0673913 0.00409466 0.000561535 0.00138236 0.986994 0.991737 -2.97118e-06 -85.6689 0.0929753 31197.4 300.359 0.983523 0.319147 0.747157 0.747152 9.99958 2.98022e-06 1.19208e-05 0.13057 0.977726 0.929655 -0.0132934 4.89276e-06 0.500564 -1.86894e-20 6.87879e-24 -1.86825e-20 0.00139501 0.997818 8.59213e-05 0.152538 2.85163 0.00139501 0.997935 0.668831 0.00104354 0.00187951 0.000859213 0.455672 0.00187951 0.434922 0.000127338 1.02 0.887364 0.534769 0.285614 1.71605e-07 3.05508e-09 2392.58 3178.13 -0.0594789 0.482113 0.277647 0.257185 -0.592652 -0.16949 0.485012 -0.268509 -0.216509 1.349 1 1.1705e-293 293.596 6.98412e-291 2.03245 1.347 0.000299971 0.880543 0.636923 0.492838 0.400683 2.03273 128.322 83.2032 18.6792 60.5202 0.00405506 0 -40 10
0.448 1.29877e-08 2.53884e-06 0.0708722 0.0708655 0.0120441 5.9035e-06 0.00115402 0.0885902 0.000656268 0.0892419 0.856135 101.883 0.246359 0.712739 4.11728 0.0536408 0.0388423 0.961158 0.0198811 0.00423612 0.0191434 0.00407853 0.0051189 0.00585656 0.204756 0.234262 57.9668 -87.8942 125.994 15.9843 145.009 0.000144017 0.267075 192.934 0.310732 0.0673913 0.00409466 0.000561535 0.00138236 0.986994 0.991737 -2.97119e-06 -85.6689 0.0929754 31197.4 300.361 0.983523 0.319147 0.747087 0.747083 9.99958 2.98022e-06 1.19208e-05 0.130571 0.977744 0.929664 -0.0132934 4.89279e-06 0.500567 -1.86902e-20 6.87913e-24 -1.86833e-20 0.00139501 0.997818 8.59213e-05 0.152538 2.85163 0.00139501 0.997934 0.668946 0.00104356 0.00187951 0.000859213 0.455671 0.00187951 0.434932 0.000127341 1.02 0.887365 0.534769 0.285615 1.71605e-07 3.0551e-09 2392.56 3177.83 -0.0594578 0.482113 0.277647 0.257166 -0.592655 -0.16949 0.485074 -0.268507 -0.216573 1.35 1 7.09945e-294 293.617 4.2368e-291 2.03265 1.348 0.000299971 0.880411 0.636985 0.492412 0.400716 2.03293 128.333 83.2065 18.6794 60.5218 0.00405492 0 -40 10
0.449 1.30167e-08 2.53884e-06 0.0709664 0.0709598 0.0120441 5.91667e-06 0.00115402 0.0887081 0.000656274 0.0893597 0.856179 101.883 0.246354 0.712801 4.11736 0.0536457 0.038843 0.961157 0.019881 0.0042362 0.0191434 0.0040786 0.00511899 0.00585665 0.20476 0.234266 57.9668 -87.8942 125.995 15.9842 145.009 0.000144004 0.267075 192.934 0.310731 0.0673913 0.00409466 0.000561536 0.00138237 0.986994 0.991737 -2.9712e-06 -85.6688 0.0929754 31197.3 300.364 0.983523 0.319147 0.747018 0.747014 9.99958 2.98023e-06 1.19208e-05 0.130572 0.977762 0.929672 -0.0132934 4.89281e-06 0.50057 -1.8691e-20 6.87947e-24 -1.86841e-20 0.00139502 0.997818 8.59214e-05 0.152538 2.85163 0.00139502 0.997933 0.669062 0.00104358 0.00187952 0.000859214 0.455671 0.00187951 0.434942 0.000127345 1.02 0.887365 0.534769 0.285617 1.71605e-07 3.05511e-09 2392.55 3177.54 -0.0594368 0.482113 0.277647 0.257148 -0.592658 -0.16949 0.485136 -0.268505 -0.216637 1.351 1 4.30603e-294 293.638 2.57018e-291 2.03285 1.349 0.000299971 0.880279 0.637047 0.491987 0.40075 2.03313 128.343 83.2099 18.6796 60.5234 0.00405477 0 -40 10
0.45 1.30456e-08 2.53884e-06 0.0710606 0.0710541 0.0120441 5.92983e-06 0.00115402 0.0888258 0.000656281 0.0894775 0.856223 101.883 0.246349 0.712862 4.11743 0.0536506 0.0388437 0.961156 0.0198809 0.00423628 0.0191433 0.00407866 0.00511909 0.00585674 0.204763 0.23427 57.9669 -87.8942 125.996 15.9842 145.009 0.00014399 0.267075 192.934 0.310731 0.0673912 0.00409466 0.000561536 0.00138237 0.986994 0.991737 -2.97122e-06 -85.6688 0.0929755 31197.3 300.366 0.983523 0.319147 0.74695 0.746945 9.99958 2.98023e-06 1.19208e-05 0.130573 0.97778 0.929681 -0.0132934 4.89283e-06 0.500573 -1.86919e-20 6.87981e-24 -1.8685e-20 0.00139502 0.997818 8.59215e-05 0.152539 2.85163 0.00139502 0.997933 0.669177 0.0010436 0.00187952 0.000859215 0.455671 0.00187952 0.434951 0.000127348 1.02 0.887366 0.534768 0.285618 1.71606e-07 3.05513e-09 2392.53 3177.25 -0.0594159 0.482113 0.277646 0.257129 -0.592662 -0.16949 0.485198 -0.268504 -0.216701 1.352 1 2.61174e-294 293.658 1.55915e-291 2.03304 1.35 0.00029997 0.880148 0.637108 0.491563 0.400783 2.03332 128.354 83.2133 18.6798 60.525 0.00405463 0 -40 10
0.451 1.30746e-08 2.53884e-06 0.0711548 0.0711482 0.012044 5.943e-06 0.00115402 0.0889435 0.000656287 0.0895951 0.856267 101.882 0.246345 0.712924 4.11751 0.0536554 0.0388444 0.961156 0.0198808 0.00423636 0.0191432 0.00407873 0.00511918 0.00585684 0.204767 0.234273 57.967 -87.8942 125.997 15.9842 145.009 0.000143977 0.267075 192.934 0.310731 0.0673912 0.00409467 0.000561537 0.00138237 0.986994 0.991737 -2.97123e-06 -85.6688 0.0929756 31197.3 300.368 0.983523 0.319147 0.746881 0.746877 9.99958 2.98023e-06 1.19208e-05 0.130573 0.977798 0.92969 -0.0132934 4.89286e-06 0.500577 -1.86927e-20 6.88015e-24 -1.86858e-20 0.00139502 0.997818 8.59215e-05 0.152539 2.85163 0.00139502 0.997932 0.669292 0.00104361 0.00187952 0.000859215 0.455671 0.00187952 0.434961 0.000127352 1.02 0.887367 0.534768 0.285619 1.71606e-07 3.05515e-09 2392.51 3176.95 -0.059395 0.482113 0.277646 0.257111 -0.592665 -0.16949 0.48526 -0.268502 -0.216764 1.353 1 1.5841e-294 293.679 9.45832e-292 2.03324 1.351 0.00029997 0.880018 0.63717 0.491141 0.400817 2.03352 128.364 83.2166 18.68 60.5267 0.00405449 0 -40 10
0.452 1.31036e-08 2.53884e-06 0.0712488 0.0712423 0.012044 5.95617e-06 0.00115402 0.089061 0.000656294 0.0897127 0.856311 101.882 0.24634 0.712986 4.11759 0.0536604 0.0388452 0.961155 0.0198807 0.00423643 0.0191431 0.00407879 0.00511928 0.00585693 0.204771 0.234277 57.967 -87.8942 125.999 15.9841 145.009 0.000143964 0.267075 192.934 0.31073 0.0673911 0.00409467 0.000561537 0.00138237 0.986994 0.991737 -2.97124e-06 -85.6688 0.0929756 31197.3 300.37 0.983523 0.319147 0.746813 0.746808 9.99958 2.98024e-06 1.19208e-05 0.130574 0.977816 0.929699 -0.0132934 4.89288e-06 0.50058 -1.86935e-20 6.88049e-24 -1.86867e-20 0.00139502 0.997818 8.59216e-05 0.152539 2.85163 0.00139502 0.997931 0.669407 0.00104363 0.00187952 0.000859216 0.455671 0.00187952 0.434971 0.000127355 1.02 0.887368 0.534768 0.28562 1.71606e-07 3.05517e-09 2392.5 3176.66 -0.0593743 0.482113 0.277646 0.257093 -0.592669 -0.16949 0.485321 -0.2685 -0.216827 1.354 1 9.60806e-295 293.699 5.73771e-292 2.03344 1.352 0.00029997 0.879888 0.637232 0.490719 0.40085 2.03372 128.375 83.22 18.6802 60.5283 0.00405436 0 -40 10
0.453 1.31325e-08 2.53884e-06 0.0713428 0.0713363 0.012044 5.96934e-06 0.00115402 0.0891785 0.000656301 0.0898302 0.856355 101.882 0.246335 0.713048 4.11766 0.0536653 0.0388459 0.961154 0.0198806 0.00423651 0.019143 0.00407886 0.00511937 0.00585703 0.204775 0.234281 57.9671 -87.8943 126 15.9841 145.009 0.000143951 0.267075 192.934 0.31073 0.0673911 0.00409467 0.000561538 0.00138237 0.986994 0.991736 -2.97125e-06 -85.6688 0.0929757 31197.3 300.372 0.983523 0.319147 0.746745 0.74674 9.99958 2.98024e-06 1.19209e-05 0.130575 0.977834 0.929707 -0.0132934 4.8929e-06 0.500583 -1.86944e-20 6.88083e-24 -1.86875e-20 0.00139502 0.997818 8.59216e-05 0.152539 2.85163 0.00139502 0.99793 0.669523 0.00104365 0.00187952 0.000859216 0.455671 0.00187952 0.434981 0.000127359 1.02 0.887369 0.534768 0.285621 1.71606e-07 3.05518e-09 2392.48 3176.37 -0.0593536 0.482113 0.277645 0.257075 -0.592672 -0.16949 0.485382 -0.268498 -0.21689 1.355 1 5.82758e-295 293.72 3.48068e-292 2.03363 1.353 0.00029997 0.879758 0.637293 0.490299 0.400883 2.03391 128.385 83.2233 18.6804 60.5299 0.00405422 0 -40 10
0.454 1.31615e-08 2.53884e-06 0.0714367 0.0714302 0.012044 5.9825e-06 0.00115402 0.0892958 0.000656307 0.0899475 0.856399 101.882 0.24633 0.71311 4.11774 0.0536702 0.0388466 0.961153 0.0198805 0.00423659 0.0191429 0.00407892 0.00511947 0.00585712 0.204779 0.234285 57.9672 -87.8943 126.001 15.984 145.009 0.000143938 0.267075 192.933 0.31073 0.0673911 0.00409467 0.000561538 0.00138237 0.986994 0.991736 -2.97126e-06 -85.6688 0.0929757 31197.3 300.374 0.983523 0.319147 0.746677 0.746673 9.99958 2.98024e-06 1.19209e-05 0.130576 0.977852 0.929716 -0.0132934 4.89293e-06 0.500586 -1.86952e-20 6.88117e-24 -1.86883e-20 0.00139502 0.997818 8.59217e-05 0.152539 2.85163 0.00139502 0.99793 0.669638 0.00104367 0.00187952 0.000859217 0.45567 0.00187952 0.434991 0.000127362 1.02 0.88737 0.534768 0.285623 1.71606e-07 3.0552e-09 2392.46 3176.09 -0.059333 0.482113 0.277645 0.257057 -0.592675 -0.16949 0.485443 -0.268497 -0.216953 1.356 1 3.53461e-295 293.74 2.11149e-292 2.03383 1.354 0.00029997 0.879629 0.637355 0.48988 0.400917 2.03411 128.396 83.2266 18.6806 60.5315 0.00405408 0 -40 10
0.455 1.31905e-08 2.53884e-06 0.0715305 0.071524 0.012044 5.99567e-06 0.00115402 0.0894131 0.000656314 0.0900648 0.856443 101.882 0.246325 0.713172 4.11782 0.0536751 0.0388474 0.961153 0.0198804 0.00423667 0.0191428 0.00407899 0.00511957 0.00585722 0.204783 0.234289 57.9672 -87.8943 126.002 15.984 145.009 0.000143925 0.267075 192.933 0.31073 0.067391 0.00409467 0.000561539 0.00138238 0.986994 0.991736 -2.97127e-06 -85.6688 0.0929758 31197.2 300.376 0.983523 0.319147 0.74661 0.746605 9.99958 2.98025e-06 1.19209e-05 0.130577 0.97787 0.929724 -0.0132934 4.89295e-06 0.50059 -1.8696e-20 6.88152e-24 -1.86892e-20 0.00139502 0.997818 8.59217e-05 0.152539 2.85163 0.00139502 0.997929 0.669753 0.00104369 0.00187952 0.000859217 0.45567 0.00187952 0.435001 0.000127366 1.02 0.887371 0.534767 0.285624 1.71607e-07 3.05522e-09 2392.45 3175.8 -0.0593124 0.482113 0.277645 0.257038 -0.592679 -0.169491 0.485504 -0.268495 -0.217015 1.357 1 2.14385e-295 293.76 1.28089e-292 2.03403 1.355 0.00029997 0.879501 0.637416 0.489462 0.40095 2.03431 128.406 83.2299 18.6807 60.5331 0.00405394 0 -40 10
0.456 1.32194e-08 2.53884e-06 0.0716242 0.0716178 0.012044 6.00884e-06 0.00115402 0.0895303 0.00065632 0.090182 0.856488 101.882 0.24632 0.713235 4.1179 0.0536801 0.0388481 0.961152 0.0198803 0.00423675 0.0191427 0.00407905 0.00511967 0.00585731 0.204787 0.234293 57.9673 -87.8943 126.003 15.984 145.009 0.000143912 0.267076 192.933 0.310729 0.067391 0.00409468 0.000561539 0.00138238 0.986994 0.991736 -2.97128e-06 -85.6688 0.0929759 31197.2 300.378 0.983523 0.319147 0.746542 0.746538 9.99958 2.98025e-06 1.19209e-05 0.130577 0.977887 0.929733 -0.0132934 4.89297e-06 0.500593 -1.86969e-20 6.88186e-24 -1.869e-20 0.00139502 0.997818 8.59218e-05 0.152539 2.85163 0.00139502 0.997928 0.669868 0.00104371 0.00187952 0.000859218 0.45567 0.00187952 0.435011 0.00012737 1.02 0.887371 0.534767 0.285625 1.71607e-07 3.05524e-09 2392.43 3175.51 -0.059292 0.482113 0.277645 0.257021 -0.592682 -0.169491 0.485564 -0.268493 -0.217078 1.358 1 1.30031e-295 293.781 7.7703e-293 2.03422 1.356 0.00029997 0.879372 0.637477 0.489045 0.400983 2.0345 128.417 83.2332 18.6809 60.5347 0.0040538 0 -40 10
0.457 1.32484e-08 2.53884e-06 0.0717179 0.0717115 0.012044 6.02201e-06 0.00115402 0.0896474 0.000656326 0.0902991 0.856532 101.882 0.246315 0.713297 4.11798 0.053685 0.0388488 0.961151 0.0198802 0.00423683 0.0191426 0.00407912 0.00511976 0.00585741 0.204791 0.234296 57.9673 -87.8943 126.005 15.9839 145.009 0.000143899 0.267076 192.933 0.310729 0.067391 0.00409468 0.00056154 0.00138238 0.986994 0.991736 -2.97129e-06 -85.6688 0.0929759 31197.2 300.381 0.983523 0.319147 0.746475 0.746471 9.99958 2.98025e-06 1.19209e-05 0.130578 0.977905 0.929742 -0.0132934 4.893e-06 0.500596 -1.86977e-20 6.8822e-24 -1.86908e-20 0.00139502 0.997818 8.59218e-05 0.152539 2.85163 0.00139502 0.997928 0.669983 0.00104373 0.00187952 0.000859218 0.45567 0.00187952 0.43502 0.000127373 1.02 0.887372 0.534767 0.285626 1.71607e-07 3.05525e-09 2392.41 3175.23 -0.0592716 0.482113 0.277644 0.257003 -0.592685 -0.169491 0.485624 -0.268491 -0.21714 1.359 1 7.88678e-296 293.801 4.7137e-293 2.03442 1.357 0.000299969 0.879245 0.637539 0.488629 0.401016 2.0347 128.427 83.2365 18.6811 60.5363 0.00405367 0 -40 10
0.458 1.32774e-08 2.53884e-06 0.0718115 0.0718051 0.0120439 6.03517e-06 0.00115402 0.0897644 0.000656333 0.0904161 0.856577 101.882 0.24631 0.71336 4.11806 0.05369 0.0388496 0.96115 0.0198801 0.00423691 0.0191425 0.00407918 0.00511986 0.00585751 0.204794 0.2343 57.9674 -87.8943 126.006 15.9839 145.009 0.000143886 0.267076 192.933 0.310729 0.0673909 0.00409468 0.00056154 0.00138238 0.986994 0.991736 -2.9713e-06 -85.6688 0.092976 31197.2 300.383 0.983523 0.319147 0.746408 0.746404 9.99958 2.98026e-06 1.19209e-05 0.130579 0.977923 0.92975 -0.0132934 4.89302e-06 0.5006 -1.86985e-20 6.88254e-24 -1.86917e-20 0.00139502 0.997818 8.59219e-05 0.152539 2.85164 0.00139502 0.997927 0.670098 0.00104375 0.00187952 0.000859219 0.45567 0.00187952 0.43503 0.000127377 1.02 0.887373 0.534767 0.285627 1.71607e-07 3.05527e-09 2392.4 3174.94 -0.0592513 0.482113 0.277644 0.256985 -0.592689 -0.169491 0.485684 -0.268489 -0.217202 1.36 1 4.78357e-296 293.821 2.85948e-293 2.03462 1.358 0.000299969 0.879118 0.6376 0.488214 0.40105 2.03489 128.438 83.2397 18.6813 60.5378 0.00405353 0 -40 10
0.459 1.33064e-08 2.53884e-06 0.071905 0.0718986 0.0120439 6.04834e-06 0.00115402 0.0898813 0.000656339 0.090533 0.856621 101.882 0.246305 0.713423 4.11813 0.053695 0.0388503 0.96115 0.01988 0.00423699 0.0191424 0.00407925 0.00511996 0.0058576 0.204798 0.234304 57.9675 -87.8943 126.007 15.9839 145.009 0.000143873 0.267076 192.933 0.310728 0.0673909 0.00409468 0.00056154 0.00138238 0.986994 0.991736 -2.97131e-06 -85.6688 0.092976 31197.2 300.385 0.983523 0.319147 0.746342 0.746337 9.99958 2.98026e-06 1.19209e-05 0.13058 0.97794 0.929759 -0.0132934 4.89304e-06 0.500603 -1.86994e-20 6.88288e-24 -1.86925e-20 0.00139502 0.997818 8.5922e-05 0.15254 2.85164 0.00139502 0.997926 0.670213 0.00104377 0.00187953 0.00085922 0.45567 0.00187952 0.43504 0.00012738 1.02 0.887374 0.534766 0.285629 1.71607e-07 3.05529e-09 2392.38 3174.66 -0.0592311 0.482114 0.277644 0.256967 -0.592692 -0.169491 0.485744 -0.268488 -0.217263 1.361 1 2.90138e-296 293.841 1.73465e-293 2.03481 1.359 0.000299969 0.878991 0.637661 0.487801 0.401083 2.03509 128.448 83.243 18.6815 60.5394 0.00405339 0 -40 10
0.46 1.33353e-08 2.53884e-06 0.0719985 0.0719921 0.0120439 6.06151e-06 0.00115402 0.0899981 0.000656346 0.0906498 0.856666 101.882 0.2463 0.713485 4.11821 0.0537 0.0388511 0.961149 0.0198799 0.00423707 0.0191423 0.00407932 0.00512006 0.0058577 0.204802 0.234308 57.9675 -87.8943 126.008 15.9838 145.009 0.00014386 0.267076 192.933 0.310728 0.0673909 0.00409469 0.000561541 0.00138238 0.986994 0.991736 -2.97132e-06 -85.6688 0.0929761 31197.2 300.387 0.983523 0.319147 0.746276 0.746271 9.99958 2.98026e-06 1.1921e-05 0.130581 0.977958 0.929767 -0.0132934 4.89307e-06 0.500606 -1.87002e-20 6.88322e-24 -1.86933e-20 0.00139502 0.997818 8.5922e-05 0.15254 2.85164 0.00139502 0.997925 0.670327 0.00104379 0.00187953 0.00085922 0.455669 0.00187953 0.43505 0.000127384 1.02 0.887375 0.534766 0.28563 1.71607e-07 3.05531e-09 2392.36 3174.37 -0.0592109 0.482114 0.277643 0.256949 -0.592695 -0.169491 0.485804 -0.268486 -0.217324 1.362 1 1.75978e-296 293.861 1.05229e-293 2.03501 1.36 0.000299969 0.878865 0.637723 0.487388 0.401116 2.03528 128.459 83.2462 18.6817 60.541 0.00405326 0 -40 10
0.461 1.33643e-08 2.53884e-06 0.0720918 0.0720855 0.0120439 6.07468e-06 0.00115402 0.0901148 0.000656352 0.0907665 0.856711 101.882 0.246295 0.713548 4.11829 0.053705 0.0388518 0.961148 0.0198798 0.00423715 0.0191422 0.00407938 0.00512016 0.0058578 0.204806 0.234312 57.9676 -87.8943 126.009 15.9838 145.009 0.000143848 0.267076 192.933 0.310728 0.0673908 0.00409469 0.000561541 0.00138238 0.986994 0.991736 -2.97133e-06 -85.6688 0.0929762 31197.1 300.389 0.983523 0.319147 0.746209 0.746205 9.99958 2.98027e-06 1.1921e-05 0.130582 0.977975 0.929775 -0.0132934 4.89309e-06 0.500609 -1.8701e-20 6.88356e-24 -1.86942e-20 0.00139502 0.997818 8.59221e-05 0.15254 2.85164 0.00139502 0.997925 0.670442 0.0010438 0.00187953 0.000859221 0.455669 0.00187953 0.43506 0.000127387 1.02 0.887376 0.534766 0.285631 1.71608e-07 3.05532e-09 2392.35 3174.09 -0.0591908 0.482114 0.277643 0.256932 -0.592699 -0.169491 0.485863 -0.268484 -0.217386 1.363 1 1.06736e-296 293.881 6.38349e-294 2.0352 1.361 0.000299969 0.878739 0.637784 0.486977 0.401149 2.03548 128.469 83.2494 18.6819 60.5425 0.00405312 0 -40 10
0.462 1.33933e-08 2.53884e-06 0.0721851 0.0721788 0.0120439 6.08784e-06 0.00115402 0.0902314 0.000656358 0.0908832 0.856756 101.882 0.24629 0.713611 4.11837 0.05371 0.0388526 0.961147 0.0198797 0.00423723 0.0191421 0.00407945 0.00512026 0.0058579 0.20481 0.234316 57.9676 -87.8943 126.011 15.9837 145.009 0.000143835 0.267076 192.933 0.310727 0.0673908 0.00409469 0.000561542 0.00138239 0.986994 0.991736 -2.97134e-06 -85.6688 0.0929762 31197.1 300.392 0.983523 0.319147 0.746144 0.746139 9.99958 2.98027e-06 1.1921e-05 0.130582 0.977992 0.929784 -0.0132934 4.89311e-06 0.500613 -1.87019e-20 6.8839e-24 -1.8695e-20 0.00139503 0.997818 8.59221e-05 0.15254 2.85164 0.00139503 0.997924 0.670557 0.00104382 0.00187953 0.000859221 0.455669 0.00187953 0.43507 0.000127391 1.02 0.887377 0.534766 0.285632 1.71608e-07 3.05534e-09 2392.33 3173.81 -0.0591708 0.482114 0.277643 0.256914 -0.592702 -0.169491 0.485922 -0.268482 -0.217446 1.364 1 6.47386e-297 293.9 3.87242e-294 2.0354 1.362 0.000299969 0.878613 0.637845 0.486567 0.401182 2.03568 128.48 83.2527 18.6821 60.5441 0.00405299 0 -40 10
0.463 1.34222e-08 2.53884e-06 0.0722783 0.072272 0.0120439 6.10101e-06 0.00115402 0.0903479 0.000656365 0.0909997 0.856801 101.882 0.246285 0.713675 4.11845 0.053715 0.0388533 0.961147 0.0198796 0.00423731 0.019142 0.00407952 0.00512036 0.00585799 0.204814 0.23432 57.9677 -87.8943 126.012 15.9837 145.01 0.000143822 0.267077 192.932 0.310727 0.0673907 0.00409469 0.000561542 0.00138239 0.986994 0.991736 -2.97136e-06 -85.6688 0.0929763 31197.1 300.394 0.983523 0.319147 0.746078 0.746074 9.99958 2.98028e-06 1.1921e-05 0.130583 0.97801 0.929792 -0.0132934 4.89314e-06 0.500616 -1.87027e-20 6.88424e-24 -1.86958e-20 0.00139503 0.997818 8.59222e-05 0.15254 2.85164 0.00139503 0.997923 0.670672 0.00104384 0.00187953 0.000859222 0.455669 0.00187953 0.435079 0.000127394 1.02 0.887378 0.534765 0.285633 1.71608e-07 3.05536e-09 2392.32 3173.53 -0.0591509 0.482114 0.277642 0.256896 -0.592705 -0.169491 0.485981 -0.26848 -0.217507 1.365 1 3.92659e-297 293.92 2.34912e-294 2.03559 1.363 0.000299969 0.878489 0.637906 0.486157 0.401215 2.03587 128.49 83.2559 18.6823 60.5456 0.00405286 0 -40 10
0.464 1.34512e-08 2.53884e-06 0.0723715 0.0723652 0.0120439 6.11418e-06 0.00115402 0.0904643 0.000656371 0.0911161 0.856846 101.881 0.24628 0.713738 4.11853 0.05372 0.0388541 0.961146 0.0198795 0.00423739 0.0191419 0.00407958 0.00512046 0.00585809 0.204818 0.234324 57.9678 -87.8943 126.013 15.9837 145.01 0.00014381 0.267077 192.932 0.310727 0.0673907 0.00409469 0.000561543 0.00138239 0.986994 0.991736 -2.97137e-06 -85.6687 0.0929763 31197.1 300.396 0.983523 0.319147 0.746013 0.746008 9.99958 2.98028e-06 1.1921e-05 0.130584 0.978027 0.929801 -0.0132934 4.89316e-06 0.50062 -1.87035e-20 6.88458e-24 -1.86967e-20 0.00139503 0.997818 8.59222e-05 0.15254 2.85164 0.00139503 0.997923 0.670786 0.00104386 0.00187953 0.000859222 0.455669 0.00187953 0.435089 0.000127398 1.02 0.887378 0.534765 0.285635 1.71608e-07 3.05538e-09 2392.3 3173.25 -0.0591311 0.482114 0.277642 0.256879 -0.592709 -0.169491 0.486039 -0.268478 -0.217567 1.366 1 2.3816e-297 293.94 1.42505e-294 2.03579 1.364 0.000299968 0.878364 0.637967 0.485749 0.401248 2.03606 128.5 83.2591 18.6824 60.5472 0.00405272 0 -40 10
0.465 1.34802e-08 2.53884e-06 0.0724645 0.0724583 0.0120439 6.12734e-06 0.00115402 0.0905807 0.000656377 0.0912325 0.856891 101.881 0.246275 0.713802 4.11862 0.053725 0.0388549 0.961145 0.0198794 0.00423748 0.0191418 0.00407965 0.00512056 0.00585819 0.204822 0.234328 57.9678 -87.8943 126.014 15.9836 145.01 0.000143797 0.267077 192.932 0.310726 0.0673907 0.0040947 0.000561543 0.00138239 0.986994 0.991736 -2.97138e-06 -85.6687 0.0929764 31197.1 300.398 0.983523 0.319147 0.745948 0.745943 9.99958 2.98028e-06 1.1921e-05 0.130585 0.978044 0.929809 -0.0132934 4.89318e-06 0.500623 -1.87044e-20 6.88491e-24 -1.86975e-20 0.00139503 0.997818 8.59223e-05 0.15254 2.85164 0.00139503 0.997922 0.670901 0.00104388 0.00187953 0.000859223 0.455669 0.00187953 0.435099 0.000127401 1.02 0.887379 0.534765 0.285636 1.71608e-07 3.05539e-09 2392.28 3172.98 -0.0591113 0.482114 0.277642 0.256861 -0.592712 -0.169491 0.486098 -0.268477 -0.217628 1.367 1 1.44451e-297 293.959 8.64475e-295 2.03598 1.365 0.000299968 0.87824 0.638028 0.485342 0.401281 2.03626 128.511 83.2622 18.6826 60.5487 0.00405259 0 -40 10
0.466 1.35091e-08 2.53884e-06 0.0725575 0.0725513 0.0120438 6.14051e-06 0.00115402 0.0906969 0.000656383 0.0913487 0.856936 101.881 0.24627 0.713865 4.1187 0.0537301 0.0388556 0.961144 0.0198793 0.00423756 0.0191417 0.00407972 0.00512066 0.00585829 0.204826 0.234332 57.9679 -87.8943 126.015 15.9836 145.01 0.000143785 0.267077 192.932 0.310726 0.0673906 0.0040947 0.000561544 0.00138239 0.986994 0.991736 -2.97139e-06 -85.6687 0.0929765 31197.1 300.4 0.983523 0.319147 0.745883 0.745878 9.99958 2.98029e-06 1.1921e-05 0.130586 0.978061 0.929817 -0.0132934 4.89321e-06 0.500626 -1.87052e-20 6.88525e-24 -1.86983e-20 0.00139503 0.997818 8.59224e-05 0.15254 2.85164 0.00139503 0.997921 0.671016 0.0010439 0.00187953 0.000859224 0.455669 0.00187953 0.435109 0.000127405 1.02 0.88738 0.534765 0.285637 1.71609e-07 3.05541e-09 2392.27 3172.7 -0.0590916 0.482114 0.277642 0.256844 -0.592715 -0.169491 0.486156 -0.268475 -0.217688 1.368 1 8.76142e-298 293.979 5.24415e-295 2.03618 1.366 0.000299968 0.878117 0.638089 0.484937 0.401314 2.03645 128.521 83.2654 18.6828 60.5503 0.00405246 0 -40 10
0.467 1.35381e-08 2.53884e-06 0.0726505 0.0726443 0.0120438 6.15368e-06 0.00115402 0.0908131 0.00065639 0.0914649 0.856981 101.881 0.246265 0.713929 4.11878 0.0537351 0.0388564 0.961144 0.0198792 0.00423764 0.0191416 0.00407979 0.00512076 0.00585839 0.20483 0.234336 57.968 -87.8943 126.016 15.9836 145.01 0.000143772 0.267077 192.932 0.310726 0.0673906 0.0040947 0.000561544 0.00138239 0.986994 0.991736 -2.9714e-06 -85.6687 0.0929765 31197.1 300.403 0.983523 0.319147 0.745818 0.745814 9.99958 2.98029e-06 1.19211e-05 0.130587 0.978078 0.929825 -0.0132934 4.89323e-06 0.50063 -1.8706e-20 6.88559e-24 -1.86991e-20 0.00139503 0.997818 8.59224e-05 0.15254 2.85164 0.00139503 0.997921 0.67113 0.00104392 0.00187953 0.000859224 0.455668 0.00187953 0.435119 0.000127408 1.02 0.887381 0.534764 0.285638 1.71609e-07 3.05543e-09 2392.25 3172.42 -0.059072 0.482114 0.277641 0.256827 -0.592718 -0.169491 0.486214 -0.268473 -0.217747 1.369 1 5.31407e-298 293.998 3.18125e-295 2.03637 1.367 0.000299968 0.877994 0.63815 0.484532 0.401347 2.03665 128.532 83.2686 18.683 60.5518 0.00405232 0 -40 10
0.468 1.35671e-08 2.53884e-06 0.0727433 0.0727371 0.0120438 6.16684e-06 0.00115402 0.0909291 0.000656396 0.0915809 0.857026 101.881 0.24626 0.713993 4.11886 0.0537402 0.0388572 0.961143 0.0198791 0.00423772 0.0191415 0.00407986 0.00512086 0.00585849 0.204835 0.23434 57.968 -87.8943 126.018 15.9835 145.01 0.00014376 0.267077 192.932 0.310726 0.0673906 0.0040947 0.000561545 0.0013824 0.986994 0.991736 -2.97141e-06 -85.6687 0.0929766 31197 300.405 0.983523 0.319147 0.745754 0.745749 9.99958 2.98029e-06 1.19211e-05 0.130587 0.978095 0.929834 -0.0132934 4.89326e-06 0.500633 -1.87069e-20 6.88593e-24 -1.87e-20 0.00139503 0.997818 8.59225e-05 0.152541 2.85164 0.00139503 0.99792 0.671245 0.00104394 0.00187954 0.000859225 0.455668 0.00187953 0.435128 0.000127412 1.02 0.887382 0.534764 0.28564 1.71609e-07 3.05545e-09 2392.23 3172.15 -0.0590525 0.482114 0.277641 0.25681 -0.592721 -0.169491 0.486271 -0.268471 -0.217807 1.37 1 3.22315e-298 294.018 1.92984e-295 2.03657 1.368 0.000299968 0.877871 0.638211 0.484128 0.40138 2.03684 128.542 83.2717 18.6832 60.5533 0.00405219 0 -40 10
0.469 1.3596e-08 2.53884e-06 0.0728361 0.0728299 0.0120438 6.18001e-06 0.00115402 0.0910451 0.000656402 0.0916969 0.857071 101.881 0.246255 0.714057 4.11894 0.0537453 0.0388579 0.961142 0.019879 0.00423781 0.0191414 0.00407992 0.00512097 0.00585859 0.204839 0.234344 57.9681 -87.8943 126.019 15.9835 145.01 0.000143747 0.267077 192.932 0.310725 0.0673905 0.00409471 0.000561545 0.0013824 0.986994 0.991736 -2.97142e-06 -85.6687 0.0929767 31197 300.407 0.983523 0.319147 0.745689 0.745685 9.99958 2.9803e-06 1.19211e-05 0.130588 0.978112 0.929842 -0.0132934 4.89328e-06 0.500637 -1.87077e-20 6.88627e-24 -1.87008e-20 0.00139503 0.997818 8.59225e-05 0.152541 2.85164 0.00139503 0.997919 0.671359 0.00104396 0.00187954 0.000859225 0.455668 0.00187954 0.435138 0.000127416 1.02 0.887383 0.534764 0.285641 1.71609e-07 3.05547e-09 2392.22 3171.88 -0.059033 0.482114 0.277641 0.256792 -0.592725 -0.169491 0.486329 -0.268469 -0.217866 1.371 1 1.95494e-298 294.037 1.1707e-295 2.03676 1.369 0.000299968 0.877749 0.638271 0.483726 0.401413 2.03704 128.552 83.2749 18.6834 60.5548 0.00405206 0 -40 10
0.47 1.3625e-08 2.53884e-06 0.0729288 0.0729226 0.0120438 6.19318e-06 0.00115402 0.091161 0.000656408 0.0918128 0.857117 101.881 0.24625 0.714121 4.11903 0.0537503 0.0388587 0.961141 0.0198789 0.00423789 0.0191413 0.00407999 0.00512107 0.00585869 0.204843 0.234348 57.9681 -87.8943 126.02 15.9834 145.01 0.000143735 0.267077 192.932 0.310725 0.0673905 0.00409471 0.000561546 0.0013824 0.986994 0.991736 -2.97143e-06 -85.6687 0.0929767 31197 300.409 0.983523 0.319147 0.745625 0.745621 9.99958 2.9803e-06 1.19211e-05 0.130589 0.978129 0.92985 -0.0132934 4.8933e-06 0.50064 -1.87085e-20 6.88661e-24 -1.87016e-20 0.00139503 0.997818 8.59226e-05 0.152541 2.85164 0.00139503 0.997919 0.671474 0.00104398 0.00187954 0.000859226 0.455668 0.00187954 0.435148 0.000127419 1.02 0.887384 0.534764 0.285642 1.71609e-07 3.05548e-09 2392.2 3171.6 -0.0590136 0.482114 0.27764 0.256775 -0.592728 -0.169491 0.486386 -0.268468 -0.217925 1.372 1 1.18573e-298 294.056 7.10177e-296 2.03695 1.37 0.000299967 0.877627 0.638332 0.483324 0.401446 2.03723 128.563 83.278 18.6836 60.5563 0.00405193 0 -40 10
0.471 1.3654e-08 2.53884e-06 0.0730214 0.0730153 0.0120438 6.20635e-06 0.00115402 0.0912768 0.000656414 0.0919286 0.857162 101.881 0.246245 0.714185 4.11911 0.0537554 0.0388595 0.96114 0.0198788 0.00423797 0.0191412 0.00408006 0.00512117 0.00585879 0.204847 0.234352 57.9682 -87.8943 126.021 15.9834 145.01 0.000143723 0.267078 192.931 0.310725 0.0673904 0.00409471 0.000561546 0.0013824 0.986994 0.991736 -2.97144e-06 -85.6687 0.0929768 31197 300.412 0.983523 0.319147 0.745562 0.745557 9.99958 2.9803e-06 1.19211e-05 0.13059 0.978146 0.929858 -0.0132934 4.89333e-06 0.500644 -1.87093e-20 6.88695e-24 -1.87025e-20 0.00139503 0.997818 8.59226e-05 0.152541 2.85164 0.00139503 0.997918 0.671588 0.001044 0.00187954 0.000859226 0.455668 0.00187954 0.435158 0.000127423 1.02 0.887385 0.534763 0.285643 1.7161e-07 3.0555e-09 2392.18 3171.33 -0.0589943 0.482114 0.27764 0.256758 -0.592731 -0.169492 0.486443 -0.268466 -0.217984 1.373 1 7.19181e-299 294.075 4.30813e-296 2.03715 1.371 0.000299967 0.877506 0.638393 0.482924 0.401479 2.03742 128.573 83.2811 18.6837 60.5578 0.0040518 0 -40 10
0.472 1.36829e-08 2.53884e-06 0.0731139 0.0731079 0.0120438 6.21951e-06 0.00115402 0.0913924 0.00065642 0.0920443 0.857208 101.881 0.246239 0.714249 4.11919 0.0537605 0.0388603 0.96114 0.0198787 0.00423806 0.0191411 0.00408013 0.00512127 0.00585889 0.204851 0.234356 57.9683 -87.8943 126.022 15.9834 145.01 0.00014371 0.267078 192.931 0.310724 0.0673904 0.00409471 0.000561547 0.0013824 0.986994 0.991736 -2.97146e-06 -85.6687 0.0929769 31197 300.414 0.983523 0.319147 0.745498 0.745494 9.99958 2.98031e-06 1.19211e-05 0.130591 0.978163 0.929866 -0.0132934 4.89335e-06 0.500647 -1.87102e-20 6.88729e-24 -1.87033e-20 0.00139503 0.997818 8.59227e-05 0.152541 2.85164 0.00139503 0.997917 0.671703 0.00104401 0.00187954 0.000859227 0.455668 0.00187954 0.435167 0.000127426 1.02 0.887385 0.534763 0.285644 1.7161e-07 3.05552e-09 2392.17 3171.06 -0.0589751 0.482114 0.27764 0.256741 -0.592734 -0.169492 0.4865 -0.268464 -0.218043 1.374 1 4.36205e-299 294.094 2.61343e-296 2.03734 1.372 0.000299967 0.877385 0.638453 0.482524 0.401512 2.03762 128.584 83.2842 18.6839 60.5593 0.00405167 0 -40 10
0.473 1.37119e-08 2.53884e-06 0.0732064 0.0732003 0.0120437 6.23268e-06 0.00115402 0.091508 0.000656426 0.0921599 0.857253 101.881 0.246234 0.714313 4.11927 0.0537656 0.0388611 0.961139 0.0198786 0.00423814 0.019141 0.0040802 0.00512138 0.005859 0.204855 0.23436 57.9683 -87.8943 126.023 15.9833 145.01 0.000143698 0.267078 192.931 0.310724 0.0673904 0.00409471 0.000561547 0.0013824 0.986993 0.991736 -2.97147e-06 -85.6687 0.0929769 31197 300.416 0.983523 0.319147 0.745435 0.74543 9.99958 2.98031e-06 1.19211e-05 0.130592 0.97818 0.929874 -0.0132934 4.89338e-06 0.500651 -1.8711e-20 6.88763e-24 -1.87041e-20 0.00139503 0.997818 8.59228e-05 0.152541 2.85165 0.00139503 0.997917 0.671817 0.00104403 0.00187954 0.000859228 0.455667 0.00187954 0.435177 0.00012743 1.02 0.887386 0.534763 0.285646 1.7161e-07 3.05554e-09 2392.15 3170.79 -0.0589559 0.482114 0.27764 0.256724 -0.592737 -0.169492 0.486556 -0.268462 -0.218101 1.375 1 2.64572e-299 294.113 1.58538e-296 2.03754 1.373 0.000299967 0.877265 0.638514 0.482126 0.401544 2.03781 128.594 83.2873 18.6841 60.5608 0.00405154 0 -40 10
0.474 1.37409e-08 2.53884e-06 0.0732988 0.0732928 0.0120437 6.24585e-06 0.00115402 0.0916235 0.000656432 0.0922754 0.857299 101.881 0.246229 0.714378 4.11936 0.0537708 0.0388619 0.961138 0.0198785 0.00423823 0.0191409 0.00408027 0.00512148 0.0058591 0.204859 0.234364 57.9684 -87.8943 126.024 15.9833 145.01 0.000143686 0.267078 192.931 0.310724 0.0673903 0.00409472 0.000561548 0.0013824 0.986993 0.991736 -2.97148e-06 -85.6687 0.092977 31196.9 300.419 0.983523 0.319147 0.745372 0.745367 9.99958 2.98031e-06 1.19212e-05 0.130593 0.978196 0.929882 -0.0132934 4.8934e-06 0.500654 -1.87118e-20 6.88796e-24 -1.87049e-20 0.00139504 0.997818 8.59228e-05 0.152541 2.85165 0.00139504 0.997916 0.671931 0.00104405 0.00187954 0.000859228 0.455667 0.00187954 0.435187 0.000127433 1.02 0.887387 0.534763 0.285647 1.7161e-07 3.05556e-09 2392.13 3170.52 -0.0589368 0.482114 0.277639 0.256707 -0.59274 -0.169492 0.486613 -0.26846 -0.218159 1.376 1 1.60471e-299 294.132 9.61734e-297 2.03773 1.374 0.000299967 0.877145 0.638575 0.481729 0.401577 2.038 128.604 83.2904 18.6843 60.5623 0.00405141 0 -40 10
0.475 1.37698e-08 2.53884e-06 0.0733911 0.0733851 0.0120437 6.25901e-06 0.00115402 0.0917389 0.000656438 0.0923908 0.857345 101.881 0.246224 0.714443 4.11944 0.0537759 0.0388627 0.961137 0.0198784 0.00423831 0.0191408 0.00408034 0.00512159 0.0058592 0.204863 0.234368 57.9685 -87.8943 126.025 15.9833 145.01 0.000143674 0.267078 192.931 0.310723 0.0673903 0.00409472 0.000561548 0.00138241 0.986993 0.991736 -2.97149e-06 -85.6687 0.092977 31196.9 300.421 0.983523 0.319147 0.745309 0.745305 9.99958 2.98032e-06 1.19212e-05 0.130593 0.978213 0.92989 -0.0132934 4.89342e-06 0.500658 -1.87126e-20 6.8883e-24 -1.87058e-20 0.00139504 0.997818 8.59229e-05 0.152541 2.85165 0.00139504 0.997915 0.672046 0.00104407 0.00187954 0.000859229 0.455667 0.00187954 0.435197 0.000127437 1.02 0.887388 0.534762 0.285648 1.7161e-07 3.05557e-09 2392.12 3170.25 -0.0589178 0.482114 0.277639 0.256691 -0.592744 -0.169492 0.486669 -0.268458 -0.218217 1.377 1 9.73306e-300 294.151 5.83414e-297 2.03792 1.375 0.000299967 0.877025 0.638635 0.481333 0.40161 2.0382 128.615 83.2935 18.6845 60.5638 0.00405129 0 -40 10
0.476 1.37988e-08 2.53884e-06 0.0734834 0.0734774 0.0120437 6.27218e-06 0.00115402 0.0918543 0.000656444 0.0925061 0.85739 101.88 0.246219 0.714507 4.11953 0.053781 0.0388635 0.961137 0.0198783 0.0042384 0.0191407 0.00408041 0.00512169 0.0058593 0.204868 0.234372 57.9685 -87.8943 126.027 15.9832 145.01 0.000143662 0.267078 192.931 0.310723 0.0673902 0.00409472 0.000561549 0.00138241 0.986993 0.991736 -2.9715e-06 -85.6687 0.0929771 31196.9 300.423 0.983523 0.319147 0.745246 0.745242 9.99958 2.98032e-06 1.19212e-05 0.130594 0.97823 0.929898 -0.0132934 4.89345e-06 0.500661 -1.87135e-20 6.88864e-24 -1.87066e-20 0.00139504 0.997818 8.59229e-05 0.152541 2.85165 0.00139504 0.997915 0.67216 0.00104409 0.00187954 0.000859229 0.455667 0.00187954 0.435206 0.00012744 1.02 0.887389 0.534762 0.285649 1.71611e-07 3.05559e-09 2392.1 3169.99 -0.0588988 0.482114 0.277639 0.256674 -0.592747 -0.169492 0.486725 -0.268457 -0.218275 1.378 1 5.9034e-300 294.17 3.53915e-297 2.03812 1.376 0.000299966 0.876906 0.638696 0.480938 0.401643 2.03839 128.625 83.2965 18.6846 60.5653 0.00405116 0 -40 10
0.477 1.38278e-08 2.53884e-06 0.0735756 0.0735696 0.0120437 6.28534e-06 0.00115402 0.0919695 0.00065645 0.0926213 0.857436 101.88 0.246214 0.714572 4.11961 0.0537862 0.0388643 0.961136 0.0198782 0.00423848 0.0191406 0.00408048 0.0051218 0.00585941 0.204872 0.234376 57.9686 -87.8943 126.028 15.9832 145.01 0.00014365 0.267078 192.931 0.310723 0.0673902 0.00409472 0.000561549 0.00138241 0.986993 0.991736 -2.97151e-06 -85.6687 0.0929772 31196.9 300.425 0.983523 0.319147 0.745184 0.74518 9.99958 2.98033e-06 1.19212e-05 0.130595 0.978246 0.929906 -0.0132934 4.89347e-06 0.500665 -1.87143e-20 6.88898e-24 -1.87074e-20 0.00139504 0.997818 8.5923e-05 0.152542 2.85165 0.00139504 0.997914 0.672274 0.00104411 0.00187955 0.00085923 0.455667 0.00187954 0.435216 0.000127444 1.02 0.88739 0.534762 0.285651 1.71611e-07 3.05561e-09 2392.08 3169.72 -0.05888 0.482115 0.277638 0.256657 -0.59275 -0.169492 0.48678 -0.268455 -0.218333 1.379 1 3.58059e-300 294.189 2.14694e-297 2.03831 1.377 0.000299966 0.876788 0.638756 0.480544 0.401675 2.03858 128.635 83.2996 18.6848 60.5668 0.00405103 0 -40 10
0.478 1.38567e-08 2.53884e-06 0.0736677 0.0736617 0.0120437 6.29851e-06 0.00115402 0.0920846 0.000656456 0.0927365 0.857482 101.88 0.246209 0.714637 4.1197 0.0537913 0.0388651 0.961135 0.0198781 0.00423857 0.0191405 0.00408055 0.0051219 0.00585951 0.204876 0.23438 57.9686 -87.8943 126.029 15.9832 145.01 0.000143638 0.267079 192.931 0.310722 0.0673902 0.00409472 0.00056155 0.00138241 0.986993 0.991736 -2.97152e-06 -85.6687 0.0929772 31196.9 300.428 0.983523 0.319147 0.745122 0.745117 9.99958 2.98033e-06 1.19212e-05 0.130596 0.978263 0.929914 -0.0132934 4.8935e-06 0.500668 -1.87151e-20 6.88932e-24 -1.87082e-20 0.00139504 0.997818 8.59231e-05 0.152542 2.85165 0.00139504 0.997914 0.672388 0.00104413 0.00187955 0.000859231 0.455667 0.00187955 0.435226 0.000127447 1.02 0.887391 0.534762 0.285652 1.71611e-07 3.05563e-09 2392.07 3169.46 -0.0588612 0.482115 0.277638 0.256641 -0.592753 -0.169492 0.486836 -0.268453 -0.21839 1.38 1 2.17174e-300 294.207 1.30239e-297 2.0385 1.378 0.000299966 0.876669 0.638816 0.480151 0.401708 2.03878 128.646 83.3026 18.685 60.5682 0.0040509 0 -40 10
0.479 1.38857e-08 2.53884e-06 0.0737597 0.0737538 0.0120437 6.31168e-06 0.00115402 0.0921996 0.000656462 0.0928515 0.857528 101.88 0.246204 0.714702 4.11978 0.0537965 0.0388659 0.961134 0.019878 0.00423865 0.0191404 0.00408062 0.00512201 0.00585961 0.20488 0.234385 57.9687 -87.8943 126.03 15.9831 145.01 0.000143626 0.267079 192.93 0.310722 0.0673901 0.00409473 0.00056155 0.00138241 0.986993 0.991736 -2.97153e-06 -85.6686 0.0929773 31196.9 300.43 0.983523 0.319147 0.74506 0.745056 9.99958 2.98033e-06 1.19212e-05 0.130597 0.978279 0.929922 -0.0132934 4.89352e-06 0.500672 -1.87159e-20 6.88965e-24 -1.8709e-20 0.00139504 0.997818 8.59231e-05 0.152542 2.85165 0.00139504 0.997913 0.672502 0.00104415 0.00187955 0.000859231 0.455666 0.00187955 0.435236 0.000127451 1.02 0.887392 0.534761 0.285653 1.71611e-07 3.05565e-09 2392.05 3169.19 -0.0588424 0.482115 0.277638 0.256624 -0.592756 -0.169492 0.486891 -0.268451 -0.218447 1.381 1 1.31723e-300 294.226 7.90065e-298 2.0387 1.379 0.000299966 0.876552 0.638877 0.479759 0.401741 2.03897 128.656 83.3057 18.6852 60.5697 0.00405078 0 -40 10
0.48 1.39147e-08 2.53884e-06 0.0738517 0.0738457 0.0120437 6.32484e-06 0.00115402 0.0923146 0.000656468 0.0929665 0.857574 101.88 0.246198 0.714768 4.11987 0.0538017 0.0388667 0.961133 0.0198779 0.00423874 0.0191403 0.00408069 0.00512211 0.00585972 0.204884 0.234389 57.9688 -87.8944 126.031 15.9831 145.01 0.000143614 0.267079 192.93 0.310722 0.0673901 0.00409473 0.000561551 0.00138241 0.986993 0.991736 -2.97155e-06 -85.6686 0.0929774 31196.8 300.432 0.983523 0.319147 0.744998 0.744994 9.99958 2.98034e-06 1.19212e-05 0.130598 0.978296 0.92993 -0.0132934 4.89354e-06 0.500675 -1.87168e-20 6.88999e-24 -1.87099e-20 0.00139504 0.997818 8.59232e-05 0.152542 2.85165 0.00139504 0.997912 0.672616 0.00104417 0.00187955 0.000859232 0.455666 0.00187955 0.435245 0.000127455 1.02 0.887393 0.534761 0.285654 1.71611e-07 3.05567e-09 2392.03 3168.93 -0.0588238 0.482115 0.277638 0.256608 -0.592759 -0.169492 0.486946 -0.268449 -0.218504 1.382 1 7.98938e-301 294.244 4.79274e-298 2.03889 1.38 0.000299966 0.876434 0.638937 0.479368 0.401773 2.03916 128.666 83.3087 18.6853 60.5712 0.00405065 0 -40 10
0.481 1.39436e-08 2.53884e-06 0.0739436 0.0739376 0.0120436 6.33801e-06 0.00115402 0.0924294 0.000656474 0.0930813 0.85762 101.88 0.246193 0.714833 4.11995 0.0538069 0.0388675 0.961133 0.0198778 0.00423883 0.0191402 0.00408077 0.00512222 0.00585982 0.204889 0.234393 57.9688 -87.8944 126.032 15.983 145.01 0.000143602 0.267079 192.93 0.310721 0.0673901 0.00409473 0.000561551 0.00138242 0.986993 0.991736 -2.97156e-06 -85.6686 0.0929774 31196.8 300.435 0.983523 0.319147 0.744937 0.744932 9.99958 2.98034e-06 1.19213e-05 0.130599 0.978312 0.929938 -0.0132934 4.89357e-06 0.500679 -1.87176e-20 6.89033e-24 -1.87107e-20 0.00139504 0.997818 8.59232e-05 0.152542 2.85165 0.00139504 0.997912 0.67273 0.00104419 0.00187955 0.000859232 0.455666 0.00187955 0.435255 0.000127458 1.02 0.887394 0.534761 0.285656 1.71612e-07 3.05568e-09 2392.02 3168.67 -0.0588052 0.482115 0.277637 0.256591 -0.592762 -0.169492 0.487001 -0.268447 -0.218561 1.383 1 4.8458e-301 294.263 2.9074e-298 2.03908 1.381 0.000299966 0.876318 0.638997 0.478978 0.401806 2.03935 128.676 83.3117 18.6855 60.5726 0.00405053 0 -40 10
0.482 1.39726e-08 2.53884e-06 0.0740354 0.0740295 0.0120436 6.35118e-06 0.00115402 0.0925442 0.00065648 0.0931961 0.857667 101.88 0.246188 0.714898 4.12004 0.053812 0.0388683 0.961132 0.0198777 0.00423891 0.0191401 0.00408084 0.00512233 0.00585993 0.204893 0.234397 57.9689 -87.8944 126.033 15.983 145.01 0.00014359 0.267079 192.93 0.310721 0.06739 0.00409473 0.000561552 0.00138242 0.986993 0.991736 -2.97157e-06 -85.6686 0.0929775 31196.8 300.437 0.983523 0.319147 0.744876 0.744871 9.99958 2.98034e-06 1.19213e-05 0.1306 0.978328 0.929946 -0.0132934 4.89359e-06 0.500682 -1.87184e-20 6.89067e-24 -1.87115e-20 0.00139504 0.997818 8.59233e-05 0.152542 2.85165 0.00139504 0.997911 0.672844 0.00104421 0.00187955 0.000859233 0.455666 0.00187955 0.435265 0.000127462 1.02 0.887394 0.534761 0.285657 1.71612e-07 3.0557e-09 2392 3168.41 -0.0587867 0.482115 0.277637 0.256575 -0.592765 -0.169492 0.487056 -0.268445 -0.218617 1.384 1 2.93913e-301 294.281 1.7637e-298 2.03927 1.382 0.000299965 0.876201 0.639058 0.478589 0.401838 2.03955 128.687 83.3147 18.6857 60.5741 0.0040504 0 -40 10
0.483 1.40016e-08 2.53884e-06 0.0741271 0.0741212 0.0120436 6.36434e-06 0.00115402 0.0926589 0.000656486 0.0933108 0.857713 101.88 0.246183 0.714964 4.12013 0.0538172 0.0388691 0.961131 0.0198776 0.004239 0.01914 0.00408091 0.00512243 0.00586003 0.204897 0.234401 57.969 -87.8944 126.034 15.983 145.01 0.000143579 0.267079 192.93 0.310721 0.06739 0.00409474 0.000561552 0.00138242 0.986993 0.991736 -2.97158e-06 -85.6686 0.0929776 31196.8 300.439 0.983523 0.319147 0.744815 0.74481 9.99958 2.98035e-06 1.19213e-05 0.130601 0.978344 0.929954 -0.0132934 4.89362e-06 0.500686 -1.87192e-20 6.891e-24 -1.87123e-20 0.00139504 0.997818 8.59234e-05 0.152542 2.85165 0.00139504 0.99791 0.672958 0.00104423 0.00187955 0.000859234 0.455666 0.00187955 0.435274 0.000127465 1.02 0.887395 0.53476 0.285658 1.71612e-07 3.05572e-09 2391.99 3168.15 -0.0587683 0.482115 0.277637 0.256558 -0.592768 -0.169492 0.48711 -0.268444 -0.218673 1.385 1 1.78267e-301 294.299 1.06991e-298 2.03946 1.383 0.000299965 0.876085 0.639118 0.478201 0.401871 2.03974 128.697 83.3177 18.6859 60.5755 0.00405028 0 -40 10
0.484 1.40305e-08 2.53884e-06 0.0742188 0.0742129 0.0120436 6.37751e-06 0.00115402 0.0927735 0.000656492 0.0934253 0.857759 101.88 0.246178 0.71503 4.12021 0.0538225 0.0388699 0.96113 0.0198775 0.00423909 0.0191399 0.00408098 0.00512254 0.00586014 0.204902 0.234406 57.969 -87.8944 126.035 15.9829 145.01 0.000143567 0.267079 192.93 0.310721 0.0673899 0.00409474 0.000561553 0.00138242 0.986993 0.991736 -2.97159e-06 -85.6686 0.0929776 31196.8 300.442 0.983523 0.319147 0.744754 0.744749 9.99958 2.98035e-06 1.19213e-05 0.130601 0.978361 0.929961 -0.0132934 4.89364e-06 0.50069 -1.872e-20 6.89134e-24 -1.87132e-20 0.00139504 0.997818 8.59234e-05 0.152542 2.85165 0.00139504 0.99791 0.673072 0.00104425 0.00187955 0.000859234 0.455666 0.00187955 0.435284 0.000127469 1.02 0.887396 0.53476 0.285659 1.71612e-07 3.05574e-09 2391.97 3167.89 -0.0587499 0.482115 0.277636 0.256542 -0.592771 -0.169492 0.487164 -0.268442 -0.218729 1.386 1 1.08124e-301 294.318 6.49033e-299 2.03966 1.384 0.000299965 0.87597 0.639178 0.477815 0.401904 2.03993 128.707 83.3206 18.686 60.5769 0.00405015 0 -40 10
0.485 1.40595e-08 2.53884e-06 0.0743104 0.0743045 0.0120436 6.39067e-06 0.00115402 0.0928879 0.000656498 0.0935398 0.857806 101.88 0.246172 0.715096 4.1203 0.0538277 0.0388707 0.961129 0.0198774 0.00423918 0.0191398 0.00408105 0.00512265 0.00586024 0.204906 0.23441 57.9691 -87.8944 126.037 15.9829 145.01 0.000143555 0.26708 192.93 0.31072 0.0673899 0.00409474 0.000561553 0.00138242 0.986993 0.991736 -2.9716e-06 -85.6686 0.0929777 31196.8 300.444 0.983523 0.319147 0.744693 0.744689 9.99958 2.98036e-06 1.19213e-05 0.130602 0.978377 0.929969 -0.0132934 4.89367e-06 0.500693 -1.87209e-20 6.89168e-24 -1.8714e-20 0.00139504 0.997818 8.59235e-05 0.152542 2.85165 0.00139504 0.997909 0.673186 0.00104426 0.00187955 0.000859235 0.455665 0.00187955 0.435294 0.000127472 1.02 0.887397 0.53476 0.285661 1.71612e-07 3.05576e-09 2391.95 3167.63 -0.0587316 0.482115 0.277636 0.256526 -0.592774 -0.169492 0.487218 -0.26844 -0.218785 1.387 1 6.55808e-302 294.336 3.9372e-299 2.03985 1.385 0.000299965 0.875855 0.639238 0.477429 0.401936 2.04012 128.718 83.3236 18.6862 60.5784 0.00405003 0 -40 10
0.486 1.40885e-08 2.53884e-06 0.0744019 0.0743961 0.0120436 6.40384e-06 0.00115402 0.0930023 0.000656504 0.0936542 0.857852 101.88 0.246167 0.715162 4.12039 0.0538329 0.0388716 0.961128 0.0198772 0.00423926 0.0191396 0.00408113 0.00512276 0.00586035 0.20491 0.234414 57.9691 -87.8944 126.038 15.9829 145.01 0.000143544 0.26708 192.93 0.31072 0.0673899 0.00409474 0.000561554 0.00138242 0.986993 0.991736 -2.97162e-06 -85.6686 0.0929778 31196.7 300.447 0.983523 0.319147 0.744633 0.744628 9.99958 2.98036e-06 1.19213e-05 0.130603 0.978393 0.929977 -0.0132934 4.89369e-06 0.500697 -1.87217e-20 6.89202e-24 -1.87148e-20 0.00139505 0.997818 8.59235e-05 0.152543 2.85165 0.00139505 0.997909 0.6733 0.00104428 0.00187956 0.000859235 0.455665 0.00187955 0.435304 0.000127476 1.02 0.887398 0.53476 0.285662 1.71613e-07 3.05578e-09 2391.94 3167.37 -0.0587134 0.482115 0.277636 0.25651 -0.592777 -0.169493 0.487272 -0.268438 -0.218841 1.388 1 3.97768e-302 294.354 2.3884e-299 2.04004 1.386 0.000299965 0.87574 0.639298 0.477044 0.401968 2.04031 128.728 83.3266 18.6864 60.5798 0.00404991 0 -40 10
0.487 1.41174e-08 2.53884e-06 0.0744933 0.0744875 0.0120436 6.41701e-06 0.00115402 0.0931166 0.000656509 0.0937685 0.857899 101.88 0.246162 0.715228 4.12047 0.0538382 0.0388724 0.961128 0.0198771 0.00423935 0.0191395 0.0040812 0.00512286 0.00586046 0.204915 0.234418 57.9692 -87.8944 126.039 15.9828 145.01 0.000143532 0.26708 192.93 0.31072 0.0673898 0.00409475 0.000561554 0.00138243 0.986993 0.991736 -2.97163e-06 -85.6686 0.0929778 31196.7 300.449 0.983523 0.319147 0.744573 0.744568 9.99958 2.98036e-06 1.19213e-05 0.130604 0.978409 0.929985 -0.0132934 4.89372e-06 0.500701 -1.87225e-20 6.89235e-24 -1.87156e-20 0.00139505 0.997818 8.59236e-05 0.152543 2.85165 0.00139505 0.997908 0.673414 0.0010443 0.00187956 0.000859236 0.455665 0.00187956 0.435313 0.000127479 1.02 0.887399 0.534759 0.285663 1.71613e-07 3.05579e-09 2391.92 3167.12 -0.0586952 0.482115 0.277636 0.256494 -0.59278 -0.169493 0.487325 -0.268436 -0.218896 1.389 1 2.41258e-302 294.372 1.44886e-299 2.04023 1.387 0.000299965 0.875626 0.639358 0.476661 0.402001 2.0405 128.738 83.3295 18.6866 60.5812 0.00404978 0 -40 10
0.488 1.41464e-08 2.53884e-06 0.0745847 0.0745789 0.0120435 6.43017e-06 0.00115402 0.0932308 0.000656515 0.0938828 0.857945 101.879 0.246157 0.715294 4.12056 0.0538434 0.0388732 0.961127 0.019877 0.00423944 0.0191394 0.00408127 0.00512297 0.00586057 0.204919 0.234423 57.9693 -87.8944 126.04 15.9828 145.01 0.000143521 0.26708 192.929 0.310719 0.0673898 0.00409475 0.000561555 0.00138243 0.986993 0.991736 -2.97164e-06 -85.6686 0.0929779 31196.7 300.451 0.983522 0.319147 0.744513 0.744508 9.99958 2.98037e-06 1.19214e-05 0.130605 0.978425 0.929992 -0.0132934 4.89374e-06 0.500704 -1.87233e-20 6.89269e-24 -1.87164e-20 0.00139505 0.997818 8.59237e-05 0.152543 2.85166 0.00139505 0.997908 0.673527 0.00104432 0.00187956 0.000859237 0.455665 0.00187956 0.435323 0.000127483 1.02 0.8874 0.534759 0.285664 1.71613e-07 3.05581e-09 2391.9 3166.86 -0.0586771 0.482115 0.277635 0.256478 -0.592783 -0.169493 0.487379 -0.268434 -0.218951 1.39 1 1.46331e-302 294.39 8.78917e-300 2.04042 1.388 0.000299964 0.875512 0.639418 0.476278 0.402033 2.0407 128.748 83.3324 18.6867 60.5826 0.00404966 0 -40 10
0.489 1.41753e-08 2.53884e-06 0.074676 0.0746702 0.0120435 6.44334e-06 0.00115402 0.093345 0.000656521 0.0939969 0.857992 101.879 0.246151 0.71536 4.12065 0.0538487 0.0388741 0.961126 0.0198769 0.00423953 0.0191393 0.00408135 0.00512308 0.00586067 0.204923 0.234427 57.9693 -87.8944 126.041 15.9827 145.01 0.000143509 0.26708 192.929 0.310719 0.0673897 0.00409475 0.000561555 0.00138243 0.986993 0.991736 -2.97165e-06 -85.6686 0.092978 31196.7 300.454 0.983522 0.319147 0.744453 0.744449 9.99958 2.98037e-06 1.19214e-05 0.130606 0.978441 0.93 -0.0132934 4.89376e-06 0.500708 -1.87242e-20 6.89303e-24 -1.87173e-20 0.00139505 0.997818 8.59237e-05 0.152543 2.85166 0.00139505 0.997907 0.673641 0.00104434 0.00187956 0.000859237 0.455665 0.00187956 0.435333 0.000127486 1.02 0.887401 0.534759 0.285666 1.71613e-07 3.05583e-09 2391.89 3166.61 -0.0586591 0.482115 0.277635 0.256462 -0.592786 -0.169493 0.487432 -0.268433 -0.219006 1.391 1 8.8754e-303 294.408 5.33173e-300 2.04062 1.389 0.000299964 0.875398 0.639478 0.475897 0.402066 2.04089 128.759 83.3354 18.6869 60.5841 0.00404954 0 -40 10
0.49 1.42043e-08 2.53884e-06 0.0747672 0.0747615 0.0120435 6.4565e-06 0.00115402 0.093459 0.000656527 0.0941109 0.858039 101.879 0.246146 0.715426 4.12074 0.0538539 0.0388749 0.961125 0.0198768 0.00423962 0.0191392 0.00408142 0.00512319 0.00586078 0.204928 0.234431 57.9694 -87.8944 126.042 15.9827 145.01 0.000143498 0.26708 192.929 0.310719 0.0673897 0.00409475 0.000561556 0.00138243 0.986993 0.991736 -2.97166e-06 -85.6686 0.092978 31196.7 300.456 0.983522 0.319147 0.744394 0.744389 9.99958 2.98037e-06 1.19214e-05 0.130607 0.978457 0.930008 -0.0132934 4.89379e-06 0.500712 -1.8725e-20 6.89336e-24 -1.87181e-20 0.00139505 0.997818 8.59238e-05 0.152543 2.85166 0.00139505 0.997906 0.673755 0.00104436 0.00187956 0.000859238 0.455664 0.00187956 0.435342 0.00012749 1.02 0.887402 0.534759 0.285667 1.71613e-07 3.05585e-09 2391.87 3166.35 -0.0586412 0.482115 0.277635 0.256446 -0.592789 -0.169493 0.487485 -0.268431 -0.219061 1.392 1 5.3832e-303 294.426 3.23435e-300 2.04081 1.39 0.000299964 0.875285 0.639538 0.475516 0.402098 2.04108 128.769 83.3383 18.6871 60.5855 0.00404942 0 -40 10
0.491 1.42333e-08 2.53885e-06 0.0748583 0.0748526 0.0120435 6.46967e-06 0.00115402 0.0935729 0.000656532 0.0942249 0.858085 101.879 0.246141 0.715493 4.12083 0.0538592 0.0388757 0.961124 0.0198767 0.00423971 0.0191391 0.00408149 0.0051233 0.00586089 0.204932 0.234436 57.9694 -87.8944 126.043 15.9827 145.01 0.000143486 0.26708 192.929 0.310718 0.0673897 0.00409475 0.000561556 0.00138243 0.986993 0.991736 -2.97167e-06 -85.6686 0.0929781 31196.7 300.459 0.983522 0.319147 0.744334 0.74433 9.99958 2.98038e-06 1.19214e-05 0.130608 0.978473 0.930015 -0.0132934 4.89381e-06 0.500715 -1.87258e-20 6.8937e-24 -1.87189e-20 0.00139505 0.997818 8.59238e-05 0.152543 2.85166 0.00139505 0.997906 0.673868 0.00104438 0.00187956 0.000859238 0.455664 0.00187956 0.435352 0.000127493 1.02 0.887403 0.534758 0.285668 1.71614e-07 3.05587e-09 2391.85 3166.1 -0.0586233 0.482115 0.277634 0.25643 -0.592792 -0.169493 0.487537 -0.268429 -0.219116 1.393 1 3.26508e-303 294.443 1.96204e-300 2.041 1.391 0.000299964 0.875173 0.639598 0.475136 0.40213 2.04127 128.779 83.3412 18.6872 60.5869 0.0040493 0 -40 10
0.492 1.42622e-08 2.53885e-06 0.0749494 0.0749437 0.0120435 6.48284e-06 0.00115402 0.0936868 0.000656538 0.0943387 0.858132 101.879 0.246136 0.71556 4.12092 0.0538645 0.0388766 0.961123 0.0198766 0.0042398 0.019139 0.00408157 0.00512341 0.005861 0.204936 0.23444 57.9695 -87.8944 126.044 15.9826 145.01 0.000143475 0.267081 192.929 0.310718 0.0673896 0.00409476 0.000561557 0.00138243 0.986993 0.991736 -2.97168e-06 -85.6686 0.0929782 31196.6 300.461 0.983522 0.319147 0.744275 0.744271 9.99958 2.98038e-06 1.19214e-05 0.130609 0.978488 0.930023 -0.0132934 4.89384e-06 0.500719 -1.87266e-20 6.89404e-24 -1.87197e-20 0.00139505 0.997818 8.59239e-05 0.152543 2.85166 0.00139505 0.997905 0.673982 0.0010444 0.00187956 0.000859239 0.455664 0.00187956 0.435362 0.000127497 1.02 0.887403 0.534758 0.285669 1.71614e-07 3.05589e-09 2391.84 3165.85 -0.0586055 0.482115 0.277634 0.256414 -0.592795 -0.169493 0.48759 -0.268427 -0.21917 1.394 1 1.98037e-303 294.461 1.19022e-300 2.04119 1.392 0.000299964 0.875061 0.639657 0.474758 0.402163 2.04146 128.789 83.3441 18.6874 60.5883 0.00404918 0 -40 10
0.493 1.42912e-08 2.53885e-06 0.0750404 0.0750347 0.0120435 6.496e-06 0.00115402 0.0938005 0.000656544 0.0944525 0.858179 101.879 0.24613 0.715626 4.12101 0.0538698 0.0388774 0.961123 0.0198765 0.00423989 0.0191389 0.00408164 0.00512352 0.00586111 0.204941 0.234444 57.9696 -87.8944 126.045 15.9826 145.01 0.000143463 0.267081 192.929 0.310718 0.0673896 0.00409476 0.000561557 0.00138244 0.986993 0.991736 -2.9717e-06 -85.6685 0.0929782 31196.6 300.464 0.983522 0.319147 0.744217 0.744212 9.99958 2.98039e-06 1.19214e-05 0.13061 0.978504 0.93003 -0.0132934 4.89386e-06 0.500723 -1.87274e-20 6.89437e-24 -1.87205e-20 0.00139505 0.997818 8.5924e-05 0.152543 2.85166 0.00139505 0.997905 0.674095 0.00104442 0.00187956 0.00085924 0.455664 0.00187956 0.435371 0.0001275 1.02 0.887404 0.534758 0.285671 1.71614e-07 3.05591e-09 2391.82 3165.6 -0.0585878 0.482115 0.277634 0.256398 -0.592798 -0.169493 0.487642 -0.268425 -0.219224 1.395 1 1.20115e-303 294.479 7.22015e-301 2.04138 1.393 0.000299964 0.874949 0.639717 0.47438 0.402195 2.04165 128.799 83.3469 18.6876 60.5896 0.00404906 0 -40 10
0.494 1.43202e-08 2.53885e-06 0.0751314 0.0751257 0.0120435 6.50917e-06 0.00115402 0.0939142 0.000656549 0.0945661 0.858226 101.879 0.246125 0.715693 4.1211 0.0538751 0.0388783 0.961122 0.0198764 0.00423998 0.0191388 0.00408172 0.00512363 0.00586122 0.204945 0.234449 57.9696 -87.8944 126.046 15.9826 145.01 0.000143452 0.267081 192.929 0.310717 0.0673895 0.00409476 0.000561558 0.00138244 0.986993 0.991736 -2.97171e-06 -85.6685 0.0929783 31196.6 300.466 0.983522 0.319147 0.744158 0.744154 9.99958 2.98039e-06 1.19214e-05 0.130611 0.97852 0.930038 -0.0132934 4.89389e-06 0.500727 -1.87282e-20 6.89471e-24 -1.87213e-20 0.00139505 0.997818 8.5924e-05 0.152543 2.85166 0.00139505 0.997904 0.674209 0.00104444 0.00187956 0.00085924 0.455664 0.00187956 0.435381 0.000127504 1.02 0.887405 0.534758 0.285672 1.71614e-07 3.05592e-09 2391.8 3165.35 -0.0585701 0.482115 0.277634 0.256383 -0.592801 -0.169493 0.487694 -0.268423 -0.219278 1.396 1 7.28537e-304 294.496 4.37991e-301 2.04157 1.394 0.000299963 0.874838 0.639777 0.474004 0.402227 2.04184 128.81 83.3498 18.6877 60.591 0.00404894 0 -40 10
0.495 1.43491e-08 2.53885e-06 0.0752222 0.0752166 0.0120435 6.52233e-06 0.00115402 0.0940278 0.000656555 0.0946797 0.858273 101.879 0.24612 0.71576 4.12119 0.0538804 0.0388791 0.961121 0.0198763 0.00424007 0.0191387 0.00408179 0.00512374 0.00586132 0.20495 0.234453 57.9697 -87.8944 126.047 15.9825 145.01 0.000143441 0.267081 192.929 0.310717 0.0673895 0.00409476 0.000561558 0.00138244 0.986993 0.991736 -2.97172e-06 -85.6685 0.0929784 31196.6 300.468 0.983522 0.319147 0.7441 0.744095 9.99958 2.98039e-06 1.19215e-05 0.130611 0.978536 0.930045 -0.0132934 4.89391e-06 0.50073 -1.87291e-20 6.89505e-24 -1.87222e-20 0.00139505 0.997818 8.59241e-05 0.152544 2.85166 0.00139505 0.997904 0.674322 0.00104446 0.00187957 0.000859241 0.455664 0.00187956 0.435391 0.000127508 1.02 0.887406 0.534757 0.285673 1.71614e-07 3.05594e-09 2391.79 3165.1 -0.0585525 0.482116 0.277633 0.256367 -0.592804 -0.169493 0.487746 -0.268421 -0.219332 1.397 1 4.4188e-304 294.514 2.65696e-301 2.04176 1.395 0.000299963 0.874727 0.639836 0.473628 0.40226 2.04203 128.82 83.3527 18.6879 60.5924 0.00404882 0 -40 10
0.496 1.43781e-08 2.53885e-06 0.075313 0.0753074 0.0120434 6.5355e-06 0.00115402 0.0941412 0.000656561 0.0947932 0.858321 101.879 0.246114 0.715827 4.12128 0.0538857 0.03888 0.96112 0.0198761 0.00424016 0.0191386 0.00408187 0.00512386 0.00586143 0.204954 0.234457 57.9698 -87.8944 126.048 15.9825 145.01 0.00014343 0.267081 192.928 0.310717 0.0673895 0.00409477 0.000561559 0.00138244 0.986993 0.991736 -2.97173e-06 -85.6685 0.0929784 31196.6 300.471 0.983522 0.319147 0.744041 0.744037 9.99958 2.9804e-06 1.19215e-05 0.130612 0.978551 0.930053 -0.0132934 4.89394e-06 0.500734 -1.87299e-20 6.89538e-24 -1.8723e-20 0.00139505 0.997818 8.59242e-05 0.152544 2.85166 0.00139505 0.997903 0.674436 0.00104448 0.00187957 0.000859242 0.455663 0.00187957 0.4354 0.000127511 1.02 0.887407 0.534757 0.285674 1.71615e-07 3.05596e-09 2391.77 3164.85 -0.058535 0.482116 0.277633 0.256351 -0.592807 -0.169493 0.487798 -0.268419 -0.219385 1.398 1 2.68014e-304 294.531 1.61177e-301 2.04195 1.396 0.000299963 0.874616 0.639896 0.473254 0.402292 2.04222 128.83 83.3555 18.6881 60.5938 0.0040487 0 -40 10
0.497 1.44071e-08 2.53885e-06 0.0754037 0.0753981 0.0120434 6.54867e-06 0.00115402 0.0942546 0.000656566 0.0949066 0.858368 101.879 0.246109 0.715894 4.12137 0.0538911 0.0388808 0.961119 0.019876 0.00424025 0.0191385 0.00408194 0.00512397 0.00586155 0.204959 0.234462 57.9698 -87.8944 126.049 15.9824 145.01 0.000143418 0.267081 192.928 0.310716 0.0673894 0.00409477 0.000561559 0.00138244 0.986993 0.991736 -2.97174e-06 -85.6685 0.0929785 31196.5 300.473 0.983522 0.319147 0.743983 0.743979 9.99958 2.9804e-06 1.19215e-05 0.130613 0.978567 0.93006 -0.0132934 4.89396e-06 0.500738 -1.87307e-20 6.89572e-24 -1.87238e-20 0.00139506 0.997818 8.59242e-05 0.152544 2.85166 0.00139506 0.997902 0.674549 0.0010445 0.00187957 0.000859242 0.455663 0.00187957 0.43541 0.000127515 1.02 0.887408 0.534757 0.285676 1.71615e-07 3.05598e-09 2391.75 3164.6 -0.0585176 0.482116 0.277633 0.256336 -0.59281 -0.169493 0.487849 -0.268418 -0.219439 1.399 1 1.62559e-304 294.549 9.77737e-302 2.04214 1.397 0.000299963 0.874506 0.639956 0.47288 0.402324 2.04241 128.84 83.3584 18.6882 60.5952 0.00404858 0 -40 10
0.498 1.4436e-08 2.53885e-06 0.0754943 0.0754888 0.0120434 6.56183e-06 0.00115402 0.0943679 0.000656572 0.0950199 0.858415 101.879 0.246104 0.715962 4.12146 0.0538964 0.0388817 0.961118 0.0198759 0.00424034 0.0191383 0.00408202 0.00512408 0.00586166 0.204963 0.234466 57.9699 -87.8944 126.05 15.9824 145.01 0.000143407 0.267082 192.928 0.310716 0.0673894 0.00409477 0.00056156 0.00138244 0.986993 0.991736 -2.97176e-06 -85.6685 0.0929786 31196.5 300.476 0.983522 0.319147 0.743926 0.743921 9.99958 2.9804e-06 1.19215e-05 0.130614 0.978582 0.930068 -0.0132934 4.89399e-06 0.500742 -1.87315e-20 6.89605e-24 -1.87246e-20 0.00139506 0.997818 8.59243e-05 0.152544 2.85166 0.00139506 0.997902 0.674663 0.00104452 0.00187957 0.000859243 0.455663 0.00187957 0.43542 0.000127518 1.02 0.887409 0.534757 0.285677 1.71615e-07 3.056e-09 2391.74 3164.36 -0.0585002 0.482116 0.277632 0.25632 -0.592813 -0.169493 0.4879 -0.268416 -0.219492 1.4 1 9.85968e-305 294.566 5.93118e-302 2.04233 1.398 0.000299963 0.874396 0.640015 0.472508 0.402356 2.0426 128.85 83.3612 18.6884 60.5965 0.00404846 0 -40 10
0.499 1.4465e-08 2.53885e-06 0.0755849 0.0755793 0.0120434 6.575e-06 0.00115402 0.0944811 0.000656578 0.0951331 0.858462 101.878 0.246098 0.716029 4.12155 0.0539017 0.0388826 0.961117 0.0198758 0.00424043 0.0191382 0.00408209 0.00512419 0.00586177 0.204968 0.234471 57.9699 -87.8944 126.051 15.9824 145.01 0.000143396 0.267082 192.928 0.310716 0.0673893 0.00409477 0.00056156 0.00138245 0.986993 0.991736 -2.97177e-06 -85.6685 0.0929786 31196.5 300.478 0.983522 0.319147 0.743868 0.743864 9.99958 2.98041e-06 1.19215e-05 0.130615 0.978598 0.930075 -0.0132934 4.89401e-06 0.500745 -1.87323e-20 6.89639e-24 -1.87254e-20 0.00139506 0.997818 8.59243e-05 0.152544 2.85166 0.00139506 0.997901 0.674776 0.00104453 0.00187957 0.000859243 0.455663 0.00187957 0.435429 0.000127522 1.02 0.88741 0.534756 0.285678 1.71615e-07 3.05602e-09 2391.72 3164.11 -0.0584829 0.482116 0.277632 0.256305 -0.592816 -0.169493 0.487951 -0.268414 -0.219545 1.401 1 5.9802e-305 294.583 3.59799e-302 2.04252 1.399 0.000299963 0.874287 0.640075 0.472136 0.402388 2.04279 128.861 83.364 18.6886 60.5979 0.00404835 0 -40 10
0.5 1.4494e-08 2.53885e-06 0.0756754 0.0756699 0.0120434 6.58816e-06 0.00115402 0.0945943 0.000656583 0.0952462 0.85851 101.878 0.246093 0.716097 4.12164 0.0539071 0.0388834 0.961117 0.0198757 0.00424053 0.0191381 0.00408217 0.00512431 0.00586188 0.204972 0.234475 57.97 -87.8944 126.052 15.9823 145.01 0.000143385 0.267082 192.928 0.310715 0.0673893 0.00409478 0.000561561 0.00138245 0.986993 0.991736 -2.97178e-06 -85.6685 0.0929787 31196.5 300.481 0.983522 0.319147 0.743811 0.743806 9.99958 2.98041e-06 1.19215e-05 0.130616 0.978613 0.930082 -0.0132934 4.89404e-06 0.500749 -1.87331e-20 6.89673e-24 -1.87262e-20 0.00139506 0.997818 8.59244e-05 0.152544 2.85166 0.00139506 0.997901 0.674889 0.00104455 0.00187957 0.000859244 0.455663 0.00187957 0.435439 0.000127525 1.02 0.887411 0.534756 0.28568 1.71615e-07 3.05604e-09 2391.7 3163.87 -0.0584656 0.482116 0.277632 0.25629 -0.592818 -0.169493 0.488002 -0.268412 -0.219597 1.402 1 3.62717e-305 294.6 2.18262e-302 2.04271 1.4 0.000299962 0.874178 0.640134 0.471766 0.402421 2.04298 128.871 83.3668 18.6887 60.5992 0.00404823 0 -40 10
0.501 1.45229e-08 2.53885e-06 0.0757658 0.0757603 0.0120434 6.60133e-06 0.00115402 0.0947073 0.000656589 0.0953593 0.858557 101.878 0.246088 0.716164 4.12174 0.0539125 0.0388843 0.961116 0.0198756 0.00424062 0.019138 0.00408225 0.00512442 0.00586199 0.204977 0.23448 57.9701 -87.8944 126.053 15.9823 145.01 0.000143374 0.267082 192.928 0.310715 0.0673893 0.00409478 0.000561561 0.00138245 0.986993 0.991736 -2.97179e-06 -85.6685 0.0929788 31196.5 300.483 0.983522 0.319147 0.743754 0.743749 9.99958 2.98042e-06 1.19216e-05 0.130617 0.978628 0.93009 -0.0132934 4.89406e-06 0.500753 -1.8734e-20 6.89706e-24 -1.87271e-20 0.00139506 0.997818 8.59245e-05 0.152544 2.85166 0.00139506 0.9979 0.675002 0.00104457 0.00187957 0.000859245 0.455663 0.00187957 0.435449 0.000127529 1.02 0.887412 0.534756 0.285681 1.71616e-07 3.05606e-09 2391.69 3163.63 -0.0584484 0.482116 0.277632 0.256274 -0.592821 -0.169494 0.488053 -0.26841 -0.21965 1.403 1 2.19999e-305 294.617 1.32403e-302 2.0429 1.401 0.000299962 0.87407 0.640193 0.471396 0.402453 2.04317 128.881 83.3696 18.6889 60.6006 0.00404811 0 -40 10
0.502 1.45519e-08 2.53885e-06 0.0758562 0.0758507 0.0120434 6.61449e-06 0.00115402 0.0948202 0.000656594 0.0954722 0.858605 101.878 0.246082 0.716232 4.12183 0.0539179 0.0388852 0.961115 0.0198755 0.00424071 0.0191379 0.00408232 0.00512453 0.0058621 0.204981 0.234484 57.9701 -87.8944 126.054 15.9823 145.01 0.000143363 0.267082 192.928 0.310715 0.0673892 0.00409478 0.000561562 0.00138245 0.986993 0.991736 -2.9718e-06 -85.6685 0.0929788 31196.5 300.486 0.983522 0.319147 0.743697 0.743692 9.99958 2.98042e-06 1.19216e-05 0.130618 0.978644 0.930097 -0.0132934 4.89409e-06 0.500757 -1.87348e-20 6.8974e-24 -1.87279e-20 0.00139506 0.997818 8.59245e-05 0.152544 2.85167 0.00139506 0.9979 0.675115 0.00104459 0.00187957 0.000859245 0.455662 0.00187957 0.435458 0.000127532 1.02 0.887413 0.534755 0.285682 1.71616e-07 3.05608e-09 2391.67 3163.38 -0.0584313 0.482116 0.277631 0.256259 -0.592824 -0.169494 0.488103 -0.268408 -0.219702 1.404 1 1.33436e-305 294.634 8.03183e-303 2.04309 1.402 0.000299962 0.873962 0.640253 0.471027 0.402485 2.04336 128.891 83.3724 18.6891 60.6019 0.004048 0 -40 10
0.503 1.45808e-08 2.53885e-06 0.0759465 0.075941 0.0120434 6.62766e-06 0.00115402 0.0949331 0.0006566 0.0955851 0.858652 101.878 0.246077 0.7163 4.12192 0.0539232 0.038886 0.961114 0.0198754 0.0042408 0.0191378 0.0040824 0.00512465 0.00586221 0.204986 0.234489 57.9702 -87.8944 126.055 15.9822 145.01 0.000143352 0.267082 192.927 0.310714 0.0673892 0.00409478 0.000561562 0.00138245 0.986993 0.991736 -2.97181e-06 -85.6685 0.0929789 31196.4 300.488 0.983522 0.319147 0.74364 0.743636 9.99958 2.98042e-06 1.19216e-05 0.130619 0.978659 0.930104 -0.0132934 4.89411e-06 0.500761 -1.87356e-20 6.89773e-24 -1.87287e-20 0.00139506 0.997818 8.59246e-05 0.152545 2.85167 0.00139506 0.997899 0.675229 0.00104461 0.00187957 0.000859246 0.455662 0.00187957 0.435468 0.000127536 1.02 0.887414 0.534755 0.285683 1.71616e-07 3.05609e-09 2391.66 3163.14 -0.0584143 0.482116 0.277631 0.256244 -0.592827 -0.169494 0.488153 -0.268406 -0.219754 1.405 1 8.09332e-306 294.651 4.87228e-303 2.04328 1.403 0.000299962 0.873854 0.640312 0.47066 0.402517 2.04355 128.901 83.3752 18.6892 60.6033 0.00404788 0 -40 10
0.504 1.46098e-08 2.53885e-06 0.0760367 0.0760312 0.0120433 6.64082e-06 0.00115402 0.0950458 0.000656605 0.0956978 0.8587 101.878 0.246071 0.716368 4.12201 0.0539286 0.0388869 0.961113 0.0198752 0.0042409 0.0191377 0.00408248 0.00512476 0.00586233 0.204991 0.234493 57.9703 -87.8944 126.056 15.9822 145.01 0.000143341 0.267082 192.927 0.310714 0.0673891 0.00409478 0.000561563 0.00138245 0.986993 0.991736 -2.97183e-06 -85.6685 0.092979 31196.4 300.491 0.983522 0.319147 0.743584 0.743579 9.99958 2.98043e-06 1.19216e-05 0.13062 0.978674 0.930112 -0.0132934 4.89414e-06 0.500765 -1.87364e-20 6.89807e-24 -1.87295e-20 0.00139506 0.997818 8.59247e-05 0.152545 2.85167 0.00139506 0.997899 0.675342 0.00104463 0.00187958 0.000859247 0.455662 0.00187957 0.435477 0.000127539 1.02 0.887415 0.534755 0.285685 1.71616e-07 3.05611e-09 2391.64 3162.9 -0.0583973 0.482116 0.277631 0.256229 -0.59283 -0.169494 0.488203 -0.268404 -0.219806 1.406 1 4.90884e-306 294.668 2.95563e-303 2.04347 1.404 0.000299962 0.873747 0.640371 0.470293 0.402549 2.04374 128.911 83.3779 18.6894 60.6046 0.00404777 0 -40 10
0.505 1.46388e-08 2.53885e-06 0.0761268 0.0761213 0.0120433 6.65399e-06 0.00115402 0.0951585 0.000656611 0.0958105 0.858748 101.878 0.246066 0.716436 4.12211 0.053934 0.0388878 0.961112 0.0198751 0.00424099 0.0191376 0.00408255 0.00512488 0.00586244 0.204995 0.234498 57.9703 -87.8944 126.057 15.9821 145.01 0.000143331 0.267083 192.927 0.310714 0.0673891 0.00409479 0.000561563 0.00138246 0.986993 0.991736 -2.97184e-06 -85.6685 0.092979 31196.4 300.493 0.983522 0.319147 0.743527 0.743523 9.99958 2.98043e-06 1.19216e-05 0.130621 0.978689 0.930119 -0.0132934 4.89416e-06 0.500769 -1.87372e-20 6.89841e-24 -1.87303e-20 0.00139506 0.997818 8.59247e-05 0.152545 2.85167 0.00139506 0.997898 0.675455 0.00104465 0.00187958 0.000859247 0.455662 0.00187958 0.435487 0.000127543 1.02 0.887415 0.534755 0.285686 1.71617e-07 3.05613e-09 2391.62 3162.66 -0.0583804 0.482116 0.27763 0.256214 -0.592833 -0.169494 0.488253 -0.268403 -0.219858 1.407 1 2.97736e-306 294.685 1.79295e-303 2.04366 1.405 0.000299961 0.87364 0.640431 0.469928 0.402581 2.04393 128.921 83.3807 18.6895 60.606 0.00404765 0 -40 10
0.506 1.46677e-08 2.53885e-06 0.0762168 0.0762114 0.0120433 6.66715e-06 0.00115402 0.095271 0.000656616 0.095923 0.858796 101.878 0.246061 0.716505 4.1222 0.0539395 0.0388887 0.961111 0.019875 0.00424108 0.0191374 0.00408263 0.00512499 0.00586255 0.205 0.234502 57.9704 -87.8945 126.058 15.9821 145.01 0.00014332 0.267083 192.927 0.310713 0.067389 0.00409479 0.000561564 0.00138246 0.986993 0.991736 -2.97185e-06 -85.6685 0.0929791 31196.4 300.496 0.983522 0.319147 0.743471 0.743467 9.99958 2.98043e-06 1.19216e-05 0.130622 0.978704 0.930126 -0.0132934 4.89419e-06 0.500772 -1.8738e-20 6.89874e-24 -1.87311e-20 0.00139506 0.997818 8.59248e-05 0.152545 2.85167 0.00139506 0.997898 0.675568 0.00104467 0.00187958 0.000859248 0.455662 0.00187958 0.435497 0.000127546 1.02 0.887416 0.534754 0.285687 1.71617e-07 3.05615e-09 2391.61 3162.42 -0.0583636 0.482116 0.27763 0.256199 -0.592835 -0.169494 0.488303 -0.268401 -0.219909 1.408 1 1.80586e-306 294.702 1.08764e-303 2.04385 1.406 0.000299961 0.873534 0.64049 0.469563 0.402613 2.04412 128.932 83.3834 18.6897 60.6073 0.00404754 0 -40 10
0.507 1.46967e-08 2.53885e-06 0.0763068 0.0763014 0.0120433 6.68032e-06 0.00115402 0.0953835 0.000656621 0.0960355 0.858844 101.878 0.246055 0.716573 4.1223 0.0539449 0.0388896 0.96111 0.0198749 0.00424118 0.0191373 0.00408271 0.00512511 0.00586267 0.205004 0.234507 57.9704 -87.8945 126.059 15.9821 145.01 0.000143309 0.267083 192.927 0.310713 0.067389 0.00409479 0.000561564 0.00138246 0.986993 0.991736 -2.97186e-06 -85.6684 0.0929792 31196.4 300.498 0.983522 0.319147 0.743416 0.743411 9.99958 2.98044e-06 1.19216e-05 0.130623 0.97872 0.930133 -0.0132934 4.89421e-06 0.500776 -1.87388e-20 6.89908e-24 -1.87319e-20 0.00139506 0.997818 8.59248e-05 0.152545 2.85167 0.00139506 0.997897 0.675681 0.00104469 0.00187958 0.000859248 0.455662 0.00187958 0.435506 0.00012755 1.02 0.887417 0.534754 0.285689 1.71617e-07 3.05617e-09 2391.59 3162.18 -0.0583468 0.482116 0.27763 0.256184 -0.592838 -0.169494 0.488352 -0.268399 -0.219961 1.409 1 1.09531e-306 294.719 6.59787e-304 2.04404 1.407 0.000299961 0.873428 0.640549 0.469199 0.402645 2.0443 128.942 83.3862 18.6899 60.6086 0.00404742 0 -40 10
0.508 1.47257e-08 2.53885e-06 0.0763967 0.0763913 0.0120433 6.69348e-06 0.00115402 0.0954958 0.000656627 0.0961478 0.858892 101.878 0.24605 0.716641 4.12239 0.0539503 0.0388905 0.96111 0.0198748 0.00424127 0.0191372 0.00408279 0.00512523 0.00586278 0.205009 0.234511 57.9705 -87.8945 126.06 15.982 145.01 0.000143298 0.267083 192.927 0.310713 0.067389 0.00409479 0.000561565 0.00138246 0.986993 0.991736 -2.97187e-06 -85.6684 0.0929792 31196.4 300.501 0.983522 0.319147 0.74336 0.743356 9.99958 2.98044e-06 1.19217e-05 0.130624 0.978735 0.93014 -0.0132934 4.89424e-06 0.50078 -1.87397e-20 6.89941e-24 -1.87328e-20 0.00139506 0.997818 8.59249e-05 0.152545 2.85167 0.00139506 0.997897 0.675794 0.00104471 0.00187958 0.000859249 0.455661 0.00187958 0.435516 0.000127553 1.02 0.887418 0.534754 0.28569 1.71617e-07 3.05619e-09 2391.57 3161.95 -0.0583301 0.482116 0.277629 0.256169 -0.592841 -0.169494 0.488401 -0.268397 -0.220012 1.41 1 6.6434e-307 294.735 4.0024e-304 2.04423 1.408 0.000299961 0.873323 0.640608 0.468837 0.402677 2.04449 128.952 83.3889 18.69 60.6099 0.00404731 0 -40 10
0.509 1.47546e-08 2.53885e-06 0.0764865 0.0764811 0.0120433 6.70665e-06 0.00115402 0.0956081 0.000656632 0.0962601 0.85894 101.878 0.246044 0.71671 4.12248 0.0539558 0.0388914 0.961109 0.0198747 0.00424137 0.0191371 0.00408287 0.00512534 0.0058629 0.205014 0.234516 57.9706 -87.8945 126.061 15.982 145.01 0.000143288 0.267083 192.927 0.310712 0.0673889 0.0040948 0.000561566 0.00138246 0.986993 0.991736 -2.97189e-06 -85.6684 0.0929793 31196.3 300.504 0.983522 0.319147 0.743305 0.7433 9.99958 2.98045e-06 1.19217e-05 0.130625 0.97875 0.930147 -0.0132934 4.89426e-06 0.500784 -1.87405e-20 6.89975e-24 -1.87336e-20 0.00139507 0.997818 8.5925e-05 0.152545 2.85167 0.00139507 0.997896 0.675907 0.00104473 0.00187958 0.00085925 0.455661 0.00187958 0.435525 0.000127557 1.02 0.887419 0.534754 0.285691 1.71617e-07 3.05621e-09 2391.56 3161.71 -0.0583135 0.482116 0.277629 0.256154 -0.592844 -0.169494 0.48845 -0.268395 -0.220062 1.411 1 4.02942e-307 294.752 2.42794e-304 2.04442 1.409 0.000299961 0.873218 0.640667 0.468476 0.402709 2.04468 128.962 83.3916 18.6902 60.6112 0.0040472 0 -40 10
0.51 1.47836e-08 2.53885e-06 0.0765763 0.0765709 0.0120433 6.71981e-06 0.00115402 0.0957203 0.000656638 0.0963723 0.858988 101.877 0.246039 0.716779 4.12258 0.0539612 0.0388923 0.961108 0.0198745 0.00424146 0.019137 0.00408294 0.00512546 0.00586301 0.205018 0.234521 57.9706 -87.8945 126.062 15.982 145.01 0.000143277 0.267083 192.927 0.310712 0.0673889 0.0040948 0.000561566 0.00138246 0.986993 0.991736 -2.9719e-06 -85.6684 0.0929794 31196.3 300.506 0.983522 0.319147 0.74325 0.743245 9.99958 2.98045e-06 1.19217e-05 0.130626 0.978764 0.930154 -0.0132934 4.89429e-06 0.500788 -1.87413e-20 6.90008e-24 -1.87344e-20 0.00139507 0.997818 8.5925e-05 0.152545 2.85167 0.00139507 0.997896 0.676019 0.00104475 0.00187958 0.00085925 0.455661 0.00187958 0.435535 0.00012756 1.02 0.88742 0.534753 0.285692 1.71618e-07 3.05623e-09 2391.54 3161.48 -0.0582969 0.482116 0.277629 0.256139 -0.592846 -0.169494 0.488499 -0.268393 -0.220113 1.412 1 2.44397e-307 294.768 1.47284e-304 2.0446 1.41 0.000299961 0.873113 0.640726 0.468115 0.402741 2.04487 128.972 83.3943 18.6903 60.6125 0.00404708 0 -40 10
0.511 1.48126e-08 2.53885e-06 0.0766659 0.0766606 0.0120432 6.73298e-06 0.00115402 0.0958324 0.000656643 0.0964845 0.859036 101.877 0.246033 0.716848 4.12267 0.0539667 0.0388932 0.961107 0.0198744 0.00424156 0.0191369 0.00408302 0.00512558 0.00586313 0.205023 0.234525 57.9707 -87.8945 126.063 15.9819 145.01 0.000143266 0.267083 192.926 0.310712 0.0673888 0.0040948 0.000561567 0.00138247 0.986993 0.991736 -2.97191e-06 -85.6684 0.0929794 31196.3 300.509 0.983522 0.319147 0.743195 0.74319 9.99958 2.98045e-06 1.19217e-05 0.130627 0.978779 0.930162 -0.0132933 4.89431e-06 0.500792 -1.87421e-20 6.90042e-24 -1.87352e-20 0.00139507 0.997818 8.59251e-05 0.152546 2.85167 0.00139507 0.997895 0.676132 0.00104477 0.00187958 0.000859251 0.455661 0.00187958 0.435545 0.000127564 1.02 0.887421 0.534753 0.285694 1.71618e-07 3.05625e-09 2391.52 3161.24 -0.0582805 0.482116 0.277629 0.256125 -0.592849 -0.169494 0.488547 -0.268391 -0.220164 1.413 1 1.48234e-307 294.785 8.93454e-305 2.04479 1.411 0.00029996 0.873009 0.640785 0.467755 0.402772 2.04506 128.982 83.397 18.6905 60.6138 0.00404697 0 -40 10
0.512 1.48415e-08 2.53885e-06 0.0767556 0.0767502 0.0120432 6.74614e-06 0.00115402 0.0959445 0.000656648 0.0965965 0.859084 101.877 0.246028 0.716916 4.12277 0.0539721 0.0388941 0.961106 0.0198743 0.00424165 0.0191368 0.0040831 0.00512569 0.00586324 0.205028 0.23453 57.9708 -87.8945 126.064 15.9819 145.011 0.000143256 0.267084 192.926 0.310711 0.0673888 0.0040948 0.000561567 0.00138247 0.986993 0.991736 -2.97192e-06 -85.6684 0.0929795 31196.3 300.511 0.983522 0.319147 0.74314 0.743135 9.99958 2.98046e-06 1.19217e-05 0.130628 0.978794 0.930169 -0.0132933 4.89434e-06 0.500796 -1.87429e-20 6.90075e-24 -1.8736e-20 0.00139507 0.997818 8.59252e-05 0.152546 2.85167 0.00139507 0.997895 0.676245 0.00104479 0.00187958 0.000859252 0.455661 0.00187958 0.435554 0.000127568 1.02 0.887422 0.534753 0.285695 1.71618e-07 3.05627e-09 2391.51 3161.01 -0.058264 0.482117 0.277628 0.25611 -0.592852 -0.169494 0.488596 -0.268389 -0.220214 1.414 1 8.99086e-308 294.801 5.41987e-305 2.04498 1.412 0.00029996 0.872905 0.640844 0.467396 0.402804 2.04525 128.992 83.3997 18.6906 60.6151 0.00404686 0 -40 10
0.513 1.48705e-08 2.53885e-06 0.0768451 0.0768398 0.0120432 6.75931e-06 0.00115402 0.0960564 0.000656654 0.0967085 0.859132 101.877 0.246022 0.716985 4.12287 0.0539776 0.038895 0.961105 0.0198742 0.00424175 0.0191366 0.00408318 0.00512581 0.00586336 0.205032 0.234534 57.9708 -87.8945 126.065 15.9818 145.011 0.000143245 0.267084 192.926 0.310711 0.0673888 0.00409481 0.000561568 0.00138247 0.986993 0.991736 -2.97193e-06 -85.6684 0.0929796 31196.3 300.514 0.983522 0.319147 0.743085 0.743081 9.99958 2.98046e-06 1.19217e-05 0.130629 0.978809 0.930176 -0.0132933 4.89436e-06 0.5008 -1.87437e-20 6.90109e-24 -1.87368e-20 0.00139507 0.997818 8.59252e-05 0.152546 2.85167 0.00139507 0.997894 0.676358 0.00104481 0.00187959 0.000859252 0.45566 0.00187959 0.435564 0.000127571 1.02 0.887423 0.534753 0.285696 1.71618e-07 3.05629e-09 2391.49 3160.77 -0.0582476 0.482117 0.277628 0.256095 -0.592855 -0.169494 0.488644 -0.268387 -0.220264 1.415 1 5.45323e-308 294.817 3.2878e-305 2.04517 1.413 0.00029996 0.872801 0.640903 0.467038 0.402836 2.04543 129.002 83.4024 18.6908 60.6164 0.00404675 0 -40 10
0.514 1.48994e-08 2.53885e-06 0.0769346 0.0769293 0.0120432 6.77247e-06 0.00115402 0.0961683 0.000656659 0.0968203 0.859181 101.877 0.246017 0.717055 4.12296 0.0539831 0.0388959 0.961104 0.0198741 0.00424185 0.0191365 0.00408326 0.00512593 0.00586348 0.205037 0.234539 57.9709 -87.8945 126.066 15.9818 145.011 0.000143235 0.267084 192.926 0.310711 0.0673887 0.00409481 0.000561568 0.00138247 0.986993 0.991736 -2.97195e-06 -85.6684 0.0929796 31196.3 300.517 0.983522 0.319147 0.743031 0.743026 9.99958 2.98047e-06 1.19218e-05 0.13063 0.978824 0.930183 -0.0132933 4.89439e-06 0.500804 -1.87445e-20 6.90142e-24 -1.87376e-20 0.00139507 0.997818 8.59253e-05 0.152546 2.85167 0.00139507 0.997894 0.676471 0.00104483 0.00187959 0.000859253 0.45566 0.00187959 0.435573 0.000127575 1.02 0.887424 0.534752 0.285698 1.71618e-07 3.0563e-09 2391.47 3160.54 -0.0582313 0.482117 0.277628 0.256081 -0.592857 -0.169494 0.488692 -0.268385 -0.220314 1.416 1 3.30755e-308 294.834 1.99445e-305 2.04536 1.414 0.00029996 0.872698 0.640962 0.466681 0.402868 2.04562 129.012 83.405 18.691 60.6177 0.00404664 0 -40 10
0.515 1.49284e-08 2.53885e-06 0.077024 0.0770187 0.0120432 6.78564e-06 0.00115402 0.09628 0.000656664 0.0969321 0.859229 101.877 0.246011 0.717124 4.12306 0.0539886 0.0388968 0.961103 0.019874 0.00424194 0.0191364 0.00408334 0.00512605 0.00586359 0.205042 0.234544 57.9709 -87.8945 126.067 15.9818 145.011 0.000143224 0.267084 192.926 0.31071 0.0673887 0.00409481 0.000561569 0.00138247 0.986993 0.991736 -2.97196e-06 -85.6684 0.0929797 31196.2 300.519 0.983522 0.319147 0.742976 0.742972 9.99958 2.98047e-06 1.19218e-05 0.130631 0.978838 0.93019 -0.0132933 4.89441e-06 0.500808 -1.87453e-20 6.90176e-24 -1.87384e-20 0.00139507 0.997818 8.59253e-05 0.152546 2.85167 0.00139507 0.997893 0.676583 0.00104484 0.00187959 0.000859253 0.45566 0.00187959 0.435583 0.000127578 1.02 0.887425 0.534752 0.285699 1.71619e-07 3.05632e-09 2391.46 3160.31 -0.0582151 0.482117 0.277627 0.256066 -0.59286 -0.169494 0.48874 -0.268384 -0.220364 1.417 1 0 294.85 0 2.04554 1.415 0.00029996 0.872595 0.641021 0.466325 0.4029 2.04581 129.022 83.4077 18.6911 60.619 0.00404653 0 -40 10
0.516 1.49574e-08 2.53885e-06 0.0771134 0.0771081 0.0120432 6.7988e-06 0.00115402 0.0963917 0.00065667 0.0970438 0.859277 101.877 0.246006 0.717193 4.12316 0.0539941 0.0388977 0.961102 0.0198738 0.00424204 0.0191363 0.00408342 0.00512617 0.00586371 0.205047 0.234548 57.971 -87.8945 126.068 15.9817 145.011 0.000143214 0.267084 192.926 0.31071 0.0673886 0.00409481 0.000561569 0.00138247 0.986993 0.991736 -2.97197e-06 -85.6684 0.0929798 31196.2 300.522 0.983522 0.319147 0.742922 0.742918 9.99958 2.98047e-06 1.19218e-05 0.130632 0.978853 0.930197 -0.0132933 4.89444e-06 0.500812 -1.87461e-20 6.90209e-24 -1.87392e-20 0.00139507 0.997818 8.59254e-05 0.152546 2.85168 0.00139507 0.997893 0.676696 0.00104486 0.00187959 0.000859254 0.45566 0.00187959 0.435592 0.000127582 1.02 0.887426 0.534752 0.2857 1.71619e-07 3.05634e-09 2391.44 3160.08 -0.0581989 0.482117 0.277627 0.256052 -0.592863 -0.169494 0.488787 -0.268382 -0.220413 1.418 1 0 294.866 0 2.04573 1.416 0.000299959 0.872493 0.641079 0.46597 0.402931 2.046 129.032 83.4103 18.6913 60.6203 0.00404642 0 -40 10
0.517 1.49863e-08 2.53885e-06 0.0772026 0.0771974 0.0120432 6.81197e-06 0.00115402 0.0965033 0.000656675 0.0971554 0.859326 101.877 0.246 0.717263 4.12325 0.0539996 0.0388986 0.961101 0.0198737 0.00424214 0.0191362 0.0040835 0.00512629 0.00586383 0.205051 0.234553 57.9711 -87.8945 126.069 15.9817 145.011 0.000143204 0.267084 192.926 0.31071 0.0673886 0.00409482 0.00056157 0.00138248 0.986993 0.991736 -2.97198e-06 -85.6684 0.0929799 31196.2 300.524 0.983522 0.319147 0.742869 0.742864 9.99958 2.98048e-06 1.19218e-05 0.130633 0.978868 0.930204 -0.0132933 4.89447e-06 0.500816 -1.8747e-20 6.90243e-24 -1.87401e-20 0.00139507 0.997818 8.59255e-05 0.152546 2.85168 0.00139507 0.997892 0.676808 0.00104488 0.00187959 0.000859255 0.45566 0.00187959 0.435602 0.000127585 1.02 0.887427 0.534752 0.285702 1.71619e-07 3.05636e-09 2391.42 3159.85 -0.0581828 0.482117 0.277627 0.256037 -0.592865 -0.169495 0.488835 -0.26838 -0.220463 1.419 1 0 294.882 0 2.04592 1.417 0.000299959 0.872391 0.641138 0.465616 0.402963 2.04619 129.042 83.413 18.6914 60.6215 0.00404631 0 -40 10
0.518 1.50153e-08 2.53885e-06 0.0772918 0.0772866 0.0120432 6.82513e-06 0.00115402 0.0966148 0.00065668 0.0972669 0.859375 101.877 0.245995 0.717332 4.12335 0.0540051 0.0388995 0.9611 0.0198736 0.00424223 0.0191361 0.00408358 0.00512641 0.00586395 0.205056 0.234558 57.9711 -87.8945 126.07 15.9817 145.011 0.000143193 0.267085 192.926 0.310709 0.0673885 0.00409482 0.00056157 0.00138248 0.986993 0.991736 -2.972e-06 -85.6684 0.0929799 31196.2 300.527 0.983522 0.319147 0.742815 0.742811 9.99958 2.98048e-06 1.19218e-05 0.130634 0.978882 0.93021 -0.0132933 4.89449e-06 0.50082 -1.87478e-20 6.90276e-24 -1.87409e-20 0.00139507 0.997818 8.59255e-05 0.152546 2.85168 0.00139507 0.997892 0.676921 0.0010449 0.00187959 0.000859255 0.45566 0.00187959 0.435611 0.000127589 1.02 0.887428 0.534751 0.285703 1.71619e-07 3.05638e-09 2391.41 3159.62 -0.0581667 0.482117 0.277627 0.256023 -0.592868 -0.169495 0.488882 -0.268378 -0.220512 1.42 1 0 294.898 0 2.04611 1.418 0.000299959 0.872289 0.641197 0.465262 0.402995 2.04637 129.052 83.4156 18.6916 60.6228 0.0040462 0 -40 10
0.519 1.50443e-08 2.53885e-06 0.0773809 0.0773757 0.0120431 6.8383e-06 0.00115402 0.0967262 0.000656685 0.0973783 0.859423 101.877 0.245989 0.717402 4.12345 0.0540107 0.0389005 0.9611 0.0198735 0.00424233 0.0191359 0.00408366 0.00512653 0.00586407 0.205061 0.234563 57.9712 -87.8945 126.071 15.9816 145.011 0.000143183 0.267085 192.925 0.310709 0.0673885 0.00409482 0.000561571 0.00138248 0.986993 0.991736 -2.97201e-06 -85.6684 0.09298 31196.2 300.53 0.983522 0.319147 0.742762 0.742757 9.99958 2.98049e-06 1.19218e-05 0.130635 0.978897 0.930217 -0.0132933 4.89452e-06 0.500824 -1.87486e-20 6.9031e-24 -1.87417e-20 0.00139507 0.997818 8.59256e-05 0.152546 2.85168 0.00139507 0.997891 0.677033 0.00104492 0.00187959 0.000859256 0.455659 0.00187959 0.435621 0.000127592 1.02 0.887429 0.534751 0.285704 1.7162e-07 3.0564e-09 2391.39 3159.4 -0.0581507 0.482117 0.277626 0.256009 -0.592871 -0.169495 0.488929 -0.268376 -0.220561 1.421 1 0 294.914 0 2.0463 1.419 0.000299959 0.872188 0.641256 0.46491 0.403027 2.04656 129.062 83.4182 18.6917 60.6241 0.00404609 0 -40 10
0.52 1.50732e-08 2.53885e-06 0.07747 0.0774648 0.0120431 6.85146e-06 0.00115402 0.0968375 0.000656691 0.0974896 0.859472 101.876 0.245984 0.717472 4.12355 0.0540162 0.0389014 0.961099 0.0198734 0.00424243 0.0191358 0.00408374 0.00512665 0.00586418 0.205066 0.234567 57.9713 -87.8945 126.072 15.9816 145.011 0.000143173 0.267085 192.925 0.310709 0.0673885 0.00409482 0.000561571 0.00138248 0.986993 0.991736 -2.97202e-06 -85.6683 0.0929801 31196.1 300.532 0.983522 0.319147 0.742708 0.742704 9.99958 2.98049e-06 1.19219e-05 0.130636 0.978911 0.930224 -0.0132933 4.89454e-06 0.500828 -1.87494e-20 6.90343e-24 -1.87425e-20 0.00139508 0.997818 8.59257e-05 0.152547 2.85168 0.00139508 0.997891 0.677146 0.00104494 0.00187959 0.000859257 0.455659 0.00187959 0.435631 0.000127596 1.02 0.88743 0.534751 0.285705 1.7162e-07 3.05642e-09 2391.37 3159.17 -0.0581348 0.482117 0.277626 0.255994 -0.592873 -0.169495 0.488976 -0.268374 -0.220609 1.422 1 0 294.93 0 2.04648 1.42 0.000299959 0.872087 0.641314 0.464559 0.403058 2.04675 129.072 83.4208 18.6919 60.6253 0.00404598 0 -40 10
0.521 1.51022e-08 2.53885e-06 0.077559 0.0775538 0.0120431 6.86463e-06 0.00115402 0.0969487 0.000656696 0.0976008 0.859521 101.876 0.245978 0.717542 4.12365 0.0540217 0.0389023 0.961098 0.0198732 0.00424253 0.0191357 0.00408383 0.00512677 0.0058643 0.205071 0.234572 57.9713 -87.8945 126.073 15.9815 145.011 0.000143162 0.267085 192.925 0.310708 0.0673884 0.00409483 0.000561572 0.00138248 0.986992 0.991736 -2.97203e-06 -85.6683 0.0929801 31196.1 300.535 0.983522 0.319147 0.742655 0.742651 9.99958 2.98049e-06 1.19219e-05 0.130637 0.978926 0.930231 -0.0132933 4.89457e-06 0.500832 -1.87502e-20 6.90377e-24 -1.87433e-20 0.00139508 0.997818 8.59257e-05 0.152547 2.85168 0.00139508 0.99789 0.677258 0.00104496 0.0018796 0.000859257 0.455659 0.00187959 0.43564 0.000127599 1.02 0.88743 0.534751 0.285707 1.7162e-07 3.05644e-09 2391.36 3158.94 -0.058119 0.482117 0.277626 0.25598 -0.592876 -0.169495 0.489023 -0.268372 -0.220658 1.423 1 0 294.946 0 2.04667 1.421 0.000299958 0.871986 0.641373 0.464208 0.40309 2.04693 129.082 83.4234 18.692 60.6266 0.00404587 0 -40 10
0.522 1.51311e-08 2.53885e-06 0.0776479 0.0776427 0.0120431 6.87779e-06 0.00115402 0.0970599 0.000656701 0.097712 0.85957 101.876 0.245973 0.717612 4.12374 0.0540273 0.0389032 0.961097 0.0198731 0.00424263 0.0191356 0.00408391 0.00512689 0.00586442 0.205076 0.234577 57.9714 -87.8945 126.074 15.9815 145.011 0.000143152 0.267085 192.925 0.310708 0.0673884 0.00409483 0.000561572 0.00138248 0.986992 0.991736 -2.97204e-06 -85.6683 0.0929802 31196.1 300.538 0.983522 0.319147 0.742603 0.742598 9.99958 2.9805e-06 1.19219e-05 0.130638 0.97894 0.930238 -0.0132933 4.89459e-06 0.500836 -1.8751e-20 6.9041e-24 -1.87441e-20 0.00139508 0.997818 8.59258e-05 0.152547 2.85168 0.00139508 0.99789 0.677371 0.00104498 0.0018796 0.000859258 0.455659 0.0018796 0.43565 0.000127603 1.02 0.887431 0.53475 0.285708 1.7162e-07 3.05646e-09 2391.34 3158.72 -0.0581032 0.482117 0.277625 0.255966 -0.592879 -0.169495 0.489069 -0.26837 -0.220706 1.424 1 0 294.962 0 2.04686 1.422 0.000299958 0.871886 0.641431 0.463858 0.403121 2.04712 129.092 83.426 18.6922 60.6278 0.00404576 0 -40 10
0.523 1.51601e-08 2.53885e-06 0.0777367 0.0777316 0.0120431 6.89096e-06 0.00115402 0.0971709 0.000656706 0.097823 0.859619 101.876 0.245967 0.717682 4.12384 0.0540329 0.0389042 0.961096 0.019873 0.00424273 0.0191355 0.00408399 0.00512701 0.00586454 0.20508 0.234582 57.9714 -87.8945 126.075 15.9815 145.011 0.000143142 0.267085 192.925 0.310707 0.0673883 0.00409483 0.000561573 0.00138249 0.986992 0.991736 -2.97206e-06 -85.6683 0.0929803 31196.1 300.54 0.983522 0.319147 0.74255 0.742546 9.99958 2.9805e-06 1.19219e-05 0.130639 0.978954 0.930245 -0.0132933 4.89462e-06 0.50084 -1.87518e-20 6.90444e-24 -1.87449e-20 0.00139508 0.997818 8.59259e-05 0.152547 2.85168 0.00139508 0.997889 0.677483 0.001045 0.0018796 0.000859259 0.455659 0.0018796 0.435659 0.000127606 1.02 0.887432 0.53475 0.285709 1.7162e-07 3.05648e-09 2391.32 3158.49 -0.0580874 0.482117 0.277625 0.255952 -0.592881 -0.169495 0.489115 -0.268368 -0.220755 1.425 1 0 294.977 0 2.04704 1.423 0.000299958 0.871787 0.64149 0.46351 0.403153 2.04731 129.102 83.4286 18.6923 60.6291 0.00404566 0 -40 10
0.524 1.51891e-08 2.53885e-06 0.0778255 0.0778204 0.0120431 6.90412e-06 0.00115402 0.0972819 0.000656711 0.097934 0.859668 101.876 0.245962 0.717752 4.12394 0.0540384 0.0389051 0.961095 0.0198729 0.00424283 0.0191353 0.00408407 0.00512713 0.00586466 0.205085 0.234586 57.9715 -87.8945 126.076 15.9814 145.011 0.000143132 0.267085 192.925 0.310707 0.0673883 0.00409483 0.000561574 0.00138249 0.986992 0.991736 -2.97207e-06 -85.6683 0.0929803 31196.1 300.543 0.983522 0.319147 0.742498 0.742493 9.99958 2.98051e-06 1.19219e-05 0.13064 0.978969 0.930251 -0.0132933 4.89464e-06 0.500845 -1.87526e-20 6.90477e-24 -1.87457e-20 0.00139508 0.997818 8.59259e-05 0.152547 2.85168 0.00139508 0.997889 0.677595 0.00104502 0.0018796 0.000859259 0.455658 0.0018796 0.435669 0.00012761 1.02 0.887433 0.53475 0.285711 1.71621e-07 3.0565e-09 2391.31 3158.27 -0.0580718 0.482117 0.277625 0.255938 -0.592884 -0.169495 0.489161 -0.268366 -0.220803 1.426 1 0 294.993 0 2.04723 1.424 0.000299958 0.871687 0.641548 0.463162 0.403185 2.04749 129.112 83.4312 18.6925 60.6303 0.00404555 0 -40 10
0.525 1.5218e-08 2.53885e-06 0.0779142 0.0779091 0.0120431 6.91728e-06 0.00115402 0.0973928 0.000656716 0.0980449 0.859717 101.876 0.245956 0.717822 4.12404 0.054044 0.0389061 0.961094 0.0198727 0.00424292 0.0191352 0.00408415 0.00512726 0.00586478 0.20509 0.234591 57.9716 -87.8945 126.077 15.9814 145.011 0.000143122 0.267086 192.925 0.310707 0.0673883 0.00409484 0.000561574 0.00138249 0.986992 0.991736 -2.97208e-06 -85.6683 0.0929804 31196.1 300.546 0.983522 0.319147 0.742445 0.742441 9.99958 2.98051e-06 1.19219e-05 0.130641 0.978983 0.930258 -0.0132933 4.89467e-06 0.500849 -1.87534e-20 6.9051e-24 -1.87465e-20 0.00139508 0.997818 8.5926e-05 0.152547 2.85168 0.00139508 0.997888 0.677708 0.00104504 0.0018796 0.00085926 0.455658 0.0018796 0.435678 0.000127613 1.02 0.887434 0.534749 0.285712 1.71621e-07 3.05652e-09 2391.29 3158.05 -0.0580562 0.482117 0.277625 0.255924 -0.592887 -0.169495 0.489207 -0.268365 -0.22085 1.427 1 0 295.009 0 2.04742 1.425 0.000299958 0.871588 0.641607 0.462815 0.403216 2.04768 129.122 83.4337 18.6926 60.6316 0.00404544 0 -40 10
0.526 1.5247e-08 2.53885e-06 0.0780028 0.0779977 0.012043 6.93045e-06 0.00115402 0.0975035 0.000656721 0.0981557 0.859766 101.876 0.24595 0.717893 4.12414 0.0540496 0.038907 0.961093 0.0198726 0.00424302 0.0191351 0.00408424 0.00512738 0.0058649 0.205095 0.234596 57.9716 -87.8945 126.078 15.9814 145.011 0.000143112 0.267086 192.924 0.310706 0.0673882 0.00409484 0.000561575 0.00138249 0.986992 0.991736 -2.97209e-06 -85.6683 0.0929805 31196 300.549 0.983522 0.319147 0.742393 0.742389 9.99958 2.98051e-06 1.19219e-05 0.130642 0.978997 0.930265 -0.0132933 4.8947e-06 0.500853 -1.87542e-20 6.90544e-24 -1.87473e-20 0.00139508 0.997818 8.59261e-05 0.152547 2.85168 0.00139508 0.997888 0.67782 0.00104506 0.0018796 0.000859261 0.455658 0.0018796 0.435688 0.000127617 1.02 0.887435 0.534749 0.285713 1.71621e-07 3.05654e-09 2391.27 3157.82 -0.0580406 0.482117 0.277624 0.25591 -0.592889 -0.169495 0.489253 -0.268363 -0.220898 1.428 1 0 295.024 0 2.0476 1.426 0.000299958 0.87149 0.641665 0.462469 0.403248 2.04787 129.132 83.4363 18.6928 60.6328 0.00404534 0 -40 10
0.527 1.52759e-08 2.53885e-06 0.0780914 0.0780863 0.012043 6.94361e-06 0.00115402 0.0976142 0.000656727 0.0982664 0.859815 101.876 0.245945 0.717963 4.12424 0.0540552 0.038908 0.961092 0.0198725 0.00424312 0.019135 0.00408432 0.0051275 0.00586502 0.2051 0.234601 57.9717 -87.8945 126.079 15.9813 145.011 0.000143102 0.267086 192.924 0.310706 0.0673882 0.00409484 0.000561575 0.00138249 0.986992 0.991736 -2.97211e-06 -85.6683 0.0929806 31196 300.551 0.983522 0.319147 0.742341 0.742337 9.99958 2.98052e-06 1.1922e-05 0.130643 0.979011 0.930272 -0.0132933 4.89472e-06 0.500857 -1.8755e-20 6.90577e-24 -1.87481e-20 0.00139508 0.997818 8.59261e-05 0.152547 2.85168 0.00139508 0.997887 0.677932 0.00104508 0.0018796 0.000859261 0.455658 0.0018796 0.435697 0.00012762 1.02 0.887436 0.534749 0.285715 1.71621e-07 3.05656e-09 2391.26 3157.6 -0.0580251 0.482117 0.277624 0.255896 -0.592892 -0.169495 0.489298 -0.268361 -0.220945 1.429 1 0 295.04 0 2.04779 1.427 0.000299957 0.871392 0.641723 0.462124 0.403279 2.04805 129.142 83.4388 18.6929 60.634 0.00404523 0 -40 10
0.528 1.53049e-08 2.53885e-06 0.0781799 0.0781748 0.012043 6.95678e-06 0.00115402 0.0977248 0.000656732 0.098377 0.859864 101.876 0.245939 0.718034 4.12434 0.0540608 0.0389089 0.961091 0.0198724 0.00424323 0.0191349 0.0040844 0.00512762 0.00586515 0.205105 0.234606 57.9718 -87.8945 126.08 15.9813 145.011 0.000143092 0.267086 192.924 0.310706 0.0673881 0.00409484 0.000561576 0.0013825 0.986992 0.991736 -2.97212e-06 -85.6683 0.0929806 31196 300.554 0.983522 0.319147 0.74229 0.742285 9.99958 2.98052e-06 1.1922e-05 0.130644 0.979025 0.930278 -0.0132933 4.89475e-06 0.500861 -1.87559e-20 6.90611e-24 -1.8749e-20 0.00139508 0.997818 8.59262e-05 0.152548 2.85168 0.00139508 0.997887 0.678044 0.0010451 0.0018796 0.000859262 0.455658 0.0018796 0.435707 0.000127624 1.02 0.887437 0.534749 0.285716 1.71621e-07 3.05658e-09 2391.24 3157.38 -0.0580097 0.482117 0.277624 0.255882 -0.592894 -0.169495 0.489344 -0.268359 -0.220993 1.43 1 0 295.055 0 2.04798 1.428 0.000299957 0.871294 0.641782 0.46178 0.403311 2.04824 129.152 83.4414 18.6931 60.6353 0.00404513 0 -40 10
0.529 1.53339e-08 2.53885e-06 0.0782683 0.0782632 0.012043 6.96994e-06 0.00115402 0.0978354 0.000656737 0.0984875 0.859913 101.876 0.245934 0.718105 4.12445 0.0540664 0.0389099 0.96109 0.0198723 0.00424333 0.0191347 0.00408449 0.00512775 0.00586527 0.20511 0.234611 57.9718 -87.8945 126.081 15.9812 145.011 0.000143082 0.267086 192.924 0.310705 0.0673881 0.00409485 0.000561576 0.0013825 0.986992 0.991736 -2.97213e-06 -85.6683 0.0929807 31196 300.557 0.983522 0.319147 0.742238 0.742234 9.99958 2.98053e-06 1.1922e-05 0.130645 0.979039 0.930285 -0.0132933 4.89477e-06 0.500865 -1.87567e-20 6.90644e-24 -1.87498e-20 0.00139508 0.997818 8.59263e-05 0.152548 2.85168 0.00139508 0.997887 0.678156 0.00104512 0.00187961 0.000859263 0.455658 0.0018796 0.435716 0.000127627 1.02 0.887438 0.534748 0.285717 1.71622e-07 3.0566e-09 2391.23 3157.16 -0.0579944 0.482118 0.277623 0.255868 -0.592897 -0.169495 0.489389 -0.268357 -0.22104 1.431 1 0 295.07 0 2.04816 1.429 0.000299957 0.871196 0.64184 0.461437 0.403342 2.04843 129.162 83.4439 18.6932 60.6365 0.00404502 0 -40 10
0.53 1.53628e-08 2.53885e-06 0.0783566 0.0783516 0.012043 6.98311e-06 0.00115402 0.0979458 0.000656742 0.0985979 0.859963 101.875 0.245928 0.718176 4.12455 0.0540721 0.0389108 0.961089 0.0198721 0.00424343 0.0191346 0.00408457 0.00512787 0.00586539 0.205115 0.234616 57.9719 -87.8945 126.082 15.9812 145.011 0.000143072 0.267086 192.924 0.310705 0.067388 0.00409485 0.000561577 0.0013825 0.986992 0.991736 -2.97214e-06 -85.6683 0.0929808 31196 300.559 0.983522 0.319147 0.742187 0.742183 9.99958 2.98053e-06 1.1922e-05 0.130646 0.979053 0.930291 -0.0132933 4.8948e-06 0.50087 -1.87575e-20 6.90678e-24 -1.87506e-20 0.00139509 0.997818 8.59263e-05 0.152548 2.85169 0.00139509 0.997886 0.678268 0.00104514 0.00187961 0.000859263 0.455657 0.00187961 0.435726 0.000127631 1.02 0.887439 0.534748 0.285719 1.71622e-07 3.05662e-09 2391.21 3156.95 -0.0579791 0.482118 0.277623 0.255855 -0.592899 -0.169495 0.489434 -0.268355 -0.221087 1.432 1 0 295.086 0 2.04835 1.43 0.000299957 0.871099 0.641898 0.461094 0.403374 2.04861 129.172 83.4464 18.6934 60.6377 0.00404492 0 -40 10
0.531 1.53918e-08 2.53885e-06 0.0784449 0.0784399 0.012043 6.99627e-06 0.00115402 0.0980561 0.000656747 0.0987083 0.860012 101.875 0.245922 0.718247 4.12465 0.0540777 0.0389118 0.961088 0.019872 0.00424353 0.0191345 0.00408465 0.005128 0.00586551 0.20512 0.234621 57.9719 -87.8945 126.082 15.9812 145.011 0.000143062 0.267087 192.924 0.310705 0.067388 0.00409485 0.000561577 0.0013825 0.986992 0.991736 -2.97216e-06 -85.6683 0.0929808 31195.9 300.562 0.983522 0.319147 0.742136 0.742132 9.99958 2.98053e-06 1.1922e-05 0.130647 0.979067 0.930298 -0.0132933 4.89482e-06 0.500874 -1.87583e-20 6.90711e-24 -1.87514e-20 0.00139509 0.997818 8.59264e-05 0.152548 2.85169 0.00139509 0.997886 0.67838 0.00104516 0.00187961 0.000859264 0.455657 0.00187961 0.435735 0.000127634 1.02 0.88744 0.534748 0.28572 1.71622e-07 3.05663e-09 2391.19 3156.73 -0.0579639 0.482118 0.277623 0.255841 -0.592902 -0.169495 0.489479 -0.268353 -0.221133 1.433 1 0 295.101 0 2.04853 1.431 0.000299957 0.871003 0.641956 0.460753 0.403405 2.0488 129.182 83.4489 18.6935 60.6389 0.00404481 0 -40 10
0.532 1.54208e-08 2.53885e-06 0.0785331 0.0785281 0.012043 7.00943e-06 0.00115402 0.0981664 0.000656752 0.0988185 0.860062 101.875 0.245917 0.718318 4.12475 0.0540834 0.0389127 0.961087 0.0198719 0.00424363 0.0191344 0.00408474 0.00512812 0.00586564 0.205125 0.234625 57.972 -87.8945 126.083 15.9811 145.011 0.000143053 0.267087 192.924 0.310704 0.067388 0.00409485 0.000561578 0.0013825 0.986992 0.991736 -2.97217e-06 -85.6683 0.0929809 31195.9 300.565 0.983522 0.319147 0.742085 0.742081 9.99958 2.98054e-06 1.1922e-05 0.130648 0.979081 0.930305 -0.0132933 4.89485e-06 0.500878 -1.87591e-20 6.90744e-24 -1.87522e-20 0.00139509 0.997818 8.59265e-05 0.152548 2.85169 0.00139509 0.997885 0.678492 0.00104518 0.00187961 0.000859265 0.455657 0.00187961 0.435745 0.000127638 1.02 0.887441 0.534748 0.285721 1.71622e-07 3.05665e-09 2391.18 3156.51 -0.0579487 0.482118 0.277623 0.255827 -0.592905 -0.169496 0.489523 -0.268351 -0.22118 1.434 1 0 295.116 0 2.04872 1.432 0.000299956 0.870906 0.642015 0.460412 0.403436 2.04898 129.192 83.4514 18.6937 60.6401 0.00404471 0 -40 10
0.533 1.54497e-08 2.53885e-06 0.0786212 0.0786162 0.012043 7.0226e-06 0.00115402 0.0982765 0.000656757 0.0989287 0.860111 101.875 0.245911 0.718389 4.12485 0.054089 0.0389137 0.961086 0.0198718 0.00424373 0.0191342 0.00408482 0.00512825 0.00586576 0.20513 0.23463 57.9721 -87.8946 126.084 15.9811 145.011 0.000143043 0.267087 192.924 0.310704 0.0673879 0.00409486 0.000561578 0.0013825 0.986992 0.991736 -2.97218e-06 -85.6682 0.092981 31195.9 300.568 0.983522 0.319147 0.742035 0.74203 9.99958 2.98054e-06 1.19221e-05 0.130649 0.979095 0.930311 -0.0132933 4.89488e-06 0.500882 -1.87599e-20 6.90778e-24 -1.8753e-20 0.00139509 0.997818 8.59265e-05 0.152548 2.85169 0.00139509 0.997885 0.678604 0.0010452 0.00187961 0.000859265 0.455657 0.00187961 0.435754 0.000127641 1.02 0.887442 0.534747 0.285723 1.71623e-07 3.05667e-09 2391.16 3156.29 -0.0579336 0.482118 0.277622 0.255814 -0.592907 -0.169496 0.489568 -0.268349 -0.221226 1.435 1 0 295.131 0 2.04891 1.433 0.000299956 0.87081 0.642073 0.460073 0.403468 2.04917 129.202 83.4539 18.6938 60.6413 0.00404461 0 -40 10
0.534 1.54787e-08 2.53885e-06 0.0787093 0.0787043 0.0120429 7.03576e-06 0.00115402 0.0983866 0.000656762 0.0990388 0.860161 101.875 0.245905 0.71846 4.12496 0.0540947 0.0389147 0.961085 0.0198716 0.00424383 0.0191341 0.00408491 0.00512837 0.00586588 0.205135 0.234635 57.9721 -87.8946 126.085 15.9811 145.011 0.000143033 0.267087 192.923 0.310704 0.0673879 0.00409486 0.000561579 0.00138251 0.986992 0.991736 -2.97219e-06 -85.6682 0.0929811 31195.9 300.57 0.983522 0.319147 0.741984 0.74198 9.99958 2.98055e-06 1.19221e-05 0.13065 0.979109 0.930318 -0.0132933 4.8949e-06 0.500886 -1.87607e-20 6.90811e-24 -1.87538e-20 0.00139509 0.997818 8.59266e-05 0.152548 2.85169 0.00139509 0.997884 0.678716 0.00104522 0.00187961 0.000859266 0.455657 0.00187961 0.435764 0.000127645 1.02 0.887443 0.534747 0.285724 1.71623e-07 3.05669e-09 2391.14 3156.08 -0.0579185 0.482118 0.277622 0.2558 -0.59291 -0.169496 0.489612 -0.268347 -0.221272 1.436 1 0 295.146 0 2.04909 1.434 0.000299956 0.870715 0.642131 0.459734 0.403499 2.04935 129.212 83.4564 18.6939 60.6425 0.0040445 0 -40 10
0.535 1.55076e-08 2.53886e-06 0.0787973 0.0787923 0.0120429 7.04893e-06 0.00115403 0.0984966 0.000656767 0.0991488 0.860211 101.875 0.2459 0.718532 4.12506 0.0541003 0.0389157 0.961084 0.0198715 0.00424394 0.019134 0.00408499 0.0051285 0.00586601 0.20514 0.23464 57.9722 -87.8946 126.086 15.981 145.011 0.000143023 0.267087 192.923 0.310703 0.0673878 0.00409486 0.00056158 0.00138251 0.986992 0.991736 -2.97221e-06 -85.6682 0.0929811 31195.9 300.573 0.983522 0.319147 0.741934 0.741929 9.99958 2.98055e-06 1.19221e-05 0.130651 0.979123 0.930324 -0.0132933 4.89493e-06 0.500891 -1.87615e-20 6.90845e-24 -1.87546e-20 0.00139509 0.997818 8.59267e-05 0.152548 2.85169 0.00139509 0.997884 0.678828 0.00104523 0.00187961 0.000859267 0.455656 0.00187961 0.435773 0.000127649 1.02 0.887444 0.534747 0.285725 1.71623e-07 3.05671e-09 2391.13 3155.86 -0.0579036 0.482118 0.277622 0.255787 -0.592912 -0.169496 0.489656 -0.268345 -0.221318 1.437 1 0 295.161 0 2.04928 1.435 0.000299956 0.870619 0.642189 0.459396 0.40353 2.04954 129.222 83.4588 18.6941 60.6437 0.0040444 0 -40 10
0.536 1.55366e-08 2.53886e-06 0.0788852 0.0788803 0.0120429 7.06209e-06 0.00115403 0.0986065 0.000656772 0.0992587 0.86026 101.875 0.245894 0.718603 4.12516 0.054106 0.0389166 0.961083 0.0198714 0.00424404 0.0191339 0.00408508 0.00512863 0.00586613 0.205145 0.234645 57.9723 -87.8946 126.087 15.981 145.011 0.000143014 0.267087 192.923 0.310703 0.0673878 0.00409486 0.00056158 0.00138251 0.986992 0.991736 -2.97222e-06 -85.6682 0.0929812 31195.8 300.576 0.983522 0.319147 0.741884 0.741879 9.99958 2.98055e-06 1.19221e-05 0.130652 0.979137 0.930331 -0.0132933 4.89495e-06 0.500895 -1.87623e-20 6.90878e-24 -1.87554e-20 0.00139509 0.997818 8.59267e-05 0.152549 2.85169 0.00139509 0.997883 0.67894 0.00104525 0.00187961 0.000859267 0.455656 0.00187961 0.435783 0.000127652 1.02 0.887445 0.534747 0.285727 1.71623e-07 3.05673e-09 2391.11 3155.65 -0.0578886 0.482118 0.277621 0.255773 -0.592915 -0.169496 0.4897 -0.268343 -0.221364 1.438 1 0 295.176 0 2.04946 1.436 0.000299956 0.870525 0.642247 0.459059 0.403562 2.04972 129.232 83.4613 18.6942 60.6449 0.0040443 0 -40 10
0.537 1.55656e-08 2.53886e-06 0.078973 0.0789681 0.0120429 7.07525e-06 0.00115403 0.0987163 0.000656777 0.0993685 0.86031 101.875 0.245888 0.718675 4.12527 0.0541117 0.0389176 0.961082 0.0198712 0.00424414 0.0191337 0.00408516 0.00512875 0.00586626 0.20515 0.23465 57.9723 -87.8946 126.088 15.9809 145.011 0.000143004 0.267087 192.923 0.310703 0.0673877 0.00409487 0.000561581 0.00138251 0.986992 0.991735 -2.97223e-06 -85.6682 0.0929813 31195.8 300.579 0.983522 0.319147 0.741834 0.741829 9.99958 2.98056e-06 1.19221e-05 0.130653 0.97915 0.930337 -0.0132933 4.89498e-06 0.500899 -1.87631e-20 6.90911e-24 -1.87562e-20 0.00139509 0.997818 8.59268e-05 0.152549 2.85169 0.00139509 0.997883 0.679052 0.00104527 0.00187962 0.000859268 0.455656 0.00187961 0.435792 0.000127656 1.02 0.887446 0.534746 0.285728 1.71623e-07 3.05675e-09 2391.09 3155.44 -0.0578738 0.482118 0.277621 0.25576 -0.592917 -0.169496 0.489743 -0.268341 -0.22141 1.439 1 0 295.191 0 2.04965 1.437 0.000299955 0.87043 0.642305 0.458723 0.403593 2.04991 129.242 83.4637 18.6944 60.6461 0.0040442 0 -40 10
0.538 1.55945e-08 2.53886e-06 0.0790608 0.0790559 0.0120429 7.08842e-06 0.00115403 0.098826 0.000656782 0.0994782 0.86036 101.875 0.245883 0.718747 4.12537 0.0541174 0.0389186 0.961081 0.0198711 0.00424425 0.0191336 0.00408525 0.00512888 0.00586638 0.205155 0.234655 57.9724 -87.8946 126.089 15.9809 145.011 0.000142995 0.267088 192.923 0.310702 0.0673877 0.00409487 0.000561581 0.00138251 0.986992 0.991735 -2.97224e-06 -85.6682 0.0929813 31195.8 300.582 0.983522 0.319147 0.741784 0.74178 9.99958 2.98056e-06 1.19221e-05 0.130654 0.979164 0.930344 -0.0132933 4.89501e-06 0.500904 -1.87639e-20 6.90945e-24 -1.8757e-20 0.00139509 0.997818 8.59269e-05 0.152549 2.85169 0.00139509 0.997883 0.679164 0.00104529 0.00187962 0.000859269 0.455656 0.00187962 0.435801 0.000127659 1.02 0.887447 0.534746 0.285729 1.71624e-07 3.05677e-09 2391.08 3155.23 -0.057859 0.482118 0.277621 0.255747 -0.59292 -0.169496 0.489787 -0.26834 -0.221455 1.44 1 0 295.206 0 2.04983 1.438 0.000299955 0.870336 0.642363 0.458387 0.403624 2.05009 129.252 83.4662 18.6945 60.6472 0.0040441 0 -40 10
0.539 1.56235e-08 2.53886e-06 0.0791485 0.0791436 0.0120429 7.10158e-06 0.00115403 0.0989357 0.000656787 0.0995879 0.86041 101.875 0.245877 0.718819 4.12548 0.0541231 0.0389196 0.96108 0.019871 0.00424435 0.0191335 0.00408533 0.00512901 0.00586651 0.20516 0.23466 57.9724 -87.8946 126.09 15.9809 145.011 0.000142985 0.267088 192.923 0.310702 0.0673876 0.00409487 0.000561582 0.00138251 0.986992 0.991735 -2.97226e-06 -85.6682 0.0929814 31195.8 300.584 0.983522 0.319147 0.741735 0.74173 9.99958 2.98057e-06 1.19222e-05 0.130655 0.979178 0.93035 -0.0132933 4.89503e-06 0.500908 -1.87647e-20 6.90978e-24 -1.87578e-20 0.00139509 0.997818 8.59269e-05 0.152549 2.85169 0.00139509 0.997882 0.679275 0.00104531 0.00187962 0.000859269 0.455656 0.00187962 0.435811 0.000127663 1.02 0.887448 0.534746 0.285731 1.71624e-07 3.05679e-09 2391.06 3155.01 -0.0578443 0.482118 0.277621 0.255733 -0.592922 -0.169496 0.48983 -0.268338 -0.2215 1.441 1 0 295.221 0 2.05002 1.439 0.000299955 0.870242 0.642421 0.458053 0.403656 2.05028 129.262 83.4686 18.6947 60.6484 0.00404399 0 -40 10
0.54 1.56524e-08 2.53886e-06 0.0792362 0.0792313 0.0120429 7.11475e-06 0.00115403 0.0990452 0.000656791 0.0996974 0.86046 101.874 0.245871 0.718891 4.12558 0.0541288 0.0389206 0.961079 0.0198709 0.00424445 0.0191334 0.00408542 0.00512913 0.00586664 0.205165 0.234665 57.9725 -87.8946 126.091 15.9808 145.011 0.000142975 0.267088 192.923 0.310702 0.0673876 0.00409487 0.000561582 0.00138252 0.986992 0.991735 -2.97227e-06 -85.6682 0.0929815 31195.8 300.587 0.983522 0.319147 0.741685 0.741681 9.99958 2.98057e-06 1.19222e-05 0.130656 0.979191 0.930356 -0.0132933 4.89506e-06 0.500912 -1.87655e-20 6.91012e-24 -1.87586e-20 0.00139509 0.997818 8.5927e-05 0.152549 2.85169 0.00139509 0.997882 0.679387 0.00104533 0.00187962 0.00085927 0.455656 0.00187962 0.43582 0.000127666 1.02 0.887449 0.534745 0.285732 1.71624e-07 3.05681e-09 2391.04 3154.8 -0.0578296 0.482118 0.27762 0.25572 -0.592925 -0.169496 0.489873 -0.268336 -0.221545 1.442 1 0 295.235 0 2.0502 1.44 0.000299955 0.870149 0.642479 0.45772 0.403687 2.05046 129.271 83.471 18.6948 60.6496 0.00404389 0 -40 10
0.541 1.56814e-08 2.53886e-06 0.0793237 0.0793189 0.0120428 7.12791e-06 0.00115403 0.0991547 0.000656796 0.0998069 0.86051 101.874 0.245865 0.718963 4.12568 0.0541345 0.0389216 0.961078 0.0198707 0.00424456 0.0191332 0.00408551 0.00512926 0.00586676 0.205171 0.23467 57.9726 -87.8946 126.091 15.9808 145.011 0.000142966 0.267088 192.922 0.310701 0.0673876 0.00409488 0.000561583 0.00138252 0.986992 0.991735 -2.97228e-06 -85.6682 0.0929816 31195.8 300.59 0.983522 0.319147 0.741636 0.741632 9.99958 2.98057e-06 1.19222e-05 0.130657 0.979205 0.930363 -0.0132933 4.89508e-06 0.500916 -1.87663e-20 6.91045e-24 -1.87594e-20 0.0013951 0.997818 8.5927e-05 0.152549 2.85169 0.0013951 0.997881 0.679499 0.00104535 0.00187962 0.00085927 0.455655 0.00187962 0.43583 0.00012767 1.02 0.88745 0.534745 0.285733 1.71624e-07 3.05683e-09 2391.03 3154.59 -0.057815 0.482118 0.27762 0.255707 -0.592927 -0.169496 0.489916 -0.268334 -0.22159 1.443 1 0 295.25 0 2.05039 1.441 0.000299955 0.870056 0.642536 0.457387 0.403718 2.05065 129.281 83.4734 18.6949 60.6507 0.00404379 0 -40 10
0.542 1.57104e-08 2.53886e-06 0.0794112 0.0794064 0.0120428 7.14107e-06 0.00115403 0.099264 0.000656801 0.0999162 0.86056 101.874 0.24586 0.719035 4.12579 0.0541403 0.0389226 0.961077 0.0198706 0.00424466 0.0191331 0.00408559 0.00512939 0.00586689 0.205176 0.234676 57.9726 -87.8946 126.092 15.9808 145.011 0.000142957 0.267088 192.922 0.310701 0.0673875 0.00409488 0.000561583 0.00138252 0.986992 0.991735 -2.97229e-06 -85.6682 0.0929816 31195.7 300.593 0.983522 0.319147 0.741587 0.741583 9.99958 2.98058e-06 1.19222e-05 0.130658 0.979218 0.930369 -0.0132933 4.89511e-06 0.500921 -1.87671e-20 6.91078e-24 -1.87602e-20 0.0013951 0.997818 8.59271e-05 0.152549 2.85169 0.0013951 0.997881 0.67961 0.00104537 0.00187962 0.000859271 0.455655 0.00187962 0.435839 0.000127673 1.02 0.887451 0.534745 0.285735 1.71625e-07 3.05685e-09 2391.01 3154.39 -0.0578004 0.482118 0.27762 0.255694 -0.592929 -0.169496 0.489959 -0.268332 -0.221635 1.444 1 0 295.265 0 2.05057 1.442 0.000299954 0.869963 0.642594 0.457055 0.403749 2.05083 129.291 83.4758 18.6951 60.6519 0.00404369 0 -40 10
0.543 1.57393e-08 2.53886e-06 0.0794987 0.0794938 0.0120428 7.15424e-06 0.00115403 0.0993733 0.000656806 0.100026 0.86061 101.874 0.245854 0.719107 4.1259 0.054146 0.0389235 0.961076 0.0198705 0.00424477 0.019133 0.00408568 0.00512952 0.00586702 0.205181 0.234681 57.9727 -87.8946 126.093 15.9807 145.011 0.000142947 0.267088 192.922 0.3107 0.0673875 0.00409488 0.000561584 0.00138252 0.986992 0.991735 -2.97231e-06 -85.6682 0.0929817 31195.7 300.596 0.983522 0.319147 0.741538 0.741534 9.99958 2.98058e-06 1.19222e-05 0.130659 0.979232 0.930375 -0.0132933 4.89514e-06 0.500925 -1.87679e-20 6.91112e-24 -1.8761e-20 0.0013951 0.997818 8.59272e-05 0.152549 2.8517 0.0013951 0.997881 0.679722 0.00104539 0.00187962 0.000859272 0.455655 0.00187962 0.435849 0.000127677 1.02 0.887451 0.534745 0.285736 1.71625e-07 3.05687e-09 2390.99 3154.18 -0.0577859 0.482118 0.277619 0.255681 -0.592932 -0.169496 0.490001 -0.26833 -0.221679 1.445 1 0 295.279 0 2.05076 1.443 0.000299954 0.869871 0.642652 0.456724 0.40378 2.05102 129.301 83.4782 18.6952 60.6531 0.00404359 0 -40 10
0.544 1.57683e-08 2.53886e-06 0.079586 0.0795812 0.0120428 7.1674e-06 0.00115403 0.0994825 0.000656811 0.100135 0.860661 101.874 0.245848 0.71918 4.126 0.0541518 0.0389245 0.961075 0.0198703 0.00424487 0.0191329 0.00408577 0.00512965 0.00586714 0.205186 0.234686 57.9728 -87.8946 126.094 15.9807 145.011 0.000142938 0.267089 192.922 0.3107 0.0673874 0.00409488 0.000561584 0.00138252 0.986992 0.991735 -2.97232e-06 -85.6682 0.0929818 31195.7 300.599 0.983522 0.319147 0.74149 0.741485 9.99958 2.98059e-06 1.19222e-05 0.130661 0.979245 0.930382 -0.0132933 4.89516e-06 0.50093 -1.87688e-20 6.91145e-24 -1.87618e-20 0.0013951 0.997818 8.59273e-05 0.15255 2.8517 0.0013951 0.99788 0.679833 0.00104541 0.00187962 0.000859273 0.455655 0.00187962 0.435858 0.00012768 1.02 0.887452 0.534744 0.285737 1.71625e-07 3.05689e-09 2390.98 3153.97 -0.0577715 0.482118 0.277619 0.255668 -0.592934 -0.169496 0.490044 -0.268328 -0.221724 1.446 1 0 295.294 0 2.05094 1.444 0.000299954 0.869779 0.64271 0.456394 0.403811 2.0512 129.311 83.4806 18.6954 60.6542 0.0040435 0 -40 10
0.545 1.57972e-08 2.53886e-06 0.0796733 0.0796685 0.0120428 7.18056e-06 0.00115403 0.0995916 0.000656816 0.100244 0.860711 101.874 0.245842 0.719252 4.12611 0.0541575 0.0389256 0.961074 0.0198702 0.00424498 0.0191327 0.00408585 0.00512978 0.00586727 0.205191 0.234691 57.9728 -87.8946 126.095 15.9806 145.011 0.000142928 0.267089 192.922 0.3107 0.0673874 0.00409489 0.000561585 0.00138253 0.986992 0.991735 -2.97233e-06 -85.6682 0.0929818 31195.7 300.601 0.983522 0.319147 0.741441 0.741437 9.99958 2.98059e-06 1.19223e-05 0.130662 0.979259 0.930388 -0.0132933 4.89519e-06 0.500934 -1.87696e-20 6.91179e-24 -1.87626e-20 0.0013951 0.997818 8.59273e-05 0.15255 2.8517 0.0013951 0.99788 0.679945 0.00104543 0.00187962 0.000859273 0.455655 0.00187962 0.435868 0.000127684 1.02 0.887453 0.534744 0.285739 1.71625e-07 3.05691e-09 2390.96 3153.76 -0.0577571 0.482119 0.277619 0.255655 -0.592937 -0.169496 0.490086 -0.268326 -0.221768 1.447 1 0 295.308 0 2.05112 1.445 0.000299954 0.869688 0.642767 0.456065 0.403843 2.05138 129.321 83.483 18.6955 60.6554 0.0040434 0 -40 10
0.546 1.58262e-08 2.53886e-06 0.0797605 0.0797557 0.0120428 7.19373e-06 0.00115403 0.0997007 0.00065682 0.100353 0.860761 101.874 0.245837 0.719325 4.12622 0.0541633 0.0389266 0.961073 0.0198701 0.00424508 0.0191326 0.00408594 0.00512991 0.0058674 0.205196 0.234696 57.9729 -87.8946 126.096 15.9806 145.011 0.000142919 0.267089 192.922 0.310699 0.0673873 0.00409489 0.000561586 0.00138253 0.986992 0.991735 -2.97234e-06 -85.6681 0.0929819 31195.7 300.604 0.983522 0.319147 0.741393 0.741389 9.99958 2.9806e-06 1.19223e-05 0.130663 0.979272 0.930394 -0.0132933 4.89521e-06 0.500938 -1.87704e-20 6.91212e-24 -1.87634e-20 0.0013951 0.997818 8.59274e-05 0.15255 2.8517 0.0013951 0.997879 0.680056 0.00104545 0.00187963 0.000859274 0.455654 0.00187963 0.435877 0.000127687 1.02 0.887454 0.534744 0.28574 1.71625e-07 3.05693e-09 2390.94 3153.56 -0.0577428 0.482119 0.277619 0.255642 -0.592939 -0.169496 0.490128 -0.268324 -0.221812 1.448 1 0 295.322 0 2.05131 1.446 0.000299953 0.869596 0.642825 0.455737 0.403874 2.05157 129.331 83.4854 18.6956 60.6565 0.0040433 0 -40 10
0.547 1.58552e-08 2.53886e-06 0.0798477 0.0798429 0.0120428 7.20689e-06 0.00115403 0.0998096 0.000656825 0.100462 0.860812 101.874 0.245831 0.719398 4.12632 0.0541691 0.0389276 0.961072 0.01987 0.00424519 0.0191325 0.00408603 0.00513004 0.00586753 0.205202 0.234701 57.9729 -87.8946 126.097 15.9806 145.011 0.00014291 0.267089 192.922 0.310699 0.0673873 0.00409489 0.000561586 0.00138253 0.986992 0.991735 -2.97236e-06 -85.6681 0.092982 31195.6 300.607 0.983522 0.319147 0.741345 0.741341 9.99958 2.9806e-06 1.19223e-05 0.130664 0.979285 0.930401 -0.0132933 4.89524e-06 0.500943 -1.87712e-20 6.91245e-24 -1.87643e-20 0.0013951 0.997818 8.59275e-05 0.15255 2.8517 0.0013951 0.997879 0.680168 0.00104547 0.00187963 0.000859275 0.455654 0.00187963 0.435886 0.000127691 1.02 0.887455 0.534744 0.285741 1.71626e-07 3.05695e-09 2390.93 3153.35 -0.0577285 0.482119 0.277618 0.255629 -0.592942 -0.169496 0.49017 -0.268322 -0.221855 1.449 1 0 295.337 0 2.05149 1.447 0.000299953 0.869506 0.642882 0.455409 0.403905 2.05175 129.34 83.4877 18.6958 60.6576 0.0040432 0 -40 10
0.548 1.58841e-08 2.53886e-06 0.0799347 0.07993 0.0120428 7.22005e-06 0.00115403 0.0999184 0.00065683 0.100571 0.860862 101.874 0.245825 0.719471 4.12643 0.0541748 0.0389286 0.961071 0.0198698 0.0042453 0.0191323 0.00408612 0.00513017 0.00586766 0.205207 0.234706 57.973 -87.8946 126.098 15.9805 145.011 0.000142901 0.267089 192.921 0.310699 0.0673873 0.00409489 0.000561587 0.00138253 0.986992 0.991735 -2.97237e-06 -85.6681 0.0929821 31195.6 300.61 0.983522 0.319147 0.741297 0.741293 9.99958 2.9806e-06 1.19223e-05 0.130665 0.979298 0.930407 -0.0132933 4.89527e-06 0.500947 -1.8772e-20 6.91279e-24 -1.87651e-20 0.0013951 0.997818 8.59275e-05 0.15255 2.8517 0.0013951 0.997879 0.680279 0.00104549 0.00187963 0.000859275 0.455654 0.00187963 0.435896 0.000127694 1.02 0.887456 0.534743 0.285743 1.71626e-07 3.05697e-09 2390.91 3153.15 -0.0577143 0.482119 0.277618 0.255616 -0.592944 -0.169497 0.490211 -0.26832 -0.221899 1.45 1 0 295.351 0 2.05168 1.448 0.000299953 0.869415 0.64294 0.455083 0.403936 2.05194 129.35 83.4901 18.6959 60.6588 0.0040431 0 -40 10
0.549 1.59131e-08 2.53886e-06 0.0800218 0.080017 0.0120427 7.23322e-06 0.00115403 0.100027 0.000656835 0.100679 0.860913 101.873 0.245819 0.719543 4.12654 0.0541806 0.0389296 0.96107 0.0198697 0.0042454 0.0191322 0.00408621 0.0051303 0.00586779 0.205212 0.234711 57.9731 -87.8946 126.098 15.9805 145.011 0.000142892 0.267089 192.921 0.310698 0.0673872 0.0040949 0.000561587 0.00138253 0.986992 0.991735 -2.97238e-06 -85.6681 0.0929821 31195.6 300.613 0.983522 0.319147 0.74125 0.741245 9.99958 2.98061e-06 1.19223e-05 0.130666 0.979312 0.930413 -0.0132933 4.89529e-06 0.500952 -1.87728e-20 6.91312e-24 -1.87659e-20 0.0013951 0.997818 8.59276e-05 0.15255 2.8517 0.0013951 0.997878 0.68039 0.00104551 0.00187963 0.000859276 0.455654 0.00187963 0.435905 0.000127698 1.02 0.887457 0.534743 0.285744 1.71626e-07 3.05699e-09 2390.89 3152.95 -0.0577002 0.482119 0.277618 0.255603 -0.592946 -0.169497 0.490253 -0.268318 -0.221943 1.451 1 0 295.365 0 2.05186 1.449 0.000299953 0.869325 0.642998 0.454757 0.403967 2.05212 129.36 83.4924 18.696 60.6599 0.00404301 0 -40 10
0.55 1.5942e-08 2.53886e-06 0.0801087 0.080104 0.0120427 7.24638e-06 0.00115403 0.100136 0.00065684 0.100788 0.860964 101.873 0.245814 0.719617 4.12665 0.0541864 0.0389306 0.961069 0.0198696 0.00424551 0.0191321 0.00408629 0.00513043 0.00586792 0.205217 0.234717 57.9731 -87.8946 126.099 15.9805 145.011 0.000142882 0.26709 192.921 0.310698 0.0673872 0.0040949 0.000561588 0.00138253 0.986992 0.991735 -2.97239e-06 -85.6681 0.0929822 31195.6 300.616 0.983521 0.319147 0.741202 0.741198 9.99958 2.98061e-06 1.19223e-05 0.130667 0.979325 0.930419 -0.0132933 4.89532e-06 0.500956 -1.87736e-20 6.91345e-24 -1.87667e-20 0.0013951 0.997818 8.59277e-05 0.15255 2.8517 0.0013951 0.997878 0.680502 0.00104553 0.00187963 0.000859277 0.455654 0.00187963 0.435915 0.000127701 1.02 0.887458 0.534743 0.285745 1.71626e-07 3.05701e-09 2390.88 3152.74 -0.0576861 0.482119 0.277617 0.255591 -0.592949 -0.169497 0.490294 -0.268316 -0.221986 1.452 1 0 295.379 0 2.05204 1.45 0.000299953 0.869235 0.643055 0.454432 0.403998 2.0523 129.37 83.4947 18.6962 60.661 0.00404291 0 -40 10
0.551 1.5971e-08 2.53886e-06 0.0801956 0.0801908 0.0120427 7.25954e-06 0.00115403 0.100244 0.000656844 0.100897 0.861014 101.873 0.245808 0.71969 4.12675 0.0541922 0.0389316 0.961068 0.0198694 0.00424562 0.019132 0.00408638 0.00513057 0.00586805 0.205223 0.234722 57.9732 -87.8946 126.1 15.9804 145.011 0.000142873 0.26709 192.921 0.310698 0.0673871 0.0040949 0.000561588 0.00138254 0.986992 0.991735 -2.97241e-06 -85.6681 0.0929823 31195.6 300.619 0.983521 0.319147 0.741155 0.74115 9.99958 2.98062e-06 1.19224e-05 0.130668 0.979338 0.930425 -0.0132933 4.89535e-06 0.500961 -1.87744e-20 6.91379e-24 -1.87675e-20 0.0013951 0.997818 8.59277e-05 0.152551 2.8517 0.0013951 0.997877 0.680613 0.00104555 0.00187963 0.000859277 0.455653 0.00187963 0.435924 0.000127705 1.02 0.887459 0.534742 0.285747 1.71627e-07 3.05703e-09 2390.86 3152.54 -0.0576721 0.482119 0.277617 0.255578 -0.592951 -0.169497 0.490335 -0.268314 -0.222029 1.453 1 0 295.393 0 2.05223 1.451 0.000299952 0.869146 0.643112 0.454108 0.404029 2.05249 129.38 83.4971 18.6963 60.6621 0.00404281 0 -40 10
0.552 1.6e-08 2.53886e-06 0.0802824 0.0802776 0.0120427 7.27271e-06 0.00115403 0.100353 0.000656849 0.101005 0.861065 101.873 0.245802 0.719763 4.12686 0.0541981 0.0389327 0.961067 0.0198693 0.00424573 0.0191318 0.00408647 0.0051307 0.00586818 0.205228 0.234727 57.9733 -87.8946 126.101 15.9804 145.011 0.000142864 0.26709 192.921 0.310697 0.0673871 0.0040949 0.000561589 0.00138254 0.986992 0.991735 -2.97242e-06 -85.6681 0.0929824 31195.5 300.622 0.983521 0.319147 0.741108 0.741103 9.99958 2.98062e-06 1.19224e-05 0.130669 0.979351 0.930431 -0.0132933 4.89537e-06 0.500965 -1.87752e-20 6.91412e-24 -1.87683e-20 0.00139511 0.997818 8.59278e-05 0.152551 2.8517 0.00139511 0.997877 0.680724 0.00104557 0.00187963 0.000859278 0.455653 0.00187963 0.435933 0.000127708 1.02 0.88746 0.534742 0.285748 1.71627e-07 3.05705e-09 2390.84 3152.34 -0.0576582 0.482119 0.277617 0.255565 -0.592953 -0.169497 0.490376 -0.268312 -0.222072 1.454 1 0 295.407 0 2.05241 1.452 0.000299952 0.869057 0.64317 0.453785 0.40406 2.05267 129.39 83.4994 18.6965 60.6633 0.00404272 0 -40 10
0.553 1.60289e-08 2.53886e-06 0.0803691 0.0803644 0.0120427 7.28587e-06 0.00115403 0.100461 0.000656854 0.101114 0.861116 101.873 0.245796 0.719836 4.12697 0.0542039 0.0389337 0.961066 0.0198692 0.00424583 0.0191317 0.00408656 0.00513083 0.00586831 0.205233 0.234732 57.9733 -87.8946 126.102 15.9804 145.011 0.000142855 0.26709 192.921 0.310697 0.067387 0.00409491 0.00056159 0.00138254 0.986992 0.991735 -2.97243e-06 -85.6681 0.0929824 31195.5 300.625 0.983521 0.319147 0.741061 0.741056 9.99958 2.98062e-06 1.19224e-05 0.13067 0.979364 0.930437 -0.0132933 4.8954e-06 0.500969 -1.8776e-20 6.91446e-24 -1.87691e-20 0.00139511 0.997818 8.59279e-05 0.152551 2.8517 0.00139511 0.997877 0.680835 0.00104559 0.00187963 0.000859279 0.455653 0.00187963 0.435943 0.000127712 1.02 0.887461 0.534742 0.285749 1.71627e-07 3.05707e-09 2390.83 3152.14 -0.0576442 0.482119 0.277617 0.255553 -0.592956 -0.169497 0.490417 -0.26831 -0.222115 1.455 1 0 295.421 0 2.05259 1.453 0.000299952 0.868968 0.643227 0.453462 0.404091 2.05285 129.399 83.5017 18.6966 60.6644 0.00404262 0 -40 10
0.554 1.60579e-08 2.53886e-06 0.0804557 0.0804511 0.0120427 7.29903e-06 0.00115403 0.10057 0.000656858 0.101222 0.861167 101.873 0.24579 0.71991 4.12708 0.0542097 0.0389347 0.961065 0.019869 0.00424594 0.0191316 0.00408665 0.00513096 0.00586844 0.205239 0.234738 57.9734 -87.8946 126.103 15.9803 145.011 0.000142846 0.26709 192.921 0.310697 0.067387 0.00409491 0.00056159 0.00138254 0.986992 0.991735 -2.97245e-06 -85.6681 0.0929825 31195.5 300.628 0.983521 0.319147 0.741014 0.74101 9.99958 2.98063e-06 1.19224e-05 0.130672 0.979377 0.930444 -0.0132933 4.89542e-06 0.500974 -1.87768e-20 6.91479e-24 -1.87699e-20 0.00139511 0.997818 8.59279e-05 0.152551 2.8517 0.00139511 0.997876 0.680947 0.00104561 0.00187964 0.000859279 0.455653 0.00187964 0.435952 0.000127715 1.02 0.887462 0.534742 0.285751 1.71627e-07 3.05709e-09 2390.81 3151.94 -0.0576304 0.482119 0.277616 0.25554 -0.592958 -0.169497 0.490458 -0.268308 -0.222157 1.456 1 0 295.435 0 2.05278 1.454 0.000299952 0.86888 0.643285 0.453141 0.404122 2.05304 129.409 83.504 18.6967 60.6655 0.00404253 0 -40 10
0.555 1.60868e-08 2.53886e-06 0.0805423 0.0805377 0.0120427 7.3122e-06 0.00115403 0.100678 0.000656863 0.10133 0.861218 101.873 0.245784 0.719983 4.12719 0.0542156 0.0389358 0.961064 0.0198689 0.00424605 0.0191314 0.00408674 0.0051311 0.00586857 0.205244 0.234743 57.9734 -87.8946 126.104 15.9803 145.011 0.000142837 0.26709 192.921 0.310696 0.0673869 0.00409491 0.000561591 0.00138254 0.986992 0.991735 -2.97246e-06 -85.6681 0.0929826 31195.5 300.631 0.983521 0.319147 0.740968 0.740963 9.99958 2.98063e-06 1.19224e-05 0.130673 0.97939 0.93045 -0.0132933 4.89545e-06 0.500978 -1.87776e-20 6.91512e-24 -1.87707e-20 0.00139511 0.997818 8.5928e-05 0.152551 2.8517 0.00139511 0.997876 0.681058 0.00104563 0.00187964 0.00085928 0.455653 0.00187964 0.435962 0.000127719 1.02 0.887463 0.534741 0.285752 1.71627e-07 3.05711e-09 2390.79 3151.74 -0.0576166 0.482119 0.277616 0.255528 -0.59296 -0.169497 0.490498 -0.268306 -0.2222 1.457 1 0 295.449 0 2.05296 1.455 0.000299952 0.868791 0.643342 0.45282 0.404153 2.05322 129.419 83.5063 18.6969 60.6666 0.00404243 0 -40 10
0.556 1.61158e-08 2.53886e-06 0.0806289 0.0806242 0.0120426 7.32536e-06 0.00115403 0.100786 0.000656868 0.101438 0.861269 101.873 0.245779 0.720057 4.1273 0.0542214 0.0389368 0.961063 0.0198688 0.00424616 0.0191313 0.00408683 0.00513123 0.0058687 0.205249 0.234748 57.9735 -87.8946 126.104 15.9802 145.011 0.000142828 0.26709 192.92 0.310696 0.0673869 0.00409491 0.000561591 0.00138255 0.986992 0.991735 -2.97247e-06 -85.6681 0.0929827 31195.5 300.633 0.983521 0.319147 0.740921 0.740917 9.99958 2.98064e-06 1.19224e-05 0.130674 0.979403 0.930456 -0.0132933 4.89548e-06 0.500983 -1.87784e-20 6.91546e-24 -1.87715e-20 0.00139511 0.997818 8.59281e-05 0.152551 2.85171 0.00139511 0.997875 0.681169 0.00104565 0.00187964 0.000859281 0.455652 0.00187964 0.435971 0.000127722 1.02 0.887464 0.534741 0.285753 1.71628e-07 3.05713e-09 2390.78 3151.54 -0.0576029 0.482119 0.277616 0.255515 -0.592963 -0.169497 0.490538 -0.268305 -0.222242 1.458 1 0 295.463 0 2.05314 1.456 0.000299951 0.868704 0.643399 0.4525 0.404183 2.0534 129.429 83.5085 18.697 60.6677 0.00404234 0 -40 10
0.557 1.61447e-08 2.53886e-06 0.0807153 0.0807107 0.0120426 7.33852e-06 0.00115403 0.100894 0.000656872 0.101546 0.86132 101.873 0.245773 0.720131 4.12741 0.0542273 0.0389378 0.961062 0.0198686 0.00424627 0.0191312 0.00408692 0.00513137 0.00586884 0.205255 0.234753 57.9736 -87.8946 126.105 15.9802 145.011 0.000142819 0.267091 192.92 0.310695 0.0673869 0.00409492 0.000561592 0.00138255 0.986992 0.991735 -2.97248e-06 -85.6681 0.0929827 31195.5 300.636 0.983521 0.319147 0.740875 0.74087 9.99958 2.98064e-06 1.19225e-05 0.130675 0.979416 0.930462 -0.0132933 4.8955e-06 0.500988 -1.87792e-20 6.91579e-24 -1.87723e-20 0.00139511 0.997818 8.59281e-05 0.152551 2.85171 0.00139511 0.997875 0.68128 0.00104567 0.00187964 0.000859281 0.455652 0.00187964 0.43598 0.000127726 1.02 0.887465 0.534741 0.285755 1.71628e-07 3.05715e-09 2390.76 3151.35 -0.0575892 0.482119 0.277615 0.255503 -0.592965 -0.169497 0.490578 -0.268303 -0.222284 1.459 1 0 295.477 0 2.05333 1.457 0.000299951 0.868616 0.643456 0.452181 0.404214 2.05358 129.439 83.5108 18.6971 60.6688 0.00404224 0 -40 10
0.558 1.61737e-08 2.53886e-06 0.0808017 0.0807971 0.0120426 7.35169e-06 0.00115403 0.101002 0.000656877 0.101654 0.861371 101.872 0.245767 0.720205 4.12752 0.0542331 0.0389389 0.961061 0.0198685 0.00424638 0.019131 0.00408701 0.0051315 0.00586897 0.20526 0.234759 57.9736 -87.8946 126.106 15.9802 145.011 0.00014281 0.267091 192.92 0.310695 0.0673868 0.00409492 0.000561592 0.00138255 0.986992 0.991735 -2.9725e-06 -85.6681 0.0929828 31195.4 300.639 0.983521 0.319147 0.740829 0.740824 9.99958 2.98064e-06 1.19225e-05 0.130676 0.979429 0.930468 -0.0132933 4.89553e-06 0.500992 -1.878e-20 6.91612e-24 -1.87731e-20 0.00139511 0.997818 8.59282e-05 0.152551 2.85171 0.00139511 0.997875 0.681391 0.00104569 0.00187964 0.000859282 0.455652 0.00187964 0.43599 0.000127729 1.02 0.887466 0.534741 0.285756 1.71628e-07 3.05717e-09 2390.74 3151.15 -0.0575756 0.482119 0.277615 0.25549 -0.592967 -0.169497 0.490618 -0.268301 -0.222326 1.46 1 0 295.49 0 2.05351 1.458 0.000299951 0.868529 0.643514 0.451863 0.404245 2.05377 129.448 83.5131 18.6973 60.6699 0.00404215 0 -40 10
0.559 1.62027e-08 2.53886e-06 0.080888 0.0808834 0.0120426 7.36485e-06 0.00115403 0.10111 0.000656882 0.101762 0.861422 101.872 0.245761 0.720279 4.12763 0.054239 0.0389399 0.96106 0.0198684 0.00424649 0.0191309 0.0040871 0.00513164 0.0058691 0.205265 0.234764 57.9737 -87.8947 126.107 15.9801 145.011 0.000142802 0.267091 192.92 0.310695 0.0673868 0.00409492 0.000561593 0.00138255 0.986992 0.991735 -2.97251e-06 -85.668 0.0929829 31195.4 300.642 0.983521 0.319147 0.740783 0.740779 9.99958 2.98065e-06 1.19225e-05 0.130677 0.979442 0.930474 -0.0132933 4.89556e-06 0.500997 -1.87808e-20 6.91646e-24 -1.87739e-20 0.00139511 0.997818 8.59283e-05 0.152552 2.85171 0.00139511 0.997874 0.681502 0.00104571 0.00187964 0.000859283 0.455652 0.00187964 0.435999 0.000127733 1.02 0.887467 0.53474 0.285758 1.71628e-07 3.05719e-09 2390.73 3150.96 -0.0575621 0.482119 0.277615 0.255478 -0.59297 -0.169497 0.490658 -0.268299 -0.222367 1.461 1 0 295.504 0 2.05369 1.459 0.000299951 0.868443 0.643571 0.451545 0.404276 2.05395 129.458 83.5153 18.6974 60.671 0.00404205 0 -40 10
0.56 1.62316e-08 2.53886e-06 0.0809742 0.0809696 0.0120426 7.37801e-06 0.00115403 0.101218 0.000656886 0.10187 0.861473 101.872 0.245755 0.720353 4.12775 0.0542449 0.038941 0.961059 0.0198682 0.0042466 0.0191308 0.00408719 0.00513177 0.00586924 0.205271 0.234769 57.9738 -87.8947 126.108 15.9801 145.011 0.000142793 0.267091 192.92 0.310694 0.0673867 0.00409492 0.000561593 0.00138255 0.986992 0.991735 -2.97252e-06 -85.668 0.0929829 31195.4 300.645 0.983521 0.319147 0.740737 0.740733 9.99958 2.98065e-06 1.19225e-05 0.130678 0.979454 0.93048 -0.0132933 4.89558e-06 0.501001 -1.87816e-20 6.91679e-24 -1.87747e-20 0.00139511 0.997818 8.59283e-05 0.152552 2.85171 0.00139511 0.997874 0.681613 0.00104572 0.00187964 0.000859283 0.455652 0.00187964 0.436008 0.000127736 1.02 0.887468 0.53474 0.285759 1.71629e-07 3.05721e-09 2390.71 3150.76 -0.0575486 0.482119 0.277615 0.255466 -0.592972 -0.169497 0.490698 -0.268297 -0.222409 1.462 1 0 295.517 0 2.05387 1.46 0.000299951 0.868357 0.643628 0.451229 0.404307 2.05413 129.468 83.5176 18.6975 60.672 0.00404196 0 -40 10
0.561 1.62606e-08 2.53886e-06 0.0810604 0.0810558 0.0120426 7.39117e-06 0.00115403 0.101326 0.000656891 0.101978 0.861525 101.872 0.245749 0.720427 4.12786 0.0542508 0.038942 0.961058 0.0198681 0.00424671 0.0191306 0.00408729 0.00513191 0.00586937 0.205276 0.234775 57.9738 -87.8947 126.108 15.9801 145.012 0.000142784 0.267091 192.92 0.310694 0.0673867 0.00409493 0.000561594 0.00138255 0.986992 0.991735 -2.97254e-06 -85.668 0.092983 31195.4 300.648 0.983521 0.319147 0.740692 0.740687 9.99958 2.98066e-06 1.19225e-05 0.130679 0.979467 0.930485 -0.0132933 4.89561e-06 0.501006 -1.87824e-20 6.91712e-24 -1.87755e-20 0.00139511 0.997818 8.59284e-05 0.152552 2.85171 0.00139511 0.997874 0.681723 0.00104574 0.00187964 0.000859284 0.455652 0.00187964 0.436018 0.00012774 1.02 0.887469 0.53474 0.28576 1.71629e-07 3.05723e-09 2390.7 3150.57 -0.0575351 0.48212 0.277614 0.255454 -0.592974 -0.169497 0.490737 -0.268295 -0.22245 1.463 1 0 295.531 0 2.05406 1.461 0.00029995 0.868271 0.643685 0.450913 0.404338 2.05431 129.478 83.5198 18.6976 60.6731 0.00404187 0 -40 10
0.562 1.62895e-08 2.53886e-06 0.0811465 0.081142 0.0120426 7.40434e-06 0.00115403 0.101433 0.000656895 0.102085 0.861576 101.872 0.245743 0.720501 4.12797 0.0542567 0.0389431 0.961057 0.019868 0.00424682 0.0191305 0.00408738 0.00513204 0.0058695 0.205282 0.23478 57.9739 -87.8947 126.109 15.98 145.012 0.000142775 0.267091 192.92 0.310694 0.0673866 0.00409493 0.000561595 0.00138256 0.986992 0.991735 -2.97255e-06 -85.668 0.0929831 31195.4 300.651 0.983521 0.319147 0.740646 0.740642 9.99958 2.98066e-06 1.19225e-05 0.13068 0.97948 0.930491 -0.0132933 4.89564e-06 0.50101 -1.87832e-20 6.91746e-24 -1.87763e-20 0.00139512 0.997818 8.59285e-05 0.152552 2.85171 0.00139512 0.997873 0.681834 0.00104576 0.00187965 0.000859285 0.455651 0.00187965 0.436027 0.000127743 1.02 0.88747 0.534739 0.285762 1.71629e-07 3.05725e-09 2390.68 3150.37 -0.0575217 0.48212 0.277614 0.255442 -0.592976 -0.169497 0.490776 -0.268293 -0.222491 1.464 1 0 295.544 0 2.05424 1.462 0.00029995 0.868185 0.643742 0.450598 0.404368 2.0545 129.487 83.522 18.6978 60.6742 0.00404178 0 -40 10
0.563 1.63185e-08 2.53886e-06 0.0812326 0.081228 0.0120426 7.4175e-06 0.00115403 0.101541 0.0006569 0.102193 0.861627 101.872 0.245737 0.720576 4.12808 0.0542626 0.0389442 0.961056 0.0198678 0.00424693 0.0191304 0.00408747 0.00513218 0.00586964 0.205287 0.234786 57.974 -87.8947 126.11 15.98 145.012 0.000142767 0.267092 192.919 0.310693 0.0673866 0.00409493 0.000561595 0.00138256 0.986992 0.991735 -2.97256e-06 -85.668 0.0929832 31195.3 300.654 0.983521 0.319147 0.740601 0.740597 9.99958 2.98067e-06 1.19226e-05 0.130682 0.979492 0.930497 -0.0132933 4.89566e-06 0.501015 -1.8784e-20 6.91779e-24 -1.87771e-20 0.00139512 0.997818 8.59285e-05 0.152552 2.85171 0.00139512 0.997873 0.681945 0.00104578 0.00187965 0.000859285 0.455651 0.00187965 0.436036 0.000127747 1.02 0.887471 0.534739 0.285763 1.71629e-07 3.05727e-09 2390.66 3150.18 -0.0575084 0.48212 0.277614 0.255429 -0.592979 -0.169498 0.490815 -0.268291 -0.222532 1.465 1 0 295.558 0 2.05442 1.463 0.00029995 0.8681 0.643799 0.450284 0.404399 2.05468 129.497 83.5242 18.6979 60.6753 0.00404168 0 -40 10
0.564 1.63475e-08 2.53886e-06 0.0813185 0.081314 0.0120425 7.43066e-06 0.00115403 0.101648 0.000656905 0.1023 0.861679 101.872 0.245731 0.72065 4.12819 0.0542685 0.0389452 0.961055 0.0198677 0.00424704 0.0191302 0.00408756 0.00513232 0.00586977 0.205293 0.234791 57.974 -87.8947 126.111 15.9799 145.012 0.000142758 0.267092 192.919 0.310693 0.0673865 0.00409493 0.000561596 0.00138256 0.986992 0.991735 -2.97257e-06 -85.668 0.0929832 31195.3 300.657 0.983521 0.319147 0.740556 0.740552 9.99958 2.98067e-06 1.19226e-05 0.130683 0.979505 0.930503 -0.0132933 4.89569e-06 0.50102 -1.87848e-20 6.91812e-24 -1.87779e-20 0.00139512 0.997818 8.59286e-05 0.152552 2.85171 0.00139512 0.997873 0.682056 0.0010458 0.00187965 0.000859286 0.455651 0.00187965 0.436046 0.00012775 1.02 0.887472 0.534739 0.285764 1.7163e-07 3.05729e-09 2390.65 3149.99 -0.0574951 0.48212 0.277613 0.255417 -0.592981 -0.169498 0.490854 -0.268289 -0.222573 1.466 1 0 295.571 0 2.0546 1.464 0.00029995 0.868015 0.643856 0.449971 0.40443 2.05486 129.507 83.5264 18.698 60.6763 0.00404159 0 -40 10
0.565 1.63764e-08 2.53886e-06 0.0814044 0.0813999 0.0120425 7.44382e-06 0.00115403 0.101756 0.000656909 0.102408 0.86173 101.872 0.245726 0.720725 4.12831 0.0542744 0.0389463 0.961054 0.0198675 0.00424715 0.0191301 0.00408765 0.00513245 0.00586991 0.205298 0.234796 57.9741 -87.8947 126.112 15.9799 145.012 0.000142749 0.267092 192.919 0.310693 0.0673865 0.00409494 0.000561596 0.00138256 0.986991 0.991735 -2.97259e-06 -85.668 0.0929833 31195.3 300.66 0.983521 0.319147 0.740512 0.740507 9.99958 2.98067e-06 1.19226e-05 0.130684 0.979518 0.930509 -0.0132933 4.89572e-06 0.501024 -1.87856e-20 6.91846e-24 -1.87787e-20 0.00139512 0.997818 8.59287e-05 0.152552 2.85171 0.00139512 0.997872 0.682166 0.00104582 0.00187965 0.000859287 0.455651 0.00187965 0.436055 0.000127754 1.02 0.887473 0.534739 0.285766 1.7163e-07 3.05731e-09 2390.63 3149.8 -0.0574819 0.48212 0.277613 0.255405 -0.592983 -0.169498 0.490893 -0.268287 -0.222614 1.467 1 0 295.584 0 2.05479 1.465 0.000299949 0.86793 0.643913 0.449658 0.404461 2.05504 129.517 83.5286 18.6982 60.6774 0.0040415 0 -40 10
0.566 1.64054e-08 2.53886e-06 0.0814903 0.0814857 0.0120425 7.45699e-06 0.00115403 0.101863 0.000656914 0.102515 0.861782 101.872 0.24572 0.7208 4.12842 0.0542804 0.0389474 0.961053 0.0198674 0.00424727 0.01913 0.00408775 0.00513259 0.00587004 0.205304 0.234802 57.9741 -87.8947 126.113 15.9799 145.012 0.000142741 0.267092 192.919 0.310692 0.0673865 0.00409494 0.000561597 0.00138256 0.986991 0.991735 -2.9726e-06 -85.668 0.0929834 31195.3 300.663 0.983521 0.319147 0.740467 0.740463 9.99958 2.98068e-06 1.19226e-05 0.130685 0.97953 0.930515 -0.0132933 4.89574e-06 0.501029 -1.87864e-20 6.91879e-24 -1.87795e-20 0.00139512 0.997818 8.59287e-05 0.152552 2.85171 0.00139512 0.997872 0.682277 0.00104584 0.00187965 0.000859287 0.455651 0.00187965 0.436064 0.000127757 1.02 0.887474 0.534738 0.285767 1.7163e-07 3.05733e-09 2390.61 3149.61 -0.0574688 0.48212 0.277613 0.255393 -0.592985 -0.169498 0.490932 -0.268285 -0.222655 1.468 1 0 295.598 0 2.05497 1.466 0.000299949 0.867846 0.64397 0.449346 0.404491 2.05522 129.526 83.5308 18.6983 60.6785 0.00404141 0 -40 10
0.567 1.64343e-08 2.53886e-06 0.081576 0.0815715 0.0120425 7.47015e-06 0.00115403 0.10197 0.000656918 0.102622 0.861834 101.871 0.245714 0.720875 4.12854 0.0542863 0.0389484 0.961052 0.0198673 0.00424738 0.0191298 0.00408784 0.00513273 0.00587018 0.205309 0.234807 57.9742 -87.8947 126.113 15.9798 145.012 0.000142732 0.267092 192.919 0.310692 0.0673864 0.00409494 0.000561597 0.00138257 0.986991 0.991735 -2.97261e-06 -85.668 0.0929835 31195.3 300.666 0.983521 0.319147 0.740422 0.740418 9.99958 2.98068e-06 1.19226e-05 0.130686 0.979543 0.930521 -0.0132933 4.89577e-06 0.501034 -1.87872e-20 6.91912e-24 -1.87803e-20 0.00139512 0.997818 8.59288e-05 0.152553 2.85171 0.00139512 0.997871 0.682388 0.00104586 0.00187965 0.000859288 0.45565 0.00187965 0.436074 0.000127761 1.02 0.887475 0.534738 0.285768 1.7163e-07 3.05735e-09 2390.6 3149.42 -0.0574557 0.48212 0.277613 0.255381 -0.592988 -0.169498 0.49097 -0.268283 -0.222695 1.469 1 0 295.611 0 2.05515 1.467 0.000299949 0.867762 0.644027 0.449036 0.404522 2.0554 129.536 83.533 18.6984 60.6795 0.00404132 0 -40 10
0.568 1.64633e-08 2.53886e-06 0.0816617 0.0816572 0.0120425 7.48331e-06 0.00115403 0.102077 0.000656923 0.102729 0.861886 101.871 0.245708 0.72095 4.12865 0.0542923 0.0389495 0.96105 0.0198671 0.00424749 0.0191297 0.00408793 0.00513287 0.00587032 0.205315 0.234813 57.9743 -87.8947 126.114 15.9798 145.012 0.000142724 0.267092 192.919 0.310691 0.0673864 0.00409494 0.000561598 0.00138257 0.986991 0.991735 -2.97263e-06 -85.668 0.0929835 31195.2 300.67 0.983521 0.319147 0.740378 0.740374 9.99958 2.98069e-06 1.19226e-05 0.130687 0.979555 0.930526 -0.0132933 4.8958e-06 0.501038 -1.8788e-20 6.91946e-24 -1.87811e-20 0.00139512 0.997818 8.59289e-05 0.152553 2.85171 0.00139512 0.997871 0.682498 0.00104588 0.00187965 0.000859289 0.45565 0.00187965 0.436083 0.000127764 1.02 0.887476 0.534738 0.28577 1.7163e-07 3.05737e-09 2390.58 3149.23 -0.0574426 0.48212 0.277612 0.25537 -0.59299 -0.169498 0.491008 -0.268281 -0.222735 1.47 1 0 295.624 0 2.05533 1.468 0.000299949 0.867678 0.644084 0.448725 0.404553 2.05559 129.546 83.5352 18.6985 60.6806 0.00404123 0 -40 10
0.569 1.64922e-08 2.53886e-06 0.0817473 0.0817428 0.0120425 7.49647e-06 0.00115403 0.102184 0.000656927 0.102836 0.861937 101.871 0.245702 0.721025 4.12876 0.0542982 0.0389506 0.961049 0.019867 0.0042476 0.0191295 0.00408803 0.00513301 0.00587045 0.20532 0.234818 57.9743 -87.8947 126.115 15.9797 145.012 0.000142715 0.267093 192.919 0.310691 0.0673863 0.00409495 0.000561599 0.00138257 0.986991 0.991735 -2.97264e-06 -85.668 0.0929836 31195.2 300.673 0.983521 0.319147 0.740334 0.74033 9.99958 2.98069e-06 1.19227e-05 0.130688 0.979567 0.930532 -0.0132933 4.89582e-06 0.501043 -1.87888e-20 6.91979e-24 -1.87819e-20 0.00139512 0.997818 8.5929e-05 0.152553 2.85172 0.00139512 0.997871 0.682609 0.0010459 0.00187966 0.00085929 0.45565 0.00187965 0.436092 0.000127768 1.02 0.887477 0.534737 0.285771 1.71631e-07 3.05739e-09 2390.56 3149.04 -0.0574296 0.48212 0.277612 0.255358 -0.592992 -0.169498 0.491046 -0.268279 -0.222775 1.471 1 0 295.637 0 2.05551 1.469 0.000299949 0.867595 0.64414 0.448416 0.404583 2.05577 129.555 83.5374 18.6987 60.6816 0.00404114 0 -40 10
0.57 1.65212e-08 2.53886e-06 0.0818329 0.0818284 0.0120425 7.50964e-06 0.00115403 0.102291 0.000656932 0.102943 0.861989 101.871 0.245696 0.7211 4.12888 0.0543042 0.0389517 0.961048 0.0198669 0.00424772 0.0191294 0.00408812 0.00513315 0.00587059 0.205326 0.234824 57.9744 -87.8947 126.116 15.9797 145.012 0.000142707 0.267093 192.918 0.310691 0.0673863 0.00409495 0.000561599 0.00138257 0.986991 0.991735 -2.97265e-06 -85.668 0.0929837 31195.2 300.676 0.983521 0.319147 0.74029 0.740286 9.99958 2.9807e-06 1.19227e-05 0.13069 0.97958 0.930538 -0.0132933 4.89585e-06 0.501048 -1.87896e-20 6.92013e-24 -1.87827e-20 0.00139512 0.997818 8.5929e-05 0.152553 2.85172 0.00139512 0.99787 0.682719 0.00104592 0.00187966 0.00085929 0.45565 0.00187966 0.436102 0.000127771 1.02 0.887478 0.534737 0.285773 1.71631e-07 3.05742e-09 2390.55 3148.85 -0.0574167 0.48212 0.277612 0.255346 -0.592994 -0.169498 0.491084 -0.268277 -0.222815 1.472 1 0 295.65 0 2.05569 1.47 0.000299948 0.867512 0.644197 0.448108 0.404614 2.05595 129.565 83.5395 18.6988 60.6826 0.00404105 0 -40 10
0.571 1.65502e-08 2.53886e-06 0.0819184 0.0819139 0.0120424 7.5228e-06 0.00115403 0.102398 0.000656936 0.10305 0.862041 101.871 0.24569 0.721175 4.12899 0.0543102 0.0389528 0.961047 0.0198667 0.00424783 0.0191293 0.00408822 0.00513328 0.00587073 0.205331 0.234829 57.9745 -87.8947 126.117 15.9797 145.012 0.000142698 0.267093 192.918 0.31069 0.0673862 0.00409495 0.0005616 0.00138257 0.986991 0.991735 -2.97267e-06 -85.6679 0.0929838 31195.2 300.679 0.983521 0.319147 0.740246 0.740242 9.99958 2.9807e-06 1.19227e-05 0.130691 0.979592 0.930544 -0.0132933 4.89588e-06 0.501052 -1.87904e-20 6.92046e-24 -1.87835e-20 0.00139512 0.997818 8.59291e-05 0.152553 2.85172 0.00139512 0.99787 0.68283 0.00104594 0.00187966 0.000859291 0.45565 0.00187966 0.436111 0.000127775 1.02 0.887479 0.534737 0.285774 1.71631e-07 3.05744e-09 2390.53 3148.67 -0.0574038 0.48212 0.277611 0.255334 -0.592996 -0.169498 0.491122 -0.268275 -0.222855 1.473 1 0 295.663 0 2.05587 1.471 0.000299948 0.86743 0.644254 0.4478 0.404644 2.05613 129.575 83.5417 18.6989 60.6837 0.00404096 0 -40 10
0.572 1.65791e-08 2.53886e-06 0.0820038 0.0819993 0.0120424 7.53596e-06 0.00115403 0.102505 0.00065694 0.103157 0.862093 101.871 0.245684 0.72125 4.12911 0.0543161 0.0389539 0.961046 0.0198666 0.00424794 0.0191291 0.00408831 0.00513342 0.00587087 0.205337 0.234835 57.9745 -87.8947 126.117 15.9796 145.012 0.00014269 0.267093 192.918 0.31069 0.0673862 0.00409495 0.0005616 0.00138258 0.986991 0.991735 -2.97268e-06 -85.6679 0.0929838 31195.2 300.682 0.983521 0.319147 0.740203 0.740198 9.99958 2.9807e-06 1.19227e-05 0.130692 0.979604 0.930549 -0.0132933 4.8959e-06 0.501057 -1.87912e-20 6.92079e-24 -1.87843e-20 0.00139513 0.997818 8.59292e-05 0.152553 2.85172 0.00139513 0.99787 0.68294 0.00104596 0.00187966 0.000859292 0.455649 0.00187966 0.43612 0.000127778 1.02 0.88748 0.534737 0.285775 1.71631e-07 3.05746e-09 2390.51 3148.48 -0.057391 0.48212 0.277611 0.255323 -0.592999 -0.169498 0.491159 -0.268273 -0.222894 1.474 1 0 295.676 0 2.05606 1.472 0.000299948 0.867347 0.644311 0.447493 0.404675 2.05631 129.585 83.5438 18.699 60.6847 0.00404087 0 -40 10
0.573 1.66081e-08 2.53887e-06 0.0820891 0.0820847 0.0120424 7.54912e-06 0.00115403 0.102611 0.000656945 0.103264 0.862145 101.871 0.245678 0.721326 4.12923 0.0543221 0.038955 0.961045 0.0198664 0.00424806 0.019129 0.0040884 0.00513357 0.00587101 0.205343 0.23484 57.9746 -87.8947 126.118 15.9796 145.012 0.000142681 0.267093 192.918 0.31069 0.0673861 0.00409496 0.000561601 0.00138258 0.986991 0.991735 -2.97269e-06 -85.6679 0.0929839 31195.1 300.685 0.983521 0.319147 0.740159 0.740155 9.99958 2.98071e-06 1.19227e-05 0.130693 0.979617 0.930555 -0.0132933 4.89593e-06 0.501062 -1.8792e-20 6.92113e-24 -1.87851e-20 0.00139513 0.997818 8.59292e-05 0.152553 2.85172 0.00139513 0.997869 0.683051 0.00104598 0.00187966 0.000859292 0.455649 0.00187966 0.43613 0.000127782 1.02 0.887481 0.534736 0.285777 1.71632e-07 3.05748e-09 2390.5 3148.29 -0.0573782 0.48212 0.277611 0.255311 -0.593001 -0.169498 0.491197 -0.268271 -0.222934 1.475 1 0 295.689 0 2.05624 1.473 0.000299948 0.867265 0.644367 0.447187 0.404705 2.05649 129.594 83.546 18.6992 60.6857 0.00404078 0 -40 10
0.574 1.6637e-08 2.53887e-06 0.0821744 0.08217 0.0120424 7.56229e-06 0.00115403 0.102718 0.000656949 0.10337 0.862197 101.871 0.245672 0.721401 4.12934 0.0543281 0.0389561 0.961044 0.0198663 0.00424817 0.0191289 0.0040885 0.00513371 0.00587115 0.205348 0.234846 57.9746 -87.8947 126.119 15.9796 145.012 0.000142673 0.267093 192.918 0.310689 0.0673861 0.00409496 0.000561602 0.00138258 0.986991 0.991735 -2.9727e-06 -85.6679 0.092984 31195.1 300.688 0.983521 0.319147 0.740116 0.740112 9.99958 2.98071e-06 1.19227e-05 0.130694 0.979629 0.930561 -0.0132933 4.89596e-06 0.501067 -1.87928e-20 6.92146e-24 -1.87859e-20 0.00139513 0.997818 8.59293e-05 0.152554 2.85172 0.00139513 0.997869 0.683161 0.001046 0.00187966 0.000859293 0.455649 0.00187966 0.436139 0.000127785 1.02 0.887482 0.534736 0.285778 1.71632e-07 3.0575e-09 2390.48 3148.11 -0.0573655 0.48212 0.277611 0.255299 -0.593003 -0.169498 0.491234 -0.268269 -0.222973 1.476 1 0 295.702 0 2.05642 1.474 0.000299947 0.867184 0.644424 0.446881 0.404736 2.05667 129.604 83.5481 18.6993 60.6868 0.00404069 0 -40 10
0.575 1.6666e-08 2.53887e-06 0.0822596 0.0822552 0.0120424 7.57545e-06 0.00115403 0.102825 0.000656954 0.103477 0.862249 101.871 0.245666 0.721477 4.12946 0.0543341 0.0389572 0.961043 0.0198662 0.00424829 0.0191287 0.00408859 0.00513385 0.00587128 0.205354 0.234851 57.9747 -87.8947 126.12 15.9795 145.012 0.000142665 0.267094 192.918 0.310689 0.067386 0.00409496 0.000561602 0.00138258 0.986991 0.991735 -2.97272e-06 -85.6679 0.0929841 31195.1 300.691 0.983521 0.319147 0.740073 0.740069 9.99958 2.98072e-06 1.19228e-05 0.130695 0.979641 0.930566 -0.0132933 4.89598e-06 0.501071 -1.87936e-20 6.92179e-24 -1.87867e-20 0.00139513 0.997818 8.59294e-05 0.152554 2.85172 0.00139513 0.997869 0.683271 0.00104602 0.00187966 0.000859294 0.455649 0.00187966 0.436148 0.000127789 1.02 0.887483 0.534736 0.285779 1.71632e-07 3.05752e-09 2390.46 3147.93 -0.0573528 0.48212 0.27761 0.255288 -0.593005 -0.169498 0.491271 -0.268267 -0.223012 1.477 1 0 295.714 0 2.0566 1.475 0.000299947 0.867103 0.644481 0.446577 0.404766 2.05685 129.614 83.5502 18.6994 60.6878 0.00404061 0 -40 10
0.576 1.66949e-08 2.53887e-06 0.0823448 0.0823404 0.0120424 7.58861e-06 0.00115403 0.102931 0.000656958 0.103583 0.862302 101.87 0.24566 0.721553 4.12958 0.0543402 0.0389583 0.961042 0.019866 0.0042484 0.0191286 0.00408869 0.00513399 0.00587142 0.20536 0.234857 57.9748 -87.8947 126.12 15.9795 145.012 0.000142656 0.267094 192.918 0.310688 0.067386 0.00409497 0.000561603 0.00138258 0.986991 0.991735 -2.97273e-06 -85.6679 0.0929841 31195.1 300.694 0.983521 0.319147 0.74003 0.740026 9.99958 2.98072e-06 1.19228e-05 0.130697 0.979653 0.930572 -0.0132933 4.89601e-06 0.501076 -1.87944e-20 6.92213e-24 -1.87875e-20 0.00139513 0.997818 8.59294e-05 0.152554 2.85172 0.00139513 0.997868 0.683382 0.00104604 0.00187966 0.000859294 0.455649 0.00187966 0.436157 0.000127792 1.02 0.887484 0.534736 0.285781 1.71632e-07 3.05754e-09 2390.45 3147.74 -0.0573402 0.482121 0.27761 0.255276 -0.593007 -0.169498 0.491308 -0.268265 -0.223051 1.478 1 0 295.727 0 2.05678 1.476 0.000299947 0.867022 0.644537 0.446273 0.404797 2.05703 129.623 83.5523 18.6995 60.6888 0.00404052 0 -40 10
0.577 1.67239e-08 2.53887e-06 0.0824298 0.0824255 0.0120424 7.60177e-06 0.00115403 0.103037 0.000656962 0.10369 0.862354 101.87 0.245654 0.721629 4.12969 0.0543462 0.0389594 0.961041 0.0198659 0.00424852 0.0191284 0.00408879 0.00513413 0.00587156 0.205365 0.234863 57.9748 -87.8947 126.121 15.9794 145.012 0.000142648 0.267094 192.917 0.310688 0.067386 0.00409497 0.000561603 0.00138258 0.986991 0.991735 -2.97274e-06 -85.6679 0.0929842 31195.1 300.697 0.983521 0.319147 0.739987 0.739983 9.99958 2.98073e-06 1.19228e-05 0.130698 0.979665 0.930577 -0.0132933 4.89604e-06 0.501081 -1.87952e-20 6.92246e-24 -1.87883e-20 0.00139513 0.997818 8.59295e-05 0.152554 2.85172 0.00139513 0.997868 0.683492 0.00104606 0.00187967 0.000859295 0.455648 0.00187966 0.436167 0.000127796 1.02 0.887485 0.534735 0.285782 1.71633e-07 3.05756e-09 2390.43 3147.56 -0.0573277 0.482121 0.27761 0.255265 -0.593009 -0.169498 0.491345 -0.268263 -0.223089 1.479 1 0 295.74 0 2.05696 1.477 0.000299947 0.866941 0.644594 0.44597 0.404827 2.05721 129.633 83.5544 18.6997 60.6898 0.00404043 0 -40 10
0.578 1.67529e-08 2.53887e-06 0.0825149 0.0825105 0.0120424 7.61494e-06 0.00115403 0.103144 0.000656967 0.103796 0.862406 101.87 0.245648 0.721705 4.12981 0.0543522 0.0389605 0.96104 0.0198657 0.00424863 0.0191283 0.00408888 0.00513427 0.0058717 0.205371 0.234868 57.9749 -87.8947 126.122 15.9794 145.012 0.00014264 0.267094 192.917 0.310688 0.0673859 0.00409497 0.000561604 0.00138259 0.986991 0.991735 -2.97276e-06 -85.6679 0.0929843 31195.1 300.701 0.983521 0.319147 0.739945 0.73994 9.99958 2.98073e-06 1.19228e-05 0.130699 0.979677 0.930583 -0.0132933 4.89606e-06 0.501086 -1.8796e-20 6.92279e-24 -1.87891e-20 0.00139513 0.997818 8.59296e-05 0.152554 2.85172 0.00139513 0.997868 0.683602 0.00104608 0.00187967 0.000859296 0.455648 0.00187967 0.436176 0.000127799 1.02 0.887486 0.534735 0.285784 1.71633e-07 3.05758e-09 2390.41 3147.38 -0.0573152 0.482121 0.277609 0.255253 -0.593012 -0.169498 0.491381 -0.268261 -0.223128 1.48 1 0 295.752 0 2.05714 1.478 0.000299947 0.866861 0.64465 0.445668 0.404858 2.05739 129.643 83.5565 18.6998 60.6908 0.00404035 0 -40 10
0.579 1.67818e-08 2.53887e-06 0.0825998 0.0825954 0.0120423 7.6281e-06 0.00115403 0.10325 0.000656971 0.103902 0.862459 101.87 0.245642 0.721781 4.12993 0.0543583 0.0389616 0.961038 0.0198656 0.00424875 0.0191282 0.00408898 0.00513441 0.00587185 0.205377 0.234874 57.975 -87.8947 126.123 15.9794 145.012 0.000142632 0.267094 192.917 0.310687 0.0673859 0.00409497 0.000561604 0.00138259 0.986991 0.991735 -2.97277e-06 -85.6679 0.0929844 31195 300.704 0.983521 0.319147 0.739902 0.739898 9.99958 2.98073e-06 1.19228e-05 0.1307 0.979689 0.930589 -0.0132933 4.89609e-06 0.501091 -1.87968e-20 6.92313e-24 -1.87899e-20 0.00139513 0.997818 8.59296e-05 0.152554 2.85172 0.00139513 0.997867 0.683712 0.0010461 0.00187967 0.000859296 0.455648 0.00187967 0.436185 0.000127803 1.02 0.887487 0.534735 0.285785 1.71633e-07 3.0576e-09 2390.4 3147.2 -0.0573027 0.482121 0.277609 0.255242 -0.593014 -0.169499 0.491418 -0.268259 -0.223166 1.481 1 0 295.765 0 2.05732 1.479 0.000299946 0.866781 0.644707 0.445366 0.404888 2.05757 129.652 83.5586 18.6999 60.6918 0.00404026 0 -40 10
0.58 1.68108e-08 2.53887e-06 0.0826847 0.0826803 0.0120423 7.64126e-06 0.00115403 0.103356 0.000656976 0.104008 0.862511 101.87 0.245636 0.721857 4.13005 0.0543643 0.0389627 0.961037 0.0198654 0.00424887 0.019128 0.00408907 0.00513456 0.00587199 0.205382 0.234879 57.975 -87.8947 126.123 15.9793 145.012 0.000142624 0.267094 192.917 0.310687 0.0673858 0.00409498 0.000561605 0.00138259 0.986991 0.991735 -2.97278e-06 -85.6679 0.0929844 31195 300.707 0.983521 0.319147 0.73986 0.739856 9.99958 2.98074e-06 1.19228e-05 0.130701 0.979701 0.930594 -0.0132933 4.89612e-06 0.501095 -1.87976e-20 6.92346e-24 -1.87907e-20 0.00139513 0.997818 8.59297e-05 0.152554 2.85172 0.00139513 0.997867 0.683822 0.00104612 0.00187967 0.000859297 0.455648 0.00187967 0.436195 0.000127806 1.02 0.887488 0.534734 0.285786 1.71633e-07 3.05762e-09 2390.38 3147.02 -0.0572903 0.482121 0.277609 0.255231 -0.593016 -0.169499 0.491454 -0.268257 -0.223205 1.482 1 0 295.778 0 2.0575 1.48 0.000299946 0.866701 0.644763 0.445066 0.404919 2.05775 129.662 83.5607 18.7 60.6928 0.00404017 0 -40 10
0.581 1.68397e-08 2.53887e-06 0.0827695 0.0827651 0.0120423 7.65442e-06 0.00115403 0.103462 0.00065698 0.104114 0.862564 101.87 0.24563 0.721933 4.13016 0.0543704 0.0389638 0.961036 0.0198653 0.00424898 0.0191279 0.00408917 0.0051347 0.00587213 0.205388 0.234885 57.9751 -87.8947 126.124 15.9793 145.012 0.000142616 0.267095 192.917 0.310687 0.0673858 0.00409498 0.000561606 0.00138259 0.986991 0.991735 -2.9728e-06 -85.6679 0.0929845 31195 300.71 0.983521 0.319147 0.739818 0.739814 9.99958 2.98074e-06 1.19229e-05 0.130703 0.979713 0.9306 -0.0132933 4.89614e-06 0.5011 -1.87984e-20 6.92379e-24 -1.87915e-20 0.00139513 0.997818 8.59298e-05 0.152554 2.85173 0.00139513 0.997867 0.683932 0.00104614 0.00187967 0.000859298 0.455648 0.00187967 0.436204 0.00012781 1.02 0.887489 0.534734 0.285788 1.71633e-07 3.05764e-09 2390.36 3146.84 -0.057278 0.482121 0.277609 0.255219 -0.593018 -0.169499 0.49149 -0.268255 -0.223243 1.483 1 0 295.79 0 2.05768 1.481 0.000299946 0.866622 0.644819 0.444766 0.404949 2.05793 129.672 83.5627 18.7001 60.6938 0.00404009 0 -40 10
0.582 1.68687e-08 2.53887e-06 0.0828542 0.0828499 0.0120423 7.66758e-06 0.00115403 0.103568 0.000656984 0.10422 0.862616 101.87 0.245624 0.72201 4.13028 0.0543764 0.0389649 0.961035 0.0198652 0.0042491 0.0191277 0.00408927 0.00513484 0.00587227 0.205394 0.234891 57.9751 -87.8947 126.125 15.9793 145.012 0.000142607 0.267095 192.917 0.310686 0.0673857 0.00409498 0.000561606 0.00138259 0.986991 0.991735 -2.97281e-06 -85.6679 0.0929846 31195 300.713 0.983521 0.319147 0.739776 0.739772 9.99958 2.98075e-06 1.19229e-05 0.130704 0.979725 0.930605 -0.0132933 4.89617e-06 0.501105 -1.87992e-20 6.92413e-24 -1.87923e-20 0.00139514 0.997818 8.59299e-05 0.152555 2.85173 0.00139514 0.997866 0.684043 0.00104616 0.00187967 0.000859299 0.455647 0.00187967 0.436213 0.000127813 1.02 0.88749 0.534734 0.285789 1.71634e-07 3.05766e-09 2390.35 3146.66 -0.0572657 0.482121 0.277608 0.255208 -0.59302 -0.169499 0.491526 -0.268253 -0.223281 1.484 1 0 295.802 0 2.05786 1.482 0.000299946 0.866543 0.644876 0.444467 0.404979 2.05811 129.681 83.5648 18.7003 60.6948 0.00404 0 -40 10
0.583 1.68976e-08 2.53887e-06 0.0829389 0.0829346 0.0120423 7.68074e-06 0.00115403 0.103674 0.000656989 0.104326 0.862669 101.87 0.245617 0.722086 4.1304 0.0543825 0.0389661 0.961034 0.019865 0.00424922 0.0191276 0.00408936 0.00513499 0.00587241 0.2054 0.234897 57.9752 -87.8947 126.126 15.9792 145.012 0.000142599 0.267095 192.917 0.310686 0.0673857 0.00409498 0.000561607 0.0013826 0.986991 0.991735 -2.97282e-06 -85.6679 0.0929847 31195 300.716 0.983521 0.319147 0.739734 0.73973 9.99958 2.98075e-06 1.19229e-05 0.130705 0.979737 0.930611 -0.0132933 4.8962e-06 0.50111 -1.88e-20 6.92446e-24 -1.87931e-20 0.00139514 0.997818 8.59299e-05 0.152555 2.85173 0.00139514 0.997866 0.684153 0.00104618 0.00187967 0.000859299 0.455647 0.00187967 0.436222 0.000127817 1.02 0.887491 0.534734 0.28579 1.71634e-07 3.05768e-09 2390.33 3146.48 -0.0572535 0.482121 0.277608 0.255197 -0.593022 -0.169499 0.491562 -0.268251 -0.223318 1.485 1 0 295.815 0 2.05804 1.483 0.000299945 0.866464 0.644932 0.444168 0.40501 2.05829 129.691 83.5668 18.7004 60.6958 0.00403992 0 -40 10
0.584 1.69266e-08 2.53887e-06 0.0830235 0.0830192 0.0120423 7.69391e-06 0.00115403 0.103779 0.000656993 0.104432 0.862722 101.869 0.245611 0.722163 4.13052 0.0543886 0.0389672 0.961033 0.0198649 0.00424933 0.0191274 0.00408946 0.00513513 0.00587256 0.205405 0.234902 57.9753 -87.8947 126.127 15.9792 145.012 0.000142591 0.267095 192.916 0.310685 0.0673856 0.00409499 0.000561607 0.0013826 0.986991 0.991735 -2.97284e-06 -85.6678 0.0929847 31194.9 300.72 0.983521 0.319147 0.739693 0.739688 9.99958 2.98076e-06 1.19229e-05 0.130706 0.979749 0.930616 -0.0132933 4.89623e-06 0.501115 -1.88008e-20 6.9248e-24 -1.87939e-20 0.00139514 0.997818 8.593e-05 0.152555 2.85173 0.00139514 0.997866 0.684263 0.0010462 0.00187967 0.0008593 0.455647 0.00187967 0.436232 0.00012782 1.02 0.887492 0.534733 0.285792 1.71634e-07 3.0577e-09 2390.31 3146.3 -0.0572413 0.482121 0.277608 0.255186 -0.593024 -0.169499 0.491597 -0.268249 -0.223356 1.486 1 0 295.827 0 2.05822 1.484 0.000299945 0.866386 0.644988 0.443871 0.40504 2.05847 129.7 83.5689 18.7005 60.6968 0.00403983 0 -40 10
0.585 1.69556e-08 2.53887e-06 0.083108 0.0831037 0.0120423 7.70707e-06 0.00115403 0.103885 0.000656997 0.104537 0.862775 101.869 0.245605 0.722239 4.13064 0.0543947 0.0389683 0.961032 0.0198647 0.00424945 0.0191273 0.00408956 0.00513528 0.0058727 0.205411 0.234908 57.9753 -87.8948 126.127 15.9791 145.012 0.000142583 0.267095 192.916 0.310685 0.0673856 0.00409499 0.000561608 0.0013826 0.986991 0.991735 -2.97285e-06 -85.6678 0.0929848 31194.9 300.723 0.983521 0.319147 0.739651 0.739647 9.99958 2.98076e-06 1.19229e-05 0.130707 0.979761 0.930621 -0.0132933 4.89625e-06 0.50112 -1.88016e-20 6.92513e-24 -1.87947e-20 0.00139514 0.997818 8.59301e-05 0.152555 2.85173 0.00139514 0.997866 0.684372 0.00104622 0.00187968 0.000859301 0.455647 0.00187967 0.436241 0.000127823 1.02 0.887493 0.534733 0.285793 1.71634e-07 3.05772e-09 2390.3 3146.13 -0.0572292 0.482121 0.277607 0.255175 -0.593026 -0.169499 0.491633 -0.268247 -0.223393 1.487 1 0 295.839 0 2.0584 1.485 0.000299945 0.866308 0.645045 0.443574 0.40507 2.05865 129.71 83.5709 18.7006 60.6978 0.00403975 0 -40 10
0.586 1.69845e-08 2.53887e-06 0.0831925 0.0831882 0.0120422 7.72023e-06 0.00115403 0.103991 0.000657001 0.104643 0.862827 101.869 0.245599 0.722316 4.13076 0.0544008 0.0389695 0.961031 0.0198646 0.00424957 0.0191272 0.00408966 0.00513542 0.00587284 0.205417 0.234914 57.9754 -87.8948 126.128 15.9791 145.012 0.000142575 0.267095 192.916 0.310685 0.0673855 0.00409499 0.000561608 0.0013826 0.986991 0.991735 -2.97286e-06 -85.6678 0.0929849 31194.9 300.726 0.983521 0.319147 0.73961 0.739606 9.99958 2.98076e-06 1.19229e-05 0.130709 0.979772 0.930627 -0.0132933 4.89628e-06 0.501125 -1.88024e-20 6.92546e-24 -1.87955e-20 0.00139514 0.997818 8.59301e-05 0.152555 2.85173 0.00139514 0.997865 0.684482 0.00104624 0.00187968 0.000859301 0.455647 0.00187968 0.43625 0.000127827 1.02 0.887494 0.534733 0.285795 1.71635e-07 3.05774e-09 2390.28 3145.95 -0.0572171 0.482121 0.277607 0.255163 -0.593028 -0.169499 0.491668 -0.268246 -0.223431 1.488 1 0 295.851 0 2.05858 1.486 0.000299945 0.86623 0.645101 0.443278 0.405101 2.05883 129.72 83.5729 18.7007 60.6988 0.00403966 0 -40 10
0.587 1.70135e-08 2.53887e-06 0.0832769 0.0832726 0.0120422 7.73339e-06 0.00115403 0.104096 0.000657006 0.104748 0.86288 101.869 0.245593 0.722393 4.13088 0.0544069 0.0389706 0.961029 0.0198644 0.00424969 0.019127 0.00408976 0.00513557 0.00587299 0.205423 0.234919 57.9755 -87.8948 126.129 15.9791 145.012 0.000142568 0.267096 192.916 0.310684 0.0673855 0.00409499 0.000561609 0.0013826 0.986991 0.991735 -2.97288e-06 -85.6678 0.092985 31194.9 300.729 0.983521 0.319147 0.739569 0.739565 9.99958 2.98077e-06 1.1923e-05 0.13071 0.979784 0.930632 -0.0132933 4.89631e-06 0.50113 -1.88032e-20 6.9258e-24 -1.87963e-20 0.00139514 0.997818 8.59302e-05 0.152555 2.85173 0.00139514 0.997865 0.684592 0.00104626 0.00187968 0.000859302 0.455646 0.00187968 0.436259 0.00012783 1.02 0.887495 0.534732 0.285796 1.71635e-07 3.05776e-09 2390.26 3145.77 -0.0572051 0.482121 0.277607 0.255152 -0.59303 -0.169499 0.491703 -0.268244 -0.223468 1.489 1 0 295.864 0 2.05876 1.487 0.000299944 0.866153 0.645157 0.442983 0.405131 2.05901 129.729 83.575 18.7009 60.6997 0.00403958 0 -40 10
0.588 1.70424e-08 2.53887e-06 0.0833612 0.0833569 0.0120422 7.74655e-06 0.00115403 0.104201 0.00065701 0.104854 0.862933 101.869 0.245587 0.72247 4.131 0.054413 0.0389717 0.961028 0.0198643 0.00424981 0.0191269 0.00408985 0.00513572 0.00587313 0.205429 0.234925 57.9755 -87.8948 126.129 15.979 145.012 0.00014256 0.267096 192.916 0.310684 0.0673855 0.004095 0.00056161 0.00138261 0.986991 0.991735 -2.97289e-06 -85.6678 0.0929851 31194.9 300.732 0.983521 0.319147 0.739528 0.739524 9.99958 2.98077e-06 1.1923e-05 0.130711 0.979796 0.930638 -0.0132933 4.89633e-06 0.501135 -1.8804e-20 6.92613e-24 -1.87971e-20 0.00139514 0.997818 8.59303e-05 0.152555 2.85173 0.00139514 0.997865 0.684702 0.00104628 0.00187968 0.000859303 0.455646 0.00187968 0.436269 0.000127834 1.02 0.887496 0.534732 0.285797 1.71635e-07 3.05778e-09 2390.25 3145.6 -0.0571931 0.482121 0.277607 0.255141 -0.593032 -0.169499 0.491738 -0.268242 -0.223505 1.49 1 0 295.876 0 2.05894 1.488 0.000299944 0.866076 0.645213 0.442688 0.405161 2.05919 129.739 83.577 18.701 60.7007 0.0040395 0 -40 10
0.589 1.70714e-08 2.53887e-06 0.0834454 0.0834412 0.0120422 7.75972e-06 0.00115403 0.104307 0.000657014 0.104959 0.862986 101.869 0.245581 0.722547 4.13113 0.0544191 0.0389729 0.961027 0.0198641 0.00424993 0.0191267 0.00408995 0.00513586 0.00587327 0.205434 0.234931 57.9756 -87.8948 126.13 15.979 145.012 0.000142552 0.267096 192.916 0.310684 0.0673854 0.004095 0.00056161 0.00138261 0.986991 0.991735 -2.9729e-06 -85.6678 0.0929851 31194.8 300.736 0.983521 0.319147 0.739487 0.739483 9.99958 2.98078e-06 1.1923e-05 0.130712 0.979808 0.930643 -0.0132933 4.89636e-06 0.50114 -1.88048e-20 6.92646e-24 -1.87979e-20 0.00139514 0.997818 8.59303e-05 0.152556 2.85173 0.00139514 0.997864 0.684812 0.0010463 0.00187968 0.000859303 0.455646 0.00187968 0.436278 0.000127837 1.02 0.887497 0.534732 0.285799 1.71635e-07 3.05781e-09 2390.23 3145.43 -0.0571812 0.482121 0.277606 0.25513 -0.593034 -0.169499 0.491773 -0.26824 -0.223541 1.491 1 0 295.888 0 2.05912 1.489 0.000299944 0.865999 0.645269 0.442394 0.405191 2.05937 129.748 83.579 18.7011 60.7017 0.00403941 0 -40 10
0.59 1.71003e-08 2.53887e-06 0.0835296 0.0835254 0.0120422 7.77288e-06 0.00115403 0.104412 0.000657018 0.105064 0.863039 101.869 0.245575 0.722624 4.13125 0.0544252 0.038974 0.961026 0.019864 0.00425005 0.0191266 0.00409005 0.00513601 0.00587342 0.20544 0.234937 57.9756 -87.8948 126.131 15.979 145.012 0.000142544 0.267096 192.916 0.310683 0.0673854 0.004095 0.000561611 0.00138261 0.986991 0.991735 -2.97292e-06 -85.6678 0.0929852 31194.8 300.739 0.983521 0.319147 0.739447 0.739442 9.99958 2.98078e-06 1.1923e-05 0.130713 0.979819 0.930648 -0.0132933 4.89639e-06 0.501145 -1.88056e-20 6.9268e-24 -1.87987e-20 0.00139514 0.997818 8.59304e-05 0.152556 2.85173 0.00139514 0.997864 0.684922 0.00104631 0.00187968 0.000859304 0.455646 0.00187968 0.436287 0.000127841 1.02 0.887498 0.534732 0.2858 1.71636e-07 3.05783e-09 2390.21 3145.25 -0.0571694 0.482121 0.277606 0.25512 -0.593036 -0.169499 0.491807 -0.268238 -0.223578 1.492 1 0 295.9 0 2.0593 1.49 0.000299944 0.865922 0.645325 0.442101 0.405222 2.05955 129.758 83.581 18.7012 60.7026 0.00403933 0 -40 10
0.591 1.71293e-08 2.53887e-06 0.0836138 0.0836096 0.0120422 7.78604e-06 0.00115403 0.104517 0.000657023 0.10517 0.863092 101.869 0.245569 0.722702 4.13137 0.0544314 0.0389752 0.961025 0.0198638 0.00425017 0.0191264 0.00409015 0.00513616 0.00587357 0.205446 0.234943 57.9757 -87.8948 126.132 15.9789 145.012 0.000142536 0.267096 192.915 0.310683 0.0673853 0.00409501 0.000561611 0.00138261 0.986991 0.991735 -2.97293e-06 -85.6678 0.0929853 31194.8 300.742 0.983521 0.319147 0.739406 0.739402 9.99958 2.98079e-06 1.1923e-05 0.130715 0.979831 0.930654 -0.0132933 4.89642e-06 0.501149 -1.88064e-20 6.92713e-24 -1.87995e-20 0.00139514 0.997818 8.59305e-05 0.152556 2.85173 0.00139514 0.997864 0.685031 0.00104633 0.00187968 0.000859305 0.455646 0.00187968 0.436296 0.000127844 1.02 0.887499 0.534731 0.285802 1.71636e-07 3.05785e-09 2390.2 3145.08 -0.0571576 0.482121 0.277606 0.255109 -0.593038 -0.169499 0.491842 -0.268236 -0.223615 1.493 1 0 295.912 0 2.05948 1.491 0.000299944 0.865846 0.645382 0.441809 0.405252 2.05973 129.768 83.583 18.7013 60.7036 0.00403925 0 -40 10
0.592 1.71582e-08 2.53887e-06 0.0836978 0.0836936 0.0120422 7.7992e-06 0.00115403 0.104622 0.000657027 0.105275 0.863146 101.869 0.245562 0.722779 4.13149 0.0544375 0.0389763 0.961024 0.0198637 0.00425029 0.0191263 0.00409025 0.0051363 0.00587371 0.205452 0.234948 57.9758 -87.8948 126.132 15.9789 145.012 0.000142528 0.267096 192.915 0.310682 0.0673853 0.00409501 0.000561612 0.00138261 0.986991 0.991735 -2.97294e-06 -85.6678 0.0929854 31194.8 300.745 0.983521 0.319147 0.739366 0.739362 9.99958 2.98079e-06 1.19231e-05 0.130716 0.979842 0.930659 -0.0132933 4.89644e-06 0.501154 -1.88072e-20 6.92747e-24 -1.88003e-20 0.00139515 0.997818 8.59306e-05 0.152556 2.85173 0.00139515 0.997863 0.685141 0.00104635 0.00187968 0.000859306 0.455645 0.00187968 0.436305 0.000127848 1.02 0.8875 0.534731 0.285803 1.71636e-07 3.05787e-09 2390.18 3144.91 -0.0571458 0.482122 0.277605 0.255098 -0.593041 -0.169499 0.491876 -0.268234 -0.223651 1.494 1 0 295.924 0 2.05966 1.492 0.000299943 0.86577 0.645438 0.441517 0.405282 2.05991 129.777 83.5849 18.7014 60.7046 0.00403917 0 -40 10
0.593 1.71872e-08 2.53887e-06 0.0837818 0.0837776 0.0120422 7.81236e-06 0.00115403 0.104727 0.000657031 0.10538 0.863199 101.868 0.245556 0.722857 4.13162 0.0544437 0.0389775 0.961022 0.0198635 0.00425041 0.0191261 0.00409035 0.00513645 0.00587386 0.205458 0.234954 57.9758 -87.8948 126.133 15.9788 145.012 0.000142521 0.267097 192.915 0.310682 0.0673852 0.00409501 0.000561613 0.00138261 0.986991 0.991735 -2.97295e-06 -85.6678 0.0929854 31194.8 300.749 0.983521 0.319147 0.739326 0.739322 9.99958 2.98079e-06 1.19231e-05 0.130717 0.979854 0.930664 -0.0132933 4.89647e-06 0.501159 -1.8808e-20 6.9278e-24 -1.88011e-20 0.00139515 0.997818 8.59306e-05 0.152556 2.85173 0.00139515 0.997863 0.685251 0.00104637 0.00187969 0.000859306 0.455645 0.00187969 0.436315 0.000127851 1.02 0.887501 0.534731 0.285804 1.71636e-07 3.05789e-09 2390.16 3144.74 -0.0571341 0.482122 0.277605 0.255087 -0.593043 -0.169499 0.491911 -0.268232 -0.223687 1.495 1 0 295.935 0 2.05983 1.493 0.000299943 0.865695 0.645494 0.441226 0.405312 2.06009 129.787 83.5869 18.7015 60.7055 0.00403908 0 -40 10
0.594 1.72161e-08 2.53887e-06 0.0838657 0.0838616 0.0120421 7.82552e-06 0.00115403 0.104832 0.000657035 0.105485 0.863252 101.868 0.24555 0.722934 4.13174 0.0544498 0.0389787 0.961021 0.0198634 0.00425053 0.019126 0.00409045 0.0051366 0.005874 0.205464 0.23496 57.9759 -87.8948 126.134 15.9788 145.012 0.000142513 0.267097 192.915 0.310682 0.0673852 0.00409501 0.000561613 0.00138262 0.986991 0.991735 -2.97297e-06 -85.6678 0.0929855 31194.7 300.752 0.983521 0.319147 0.739286 0.739282 9.99958 2.9808e-06 1.19231e-05 0.130718 0.979865 0.93067 -0.0132932 4.8965e-06 0.501165 -1.88088e-20 6.92813e-24 -1.88019e-20 0.00139515 0.997818 8.59307e-05 0.152556 2.85174 0.00139515 0.997863 0.68536 0.00104639 0.00187969 0.000859307 0.455645 0.00187969 0.436324 0.000127855 1.02 0.887502 0.53473 0.285806 1.71637e-07 3.05791e-09 2390.15 3144.57 -0.0571224 0.482122 0.277605 0.255076 -0.593045 -0.1695 0.491945 -0.26823 -0.223723 1.496 1 0 295.947 0 2.06001 1.494 0.000299943 0.86562 0.64555 0.440936 0.405342 2.06026 129.796 83.5889 18.7017 60.7065 0.004039 0 -40 10
0.595 1.72451e-08 2.53887e-06 0.0839496 0.0839454 0.0120421 7.83868e-06 0.00115403 0.104937 0.000657039 0.105589 0.863306 101.868 0.245544 0.723012 4.13186 0.054456 0.0389798 0.96102 0.0198633 0.00425065 0.0191258 0.00409055 0.00513675 0.00587415 0.20547 0.234966 57.976 -87.8948 126.135 15.9788 145.012 0.000142505 0.267097 192.915 0.310681 0.0673851 0.00409502 0.000561614 0.00138262 0.986991 0.991735 -2.97298e-06 -85.6678 0.0929856 31194.7 300.755 0.983521 0.319147 0.739246 0.739242 9.99958 2.9808e-06 1.19231e-05 0.13072 0.979877 0.930675 -0.0132932 4.89652e-06 0.50117 -1.88096e-20 6.92847e-24 -1.88027e-20 0.00139515 0.997818 8.59308e-05 0.152556 2.85174 0.00139515 0.997863 0.68547 0.00104641 0.00187969 0.000859308 0.455645 0.00187969 0.436333 0.000127858 1.02 0.887503 0.53473 0.285807 1.71637e-07 3.05793e-09 2390.13 3144.4 -0.0571108 0.482122 0.277605 0.255066 -0.593047 -0.1695 0.491978 -0.268228 -0.223759 1.497 1 0 295.959 0 2.06019 1.495 0.000299943 0.865545 0.645605 0.440647 0.405372 2.06044 129.806 83.5908 18.7018 60.7074 0.00403892 0 -40 10
0.596 1.72741e-08 2.53887e-06 0.0840334 0.0840292 0.0120421 7.85185e-06 0.00115403 0.105042 0.000657043 0.105694 0.863359 101.868 0.245538 0.72309 4.13199 0.0544622 0.038981 0.961019 0.0198631 0.00425077 0.0191257 0.00409065 0.0051369 0.0058743 0.205476 0.234972 57.976 -87.8948 126.135 15.9787 145.012 0.000142498 0.267097 192.915 0.310681 0.0673851 0.00409502 0.000561614 0.00138262 0.986991 0.991735 -2.97299e-06 -85.6677 0.0929857 31194.7 300.758 0.983521 0.319147 0.739207 0.739202 9.99958 2.98081e-06 1.19231e-05 0.130721 0.979888 0.93068 -0.0132932 4.89655e-06 0.501175 -1.88104e-20 6.9288e-24 -1.88035e-20 0.00139515 0.997818 8.59308e-05 0.152556 2.85174 0.00139515 0.997862 0.685579 0.00104643 0.00187969 0.000859308 0.455645 0.00187969 0.436342 0.000127862 1.02 0.887504 0.53473 0.285809 1.71637e-07 3.05795e-09 2390.11 3144.23 -0.0570993 0.482122 0.277604 0.255055 -0.593048 -0.1695 0.492012 -0.268226 -0.223795 1.498 1 0 295.971 0 2.06037 1.496 0.000299942 0.86547 0.645661 0.440358 0.405402 2.06062 129.815 83.5928 18.7019 60.7083 0.00403884 0 -40 10
0.597 1.7303e-08 2.53887e-06 0.0841171 0.084113 0.0120421 7.86501e-06 0.00115403 0.105146 0.000657047 0.105799 0.863412 101.868 0.245532 0.723168 4.13211 0.0544684 0.0389822 0.961018 0.019863 0.00425089 0.0191256 0.00409075 0.00513705 0.00587445 0.205482 0.234978 57.9761 -87.8948 126.136 15.9787 145.012 0.00014249 0.267097 192.915 0.310681 0.067385 0.00409502 0.000561615 0.00138262 0.986991 0.991735 -2.97301e-06 -85.6677 0.0929857 31194.7 300.762 0.983521 0.319147 0.739167 0.739163 9.99958 2.98081e-06 1.19231e-05 0.130722 0.979899 0.930685 -0.0132932 4.89658e-06 0.50118 -1.88112e-20 6.92914e-24 -1.88043e-20 0.00139515 0.997818 8.59309e-05 0.152557 2.85174 0.00139515 0.997862 0.685689 0.00104645 0.00187969 0.000859309 0.455644 0.00187969 0.436351 0.000127865 1.02 0.887505 0.53473 0.28581 1.71637e-07 3.05797e-09 2390.1 3144.06 -0.0570878 0.482122 0.277604 0.255045 -0.59305 -0.1695 0.492046 -0.268224 -0.22383 1.499 1 0 295.982 0 2.06055 1.497 0.000299942 0.865396 0.645717 0.44007 0.405433 2.0608 129.825 83.5947 18.702 60.7093 0.00403876 0 -40 10
0.598 1.7332e-08 2.53887e-06 0.0842008 0.0841966 0.0120421 7.87817e-06 0.00115403 0.105251 0.000657052 0.105903 0.863466 101.868 0.245525 0.723246 4.13223 0.0544746 0.0389833 0.961017 0.0198628 0.00425101 0.0191254 0.00409085 0.0051372 0.00587459 0.205488 0.234984 57.9761 -87.8948 126.137 15.9787 145.012 0.000142482 0.267097 192.914 0.31068 0.067385 0.00409502 0.000561616 0.00138262 0.986991 0.991735 -2.97302e-06 -85.6677 0.0929858 31194.7 300.765 0.983521 0.319147 0.739128 0.739123 9.99958 2.98082e-06 1.19232e-05 0.130723 0.979911 0.93069 -0.0132932 4.89661e-06 0.501185 -1.8812e-20 6.92947e-24 -1.88051e-20 0.00139515 0.997818 8.5931e-05 0.152557 2.85174 0.00139515 0.997862 0.685798 0.00104647 0.00187969 0.00085931 0.455644 0.00187969 0.436361 0.000127869 1.02 0.887506 0.534729 0.285811 1.71638e-07 3.05799e-09 2390.08 3143.89 -0.0570764 0.482122 0.277604 0.255034 -0.593052 -0.1695 0.492079 -0.268222 -0.223866 1.5 1 0 295.994 0 2.06073 1.498 0.000299942 0.865322 0.645773 0.439783 0.405463 2.06098 129.835 83.5967 18.7021 60.7102 0.00403868 0 -40 10
0.599 1.73609e-08 2.53887e-06 0.0842843 0.0842802 0.0120421 7.89133e-06 0.00115403 0.105355 0.000657056 0.106008 0.86352 101.868 0.245519 0.723324 4.13236 0.0544808 0.0389845 0.961015 0.0198627 0.00425113 0.0191253 0.00409096 0.00513735 0.00587474 0.205494 0.23499 57.9762 -87.8948 126.137 15.9786 145.012 0.000142475 0.267098 192.914 0.31068 0.0673849 0.00409503 0.000561616 0.00138263 0.986991 0.991735 -2.97303e-06 -85.6677 0.0929859 31194.6 300.768 0.983521 0.319147 0.739089 0.739084 9.99958 2.98082e-06 1.19232e-05 0.130725 0.979922 0.930696 -0.0132932 4.89663e-06 0.50119 -1.88128e-20 6.9298e-24 -1.88059e-20 0.00139515 0.997818 8.59311e-05 0.152557 2.85174 0.00139515 0.997861 0.685907 0.00104649 0.00187969 0.000859311 0.455644 0.00187969 0.43637 0.000127872 1.02 0.887507 0.534729 0.285813 1.71638e-07 3.05801e-09 2390.06 3143.72 -0.057065 0.482122 0.277603 0.255023 -0.593054 -0.1695 0.492112 -0.26822 -0.223901 1.501 1 0 296.005 0 2.06091 1.499 0.000299942 0.865248 0.645829 0.439497 0.405493 2.06116 129.844 83.5986 18.7022 60.7111 0.0040386 0 -40 10
0.6 1.73899e-08 2.53887e-06 0.0843679 0.0843638 0.0120421 7.90449e-06 0.00115403 0.10546 0.00065706 0.106112 0.863573 101.868 0.245513 0.723402 4.13248 0.054487 0.0389857 0.961014 0.0198625 0.00425126 0.0191251 0.00409106 0.0051375 0.00587489 0.2055 0.234996 57.9763 -87.8948 126.138 15.9786 145.012 0.000142467 0.267098 192.914 0.310679 0.0673849 0.00409503 0.000561617 0.00138263 0.986991 0.991735 -2.97305e-06 -85.6677 0.092986 31194.6 300.772 0.983521 0.319147 0.73905 0.739045 9.99958 2.98083e-06 1.19232e-05 0.130726 0.979933 0.930701 -0.0132932 4.89666e-06 0.501195 -1.88136e-20 6.93014e-24 -1.88067e-20 0.00139515 0.997818 8.59311e-05 0.152557 2.85174 0.00139515 0.997861 0.686017 0.00104651 0.0018797 0.000859311 0.455644 0.00187969 0.436379 0.000127876 1.02 0.887508 0.534729 0.285814 1.71638e-07 3.05803e-09 2390.05 3143.56 -0.0570536 0.482122 0.277603 0.255013 -0.593056 -0.1695 0.492145 -0.268218 -0.223936 1.502 1 0 296.017 0 2.06108 1.5 0.000299941 0.865175 0.645885 0.439211 0.405523 2.06133 129.854 83.6005 18.7023 60.7121 0.00403852 0 -40 10
0.601 1.74188e-08 2.53887e-06 0.0844513 0.0844472 0.012042 7.91765e-06 0.00115403 0.105564 0.000657064 0.106217 0.863627 101.867 0.245507 0.72348 4.13261 0.0544932 0.0389869 0.961013 0.0198624 0.00425138 0.019125 0.00409116 0.00513765 0.00587504 0.205506 0.235002 57.9763 -87.8948 126.139 15.9785 145.012 0.00014246 0.267098 192.914 0.310679 0.0673848 0.00409503 0.000561617 0.00138263 0.986991 0.991735 -2.97306e-06 -85.6677 0.0929861 31194.6 300.775 0.983521 0.319147 0.739011 0.739006 9.99958 2.98083e-06 1.19232e-05 0.130727 0.979945 0.930706 -0.0132932 4.89669e-06 0.5012 -1.88144e-20 6.93047e-24 -1.88075e-20 0.00139515 0.997818 8.59312e-05 0.152557 2.85174 0.00139515 0.997861 0.686126 0.00104653 0.0018797 0.000859312 0.455644 0.0018797 0.436388 0.000127879 1.02 0.887509 0.534729 0.285815 1.71638e-07 3.05805e-09 2390.03 3143.39 -0.0570423 0.482122 0.277603 0.255003 -0.593058 -0.1695 0.492178 -0.268216 -0.223971 1.503 1 0 296.028 0 2.06126 1.501 0.000299941 0.865102 0.64594 0.438926 0.405553 2.06151 129.863 83.6024 18.7024 60.713 0.00403844 0 -40 10
0.602 1.74478e-08 2.53887e-06 0.0845347 0.0845306 0.012042 7.93081e-06 0.00115403 0.105668 0.000657068 0.106321 0.863681 101.867 0.245501 0.723559 4.13274 0.0544994 0.0389881 0.961012 0.0198622 0.0042515 0.0191248 0.00409126 0.0051378 0.00587519 0.205512 0.235008 57.9764 -87.8948 126.14 15.9785 145.012 0.000142452 0.267098 192.914 0.310679 0.0673848 0.00409503 0.000561618 0.00138263 0.986991 0.991735 -2.97307e-06 -85.6677 0.0929861 31194.6 300.778 0.983521 0.319147 0.738972 0.738968 9.99958 2.98083e-06 1.19232e-05 0.130728 0.979956 0.930711 -0.0132932 4.89671e-06 0.501205 -1.88152e-20 6.93081e-24 -1.88083e-20 0.00139516 0.997818 8.59313e-05 0.152557 2.85174 0.00139516 0.997861 0.686235 0.00104655 0.0018797 0.000859313 0.455643 0.0018797 0.436397 0.000127883 1.02 0.88751 0.534728 0.285817 1.71638e-07 3.05807e-09 2390.01 3143.23 -0.0570311 0.482122 0.277602 0.254992 -0.59306 -0.1695 0.492211 -0.268214 -0.224006 1.504 1 0 296.04 0 2.06144 1.502 0.000299941 0.865029 0.645996 0.438642 0.405583 2.06169 129.873 83.6043 18.7026 60.7139 0.00403836 0 -40 10
0.603 1.74767e-08 2.53887e-06 0.084618 0.084614 0.012042 7.94397e-06 0.00115403 0.105773 0.000657072 0.106425 0.863735 101.867 0.245494 0.723637 4.13286 0.0545057 0.0389893 0.961011 0.019862 0.00425163 0.0191247 0.00409136 0.00513795 0.00587534 0.205518 0.235014 57.9765 -87.8948 126.14 15.9785 145.012 0.000142445 0.267098 192.914 0.310678 0.0673848 0.00409504 0.000561618 0.00138263 0.986991 0.991735 -2.97309e-06 -85.6677 0.0929862 31194.6 300.782 0.983521 0.319147 0.738934 0.738929 9.99958 2.98084e-06 1.19232e-05 0.13073 0.979967 0.930716 -0.0132932 4.89674e-06 0.50121 -1.8816e-20 6.93114e-24 -1.88091e-20 0.00139516 0.997818 8.59313e-05 0.152557 2.85174 0.00139516 0.99786 0.686345 0.00104657 0.0018797 0.000859313 0.455643 0.0018797 0.436406 0.000127886 1.02 0.887511 0.534728 0.285818 1.71639e-07 3.0581e-09 2390 3143.06 -0.0570199 0.482122 0.277602 0.254982 -0.593062 -0.1695 0.492244 -0.268212 -0.224041 1.505 1 0 296.051 0 2.06162 1.503 0.000299941 0.864957 0.646052 0.438359 0.405613 2.06187 129.882 83.6062 18.7027 60.7148 0.00403828 0 -40 10
0.604 1.75057e-08 2.53887e-06 0.0847013 0.0846972 0.012042 7.95713e-06 0.00115403 0.105877 0.000657076 0.106529 0.863788 101.867 0.245488 0.723716 4.13299 0.0545119 0.0389905 0.96101 0.0198619 0.00425175 0.0191245 0.00409147 0.0051381 0.00587549 0.205524 0.23502 57.9765 -87.8948 126.141 15.9784 145.012 0.000142438 0.267098 192.914 0.310678 0.0673847 0.00409504 0.000561619 0.00138264 0.986991 0.991735 -2.9731e-06 -85.6677 0.0929863 31194.5 300.785 0.983521 0.319147 0.738895 0.738891 9.99958 2.98084e-06 1.19233e-05 0.130731 0.979978 0.930721 -0.0132932 4.89677e-06 0.501215 -1.88168e-20 6.93147e-24 -1.88099e-20 0.00139516 0.997818 8.59314e-05 0.152558 2.85174 0.00139516 0.99786 0.686454 0.00104659 0.0018797 0.000859314 0.455643 0.0018797 0.436416 0.00012789 1.02 0.887512 0.534728 0.28582 1.71639e-07 3.05812e-09 2389.98 3142.9 -0.0570087 0.482122 0.277602 0.254971 -0.593064 -0.1695 0.492276 -0.26821 -0.224075 1.506 1 0 296.062 0 2.0618 1.504 0.00029994 0.864884 0.646107 0.438076 0.405643 2.06205 129.892 83.6081 18.7028 60.7157 0.00403821 0 -40 10
0.605 1.75346e-08 2.53887e-06 0.0847845 0.0847804 0.012042 7.9703e-06 0.00115403 0.105981 0.00065708 0.106633 0.863842 101.867 0.245482 0.723794 4.13312 0.0545182 0.0389917 0.961008 0.0198617 0.00425187 0.0191244 0.00409157 0.00513826 0.00587564 0.20553 0.235026 57.9766 -87.8948 126.142 15.9784 145.012 0.00014243 0.267099 192.913 0.310678 0.0673847 0.00409504 0.00056162 0.00138264 0.986991 0.991735 -2.97312e-06 -85.6677 0.0929864 31194.5 300.788 0.983521 0.319147 0.738857 0.738853 9.99958 2.98085e-06 1.19233e-05 0.130732 0.979989 0.930726 -0.0132932 4.8968e-06 0.501221 -1.88176e-20 6.93181e-24 -1.88107e-20 0.00139516 0.997818 8.59315e-05 0.152558 2.85174 0.00139516 0.99786 0.686563 0.00104661 0.0018797 0.000859315 0.455643 0.0018797 0.436425 0.000127893 1.02 0.887513 0.534727 0.285821 1.71639e-07 3.05814e-09 2389.96 3142.73 -0.0569976 0.482122 0.277602 0.254961 -0.593066 -0.1695 0.492309 -0.268208 -0.224109 1.507 1 0 296.074 0 2.06197 1.505 0.00029994 0.864813 0.646163 0.437794 0.405673 2.06222 129.901 83.61 18.7029 60.7166 0.00403813 0 -40 10
0.606 1.75636e-08 2.53887e-06 0.0848676 0.0848636 0.012042 7.98346e-06 0.00115403 0.106084 0.000657084 0.106737 0.863896 101.867 0.245476 0.723873 4.13324 0.0545244 0.0389929 0.961007 0.0198616 0.004252 0.0191242 0.00409167 0.00513841 0.00587579 0.205536 0.235032 57.9767 -87.8948 126.142 15.9784 145.012 0.000142423 0.267099 192.913 0.310677 0.0673846 0.00409505 0.00056162 0.00138264 0.986991 0.991735 -2.97313e-06 -85.6677 0.0929864 31194.5 300.792 0.983521 0.319147 0.738819 0.738815 9.99958 2.98085e-06 1.19233e-05 0.130733 0.98 0.930731 -0.0132932 4.89682e-06 0.501226 -1.88184e-20 6.93214e-24 -1.88115e-20 0.00139516 0.997818 8.59316e-05 0.152558 2.85175 0.00139516 0.997859 0.686672 0.00104663 0.0018797 0.000859316 0.455643 0.0018797 0.436434 0.000127896 1.02 0.887514 0.534727 0.285823 1.71639e-07 3.05816e-09 2389.95 3142.57 -0.0569866 0.482122 0.277601 0.254951 -0.593068 -0.1695 0.492341 -0.268206 -0.224144 1.508 1 0 296.085 0 2.06215 1.506 0.00029994 0.864741 0.646219 0.437512 0.405702 2.0624 129.911 83.6119 18.703 60.7175 0.00403805 0 -40 10
0.607 1.75926e-08 2.53888e-06 0.0849506 0.0849466 0.012042 7.99662e-06 0.00115403 0.106188 0.000657088 0.106841 0.86395 101.867 0.245469 0.723952 4.13337 0.0545307 0.0389941 0.961006 0.0198614 0.00425212 0.0191241 0.00409178 0.00513856 0.00587594 0.205542 0.235038 57.9767 -87.8948 126.143 15.9783 145.012 0.000142416 0.267099 192.913 0.310677 0.0673846 0.00409505 0.000561621 0.00138264 0.986991 0.991735 -2.97314e-06 -85.6677 0.0929865 31194.5 300.795 0.98352 0.319147 0.738781 0.738777 9.99958 2.98086e-06 1.19233e-05 0.130735 0.980011 0.930736 -0.0132932 4.89685e-06 0.501231 -1.88192e-20 6.93248e-24 -1.88123e-20 0.00139516 0.997818 8.59316e-05 0.152558 2.85175 0.00139516 0.997859 0.686781 0.00104665 0.0018797 0.000859316 0.455642 0.0018797 0.436443 0.0001279 1.02 0.887515 0.534727 0.285824 1.7164e-07 3.05818e-09 2389.93 3142.41 -0.0569756 0.482123 0.277601 0.254941 -0.59307 -0.1695 0.492373 -0.268204 -0.224178 1.509 1 0 296.096 0 2.06233 1.507 0.00029994 0.86467 0.646274 0.437232 0.405732 2.06258 129.92 83.6137 18.7031 60.7184 0.00403797 0 -40 10
0.608 1.76215e-08 2.53888e-06 0.0850336 0.0850296 0.012042 8.00978e-06 0.00115403 0.106292 0.000657092 0.106945 0.864005 101.867 0.245463 0.724031 4.1335 0.054537 0.0389953 0.961005 0.0198613 0.00425225 0.0191239 0.00409188 0.00513872 0.0058761 0.205549 0.235044 57.9768 -87.8948 126.144 15.9783 145.012 0.000142408 0.267099 192.913 0.310676 0.0673845 0.00409505 0.000561621 0.00138264 0.98699 0.991735 -2.97316e-06 -85.6676 0.0929866 31194.5 300.798 0.98352 0.319147 0.738743 0.738739 9.99958 2.98086e-06 1.19233e-05 0.130736 0.980022 0.930741 -0.0132932 4.89688e-06 0.501236 -1.882e-20 6.93281e-24 -1.88131e-20 0.00139516 0.997818 8.59317e-05 0.152558 2.85175 0.00139516 0.997859 0.68689 0.00104667 0.00187971 0.000859317 0.455642 0.0018797 0.436452 0.000127903 1.02 0.887516 0.534727 0.285825 1.7164e-07 3.0582e-09 2389.91 3142.25 -0.0569647 0.482123 0.277601 0.254931 -0.593072 -0.1695 0.492405 -0.268202 -0.224212 1.51 1 0 296.107 0 2.06251 1.508 0.000299939 0.864599 0.64633 0.436952 0.405762 2.06275 129.93 83.6156 18.7032 60.7193 0.0040379 0 -40 10
0.609 1.76505e-08 2.53888e-06 0.0851165 0.0851125 0.0120419 8.02294e-06 0.00115403 0.106396 0.000657096 0.107048 0.864059 101.866 0.245457 0.72411 4.13363 0.0545432 0.0389965 0.961004 0.0198611 0.00425237 0.0191238 0.00409198 0.00513887 0.00587625 0.205555 0.23505 57.9768 -87.8948 126.144 15.9782 145.013 0.000142401 0.267099 192.913 0.310676 0.0673845 0.00409505 0.000561622 0.00138265 0.98699 0.991735 -2.97317e-06 -85.6676 0.0929867 31194.4 300.802 0.98352 0.319147 0.738706 0.738701 9.99958 2.98086e-06 1.19234e-05 0.130737 0.980033 0.930746 -0.0132932 4.89691e-06 0.501241 -1.88208e-20 6.93315e-24 -1.88139e-20 0.00139516 0.997818 8.59318e-05 0.152558 2.85175 0.00139516 0.997859 0.686999 0.00104669 0.00187971 0.000859318 0.455642 0.00187971 0.436461 0.000127907 1.02 0.887517 0.534726 0.285827 1.7164e-07 3.05822e-09 2389.9 3142.09 -0.0569538 0.482123 0.2776 0.254921 -0.593074 -0.1695 0.492437 -0.2682 -0.224245 1.511 1 0 296.118 0 2.06268 1.509 0.000299939 0.864528 0.646385 0.436672 0.405792 2.06293 129.939 83.6174 18.7033 60.7202 0.00403782 0 -40 10
0.61 1.76794e-08 2.53888e-06 0.0851994 0.0851954 0.0120419 8.0361e-06 0.00115403 0.106499 0.0006571 0.107152 0.864113 101.866 0.24545 0.724189 4.13376 0.0545495 0.0389977 0.961002 0.019861 0.0042525 0.0191236 0.00409209 0.00513902 0.0058764 0.205561 0.235056 57.9769 -87.8948 126.145 15.9782 145.013 0.000142394 0.267099 192.913 0.310676 0.0673844 0.00409506 0.000561623 0.00138265 0.98699 0.991734 -2.97318e-06 -85.6676 0.0929868 31194.4 300.805 0.98352 0.319147 0.738668 0.738664 9.99958 2.98087e-06 1.19234e-05 0.130739 0.980044 0.930751 -0.0132932 4.89693e-06 0.501247 -1.88216e-20 6.93348e-24 -1.88147e-20 0.00139516 0.997818 8.59318e-05 0.152558 2.85175 0.00139516 0.997858 0.687108 0.00104671 0.00187971 0.000859318 0.455642 0.00187971 0.43647 0.00012791 1.02 0.887518 0.534726 0.285828 1.7164e-07 3.05824e-09 2389.88 3141.93 -0.0569429 0.482123 0.2776 0.254911 -0.593075 -0.169501 0.492468 -0.268198 -0.224279 1.512 1 0 296.129 0 2.06286 1.51 0.000299939 0.864458 0.646441 0.436394 0.405822 2.06311 129.949 83.6193 18.7034 60.7211 0.00403774 0 -40 10
0.611 1.77084e-08 2.53888e-06 0.0852822 0.0852782 0.0120419 8.04926e-06 0.00115403 0.106603 0.000657104 0.107255 0.864167 101.866 0.245444 0.724269 4.13389 0.0545558 0.0389989 0.961001 0.0198608 0.00425263 0.0191234 0.00409219 0.00513918 0.00587655 0.205567 0.235062 57.977 -87.8948 126.146 15.9782 145.013 0.000142387 0.2671 192.913 0.310675 0.0673844 0.00409506 0.000561623 0.00138265 0.98699 0.991734 -2.9732e-06 -85.6676 0.0929868 31194.4 300.809 0.98352 0.319147 0.738631 0.738627 9.99958 2.98087e-06 1.19234e-05 0.13074 0.980055 0.930756 -0.0132932 4.89696e-06 0.501252 -1.88224e-20 6.93382e-24 -1.88155e-20 0.00139516 0.997818 8.59319e-05 0.152559 2.85175 0.00139516 0.997858 0.687217 0.00104673 0.00187971 0.000859319 0.455642 0.00187971 0.43648 0.000127914 1.02 0.887519 0.534726 0.28583 1.71641e-07 3.05826e-09 2389.86 3141.77 -0.0569321 0.482123 0.2776 0.254901 -0.593077 -0.169501 0.4925 -0.268196 -0.224313 1.513 1 0 296.14 0 2.06304 1.511 0.000299939 0.864388 0.646496 0.436116 0.405852 2.06329 129.958 83.6211 18.7035 60.722 0.00403767 0 -40 10
0.612 1.77373e-08 2.53888e-06 0.0853649 0.0853609 0.0120419 8.06242e-06 0.00115403 0.106706 0.000657108 0.107359 0.864222 101.866 0.245438 0.724348 4.13402 0.0545621 0.0390001 0.961 0.0198607 0.00425275 0.0191233 0.0040923 0.00513933 0.00587671 0.205573 0.235068 57.977 -87.8949 126.146 15.9781 145.013 0.00014238 0.2671 192.912 0.310675 0.0673843 0.00409506 0.000561624 0.00138265 0.98699 0.991734 -2.97321e-06 -85.6676 0.0929869 31194.4 300.812 0.98352 0.319147 0.738594 0.738589 9.99958 2.98088e-06 1.19234e-05 0.130741 0.980066 0.930761 -0.0132932 4.89699e-06 0.501257 -1.88232e-20 6.93415e-24 -1.88163e-20 0.00139517 0.997818 8.5932e-05 0.152559 2.85175 0.00139517 0.997858 0.687326 0.00104675 0.00187971 0.00085932 0.455641 0.00187971 0.436489 0.000127917 1.02 0.88752 0.534725 0.285831 1.71641e-07 3.05828e-09 2389.85 3141.61 -0.0569214 0.482123 0.2776 0.254891 -0.593079 -0.169501 0.492531 -0.268194 -0.224346 1.514 1 0 296.151 0 2.06321 1.512 0.000299938 0.864318 0.646551 0.435839 0.405882 2.06346 129.968 83.6229 18.7036 60.7229 0.00403759 0 -40 10
0.613 1.77663e-08 2.53888e-06 0.0854476 0.0854436 0.0120419 8.07558e-06 0.00115403 0.106809 0.000657112 0.107462 0.864276 101.866 0.245432 0.724427 4.13415 0.0545684 0.0390014 0.960999 0.0198605 0.00425288 0.0191231 0.0040924 0.00513949 0.00587686 0.20558 0.235074 57.9771 -87.8949 126.147 15.9781 145.013 0.000142372 0.2671 192.912 0.310675 0.0673843 0.00409506 0.000561624 0.00138265 0.98699 0.991734 -2.97322e-06 -85.6676 0.092987 31194.4 300.816 0.98352 0.319147 0.738557 0.738552 9.99958 2.98088e-06 1.19234e-05 0.130742 0.980077 0.930766 -0.0132932 4.89702e-06 0.501262 -1.88241e-20 6.93448e-24 -1.88171e-20 0.00139517 0.997818 8.59321e-05 0.152559 2.85175 0.00139517 0.997858 0.687435 0.00104677 0.00187971 0.000859321 0.455641 0.00187971 0.436498 0.000127921 1.02 0.887521 0.534725 0.285832 1.71641e-07 3.05831e-09 2389.83 3141.45 -0.0569107 0.482123 0.277599 0.254881 -0.593081 -0.169501 0.492562 -0.268192 -0.224379 1.515 1 0 296.162 0 2.06339 1.513 0.000299938 0.864249 0.646607 0.435563 0.405911 2.06364 129.977 83.6248 18.7037 60.7238 0.00403752 0 -40 10
0.614 1.77952e-08 2.53888e-06 0.0855301 0.0855262 0.0120419 8.08874e-06 0.00115404 0.106913 0.000657116 0.107565 0.864331 101.866 0.245425 0.724507 4.13428 0.0545748 0.0390026 0.960997 0.0198604 0.00425301 0.019123 0.00409251 0.00513965 0.00587702 0.205586 0.235081 57.9772 -87.8949 126.148 15.9781 145.013 0.000142365 0.2671 192.912 0.310674 0.0673842 0.00409507 0.000561625 0.00138265 0.98699 0.991734 -2.97324e-06 -85.6676 0.0929871 31194.3 300.819 0.98352 0.319147 0.73852 0.738516 9.99958 2.98089e-06 1.19234e-05 0.130744 0.980087 0.930771 -0.0132932 4.89704e-06 0.501268 -1.88249e-20 6.93482e-24 -1.88179e-20 0.00139517 0.997818 8.59321e-05 0.152559 2.85175 0.00139517 0.997857 0.687544 0.00104679 0.00187971 0.000859321 0.455641 0.00187971 0.436507 0.000127924 1.02 0.887522 0.534725 0.285834 1.71641e-07 3.05833e-09 2389.81 3141.29 -0.0569 0.482123 0.277599 0.254871 -0.593083 -0.169501 0.492593 -0.26819 -0.224412 1.516 1 0 296.173 0 2.06357 1.514 0.000299938 0.864179 0.646662 0.435287 0.405941 2.06382 129.986 83.6266 18.7038 60.7246 0.00403744 0 -40 10
0.615 1.78242e-08 2.53888e-06 0.0856127 0.0856087 0.0120419 8.1019e-06 0.00115404 0.107016 0.00065712 0.107668 0.864385 101.866 0.245419 0.724587 4.13441 0.0545811 0.0390038 0.960996 0.0198602 0.00425313 0.0191228 0.00409261 0.0051398 0.00587717 0.205592 0.235087 57.9772 -87.8949 126.148 15.978 145.013 0.000142358 0.2671 192.912 0.310674 0.0673842 0.00409507 0.000561626 0.00138266 0.98699 0.991734 -2.97325e-06 -85.6676 0.0929871 31194.3 300.822 0.98352 0.319147 0.738483 0.738479 9.99958 2.98089e-06 1.19235e-05 0.130745 0.980098 0.930776 -0.0132932 4.89707e-06 0.501273 -1.88257e-20 6.93515e-24 -1.88187e-20 0.00139517 0.997818 8.59322e-05 0.152559 2.85175 0.00139517 0.997857 0.687653 0.00104681 0.00187972 0.000859322 0.455641 0.00187971 0.436516 0.000127928 1.02 0.887523 0.534725 0.285835 1.71642e-07 3.05835e-09 2389.8 3141.14 -0.0568894 0.482123 0.277599 0.254861 -0.593085 -0.169501 0.492624 -0.268188 -0.224445 1.517 1 0 296.183 0 2.06374 1.515 0.000299938 0.864111 0.646717 0.435012 0.405971 2.06399 129.996 83.6284 18.704 60.7255 0.00403737 0 -40 10
0.616 1.78531e-08 2.53888e-06 0.0856951 0.0856912 0.0120418 8.11506e-06 0.00115404 0.107119 0.000657124 0.107771 0.86444 101.865 0.245413 0.724666 4.13454 0.0545874 0.0390051 0.960995 0.01986 0.00425326 0.0191227 0.00409272 0.00513996 0.00587733 0.205598 0.235093 57.9773 -87.8949 126.149 15.978 145.013 0.000142351 0.2671 192.912 0.310673 0.0673841 0.00409507 0.000561626 0.00138266 0.98699 0.991734 -2.97326e-06 -85.6676 0.0929872 31194.3 300.826 0.98352 0.319147 0.738447 0.738442 9.99958 2.9809e-06 1.19235e-05 0.130746 0.980109 0.93078 -0.0132932 4.8971e-06 0.501278 -1.88265e-20 6.93549e-24 -1.88195e-20 0.00139517 0.997818 8.59323e-05 0.152559 2.85175 0.00139517 0.997857 0.687761 0.00104683 0.00187972 0.000859323 0.455641 0.00187972 0.436525 0.000127931 1.02 0.887524 0.534724 0.285837 1.71642e-07 3.05837e-09 2389.78 3140.98 -0.0568789 0.482123 0.277598 0.254851 -0.593086 -0.169501 0.492655 -0.268186 -0.224478 1.518 1 0 296.194 0 2.06392 1.516 0.000299937 0.864042 0.646773 0.434738 0.406001 2.06417 130.005 83.6302 18.7041 60.7264 0.00403729 0 -40 10
0.617 1.78821e-08 2.53888e-06 0.0857775 0.0857736 0.0120418 8.12822e-06 0.00115404 0.107222 0.000657128 0.107874 0.864494 101.865 0.245406 0.724746 4.13467 0.0545938 0.0390063 0.960994 0.0198599 0.00425339 0.0191225 0.00409283 0.00514012 0.00587748 0.205605 0.235099 57.9773 -87.8949 126.15 15.9779 145.013 0.000142344 0.267101 192.912 0.310673 0.0673841 0.00409508 0.000561627 0.00138266 0.98699 0.991734 -2.97328e-06 -85.6676 0.0929873 31194.3 300.829 0.98352 0.319147 0.73841 0.738406 9.99958 2.9809e-06 1.19235e-05 0.130748 0.980119 0.930785 -0.0132932 4.89713e-06 0.501284 -1.88273e-20 6.93582e-24 -1.88203e-20 0.00139517 0.997818 8.59323e-05 0.152559 2.85175 0.00139517 0.997857 0.68787 0.00104685 0.00187972 0.000859323 0.45564 0.00187972 0.436534 0.000127935 1.02 0.887525 0.534724 0.285838 1.71642e-07 3.05839e-09 2389.76 3140.83 -0.0568684 0.482123 0.277598 0.254841 -0.593088 -0.169501 0.492686 -0.268184 -0.22451 1.519 1 0 296.205 0 2.0641 1.517 0.000299937 0.863974 0.646828 0.434464 0.40603 2.06434 130.015 83.632 18.7042 60.7272 0.00403722 0 -40 10
0.618 1.7911e-08 2.53888e-06 0.0858598 0.0858559 0.0120418 8.14138e-06 0.00115404 0.107325 0.000657132 0.107977 0.864549 101.865 0.2454 0.724826 4.1348 0.0546001 0.0390075 0.960992 0.0198597 0.00425352 0.0191224 0.00409293 0.00514027 0.00587764 0.205611 0.235105 57.9774 -87.8949 126.15 15.9779 145.013 0.000142337 0.267101 192.911 0.310673 0.067384 0.00409508 0.000561627 0.00138266 0.98699 0.991734 -2.97329e-06 -85.6676 0.0929874 31194.3 300.833 0.98352 0.319147 0.738374 0.73837 9.99958 2.9809e-06 1.19235e-05 0.130749 0.98013 0.93079 -0.0132932 4.89715e-06 0.501289 -1.88281e-20 6.93616e-24 -1.88211e-20 0.00139517 0.997818 8.59324e-05 0.152559 2.85176 0.00139517 0.997856 0.687979 0.00104687 0.00187972 0.000859324 0.45564 0.00187972 0.436543 0.000127938 1.02 0.887526 0.534724 0.285839 1.71642e-07 3.05841e-09 2389.75 3140.67 -0.0568579 0.482123 0.277598 0.254832 -0.59309 -0.169501 0.492716 -0.268182 -0.224543 1.52 1 0 296.215 0 2.06427 1.518 0.000299937 0.863906 0.646883 0.434191 0.40606 2.06452 130.024 83.6337 18.7043 60.7281 0.00403714 0 -40 10
0.619 1.794e-08 2.53888e-06 0.0859421 0.0859382 0.0120418 8.15454e-06 0.00115404 0.107428 0.000657136 0.10808 0.864604 101.865 0.245394 0.724906 4.13493 0.0546065 0.0390088 0.960991 0.0198596 0.00425365 0.0191222 0.00409304 0.00514043 0.00587779 0.205617 0.235112 57.9775 -87.8949 126.151 15.9779 145.013 0.00014233 0.267101 192.911 0.310672 0.067384 0.00409508 0.000561628 0.00138266 0.98699 0.991734 -2.9733e-06 -85.6676 0.0929875 31194.2 300.836 0.98352 0.319147 0.738338 0.738334 9.99958 2.98091e-06 1.19235e-05 0.13075 0.980141 0.930795 -0.0132932 4.89718e-06 0.501294 -1.88289e-20 6.93649e-24 -1.88219e-20 0.00139517 0.997818 8.59325e-05 0.15256 2.85176 0.00139517 0.997856 0.688087 0.00104689 0.00187972 0.000859325 0.45564 0.00187972 0.436552 0.000127941 1.02 0.887527 0.534723 0.285841 1.71643e-07 3.05843e-09 2389.73 3140.52 -0.0568475 0.482123 0.277598 0.254822 -0.593092 -0.169501 0.492746 -0.26818 -0.224575 1.521 1 0 296.226 0 2.06445 1.519 0.000299937 0.863838 0.646938 0.433919 0.40609 2.0647 130.034 83.6355 18.7044 60.729 0.00403707 0 -40 10
0.62 1.79689e-08 2.53888e-06 0.0860243 0.0860204 0.0120418 8.1677e-06 0.00115404 0.10753 0.000657139 0.108183 0.864659 101.865 0.245387 0.724986 4.13506 0.0546129 0.03901 0.96099 0.0198594 0.00425377 0.0191221 0.00409315 0.00514059 0.00587795 0.205624 0.235118 57.9775 -87.8949 126.152 15.9778 145.013 0.000142323 0.267101 192.911 0.310672 0.067384 0.00409508 0.000561629 0.00138267 0.98699 0.991734 -2.97332e-06 -85.6675 0.0929875 31194.2 300.84 0.98352 0.319147 0.738302 0.738298 9.99958 2.98091e-06 1.19235e-05 0.130752 0.980151 0.9308 -0.0132932 4.89721e-06 0.5013 -1.88297e-20 6.93683e-24 -1.88227e-20 0.00139517 0.997818 8.59326e-05 0.15256 2.85176 0.00139517 0.997856 0.688196 0.00104691 0.00187972 0.000859326 0.45564 0.00187972 0.436562 0.000127945 1.02 0.887528 0.534723 0.285842 1.71643e-07 3.05845e-09 2389.72 3140.36 -0.0568372 0.482123 0.277597 0.254812 -0.593094 -0.169501 0.492776 -0.268178 -0.224607 1.522 1 0 296.237 0 2.06463 1.52 0.000299936 0.86377 0.646994 0.433647 0.406119 2.06487 130.043 83.6373 18.7045 60.7298 0.004037 0 -40 10
0.621 1.79979e-08 2.53888e-06 0.0861064 0.0861025 0.0120418 8.18086e-06 0.00115404 0.107633 0.000657143 0.108286 0.864714 101.865 0.245381 0.725067 4.1352 0.0546192 0.0390113 0.960989 0.0198593 0.0042539 0.0191219 0.00409325 0.00514075 0.00587811 0.20563 0.235124 57.9776 -87.8949 126.152 15.9778 145.013 0.000142316 0.267101 192.911 0.310671 0.0673839 0.00409509 0.000561629 0.00138267 0.98699 0.991734 -2.97333e-06 -85.6675 0.0929876 31194.2 300.843 0.98352 0.319147 0.738266 0.738262 9.99958 2.98092e-06 1.19236e-05 0.130753 0.980162 0.930804 -0.0132932 4.89724e-06 0.501305 -1.88305e-20 6.93716e-24 -1.88235e-20 0.00139517 0.997818 8.59326e-05 0.15256 2.85176 0.00139517 0.997856 0.688304 0.00104693 0.00187972 0.000859326 0.45564 0.00187972 0.436571 0.000127948 1.02 0.887529 0.534723 0.285844 1.71643e-07 3.05847e-09 2389.7 3140.21 -0.0568268 0.482123 0.277597 0.254803 -0.593095 -0.169501 0.492806 -0.268176 -0.224639 1.523 1 0 296.247 0 2.0648 1.521 0.000299936 0.863703 0.647049 0.433376 0.406149 2.06505 130.053 83.6391 18.7046 60.7307 0.00403692 0 -40 10
0.622 1.80269e-08 2.53888e-06 0.0861885 0.0861846 0.0120418 8.19402e-06 0.00115404 0.107736 0.000657147 0.108388 0.864768 101.865 0.245374 0.725147 4.13533 0.0546256 0.0390125 0.960987 0.0198591 0.00425403 0.0191217 0.00409336 0.00514091 0.00587826 0.205636 0.235131 57.9777 -87.8949 126.153 15.9778 145.013 0.00014231 0.267102 192.911 0.310671 0.0673839 0.00409509 0.00056163 0.00138267 0.98699 0.991734 -2.97334e-06 -85.6675 0.0929877 31194.2 300.847 0.98352 0.319147 0.738231 0.738226 9.99958 2.98092e-06 1.19236e-05 0.130754 0.980172 0.930809 -0.0132932 4.89726e-06 0.50131 -1.88313e-20 6.9375e-24 -1.88243e-20 0.00139518 0.997818 8.59327e-05 0.15256 2.85176 0.00139518 0.997855 0.688413 0.00104695 0.00187972 0.000859327 0.455639 0.00187972 0.43658 0.000127952 1.02 0.88753 0.534723 0.285845 1.71643e-07 3.05849e-09 2389.68 3140.06 -0.0568166 0.482124 0.277597 0.254793 -0.593097 -0.169501 0.492836 -0.268174 -0.224671 1.524 1 0 296.258 0 2.06498 1.522 0.000299936 0.863636 0.647104 0.433106 0.406179 2.06522 130.062 83.6408 18.7047 60.7315 0.00403685 0 -40 10
0.623 1.80558e-08 2.53888e-06 0.0862705 0.0862666 0.0120418 8.20718e-06 0.00115404 0.107838 0.000657151 0.108491 0.864823 101.865 0.245368 0.725227 4.13546 0.054632 0.0390138 0.960986 0.0198589 0.00425416 0.0191216 0.00409347 0.00514107 0.00587842 0.205643 0.235137 57.9777 -87.8949 126.154 15.9777 145.013 0.000142303 0.267102 192.911 0.310671 0.0673838 0.00409509 0.00056163 0.00138267 0.98699 0.991734 -2.97336e-06 -85.6675 0.0929878 31194.2 300.85 0.98352 0.319147 0.738195 0.738191 9.99958 2.98093e-06 1.19236e-05 0.130756 0.980183 0.930814 -0.0132932 4.89729e-06 0.501316 -1.88321e-20 6.93783e-24 -1.88251e-20 0.00139518 0.997818 8.59328e-05 0.15256 2.85176 0.00139518 0.997855 0.688521 0.00104697 0.00187973 0.000859328 0.455639 0.00187972 0.436589 0.000127955 1.02 0.887531 0.534722 0.285846 1.71644e-07 3.05852e-09 2389.67 3139.91 -0.0568064 0.482124 0.277596 0.254783 -0.593099 -0.169501 0.492866 -0.268172 -0.224703 1.525 1 0 296.268 0 2.06515 1.523 0.000299936 0.86357 0.647159 0.432837 0.406208 2.0654 130.071 83.6426 18.7048 60.7323 0.00403678 0 -40 10
0.624 1.80848e-08 2.53888e-06 0.0863524 0.0863486 0.0120417 8.22034e-06 0.00115404 0.10794 0.000657155 0.108593 0.864878 101.864 0.245362 0.725308 4.1356 0.0546384 0.0390151 0.960985 0.0198588 0.00425429 0.0191214 0.00409358 0.00514123 0.00587858 0.205649 0.235143 57.9778 -87.8949 126.154 15.9777 145.013 0.000142296 0.267102 192.911 0.31067 0.0673838 0.00409509 0.000561631 0.00138267 0.98699 0.991734 -2.97337e-06 -85.6675 0.0929878 31194.1 300.854 0.98352 0.319147 0.73816 0.738155 9.99958 2.98093e-06 1.19236e-05 0.130757 0.980193 0.930819 -0.0132932 4.89732e-06 0.501321 -1.88329e-20 6.93817e-24 -1.88259e-20 0.00139518 0.997818 8.59329e-05 0.15256 2.85176 0.00139518 0.997855 0.68863 0.00104699 0.00187973 0.000859329 0.455639 0.00187973 0.436598 0.000127959 1.02 0.887532 0.534722 0.285848 1.71644e-07 3.05854e-09 2389.65 3139.76 -0.0567962 0.482124 0.277596 0.254774 -0.593101 -0.169501 0.492896 -0.26817 -0.224735 1.526 1 0 296.278 0 2.06533 1.524 0.000299935 0.863504 0.647214 0.432568 0.406238 2.06558 130.081 83.6443 18.7049 60.7332 0.00403671 0 -40 10
0.625 1.81137e-08 2.53888e-06 0.0864343 0.0864304 0.0120417 8.2335e-06 0.00115404 0.108043 0.000657159 0.108695 0.864934 101.864 0.245355 0.725389 4.13573 0.0546448 0.0390163 0.960984 0.0198586 0.00425442 0.0191213 0.00409369 0.00514139 0.00587874 0.205656 0.23515 57.9778 -87.8949 126.155 15.9776 145.013 0.000142289 0.267102 192.91 0.31067 0.0673837 0.0040951 0.000561632 0.00138268 0.98699 0.991734 -2.97339e-06 -85.6675 0.0929879 31194.1 300.857 0.98352 0.319147 0.738125 0.73812 9.99958 2.98094e-06 1.19236e-05 0.130758 0.980204 0.930823 -0.0132932 4.89735e-06 0.501327 -1.88337e-20 6.9385e-24 -1.88267e-20 0.00139518 0.997818 8.59329e-05 0.15256 2.85176 0.00139518 0.997855 0.688738 0.00104701 0.00187973 0.000859329 0.455639 0.00187973 0.436607 0.000127962 1.02 0.887533 0.534722 0.285849 1.71644e-07 3.05856e-09 2389.63 3139.61 -0.0567861 0.482124 0.277596 0.254764 -0.593103 -0.169502 0.492925 -0.268168 -0.224766 1.527 1 0 296.289 0 2.06551 1.525 0.000299935 0.863438 0.647269 0.4323 0.406267 2.06575 130.09 83.646 18.705 60.734 0.00403664 0 -40 10
0.626 1.81427e-08 2.53888e-06 0.0865161 0.0865122 0.0120417 8.24666e-06 0.00115404 0.108145 0.000657163 0.108798 0.864989 101.864 0.245349 0.725469 4.13587 0.0546512 0.0390176 0.960982 0.0198585 0.00425455 0.0191211 0.00409379 0.00514155 0.0058789 0.205662 0.235156 57.9779 -87.8949 126.155 15.9776 145.013 0.000142282 0.267102 192.91 0.31067 0.0673837 0.0040951 0.000561632 0.00138268 0.98699 0.991734 -2.9734e-06 -85.6675 0.092988 31194.1 300.861 0.98352 0.319147 0.73809 0.738085 9.99958 2.98094e-06 1.19237e-05 0.13076 0.980214 0.930828 -0.0132932 4.89737e-06 0.501332 -1.88345e-20 6.93884e-24 -1.88275e-20 0.00139518 0.997818 8.5933e-05 0.152561 2.85176 0.00139518 0.997854 0.688847 0.00104702 0.00187973 0.00085933 0.455639 0.00187973 0.436616 0.000127966 1.02 0.887534 0.534721 0.285851 1.71644e-07 3.05858e-09 2389.62 3139.46 -0.056776 0.482124 0.277596 0.254755 -0.593104 -0.169502 0.492954 -0.268166 -0.224797 1.528 1 0 296.299 0 2.06568 1.526 0.000299935 0.863372 0.647324 0.432032 0.406297 2.06593 130.1 83.6478 18.7051 60.7349 0.00403656 0 -40 10
0.627 1.81716e-08 2.53888e-06 0.0865978 0.086594 0.0120417 8.25982e-06 0.00115404 0.108247 0.000657166 0.1089 0.865044 101.864 0.245342 0.72555 4.136 0.0546576 0.0390189 0.960981 0.0198583 0.00425468 0.0191209 0.0040939 0.00514171 0.00587906 0.205668 0.235162 57.978 -87.8949 126.156 15.9776 145.013 0.000142276 0.267102 192.91 0.310669 0.0673836 0.0040951 0.000561633 0.00138268 0.98699 0.991734 -2.97341e-06 -85.6675 0.0929881 31194.1 300.864 0.98352 0.319147 0.738055 0.73805 9.99958 2.98094e-06 1.19237e-05 0.130761 0.980224 0.930833 -0.0132932 4.8974e-06 0.501338 -1.88353e-20 6.93918e-24 -1.88283e-20 0.00139518 0.997818 8.59331e-05 0.152561 2.85176 0.00139518 0.997854 0.688955 0.00104704 0.00187973 0.000859331 0.455638 0.00187973 0.436625 0.000127969 1.02 0.887535 0.534721 0.285852 1.71644e-07 3.0586e-09 2389.6 3139.31 -0.056766 0.482124 0.277595 0.254746 -0.593106 -0.169502 0.492984 -0.268164 -0.224828 1.529 1 0 296.309 0 2.06586 1.527 0.000299935 0.863306 0.647379 0.431765 0.406327 2.0661 130.109 83.6495 18.7052 60.7357 0.00403649 0 -40 10
0.628 1.82006e-08 2.53888e-06 0.0866794 0.0866757 0.0120417 8.27298e-06 0.00115404 0.108349 0.00065717 0.109002 0.865099 101.864 0.245336 0.725631 4.13614 0.0546641 0.0390201 0.96098 0.0198581 0.00425482 0.0191208 0.00409401 0.00514187 0.00587922 0.205675 0.235169 57.978 -87.8949 126.157 15.9775 145.013 0.000142269 0.267103 192.91 0.310669 0.0673836 0.00409511 0.000561633 0.00138268 0.98699 0.991734 -2.97343e-06 -85.6675 0.0929882 31194.1 300.868 0.98352 0.319147 0.73802 0.738015 9.99958 2.98095e-06 1.19237e-05 0.130762 0.980235 0.930837 -0.0132932 4.89743e-06 0.501343 -1.88361e-20 6.93951e-24 -1.88291e-20 0.00139518 0.997818 8.59331e-05 0.152561 2.85176 0.00139518 0.997854 0.689063 0.00104706 0.00187973 0.000859331 0.455638 0.00187973 0.436634 0.000127973 1.02 0.887536 0.534721 0.285854 1.71645e-07 3.05862e-09 2389.58 3139.16 -0.056756 0.482124 0.277595 0.254736 -0.593108 -0.169502 0.493013 -0.268162 -0.22486 1.53 1 0 296.319 0 2.06603 1.528 0.000299934 0.863241 0.647434 0.431499 0.406356 2.06628 130.118 83.6512 18.7053 60.7365 0.00403642 0 -40 10
0.629 1.82295e-08 2.53888e-06 0.086761 0.0867573 0.0120417 8.28614e-06 0.00115404 0.108451 0.000657174 0.109104 0.865155 101.864 0.245329 0.725712 4.13627 0.0546705 0.0390214 0.960979 0.019858 0.00425495 0.0191206 0.00409412 0.00514203 0.00587938 0.205681 0.235175 57.9781 -87.8949 126.157 15.9775 145.013 0.000142262 0.267103 192.91 0.310668 0.0673835 0.00409511 0.000561634 0.00138268 0.98699 0.991734 -2.97344e-06 -85.6675 0.0929882 31194 300.872 0.98352 0.319147 0.737985 0.737981 9.99958 2.98095e-06 1.19237e-05 0.130764 0.980245 0.930842 -0.0132932 4.89746e-06 0.501349 -1.88369e-20 6.93985e-24 -1.88299e-20 0.00139518 0.997818 8.59332e-05 0.152561 2.85176 0.00139518 0.997854 0.689172 0.00104708 0.00187973 0.000859332 0.455638 0.00187973 0.436643 0.000127976 1.02 0.887537 0.534721 0.285855 1.71645e-07 3.05864e-09 2389.57 3139.01 -0.056746 0.482124 0.277595 0.254727 -0.59311 -0.169502 0.493041 -0.268159 -0.22489 1.531 1 0 296.329 0 2.06621 1.529 0.000299934 0.863176 0.647488 0.431234 0.406386 2.06645 130.128 83.6529 18.7054 60.7373 0.00403635 0 -40 10
0.63 1.82585e-08 2.53888e-06 0.0868426 0.0868388 0.0120417 8.2993e-06 0.00115404 0.108553 0.000657178 0.109206 0.86521 101.864 0.245323 0.725793 4.13641 0.0546769 0.0390227 0.960977 0.0198578 0.00425508 0.0191205 0.00409423 0.0051422 0.00587954 0.205688 0.235181 57.9782 -87.8949 126.158 15.9775 145.013 0.000142256 0.267103 192.91 0.310668 0.0673835 0.00409511 0.000561635 0.00138269 0.98699 0.991734 -2.97345e-06 -85.6675 0.0929883 31194 300.875 0.98352 0.319147 0.737951 0.737946 9.99958 2.98096e-06 1.19237e-05 0.130765 0.980255 0.930846 -0.0132932 4.89748e-06 0.501354 -1.88377e-20 6.94018e-24 -1.88307e-20 0.00139518 0.997818 8.59333e-05 0.152561 2.85177 0.00139518 0.997853 0.68928 0.0010471 0.00187974 0.000859333 0.455638 0.00187973 0.436652 0.000127979 1.02 0.887538 0.53472 0.285856 1.71645e-07 3.05866e-09 2389.55 3138.86 -0.0567362 0.482124 0.277594 0.254718 -0.593111 -0.169502 0.49307 -0.268157 -0.224921 1.532 1 0 296.339 0 2.06638 1.53 0.000299934 0.863112 0.647543 0.430969 0.406415 2.06663 130.137 83.6546 18.7055 60.7381 0.00403628 0 -40 10
0.631 1.82874e-08 2.53888e-06 0.0869241 0.0869203 0.0120417 8.31246e-06 0.00115404 0.108655 0.000657181 0.109308 0.865265 101.863 0.245317 0.725874 4.13654 0.0546834 0.039024 0.960976 0.0198576 0.00425521 0.0191203 0.00409434 0.00514236 0.0058797 0.205694 0.235188 57.9782 -87.8949 126.159 15.9774 145.013 0.000142249 0.267103 192.91 0.310668 0.0673834 0.00409511 0.000561635 0.00138269 0.98699 0.991734 -2.97347e-06 -85.6675 0.0929884 31194 300.879 0.98352 0.319147 0.737916 0.737912 9.99958 2.98096e-06 1.19237e-05 0.130766 0.980265 0.930851 -0.0132932 4.89751e-06 0.50136 -1.88385e-20 6.94052e-24 -1.88315e-20 0.00139519 0.997818 8.59334e-05 0.152561 2.85177 0.00139519 0.997853 0.689388 0.00104712 0.00187974 0.000859334 0.455638 0.00187974 0.436661 0.000127983 1.02 0.887539 0.53472 0.285858 1.71645e-07 3.05869e-09 2389.53 3138.72 -0.0567263 0.482124 0.277594 0.254709 -0.593113 -0.169502 0.493099 -0.268155 -0.224952 1.533 1 0 296.349 0 2.06656 1.531 0.000299933 0.863047 0.647598 0.430705 0.406445 2.0668 130.146 83.6563 18.7056 60.739 0.00403621 0 -40 10
0.632 1.83164e-08 2.53888e-06 0.0870055 0.0870017 0.0120416 8.32562e-06 0.00115404 0.108757 0.000657185 0.109409 0.865321 101.863 0.24531 0.725956 4.13668 0.0546899 0.0390253 0.960975 0.0198575 0.00425534 0.0191201 0.00409445 0.00514252 0.00587986 0.205701 0.235194 57.9783 -87.8949 126.159 15.9774 145.013 0.000142242 0.267103 192.909 0.310667 0.0673834 0.00409512 0.000561636 0.00138269 0.98699 0.991734 -2.97348e-06 -85.6674 0.0929885 31194 300.882 0.98352 0.319147 0.737882 0.737878 9.99958 2.98097e-06 1.19238e-05 0.130768 0.980276 0.930856 -0.0132932 4.89754e-06 0.501365 -1.88393e-20 6.94085e-24 -1.88323e-20 0.00139519 0.997818 8.59334e-05 0.152561 2.85177 0.00139519 0.997853 0.689496 0.00104714 0.00187974 0.000859334 0.455637 0.00187974 0.43667 0.000127986 1.02 0.88754 0.53472 0.285859 1.71646e-07 3.05871e-09 2389.52 3138.57 -0.0567165 0.482124 0.277594 0.254699 -0.593115 -0.169502 0.493127 -0.268153 -0.224982 1.534 1 0 296.359 0 2.06673 1.532 0.000299933 0.862983 0.647653 0.430441 0.406474 2.06698 130.156 83.658 18.7057 60.7398 0.00403614 0 -40 10
0.633 1.83453e-08 2.53888e-06 0.0870868 0.0870831 0.0120416 8.33878e-06 0.00115404 0.108858 0.000657189 0.109511 0.865376 101.863 0.245304 0.726037 4.13682 0.0546963 0.0390266 0.960973 0.0198573 0.00425548 0.01912 0.00409456 0.00514268 0.00588002 0.205707 0.235201 57.9784 -87.8949 126.16 15.9773 145.013 0.000142236 0.267103 192.909 0.310667 0.0673833 0.00409512 0.000561637 0.00138269 0.98699 0.991734 -2.97349e-06 -85.6674 0.0929886 31194 300.886 0.98352 0.319147 0.737848 0.737844 9.99958 2.98097e-06 1.19238e-05 0.130769 0.980286 0.93086 -0.0132932 4.89757e-06 0.501371 -1.88401e-20 6.94119e-24 -1.88331e-20 0.00139519 0.997818 8.59335e-05 0.152562 2.85177 0.00139519 0.997853 0.689604 0.00104716 0.00187974 0.000859335 0.455637 0.00187974 0.436679 0.00012799 1.02 0.887541 0.534719 0.285861 1.71646e-07 3.05873e-09 2389.5 3138.42 -0.0567068 0.482124 0.277594 0.25469 -0.593116 -0.169502 0.493156 -0.268151 -0.225013 1.535 1 0 296.369 0 2.06691 1.533 0.000299933 0.862919 0.647708 0.430178 0.406503 2.06715 130.165 83.6596 18.7058 60.7406 0.00403607 0 -40 10
0.634 1.83743e-08 2.53888e-06 0.0871681 0.0871643 0.0120416 8.35194e-06 0.00115404 0.10896 0.000657193 0.109613 0.865432 101.863 0.245297 0.726118 4.13695 0.0547028 0.0390279 0.960972 0.0198572 0.00425561 0.0191198 0.00409467 0.00514285 0.00588018 0.205714 0.235207 57.9784 -87.8949 126.16 15.9773 145.013 0.000142229 0.267104 192.909 0.310666 0.0673833 0.00409512 0.000561637 0.00138269 0.98699 0.991734 -2.97351e-06 -85.6674 0.0929886 31193.9 300.89 0.98352 0.319147 0.737814 0.73781 9.99958 2.98098e-06 1.19238e-05 0.13077 0.980296 0.930865 -0.0132932 4.8976e-06 0.501376 -1.88409e-20 6.94152e-24 -1.88339e-20 0.00139519 0.997818 8.59336e-05 0.152562 2.85177 0.00139519 0.997852 0.689712 0.00104718 0.00187974 0.000859336 0.455637 0.00187974 0.436688 0.000127993 1.02 0.887543 0.534719 0.285862 1.71646e-07 3.05875e-09 2389.48 3138.28 -0.0566971 0.482124 0.277593 0.254681 -0.593118 -0.169502 0.493184 -0.268149 -0.225043 1.536 1 0 296.379 0 2.06708 1.534 0.000299933 0.862856 0.647762 0.429916 0.406533 2.06733 130.175 83.6613 18.7059 60.7414 0.004036 0 -40 10
0.635 1.84032e-08 2.53888e-06 0.0872493 0.0872456 0.0120416 8.3651e-06 0.00115404 0.109062 0.000657196 0.109714 0.865488 101.863 0.245291 0.7262 4.13709 0.0547093 0.0390292 0.960971 0.019857 0.00425574 0.0191197 0.00409478 0.00514301 0.00588035 0.20572 0.235214 57.9785 -87.8949 126.161 15.9773 145.013 0.000142223 0.267104 192.909 0.310666 0.0673832 0.00409512 0.000561638 0.0013827 0.98699 0.991734 -2.97352e-06 -85.6674 0.0929887 31193.9 300.893 0.98352 0.319147 0.73778 0.737776 9.99958 2.98098e-06 1.19238e-05 0.130772 0.980306 0.930869 -0.0132932 4.89762e-06 0.501382 -1.88417e-20 6.94186e-24 -1.88348e-20 0.00139519 0.997818 8.59337e-05 0.152562 2.85177 0.00139519 0.997852 0.68982 0.0010472 0.00187974 0.000859337 0.455637 0.00187974 0.436697 0.000127997 1.02 0.887544 0.534719 0.285864 1.71646e-07 3.05877e-09 2389.47 3138.14 -0.0566874 0.482124 0.277593 0.254672 -0.59312 -0.169502 0.493212 -0.268147 -0.225073 1.537 1 0 296.389 0 2.06726 1.535 0.000299932 0.862793 0.647817 0.429655 0.406562 2.0675 130.184 83.663 18.706 60.7422 0.00403593 0 -40 10
0.636 1.84322e-08 2.53888e-06 0.0873304 0.0873267 0.0120416 8.37826e-06 0.00115404 0.109163 0.0006572 0.109816 0.865543 101.863 0.245284 0.726282 4.13723 0.0547158 0.0390305 0.96097 0.0198568 0.00425588 0.0191195 0.00409489 0.00514318 0.00588051 0.205727 0.23522 57.9785 -87.8949 126.162 15.9772 145.013 0.000142216 0.267104 192.909 0.310666 0.0673832 0.00409513 0.000561638 0.0013827 0.98699 0.991734 -2.97354e-06 -85.6674 0.0929888 31193.9 300.897 0.98352 0.319147 0.737747 0.737742 9.99958 2.98098e-06 1.19238e-05 0.130773 0.980316 0.930874 -0.0132932 4.89765e-06 0.501387 -1.88425e-20 6.9422e-24 -1.88356e-20 0.00139519 0.997818 8.59337e-05 0.152562 2.85177 0.00139519 0.997852 0.689928 0.00104722 0.00187974 0.000859337 0.455637 0.00187974 0.436706 0.000128 1.02 0.887545 0.534719 0.285865 1.71647e-07 3.05879e-09 2389.45 3137.99 -0.0566778 0.482125 0.277593 0.254663 -0.593121 -0.169502 0.49324 -0.268145 -0.225103 1.538 1 0 296.399 0 2.06743 1.536 0.000299932 0.86273 0.647872 0.429394 0.406592 2.06768 130.193 83.6646 18.7061 60.743 0.00403587 0 -40 10
0.637 1.84611e-08 2.53888e-06 0.0874115 0.0874078 0.0120416 8.39142e-06 0.00115404 0.109264 0.000657204 0.109917 0.865599 101.863 0.245278 0.726363 4.13737 0.0547223 0.0390318 0.960968 0.0198567 0.00425601 0.0191193 0.00409501 0.00514334 0.00588067 0.205734 0.235227 57.9786 -87.8949 126.162 15.9772 145.013 0.00014221 0.267104 192.909 0.310665 0.0673831 0.00409513 0.000561639 0.0013827 0.98699 0.991734 -2.97355e-06 -85.6674 0.0929889 31193.9 300.9 0.98352 0.319147 0.737713 0.737709 9.99958 2.98099e-06 1.19239e-05 0.130774 0.980326 0.930878 -0.0132932 4.89768e-06 0.501393 -1.88433e-20 6.94253e-24 -1.88364e-20 0.00139519 0.997818 8.59338e-05 0.152562 2.85177 0.00139519 0.997852 0.690036 0.00104724 0.00187974 0.000859338 0.455636 0.00187974 0.436715 0.000128004 1.02 0.887546 0.534718 0.285866 1.71647e-07 3.05881e-09 2389.43 3137.85 -0.0566682 0.482125 0.277592 0.254654 -0.593123 -0.169502 0.493268 -0.268143 -0.225133 1.539 1 0 296.409 0 2.06761 1.537 0.000299932 0.862667 0.647926 0.429133 0.406621 2.06785 130.203 83.6663 18.7062 60.7438 0.0040358 0 -40 10
0.638 1.84901e-08 2.53888e-06 0.0874925 0.0874888 0.0120416 8.40458e-06 0.00115404 0.109366 0.000657207 0.110018 0.865655 101.862 0.245271 0.726445 4.13751 0.0547288 0.0390331 0.960967 0.0198565 0.00425615 0.0191192 0.00409512 0.00514351 0.00588084 0.20574 0.235233 57.9787 -87.895 126.163 15.9772 145.013 0.000142203 0.267104 192.909 0.310665 0.0673831 0.00409513 0.00056164 0.0013827 0.98699 0.991734 -2.97356e-06 -85.6674 0.092989 31193.8 300.904 0.98352 0.319147 0.73768 0.737676 9.99958 2.98099e-06 1.19239e-05 0.130776 0.980336 0.930883 -0.0132932 4.89771e-06 0.501398 -1.88441e-20 6.94287e-24 -1.88372e-20 0.00139519 0.997818 8.59339e-05 0.152562 2.85177 0.00139519 0.997852 0.690144 0.00104726 0.00187975 0.000859339 0.455636 0.00187975 0.436724 0.000128007 1.02 0.887547 0.534718 0.285868 1.71647e-07 3.05883e-09 2389.42 3137.71 -0.0566587 0.482125 0.277592 0.254645 -0.593125 -0.169502 0.493295 -0.268141 -0.225162 1.54 1 0 296.418 0 2.06778 1.538 0.000299932 0.862605 0.647981 0.428874 0.40665 2.06802 130.212 83.6679 18.7063 60.7446 0.00403573 0 -40 10
0.639 1.8519e-08 2.53889e-06 0.0875735 0.0875698 0.0120415 8.41774e-06 0.00115404 0.109467 0.000657211 0.110119 0.865711 101.862 0.245265 0.726527 4.13765 0.0547353 0.0390344 0.960966 0.0198563 0.00425628 0.019119 0.00409523 0.00514367 0.005881 0.205747 0.23524 57.9787 -87.895 126.163 15.9771 145.013 0.000142197 0.267104 192.908 0.310664 0.067383 0.00409514 0.00056164 0.0013827 0.98699 0.991734 -2.97358e-06 -85.6674 0.092989 31193.8 300.908 0.98352 0.319147 0.737647 0.737642 9.99958 2.981e-06 1.19239e-05 0.130777 0.980346 0.930887 -0.0132932 4.89773e-06 0.501404 -1.88449e-20 6.94321e-24 -1.8838e-20 0.00139519 0.997818 8.59339e-05 0.152562 2.85177 0.00139519 0.997851 0.690252 0.00104728 0.00187975 0.000859339 0.455636 0.00187975 0.436733 0.00012801 1.02 0.887548 0.534718 0.285869 1.71647e-07 3.05886e-09 2389.4 3137.56 -0.0566492 0.482125 0.277592 0.254636 -0.593126 -0.169502 0.493323 -0.268139 -0.225192 1.541 1 0 296.428 0 2.06795 1.539 0.000299931 0.862543 0.648036 0.428615 0.40668 2.0682 130.221 83.6696 18.7063 60.7454 0.00403566 0 -40 10
0.64 1.8548e-08 2.53889e-06 0.0876543 0.0876507 0.0120415 8.4309e-06 0.00115404 0.109568 0.000657215 0.110221 0.865767 101.862 0.245258 0.726609 4.13779 0.0547418 0.0390357 0.960964 0.0198562 0.00425642 0.0191188 0.00409534 0.00514384 0.00588116 0.205754 0.235247 57.9788 -87.895 126.164 15.9771 145.013 0.000142191 0.267105 192.908 0.310664 0.067383 0.00409514 0.000561641 0.00138271 0.98699 0.991734 -2.97359e-06 -85.6674 0.0929891 31193.8 300.911 0.98352 0.319147 0.737614 0.737609 9.99958 2.981e-06 1.19239e-05 0.130779 0.980356 0.930892 -0.0132932 4.89776e-06 0.50141 -1.88457e-20 6.94354e-24 -1.88388e-20 0.00139519 0.997818 8.5934e-05 0.152563 2.85177 0.00139519 0.997851 0.69036 0.0010473 0.00187975 0.00085934 0.455636 0.00187975 0.436742 0.000128014 1.02 0.887549 0.534717 0.285871 1.71648e-07 3.05888e-09 2389.38 3137.42 -0.0566398 0.482125 0.277592 0.254627 -0.593128 -0.169502 0.49335 -0.268137 -0.225221 1.542 1 0 296.438 0 2.06813 1.54 0.000299931 0.862481 0.64809 0.428357 0.406709 2.06837 130.231 83.6712 18.7064 60.7462 0.00403559 0 -40 10
0.641 1.85769e-08 2.53889e-06 0.0877352 0.0877315 0.0120415 8.44406e-06 0.00115404 0.109669 0.000657218 0.110322 0.865823 101.862 0.245252 0.726691 4.13793 0.0547483 0.039037 0.960963 0.019856 0.00425655 0.0191187 0.00409545 0.00514401 0.00588133 0.20576 0.235253 57.9789 -87.895 126.165 15.977 145.013 0.000142184 0.267105 192.908 0.310664 0.067383 0.00409514 0.000561641 0.00138271 0.98699 0.991734 -2.9736e-06 -85.6674 0.0929892 31193.8 300.915 0.98352 0.319147 0.737581 0.737576 9.99958 2.98101e-06 1.19239e-05 0.13078 0.980366 0.930896 -0.0132932 4.89779e-06 0.501415 -1.88465e-20 6.94388e-24 -1.88396e-20 0.0013952 0.997818 8.59341e-05 0.152563 2.85177 0.0013952 0.997851 0.690468 0.00104732 0.00187975 0.000859341 0.455636 0.00187975 0.436751 0.000128017 1.02 0.88755 0.534717 0.285872 1.71648e-07 3.0589e-09 2389.37 3137.28 -0.0566304 0.482125 0.277591 0.254618 -0.59313 -0.169503 0.493377 -0.268135 -0.225251 1.543 1 0 296.447 0 2.0683 1.541 0.000299931 0.862419 0.648145 0.428099 0.406738 2.06855 130.24 83.6728 18.7065 60.7469 0.00403553 0 -40 10
0.642 1.86059e-08 2.53889e-06 0.0878159 0.0878123 0.0120415 8.45722e-06 0.00115404 0.10977 0.000657222 0.110423 0.865879 101.862 0.245245 0.726774 4.13807 0.0547549 0.0390384 0.960962 0.0198558 0.00425669 0.0191185 0.00409557 0.00514417 0.00588149 0.205767 0.23526 57.9789 -87.895 126.165 15.977 145.013 0.000142178 0.267105 192.908 0.310663 0.0673829 0.00409514 0.000561642 0.00138271 0.98699 0.991734 -2.97362e-06 -85.6674 0.0929893 31193.8 300.919 0.98352 0.319147 0.737548 0.737544 9.99958 2.98101e-06 1.19239e-05 0.130781 0.980376 0.9309 -0.0132932 4.89782e-06 0.501421 -1.88473e-20 6.94421e-24 -1.88404e-20 0.0013952 0.997818 8.59342e-05 0.152563 2.85178 0.0013952 0.997851 0.690575 0.00104734 0.00187975 0.000859342 0.455635 0.00187975 0.43676 0.000128021 1.02 0.887551 0.534717 0.285874 1.71648e-07 3.05892e-09 2389.35 3137.14 -0.0566211 0.482125 0.277591 0.25461 -0.593131 -0.169503 0.493404 -0.268133 -0.22528 1.544 1 0 296.457 0 2.06848 1.542 0.000299931 0.862358 0.648199 0.427842 0.406768 2.06872 130.249 83.6744 18.7066 60.7477 0.00403546 0 -40 10
0.643 1.86348e-08 2.53889e-06 0.0878966 0.087893 0.0120415 8.47038e-06 0.00115404 0.109871 0.000657226 0.110523 0.865935 101.862 0.245239 0.726856 4.13821 0.0547614 0.0390397 0.96096 0.0198557 0.00425682 0.0191183 0.00409568 0.00514434 0.00588166 0.205774 0.235266 57.979 -87.895 126.166 15.977 145.013 0.000142172 0.267105 192.908 0.310663 0.0673829 0.00409515 0.000561643 0.00138271 0.98699 0.991734 -2.97363e-06 -85.6673 0.0929894 31193.7 300.922 0.98352 0.319147 0.737515 0.737511 9.99958 2.98102e-06 1.1924e-05 0.130783 0.980385 0.930905 -0.0132932 4.89785e-06 0.501427 -1.88481e-20 6.94455e-24 -1.88412e-20 0.0013952 0.997818 8.59342e-05 0.152563 2.85178 0.0013952 0.997851 0.690683 0.00104736 0.00187975 0.000859342 0.455635 0.00187975 0.436769 0.000128024 1.02 0.887552 0.534716 0.285875 1.71648e-07 3.05894e-09 2389.33 3137 -0.0566118 0.482125 0.277591 0.254601 -0.593133 -0.169503 0.493431 -0.268131 -0.225309 1.545 1 0 296.466 0 2.06865 1.543 0.00029993 0.862297 0.648254 0.427586 0.406797 2.06889 130.259 83.676 18.7067 60.7485 0.00403539 0 -40 10
0.644 1.86638e-08 2.53889e-06 0.0879772 0.0879736 0.0120415 8.48354e-06 0.00115404 0.109972 0.000657229 0.110624 0.865991 101.862 0.245232 0.726938 4.13835 0.054768 0.039041 0.960959 0.0198555 0.00425696 0.0191182 0.00409579 0.00514451 0.00588183 0.20578 0.235273 57.979 -87.895 126.166 15.9769 145.013 0.000142165 0.267105 192.908 0.310662 0.0673828 0.00409515 0.000561643 0.00138271 0.98699 0.991734 -2.97365e-06 -85.6673 0.0929894 31193.7 300.926 0.98352 0.319147 0.737483 0.737478 9.99958 2.98102e-06 1.1924e-05 0.130784 0.980395 0.930909 -0.0132932 4.89787e-06 0.501432 -1.88489e-20 6.94489e-24 -1.8842e-20 0.0013952 0.997818 8.59343e-05 0.152563 2.85178 0.0013952 0.99785 0.690791 0.00104738 0.00187975 0.000859343 0.455635 0.00187975 0.436778 0.000128028 1.02 0.887553 0.534716 0.285876 1.71649e-07 3.05896e-09 2389.32 3136.86 -0.0566025 0.482125 0.27759 0.254592 -0.593135 -0.169503 0.493458 -0.268129 -0.225338 1.546 1 0 296.476 0 2.06882 1.544 0.00029993 0.862236 0.648308 0.42733 0.406826 2.06907 130.268 83.6776 18.7068 60.7493 0.00403533 0 -40 10
0.645 1.86927e-08 2.53889e-06 0.0880578 0.0880542 0.0120415 8.4967e-06 0.00115404 0.110072 0.000657233 0.110725 0.866048 101.862 0.245225 0.727021 4.13849 0.0547745 0.0390423 0.960958 0.0198553 0.0042571 0.019118 0.00409591 0.00514468 0.00588199 0.205787 0.23528 57.9791 -87.895 126.167 15.9769 145.013 0.000142159 0.267105 192.907 0.310662 0.0673828 0.00409515 0.000561644 0.00138272 0.98699 0.991734 -2.97366e-06 -85.6673 0.0929895 31193.7 300.93 0.98352 0.319147 0.737451 0.737446 9.99958 2.98103e-06 1.1924e-05 0.130786 0.980405 0.930913 -0.0132932 4.8979e-06 0.501438 -1.88497e-20 6.94522e-24 -1.88428e-20 0.0013952 0.997818 8.59344e-05 0.152563 2.85178 0.0013952 0.99785 0.690898 0.0010474 0.00187976 0.000859344 0.455635 0.00187975 0.436787 0.000128031 1.02 0.887554 0.534716 0.285878 1.71649e-07 3.05898e-09 2389.3 3136.73 -0.0565933 0.482125 0.27759 0.254583 -0.593136 -0.169503 0.493485 -0.268127 -0.225366 1.547 1 0 296.485 0 2.069 1.545 0.00029993 0.862175 0.648363 0.427075 0.406855 2.06924 130.277 83.6792 18.7069 60.75 0.00403526 0 -40 10
0.646 1.87217e-08 2.53889e-06 0.0881383 0.0881347 0.0120415 8.50986e-06 0.00115404 0.110173 0.000657237 0.110825 0.866104 101.861 0.245219 0.727104 4.13863 0.0547811 0.0390437 0.960956 0.0198552 0.00425723 0.0191178 0.00409602 0.00514484 0.00588216 0.205794 0.235286 57.9792 -87.895 126.168 15.9769 145.013 0.000142153 0.267106 192.907 0.310662 0.0673827 0.00409515 0.000561644 0.00138272 0.98699 0.991734 -2.97367e-06 -85.6673 0.0929896 31193.7 300.934 0.98352 0.319147 0.737418 0.737414 9.99958 2.98103e-06 1.1924e-05 0.130787 0.980415 0.930918 -0.0132932 4.89793e-06 0.501444 -1.88505e-20 6.94556e-24 -1.88436e-20 0.0013952 0.997818 8.59345e-05 0.152563 2.85178 0.0013952 0.99785 0.691006 0.00104742 0.00187976 0.000859345 0.455635 0.00187976 0.436796 0.000128034 1.02 0.887555 0.534716 0.285879 1.71649e-07 3.059e-09 2389.28 3136.59 -0.0565841 0.482125 0.27759 0.254575 -0.593138 -0.169503 0.493511 -0.268125 -0.225395 1.548 1 0 296.495 0 2.06917 1.546 0.000299929 0.862115 0.648417 0.426821 0.406885 2.06942 130.286 83.6808 18.707 60.7508 0.0040352 0 -40 10
0.647 1.87506e-08 2.53889e-06 0.0882187 0.0882151 0.0120414 8.52301e-06 0.00115404 0.110273 0.00065724 0.110926 0.86616 101.861 0.245212 0.727186 4.13877 0.0547877 0.039045 0.960955 0.019855 0.00425737 0.0191177 0.00409614 0.00514501 0.00588233 0.205801 0.235293 57.9792 -87.895 126.168 15.9768 145.013 0.000142147 0.267106 192.907 0.310661 0.0673827 0.00409516 0.000561645 0.00138272 0.98699 0.991734 -2.97369e-06 -85.6673 0.0929897 31193.7 300.937 0.98352 0.319147 0.737386 0.737382 9.99958 2.98103e-06 1.1924e-05 0.130788 0.980425 0.930922 -0.0132932 4.89796e-06 0.50145 -1.88513e-20 6.9459e-24 -1.88444e-20 0.0013952 0.997818 8.59345e-05 0.152564 2.85178 0.0013952 0.99785 0.691114 0.00104744 0.00187976 0.000859345 0.455634 0.00187976 0.436805 0.000128038 1.02 0.887556 0.534715 0.285881 1.71649e-07 3.05903e-09 2389.27 3136.45 -0.056575 0.482125 0.27759 0.254566 -0.593139 -0.169503 0.493538 -0.268123 -0.225423 1.549 1 0 296.504 0 2.06935 1.547 0.000299929 0.862055 0.648471 0.426567 0.406914 2.06959 130.296 83.6824 18.7071 60.7516 0.00403513 0 -40 10
0.648 1.87796e-08 2.53889e-06 0.0882991 0.0882955 0.0120414 8.53617e-06 0.00115404 0.110374 0.000657244 0.111026 0.866217 101.861 0.245206 0.727269 4.13892 0.0547942 0.0390464 0.960954 0.0198548 0.00425751 0.0191175 0.00409625 0.00514518 0.00588249 0.205807 0.2353 57.9793 -87.895 126.169 15.9768 145.013 0.000142141 0.267106 192.907 0.310661 0.0673826 0.00409516 0.000561646 0.00138272 0.986989 0.991734 -2.9737e-06 -85.6673 0.0929898 31193.6 300.941 0.98352 0.319147 0.737354 0.73735 9.99958 2.98104e-06 1.1924e-05 0.13079 0.980434 0.930926 -0.0132932 4.89799e-06 0.501455 -1.88521e-20 6.94623e-24 -1.88452e-20 0.0013952 0.997818 8.59346e-05 0.152564 2.85178 0.0013952 0.997849 0.691221 0.00104746 0.00187976 0.000859346 0.455634 0.00187976 0.436814 0.000128041 1.02 0.887557 0.534715 0.285882 1.7165e-07 3.05905e-09 2389.25 3136.31 -0.056566 0.482125 0.277589 0.254557 -0.593141 -0.169503 0.493564 -0.268121 -0.225452 1.55 1 0 296.513 0 2.06952 1.548 0.000299929 0.861996 0.648526 0.426314 0.406943 2.06976 130.305 83.684 18.7072 60.7523 0.00403507 0 -40 10
0.649 1.88085e-08 2.53889e-06 0.0883794 0.0883758 0.0120414 8.54933e-06 0.00115404 0.110474 0.000657247 0.111127 0.866273 101.861 0.245199 0.727352 4.13906 0.0548008 0.0390477 0.960952 0.0198546 0.00425765 0.0191173 0.00409636 0.00514535 0.00588266 0.205814 0.235306 57.9794 -87.895 126.169 15.9767 145.013 0.000142134 0.267106 192.907 0.310661 0.0673826 0.00409516 0.000561646 0.00138272 0.986989 0.991734 -2.97372e-06 -85.6673 0.0929898 31193.6 300.945 0.98352 0.319147 0.737322 0.737318 9.99958 2.98104e-06 1.19241e-05 0.130791 0.980444 0.930931 -0.0132932 4.89801e-06 0.501461 -1.8853e-20 6.94657e-24 -1.8846e-20 0.0013952 0.997818 8.59347e-05 0.152564 2.85178 0.0013952 0.997849 0.691329 0.00104748 0.00187976 0.000859347 0.455634 0.00187976 0.436823 0.000128045 1.02 0.887558 0.534715 0.285884 1.7165e-07 3.05907e-09 2389.23 3136.18 -0.0565569 0.482125 0.277589 0.254549 -0.593143 -0.169503 0.49359 -0.268119 -0.22548 1.551 1 0 296.523 0 2.06969 1.549 0.000299929 0.861936 0.64858 0.426061 0.406972 2.06994 130.314 83.6855 18.7073 60.7531 0.004035 0 -40 10
0.65 1.88375e-08 2.53889e-06 0.0884596 0.0884561 0.0120414 8.56249e-06 0.00115404 0.110575 0.000657251 0.111227 0.866329 101.861 0.245193 0.727435 4.1392 0.0548074 0.0390491 0.960951 0.0198545 0.00425779 0.0191172 0.00409648 0.00514552 0.00588283 0.205821 0.235313 57.9794 -87.895 126.17 15.9767 145.013 0.000142128 0.267106 192.907 0.31066 0.0673825 0.00409517 0.000561647 0.00138273 0.986989 0.991734 -2.97373e-06 -85.6673 0.0929899 31193.6 300.949 0.98352 0.319147 0.737291 0.737286 9.99958 2.98105e-06 1.19241e-05 0.130793 0.980453 0.930935 -0.0132932 4.89804e-06 0.501467 -1.88538e-20 6.94691e-24 -1.88468e-20 0.00139521 0.997818 8.59348e-05 0.152564 2.85178 0.0013952 0.997849 0.691436 0.0010475 0.00187976 0.000859348 0.455634 0.00187976 0.436832 0.000128048 1.02 0.887559 0.534714 0.285885 1.7165e-07 3.05909e-09 2389.22 3136.04 -0.0565479 0.482125 0.277589 0.25454 -0.593144 -0.169503 0.493616 -0.268117 -0.225508 1.552 1 0 296.532 0 2.06987 1.55 0.000299928 0.861877 0.648634 0.425809 0.407001 2.07011 130.324 83.6871 18.7074 60.7538 0.00403494 0 -40 10
0.651 1.88664e-08 2.53889e-06 0.0885398 0.0885362 0.0120414 8.57565e-06 0.00115404 0.110675 0.000657255 0.111327 0.866386 101.861 0.245186 0.727518 4.13934 0.054814 0.0390504 0.96095 0.0198543 0.00425792 0.019117 0.0040966 0.00514569 0.005883 0.205828 0.23532 57.9795 -87.895 126.171 15.9767 145.013 0.000142122 0.267107 192.907 0.31066 0.0673825 0.00409517 0.000561648 0.00138273 0.986989 0.991734 -2.97374e-06 -85.6673 0.09299 31193.6 300.952 0.98352 0.319147 0.737259 0.737255 9.99958 2.98105e-06 1.19241e-05 0.130794 0.980463 0.930939 -0.0132932 4.89807e-06 0.501473 -1.88546e-20 6.94725e-24 -1.88476e-20 0.00139521 0.997818 8.59348e-05 0.152564 2.85178 0.00139521 0.997849 0.691543 0.00104752 0.00187976 0.000859348 0.455633 0.00187976 0.436841 0.000128052 1.02 0.88756 0.534714 0.285886 1.7165e-07 3.05911e-09 2389.2 3135.91 -0.056539 0.482126 0.277588 0.254532 -0.593146 -0.169503 0.493642 -0.268115 -0.225536 1.553 1 0 296.541 0 2.07004 1.551 0.000299928 0.861818 0.648688 0.425558 0.40703 2.07028 130.333 83.6887 18.7075 60.7546 0.00403487 0 -40 10
0.652 1.88954e-08 2.53889e-06 0.0886199 0.0886164 0.0120414 8.58881e-06 0.00115404 0.110775 0.000657258 0.111428 0.866443 101.861 0.245179 0.727601 4.13949 0.0548206 0.0390518 0.960948 0.0198541 0.00425806 0.0191168 0.00409671 0.00514586 0.00588317 0.205835 0.235327 57.9795 -87.895 126.171 15.9766 145.013 0.000142116 0.267107 192.906 0.310659 0.0673824 0.00409517 0.000561648 0.00138273 0.986989 0.991734 -2.97376e-06 -85.6673 0.0929901 31193.6 300.956 0.98352 0.319147 0.737228 0.737223 9.99958 2.98106e-06 1.19241e-05 0.130795 0.980473 0.930943 -0.0132932 4.8981e-06 0.501478 -1.88554e-20 6.94758e-24 -1.88484e-20 0.00139521 0.997818 8.59349e-05 0.152564 2.85178 0.00139521 0.997849 0.691651 0.00104754 0.00187977 0.000859349 0.455633 0.00187976 0.43685 0.000128055 1.02 0.887561 0.534714 0.285888 1.71651e-07 3.05913e-09 2389.18 3135.77 -0.0565301 0.482126 0.277588 0.254523 -0.593147 -0.169503 0.493668 -0.268113 -0.225564 1.554 1 0 296.55 0 2.07021 1.552 0.000299928 0.861759 0.648743 0.425307 0.40706 2.07046 130.342 83.6902 18.7075 60.7553 0.00403481 0 -40 10
0.653 1.89243e-08 2.53889e-06 0.0886999 0.0886964 0.0120414 8.60197e-06 0.00115404 0.110875 0.000657262 0.111528 0.866499 101.86 0.245173 0.727684 4.13963 0.0548272 0.0390531 0.960947 0.019854 0.0042582 0.0191167 0.00409683 0.00514603 0.00588334 0.205841 0.235334 57.9796 -87.895 126.172 15.9766 145.013 0.00014211 0.267107 192.906 0.310659 0.0673824 0.00409517 0.000561649 0.00138273 0.986989 0.991734 -2.97377e-06 -85.6673 0.0929902 31193.5 300.96 0.98352 0.319147 0.737196 0.737192 9.99958 2.98106e-06 1.19241e-05 0.130797 0.980482 0.930948 -0.0132932 4.89813e-06 0.501484 -1.88562e-20 6.94792e-24 -1.88492e-20 0.00139521 0.997818 8.5935e-05 0.152564 2.85178 0.00139521 0.997848 0.691758 0.00104756 0.00187977 0.00085935 0.455633 0.00187977 0.436859 0.000128058 1.02 0.887562 0.534714 0.285889 1.71651e-07 3.05915e-09 2389.17 3135.64 -0.0565212 0.482126 0.277588 0.254515 -0.593149 -0.169503 0.493694 -0.268111 -0.225591 1.555 1 0 296.559 0 2.07039 1.553 0.000299928 0.861701 0.648797 0.425057 0.407089 2.07063 130.351 83.6917 18.7076 60.7561 0.00403474 0 -40 10
0.654 1.89533e-08 2.53889e-06 0.0887799 0.0887764 0.0120413 8.61513e-06 0.00115404 0.110975 0.000657265 0.111628 0.866556 101.86 0.245166 0.727768 4.13978 0.0548339 0.0390545 0.960945 0.0198538 0.00425834 0.0191165 0.00409694 0.00514621 0.00588351 0.205848 0.23534 57.9797 -87.895 126.172 15.9766 145.013 0.000142104 0.267107 192.906 0.310659 0.0673823 0.00409518 0.000561649 0.00138273 0.986989 0.991734 -2.97378e-06 -85.6673 0.0929902 31193.5 300.964 0.98352 0.319147 0.737165 0.737161 9.99958 2.98107e-06 1.19242e-05 0.130798 0.980492 0.930952 -0.0132932 4.89815e-06 0.50149 -1.8857e-20 6.94826e-24 -1.885e-20 0.00139521 0.997818 8.59351e-05 0.152565 2.85179 0.00139521 0.997848 0.691865 0.00104758 0.00187977 0.000859351 0.455633 0.00187977 0.436868 0.000128062 1.02 0.887563 0.534713 0.285891 1.71651e-07 3.05918e-09 2389.15 3135.51 -0.0565124 0.482126 0.277588 0.254507 -0.593151 -0.169503 0.493719 -0.268109 -0.225619 1.556 1 0 296.568 0 2.07056 1.554 0.000299927 0.861643 0.648851 0.424808 0.407118 2.0708 130.361 83.6933 18.7077 60.7568 0.00403468 0 -40 10
0.655 1.89822e-08 2.53889e-06 0.0888598 0.0888563 0.0120413 8.62829e-06 0.00115404 0.111075 0.000657269 0.111727 0.866613 101.86 0.24516 0.727851 4.13992 0.0548405 0.0390559 0.960944 0.0198536 0.00425848 0.0191163 0.00409706 0.00514638 0.00588368 0.205855 0.235347 57.9797 -87.895 126.173 15.9765 145.013 0.000142098 0.267107 192.906 0.310658 0.0673823 0.00409518 0.00056165 0.00138274 0.986989 0.991734 -2.9738e-06 -85.6672 0.0929903 31193.5 300.967 0.98352 0.319147 0.737134 0.73713 9.99958 2.98107e-06 1.19242e-05 0.1308 0.980501 0.930956 -0.0132932 4.89818e-06 0.501496 -1.88578e-20 6.94859e-24 -1.88508e-20 0.00139521 0.997818 8.59351e-05 0.152565 2.85179 0.00139521 0.997848 0.691973 0.0010476 0.00187977 0.000859351 0.455633 0.00187977 0.436877 0.000128065 1.02 0.887564 0.534713 0.285892 1.71651e-07 3.0592e-09 2389.13 3135.37 -0.0565037 0.482126 0.277587 0.254498 -0.593152 -0.169503 0.493745 -0.268107 -0.225646 1.557 1 0 296.577 0 2.07073 1.555 0.000299927 0.861585 0.648905 0.424559 0.407147 2.07097 130.37 83.6948 18.7078 60.7575 0.00403462 0 -40 10
0.656 1.90112e-08 2.53889e-06 0.0889397 0.0889362 0.0120413 8.64144e-06 0.00115404 0.111175 0.000657272 0.111827 0.86667 101.86 0.245153 0.727935 4.14007 0.0548471 0.0390572 0.960943 0.0198534 0.00425862 0.0191162 0.00409718 0.00514655 0.00588385 0.205862 0.235354 57.9798 -87.895 126.173 15.9765 145.013 0.000142092 0.267107 192.906 0.310658 0.0673822 0.00409518 0.000561651 0.00138274 0.986989 0.991734 -2.97381e-06 -85.6672 0.0929904 31193.5 300.971 0.98352 0.319147 0.737103 0.737099 9.99958 2.98108e-06 1.19242e-05 0.130801 0.980511 0.93096 -0.0132932 4.89821e-06 0.501502 -1.88586e-20 6.94893e-24 -1.88516e-20 0.00139521 0.997818 8.59352e-05 0.152565 2.85179 0.00139521 0.997848 0.69208 0.00104762 0.00187977 0.000859352 0.455632 0.00187977 0.436886 0.000128069 1.02 0.887565 0.534713 0.285894 1.71652e-07 3.05922e-09 2389.12 3135.24 -0.0564949 0.482126 0.277587 0.25449 -0.593154 -0.169504 0.49377 -0.268105 -0.225674 1.558 1 0 296.586 0 2.0709 1.556 0.000299927 0.861527 0.648959 0.424311 0.407176 2.07115 130.379 83.6963 18.7079 60.7583 0.00403455 0 -40 10
0.657 1.90401e-08 2.53889e-06 0.0890195 0.089016 0.0120413 8.6546e-06 0.00115404 0.111274 0.000657276 0.111927 0.866727 101.86 0.245146 0.728018 4.14021 0.0548538 0.0390586 0.960941 0.0198533 0.00425876 0.019116 0.00409729 0.00514672 0.00588402 0.205869 0.235361 57.9799 -87.895 126.174 15.9764 145.013 0.000142086 0.267108 192.906 0.310657 0.0673822 0.00409519 0.000561651 0.00138274 0.986989 0.991734 -2.97383e-06 -85.6672 0.0929905 31193.5 300.975 0.98352 0.319147 0.737073 0.737068 9.99958 2.98108e-06 1.19242e-05 0.130803 0.98052 0.930964 -0.0132932 4.89824e-06 0.501508 -1.88594e-20 6.94927e-24 -1.88524e-20 0.00139521 0.997818 8.59353e-05 0.152565 2.85179 0.00139521 0.997848 0.692187 0.00104764 0.00187977 0.000859353 0.455632 0.00187977 0.436895 0.000128072 1.02 0.887566 0.534712 0.285895 1.71652e-07 3.05924e-09 2389.1 3135.11 -0.0564862 0.482126 0.277587 0.254482 -0.593155 -0.169504 0.493795 -0.268103 -0.225701 1.559 1 0 296.595 0 2.07108 1.557 0.000299926 0.86147 0.649013 0.424063 0.407205 2.07132 130.388 83.6978 18.708 60.759 0.00403449 0 -40 10
0.658 1.90691e-08 2.53889e-06 0.0890992 0.0890957 0.0120413 8.66776e-06 0.00115404 0.111374 0.000657279 0.112027 0.866783 101.86 0.24514 0.728102 4.14036 0.0548604 0.03906 0.96094 0.0198531 0.0042589 0.0191158 0.00409741 0.0051469 0.00588419 0.205876 0.235368 57.9799 -87.895 126.174 15.9764 145.014 0.00014208 0.267108 192.905 0.310657 0.0673821 0.00409519 0.000561652 0.00138274 0.986989 0.991734 -2.97384e-06 -85.6672 0.0929906 31193.4 300.979 0.98352 0.319147 0.737042 0.737038 9.99958 2.98108e-06 1.19242e-05 0.130804 0.980529 0.930968 -0.0132932 4.89827e-06 0.501513 -1.88602e-20 6.94961e-24 -1.88533e-20 0.00139521 0.997818 8.59354e-05 0.152565 2.85179 0.00139521 0.997847 0.692294 0.00104766 0.00187977 0.000859354 0.455632 0.00187977 0.436904 0.000128076 1.02 0.887567 0.534712 0.285896 1.71652e-07 3.05926e-09 2389.08 3134.98 -0.0564776 0.482126 0.277586 0.254474 -0.593157 -0.169504 0.49382 -0.268101 -0.225728 1.56 1 0 296.604 0 2.07125 1.558 0.000299926 0.861413 0.649067 0.423816 0.407234 2.07149 130.398 83.6993 18.7081 60.7597 0.00403443 0 -40 10
0.659 1.9098e-08 2.53889e-06 0.0891789 0.0891754 0.0120413 8.68092e-06 0.00115404 0.111474 0.000657283 0.112126 0.86684 101.859 0.245133 0.728186 4.14051 0.0548671 0.0390614 0.960939 0.0198529 0.00425905 0.0191156 0.00409753 0.00514707 0.00588436 0.205883 0.235375 57.98 -87.895 126.175 15.9764 145.014 0.000142075 0.267108 192.905 0.310657 0.0673821 0.00409519 0.000561652 0.00138274 0.986989 0.991734 -2.97385e-06 -85.6672 0.0929906 31193.4 300.983 0.98352 0.319147 0.737012 0.737007 9.99958 2.98109e-06 1.19242e-05 0.130806 0.980539 0.930973 -0.0132932 4.89829e-06 0.501519 -1.8861e-20 6.94995e-24 -1.88541e-20 0.00139521 0.997818 8.59354e-05 0.152565 2.85179 0.00139521 0.997847 0.692401 0.00104768 0.00187977 0.000859354 0.455632 0.00187977 0.436912 0.000128079 1.02 0.887568 0.534712 0.285898 1.71652e-07 3.05928e-09 2389.07 3134.85 -0.056469 0.482126 0.277586 0.254465 -0.593158 -0.169504 0.493845 -0.268099 -0.225755 1.561 1 0 296.613 0 2.07142 1.559 0.000299926 0.861356 0.649121 0.42357 0.407263 2.07166 130.407 83.7008 18.7082 60.7605 0.00403437 0 -40 10
0.66 1.9127e-08 2.53889e-06 0.0892585 0.089255 0.0120413 8.69408e-06 0.00115404 0.111573 0.000657286 0.112226 0.866898 101.859 0.245126 0.72827 4.14065 0.0548738 0.0390628 0.960937 0.0198528 0.00425919 0.0191155 0.00409764 0.00514724 0.00588454 0.20589 0.235381 57.9801 -87.895 126.176 15.9763 145.014 0.000142069 0.267108 192.905 0.310656 0.067382 0.00409519 0.000561653 0.00138275 0.986989 0.991734 -2.97387e-06 -85.6672 0.0929907 31193.4 300.987 0.98352 0.319147 0.736981 0.736977 9.99958 2.98109e-06 1.19243e-05 0.130807 0.980548 0.930977 -0.0132932 4.89832e-06 0.501525 -1.88618e-20 6.95028e-24 -1.88549e-20 0.00139522 0.997818 8.59355e-05 0.152565 2.85179 0.00139522 0.997847 0.692508 0.0010477 0.00187978 0.000859355 0.455632 0.00187978 0.436921 0.000128082 1.02 0.887569 0.534712 0.285899 1.71653e-07 3.05931e-09 2389.05 3134.72 -0.0564604 0.482126 0.277586 0.254457 -0.59316 -0.169504 0.49387 -0.268097 -0.225782 1.562 1 0 296.621 0 2.0716 1.56 0.000299926 0.861299 0.649175 0.423324 0.407292 2.07184 130.416 83.7023 18.7082 60.7612 0.00403431 0 -40 10
0.661 1.91559e-08 2.53889e-06 0.089338 0.0893345 0.0120413 8.70724e-06 0.00115404 0.111673 0.00065729 0.112325 0.866955 101.859 0.24512 0.728354 4.1408 0.0548804 0.0390642 0.960936 0.0198526 0.00425933 0.0191153 0.00409776 0.00514742 0.00588471 0.205897 0.235388 57.9801 -87.895 126.176 15.9763 145.014 0.000142063 0.267108 192.905 0.310656 0.067382 0.0040952 0.000561654 0.00138275 0.986989 0.991734 -2.97388e-06 -85.6672 0.0929908 31193.4 300.99 0.983519 0.319147 0.736951 0.736947 9.99958 2.9811e-06 1.19243e-05 0.130808 0.980557 0.930981 -0.0132932 4.89835e-06 0.501531 -1.88626e-20 6.95062e-24 -1.88557e-20 0.00139522 0.997818 8.59356e-05 0.152566 2.85179 0.00139522 0.997847 0.692616 0.00104772 0.00187978 0.000859356 0.455631 0.00187978 0.43693 0.000128086 1.02 0.88757 0.534711 0.285901 1.71653e-07 3.05933e-09 2389.03 3134.59 -0.0564519 0.482126 0.277586 0.254449 -0.593161 -0.169504 0.493894 -0.268095 -0.225808 1.563 1 0 296.63 0 2.07177 1.561 0.000299925 0.861243 0.649229 0.423079 0.407321 2.07201 130.425 83.7038 18.7083 60.7619 0.00403424 0 -40 10
0.662 1.91849e-08 2.53889e-06 0.0894175 0.089414 0.0120412 8.7204e-06 0.00115404 0.111772 0.000657293 0.112425 0.867012 101.859 0.245113 0.728438 4.14095 0.0548871 0.0390655 0.960934 0.0198524 0.00425947 0.0191151 0.00409788 0.00514759 0.00588488 0.205904 0.235395 57.9802 -87.895 126.177 15.9762 145.014 0.000142057 0.267108 192.905 0.310655 0.0673819 0.0040952 0.000561654 0.00138275 0.986989 0.991734 -2.9739e-06 -85.6672 0.0929909 31193.4 300.994 0.983519 0.319147 0.736921 0.736917 9.99958 2.9811e-06 1.19243e-05 0.13081 0.980567 0.930985 -0.0132932 4.89838e-06 0.501537 -1.88634e-20 6.95096e-24 -1.88565e-20 0.00139522 0.997818 8.59356e-05 0.152566 2.85179 0.00139522 0.997847 0.692723 0.00104774 0.00187978 0.000859356 0.455631 0.00187978 0.436939 0.000128089 1.02 0.887571 0.534711 0.285902 1.71653e-07 3.05935e-09 2389.02 3134.46 -0.0564435 0.482126 0.277585 0.254441 -0.593163 -0.169504 0.493919 -0.268093 -0.225835 1.564 1 0 296.639 0 2.07194 1.562 0.000299925 0.861187 0.649283 0.422834 0.40735 2.07218 130.435 83.7053 18.7084 60.7626 0.00403418 0 -40 10
0.663 1.92138e-08 2.53889e-06 0.0894969 0.0894934 0.0120412 8.73355e-06 0.00115404 0.111871 0.000657297 0.112524 0.867069 101.859 0.245106 0.728522 4.1411 0.0548938 0.0390669 0.960933 0.0198522 0.00425961 0.0191149 0.004098 0.00514777 0.00588506 0.205911 0.235402 57.9802 -87.895 126.177 15.9762 145.014 0.000142051 0.267109 192.905 0.310655 0.0673819 0.0040952 0.000561655 0.00138275 0.986989 0.991734 -2.97391e-06 -85.6672 0.092991 31193.3 300.998 0.983519 0.319147 0.736891 0.736887 9.99958 2.98111e-06 1.19243e-05 0.130811 0.980576 0.930989 -0.0132932 4.89841e-06 0.501543 -1.88642e-20 6.9513e-24 -1.88573e-20 0.00139522 0.997818 8.59357e-05 0.152566 2.85179 0.00139522 0.997847 0.692829 0.00104776 0.00187978 0.000859357 0.455631 0.00187978 0.436948 0.000128093 1.02 0.887573 0.534711 0.285904 1.71653e-07 3.05937e-09 2389 3134.33 -0.056435 0.482126 0.277585 0.254433 -0.593164 -0.169504 0.493943 -0.268091 -0.225861 1.565 1 0 296.648 0 2.07211 1.563 0.000299925 0.861131 0.649337 0.42259 0.407379 2.07235 130.444 83.7068 18.7085 60.7633 0.00403412 0 -40 10
0.664 1.92428e-08 2.53889e-06 0.0895762 0.0895728 0.0120412 8.74671e-06 0.00115404 0.11197 0.0006573 0.112623 0.867126 101.859 0.245099 0.728606 4.14124 0.0549005 0.0390683 0.960932 0.0198521 0.00425976 0.0191148 0.00409812 0.00514794 0.00588523 0.205918 0.235409 57.9803 -87.895 126.178 15.9762 145.014 0.000142046 0.267109 192.905 0.310655 0.0673818 0.00409521 0.000561656 0.00138275 0.986989 0.991734 -2.97392e-06 -85.6672 0.092991 31193.3 301.002 0.983519 0.319147 0.736861 0.736857 9.99958 2.98111e-06 1.19243e-05 0.130813 0.980585 0.930993 -0.0132932 4.89843e-06 0.501549 -1.8865e-20 6.95164e-24 -1.88581e-20 0.00139522 0.997818 8.59358e-05 0.152566 2.85179 0.00139522 0.997846 0.692936 0.00104778 0.00187978 0.000859358 0.455631 0.00187978 0.436957 0.000128096 1.02 0.887574 0.53471 0.285905 1.71654e-07 3.05939e-09 2388.98 3134.21 -0.0564266 0.482126 0.277585 0.254425 -0.593166 -0.169504 0.493967 -0.268089 -0.225888 1.566 1 0 296.656 0 2.07228 1.564 0.000299924 0.861075 0.649391 0.422347 0.407408 2.07252 130.453 83.7083 18.7086 60.764 0.00403406 0 -40 10
0.665 1.92717e-08 2.53889e-06 0.0896555 0.0896521 0.0120412 8.75987e-06 0.00115404 0.112069 0.000657304 0.112722 0.867184 101.859 0.245093 0.728691 4.14139 0.0549072 0.0390697 0.96093 0.0198519 0.0042599 0.0191146 0.00409824 0.00514812 0.0058854 0.205925 0.235416 57.9804 -87.8951 126.178 15.9761 145.014 0.00014204 0.267109 192.904 0.310654 0.0673818 0.00409521 0.000561656 0.00138276 0.986989 0.991734 -2.97394e-06 -85.6672 0.0929911 31193.3 301.006 0.983519 0.319147 0.736832 0.736827 9.99958 2.98112e-06 1.19244e-05 0.130814 0.980594 0.930997 -0.0132932 4.89846e-06 0.501555 -1.88659e-20 6.95197e-24 -1.88589e-20 0.00139522 0.997818 8.59359e-05 0.152566 2.85179 0.00139522 0.997846 0.693043 0.00104779 0.00187978 0.000859359 0.455631 0.00187978 0.436966 0.0001281 1.02 0.887575 0.53471 0.285907 1.71654e-07 3.05941e-09 2388.97 3134.08 -0.0564183 0.482127 0.277584 0.254417 -0.593167 -0.169504 0.493991 -0.268086 -0.225914 1.567 1 0 296.665 0 2.07246 1.565 0.000299924 0.86102 0.649445 0.422104 0.407437 2.0727 130.462 83.7097 18.7087 60.7647 0.004034 0 -40 10
0.666 1.93007e-08 2.53889e-06 0.0897347 0.0897313 0.0120412 8.77303e-06 0.00115404 0.112168 0.000657307 0.112821 0.867241 101.858 0.245086 0.728775 4.14154 0.0549139 0.0390711 0.960929 0.0198517 0.00426004 0.0191144 0.00409836 0.0051483 0.00588558 0.205932 0.235423 57.9804 -87.8951 126.179 15.9761 145.014 0.000142034 0.267109 192.904 0.310654 0.0673817 0.00409521 0.000561657 0.00138276 0.986989 0.991734 -2.97395e-06 -85.6671 0.0929912 31193.3 301.01 0.983519 0.319147 0.736802 0.736798 9.99958 2.98112e-06 1.19244e-05 0.130816 0.980603 0.931001 -0.0132932 4.89849e-06 0.501561 -1.88667e-20 6.95231e-24 -1.88597e-20 0.00139522 0.997818 8.59359e-05 0.152566 2.8518 0.00139522 0.997846 0.69315 0.00104781 0.00187978 0.000859359 0.45563 0.00187978 0.436975 0.000128103 1.02 0.887576 0.53471 0.285908 1.71654e-07 3.05943e-09 2388.95 3133.95 -0.05641 0.482127 0.277584 0.254409 -0.593169 -0.169504 0.494015 -0.268084 -0.22594 1.568 1 0 296.673 0 2.07263 1.566 0.000299924 0.860965 0.649499 0.421862 0.407466 2.07287 130.471 83.7112 18.7088 60.7654 0.00403394 0 -40 10
0.667 1.93296e-08 2.53889e-06 0.0898139 0.0898104 0.0120412 8.78619e-06 0.00115404 0.112267 0.00065731 0.11292 0.867298 101.858 0.245079 0.72886 4.14169 0.0549206 0.0390726 0.960927 0.0198515 0.00426019 0.0191142 0.00409848 0.00514847 0.00588575 0.205939 0.23543 57.9805 -87.8951 126.179 15.9761 145.014 0.000142028 0.267109 192.904 0.310653 0.0673817 0.00409521 0.000561657 0.00138276 0.986989 0.991734 -2.97397e-06 -85.6671 0.0929913 31193.2 301.014 0.983519 0.319147 0.736773 0.736768 9.99958 2.98113e-06 1.19244e-05 0.130817 0.980613 0.931005 -0.0132932 4.89852e-06 0.501567 -1.88675e-20 6.95265e-24 -1.88605e-20 0.00139522 0.997818 8.5936e-05 0.152566 2.8518 0.00139522 0.997846 0.693257 0.00104783 0.00187979 0.00085936 0.45563 0.00187978 0.436984 0.000128106 1.02 0.887577 0.53471 0.285909 1.71654e-07 3.05946e-09 2388.93 3133.83 -0.0564017 0.482127 0.277584 0.254401 -0.59317 -0.169504 0.494039 -0.268082 -0.225966 1.569 1 0 296.682 0 2.0728 1.567 0.000299924 0.86091 0.649553 0.421621 0.407495 2.07304 130.481 83.7126 18.7088 60.7661 0.00403388 0 -40 10
0.668 1.93586e-08 2.5389e-06 0.0898929 0.0898895 0.0120412 8.79934e-06 0.00115404 0.112366 0.000657314 0.113019 0.867356 101.858 0.245073 0.728944 4.14184 0.0549274 0.039074 0.960926 0.0198513 0.00426033 0.0191141 0.0040986 0.00514865 0.00588593 0.205946 0.235437 57.9806 -87.8951 126.18 15.976 145.014 0.000142023 0.26711 192.904 0.310653 0.0673816 0.00409522 0.000561658 0.00138276 0.986989 0.991734 -2.97398e-06 -85.6671 0.0929914 31193.2 301.018 0.983519 0.319147 0.736743 0.736739 9.99958 2.98113e-06 1.19244e-05 0.130819 0.980622 0.931009 -0.0132932 4.89855e-06 0.501573 -1.88683e-20 6.95299e-24 -1.88613e-20 0.00139522 0.997818 8.59361e-05 0.152566 2.8518 0.00139522 0.997846 0.693364 0.00104785 0.00187979 0.000859361 0.45563 0.00187979 0.436993 0.00012811 1.02 0.887578 0.534709 0.285911 1.71655e-07 3.05948e-09 2388.92 3133.7 -0.0563935 0.482127 0.277584 0.254393 -0.593172 -0.169504 0.494063 -0.26808 -0.225991 1.57 1 0 296.69 0 2.07297 1.568 0.000299923 0.860856 0.649606 0.42138 0.407523 2.07321 130.49 83.7141 18.7089 60.7668 0.00403382 0 -40 10
0.669 1.93875e-08 2.5389e-06 0.089972 0.0899686 0.0120411 8.8125e-06 0.00115404 0.112465 0.000657317 0.113118 0.867413 101.858 0.245066 0.729029 4.14199 0.0549341 0.0390754 0.960925 0.0198512 0.00426048 0.0191139 0.00409872 0.00514883 0.00588611 0.205953 0.235444 57.9806 -87.8951 126.18 15.976 145.014 0.000142017 0.26711 192.904 0.310653 0.0673816 0.00409522 0.000561659 0.00138276 0.986989 0.991734 -2.97399e-06 -85.6671 0.0929914 31193.2 301.021 0.983519 0.319147 0.736714 0.73671 9.99958 2.98114e-06 1.19244e-05 0.13082 0.980631 0.931013 -0.0132932 4.89858e-06 0.501579 -1.88691e-20 6.95333e-24 -1.88621e-20 0.00139523 0.997818 8.59362e-05 0.152567 2.8518 0.00139523 0.997845 0.69347 0.00104787 0.00187979 0.000859362 0.45563 0.00187979 0.437001 0.000128113 1.02 0.887579 0.534709 0.285912 1.71655e-07 3.0595e-09 2388.9 3133.58 -0.0563853 0.482127 0.277583 0.254385 -0.593173 -0.169504 0.494087 -0.268078 -0.226017 1.571 1 0 296.699 0 2.07314 1.569 0.000299923 0.860801 0.64966 0.421139 0.407552 2.07338 130.499 83.7155 18.709 60.7675 0.00403376 0 -40 10
0.67 1.94165e-08 2.5389e-06 0.0900509 0.0900475 0.0120411 8.82566e-06 0.00115404 0.112564 0.000657321 0.113216 0.867471 101.858 0.245059 0.729114 4.14214 0.0549408 0.0390768 0.960923 0.019851 0.00426062 0.0191137 0.00409884 0.00514901 0.00588628 0.20596 0.235451 57.9807 -87.8951 126.181 15.9759 145.014 0.000142012 0.26711 192.904 0.310652 0.0673815 0.00409522 0.000561659 0.00138277 0.986989 0.991734 -2.97401e-06 -85.6671 0.0929915 31193.2 301.025 0.983519 0.319147 0.736685 0.736681 9.99958 2.98114e-06 1.19245e-05 0.130822 0.98064 0.931017 -0.0132932 4.8986e-06 0.501585 -1.88699e-20 6.95367e-24 -1.88629e-20 0.00139523 0.997818 8.59362e-05 0.152567 2.8518 0.00139523 0.997845 0.693577 0.00104789 0.00187979 0.000859362 0.45563 0.00187979 0.43701 0.000128117 1.02 0.88758 0.534709 0.285914 1.71655e-07 3.05952e-09 2388.88 3133.45 -0.0563772 0.482127 0.277583 0.254378 -0.593175 -0.169504 0.49411 -0.268076 -0.226043 1.572 1 0 296.707 0 2.07331 1.57 0.000299923 0.860747 0.649714 0.4209 0.407581 2.07355 130.508 83.7169 18.7091 60.7682 0.0040337 0 -40 10
0.671 1.94454e-08 2.5389e-06 0.0901298 0.0901264 0.0120411 8.83882e-06 0.00115404 0.112662 0.000657324 0.113315 0.867529 101.858 0.245052 0.729199 4.14229 0.0549476 0.0390782 0.960922 0.0198508 0.00426076 0.0191135 0.00409896 0.00514918 0.00588646 0.205967 0.235458 57.9807 -87.8951 126.181 15.9759 145.014 0.000142006 0.26711 192.904 0.310652 0.0673815 0.00409522 0.00056166 0.00138277 0.986989 0.991734 -2.97402e-06 -85.6671 0.0929916 31193.2 301.029 0.983519 0.319147 0.736656 0.736652 9.99958 2.98114e-06 1.19245e-05 0.130823 0.980649 0.931021 -0.0132931 4.89863e-06 0.501591 -1.88707e-20 6.95401e-24 -1.88638e-20 0.00139523 0.997818 8.59363e-05 0.152567 2.8518 0.00139523 0.997845 0.693684 0.00104791 0.00187979 0.000859363 0.455629 0.00187979 0.437019 0.00012812 1.02 0.887581 0.534708 0.285915 1.71655e-07 3.05954e-09 2388.87 3133.33 -0.0563691 0.482127 0.277583 0.25437 -0.593176 -0.169504 0.494134 -0.268074 -0.226068 1.573 1 0 296.715 0 2.07349 1.571 0.000299922 0.860693 0.649768 0.420661 0.40761 2.07373 130.517 83.7184 18.7092 60.7689 0.00403364 0 -40 10
0.672 1.94743e-08 2.5389e-06 0.0902087 0.0902053 0.0120411 8.85198e-06 0.00115404 0.112761 0.000657327 0.113414 0.867586 101.858 0.245046 0.729284 4.14244 0.0549543 0.0390797 0.96092 0.0198506 0.00426091 0.0191134 0.00409908 0.00514936 0.00588664 0.205975 0.235465 57.9808 -87.8951 126.182 15.9759 145.014 0.000142 0.26711 192.903 0.310651 0.0673814 0.00409523 0.000561661 0.00138277 0.986989 0.991734 -2.97404e-06 -85.6671 0.0929917 31193.1 301.033 0.983519 0.319147 0.736627 0.736623 9.99958 2.98115e-06 1.19245e-05 0.130825 0.980658 0.931025 -0.0132931 4.89866e-06 0.501597 -1.88715e-20 6.95435e-24 -1.88646e-20 0.00139523 0.997818 8.59364e-05 0.152567 2.8518 0.00139523 0.997845 0.69379 0.00104793 0.00187979 0.000859364 0.455629 0.00187979 0.437028 0.000128123 1.02 0.887582 0.534708 0.285917 1.71656e-07 3.05956e-09 2388.85 3133.21 -0.056361 0.482127 0.277582 0.254362 -0.593177 -0.169505 0.494157 -0.268072 -0.226093 1.574 1 0 296.724 0 2.07366 1.572 0.000299922 0.86064 0.649821 0.420422 0.407639 2.0739 130.527 83.7198 18.7093 60.7696 0.00403358 0 -40 10
0.673 1.95033e-08 2.5389e-06 0.0902874 0.0902841 0.0120411 8.86514e-06 0.00115404 0.112859 0.000657331 0.113512 0.867644 101.857 0.245039 0.729369 4.1426 0.0549611 0.0390811 0.960919 0.0198505 0.00426106 0.0191132 0.0040992 0.00514954 0.00588681 0.205982 0.235473 57.9809 -87.8951 126.182 15.9758 145.014 0.000141995 0.26711 192.903 0.310651 0.0673814 0.00409523 0.000561661 0.00138277 0.986989 0.991734 -2.97405e-06 -85.6671 0.0929918 31193.1 301.037 0.983519 0.319147 0.736599 0.736594 9.99958 2.98115e-06 1.19245e-05 0.130826 0.980667 0.931029 -0.0132931 4.89869e-06 0.501603 -1.88723e-20 6.95468e-24 -1.88654e-20 0.00139523 0.997818 8.59365e-05 0.152567 2.8518 0.00139523 0.997845 0.693897 0.00104795 0.00187979 0.000859365 0.455629 0.00187979 0.437037 0.000128127 1.02 0.887583 0.534708 0.285918 1.71656e-07 3.05959e-09 2388.83 3133.08 -0.056353 0.482127 0.277582 0.254354 -0.593179 -0.169505 0.49418 -0.26807 -0.226118 1.575 1 0 296.732 0 2.07383 1.573 0.000299922 0.860586 0.649875 0.420184 0.407668 2.07407 130.536 83.7212 18.7093 60.7703 0.00403353 0 -40 10
0.674 1.95322e-08 2.5389e-06 0.0903661 0.0903628 0.0120411 8.87829e-06 0.00115404 0.112958 0.000657334 0.11361 0.867702 101.857 0.245032 0.729454 4.14275 0.0549679 0.0390825 0.960917 0.0198503 0.0042612 0.019113 0.00409932 0.00514972 0.00588699 0.205989 0.23548 57.9809 -87.8951 126.183 15.9758 145.014 0.000141989 0.267111 192.903 0.310651 0.0673814 0.00409523 0.000561662 0.00138277 0.986989 0.991734 -2.97406e-06 -85.6671 0.0929918 31193.1 301.041 0.983519 0.319147 0.73657 0.736566 9.99958 2.98116e-06 1.19245e-05 0.130828 0.980676 0.931032 -0.0132931 4.89872e-06 0.501609 -1.88731e-20 6.95502e-24 -1.88662e-20 0.00139523 0.997818 8.59365e-05 0.152567 2.8518 0.00139523 0.997845 0.694004 0.00104797 0.0018798 0.000859365 0.455629 0.00187979 0.437046 0.00012813 1.02 0.887584 0.534707 0.28592 1.71656e-07 3.05961e-09 2388.82 3132.96 -0.0563451 0.482127 0.277582 0.254347 -0.59318 -0.169505 0.494203 -0.268068 -0.226144 1.576 1 0 296.74 0 2.074 1.574 0.000299921 0.860533 0.649928 0.419947 0.407696 2.07424 130.545 83.7226 18.7094 60.7709 0.00403347 0 -40 10
0.675 1.95612e-08 2.5389e-06 0.0904448 0.0904414 0.0120411 8.89145e-06 0.00115404 0.113056 0.000657337 0.113709 0.86776 101.857 0.245025 0.729539 4.1429 0.0549747 0.039084 0.960916 0.0198501 0.00426135 0.0191128 0.00409944 0.0051499 0.00588717 0.205996 0.235487 57.981 -87.8951 126.184 15.9758 145.014 0.000141984 0.267111 192.903 0.31065 0.0673813 0.00409524 0.000561662 0.00138278 0.986989 0.991734 -2.97408e-06 -85.6671 0.0929919 31193.1 301.045 0.983519 0.319147 0.736542 0.736537 9.99958 2.98116e-06 1.19245e-05 0.130829 0.980684 0.931036 -0.0132931 4.89874e-06 0.501615 -1.88739e-20 6.95536e-24 -1.8867e-20 0.00139523 0.997818 8.59366e-05 0.152567 2.8518 0.00139523 0.997844 0.69411 0.00104799 0.0018798 0.000859366 0.455628 0.0018798 0.437055 0.000128134 1.02 0.887585 0.534707 0.285921 1.71656e-07 3.05963e-09 2388.8 3132.84 -0.0563371 0.482127 0.277582 0.254339 -0.593182 -0.169505 0.494226 -0.268066 -0.226168 1.577 1 0 296.748 0 2.07417 1.575 0.000299921 0.860481 0.649982 0.41971 0.407725 2.07441 130.554 83.724 18.7095 60.7716 0.00403341 0 -40 10
0.676 1.95901e-08 2.5389e-06 0.0905234 0.09052 0.0120411 8.90461e-06 0.00115404 0.113154 0.000657341 0.113807 0.867818 101.857 0.245019 0.729624 4.14305 0.0549814 0.0390854 0.960915 0.0198499 0.00426149 0.0191127 0.00409957 0.00515008 0.00588735 0.206003 0.235494 57.9811 -87.8951 126.184 15.9757 145.014 0.000141978 0.267111 192.903 0.31065 0.0673813 0.00409524 0.000561663 0.00138278 0.986989 0.991734 -2.97409e-06 -85.6671 0.092992 31193.1 301.049 0.983519 0.319147 0.736513 0.736509 9.99958 2.98117e-06 1.19246e-05 0.130831 0.980693 0.93104 -0.0132931 4.89877e-06 0.501622 -1.88748e-20 6.9557e-24 -1.88678e-20 0.00139523 0.997818 8.59367e-05 0.152568 2.8518 0.00139523 0.997844 0.694217 0.00104801 0.0018798 0.000859367 0.455628 0.0018798 0.437063 0.000128137 1.02 0.887586 0.534707 0.285922 1.71657e-07 3.05965e-09 2388.78 3132.72 -0.0563292 0.482127 0.277581 0.254331 -0.593183 -0.169505 0.494249 -0.268064 -0.226193 1.578 1 0 296.756 0 2.07434 1.576 0.000299921 0.860428 0.650036 0.419474 0.407754 2.07458 130.563 83.7254 18.7096 60.7723 0.00403335 0 -40 10
0.677 1.96191e-08 2.5389e-06 0.0906019 0.0905986 0.012041 8.91777e-06 0.00115404 0.113252 0.000657344 0.113905 0.867876 101.857 0.245012 0.72971 4.14321 0.0549882 0.0390868 0.960913 0.0198497 0.00426164 0.0191125 0.00409969 0.00515026 0.00588753 0.20601 0.235501 57.9811 -87.8951 126.185 15.9757 145.014 0.000141973 0.267111 192.903 0.310649 0.0673812 0.00409524 0.000561664 0.00138278 0.986989 0.991734 -2.97411e-06 -85.6671 0.0929921 31193 301.053 0.983519 0.319147 0.736485 0.736481 9.99958 2.98117e-06 1.19246e-05 0.130832 0.980702 0.931044 -0.0132931 4.8988e-06 0.501628 -1.88756e-20 6.95604e-24 -1.88686e-20 0.00139523 0.997818 8.59368e-05 0.152568 2.85181 0.00139523 0.997844 0.694323 0.00104803 0.0018798 0.000859368 0.455628 0.0018798 0.437072 0.00012814 1.02 0.887587 0.534707 0.285924 1.71657e-07 3.05967e-09 2388.77 3132.6 -0.0563214 0.482127 0.277581 0.254324 -0.593184 -0.169505 0.494271 -0.268062 -0.226218 1.579 1 0 296.765 0 2.07451 1.577 0.000299921 0.860376 0.650089 0.419238 0.407783 2.07475 130.572 83.7268 18.7097 60.773 0.0040333 0 -40 10
0.678 1.9648e-08 2.5389e-06 0.0906803 0.090677 0.012041 8.93092e-06 0.00115404 0.11335 0.000657347 0.114003 0.867934 101.857 0.245005 0.729795 4.14336 0.054995 0.0390883 0.960912 0.0198496 0.00426179 0.0191123 0.00409981 0.00515044 0.00588771 0.206018 0.235508 57.9812 -87.8951 126.185 15.9756 145.014 0.000141968 0.267111 192.902 0.310649 0.0673812 0.00409524 0.000561664 0.00138278 0.986989 0.991734 -2.97412e-06 -85.667 0.0929922 31193 301.057 0.983519 0.319147 0.736457 0.736453 9.99958 2.98118e-06 1.19246e-05 0.130834 0.980711 0.931048 -0.0132931 4.89883e-06 0.501634 -1.88764e-20 6.95638e-24 -1.88694e-20 0.00139523 0.997818 8.59368e-05 0.152568 2.85181 0.00139523 0.997844 0.694429 0.00104805 0.0018798 0.000859368 0.455628 0.0018798 0.437081 0.000128144 1.02 0.887588 0.534706 0.285925 1.71657e-07 3.05969e-09 2388.75 3132.48 -0.0563136 0.482127 0.277581 0.254316 -0.593186 -0.169505 0.494294 -0.26806 -0.226243 1.58 1 0 296.773 0 2.07468 1.578 0.00029992 0.860323 0.650143 0.419003 0.407811 2.07492 130.581 83.7282 18.7097 60.7736 0.00403324 0 -40 10
0.679 1.9677e-08 2.5389e-06 0.0907587 0.0907554 0.012041 8.94408e-06 0.00115405 0.113448 0.000657351 0.114101 0.867992 101.856 0.244998 0.729881 4.14351 0.0550018 0.0390897 0.96091 0.0198494 0.00426194 0.0191121 0.00409993 0.00515062 0.00588789 0.206025 0.235515 57.9813 -87.8951 126.186 15.9756 145.014 0.000141962 0.267112 192.902 0.310649 0.0673811 0.00409525 0.000561665 0.00138278 0.986989 0.991733 -2.97413e-06 -85.667 0.0929923 31193 301.061 0.983519 0.319147 0.736429 0.736425 9.99958 2.98118e-06 1.19246e-05 0.130835 0.98072 0.931052 -0.0132931 4.89886e-06 0.50164 -1.88772e-20 6.95672e-24 -1.88702e-20 0.00139524 0.997818 8.59369e-05 0.152568 2.85181 0.00139524 0.997844 0.694536 0.00104807 0.0018798 0.000859369 0.455628 0.0018798 0.43709 0.000128147 1.02 0.887589 0.534706 0.285927 1.71657e-07 3.05972e-09 2388.73 3132.36 -0.0563058 0.482127 0.27758 0.254309 -0.593187 -0.169505 0.494316 -0.268058 -0.226267 1.581 1 0 296.781 0 2.07486 1.579 0.00029992 0.860272 0.650196 0.418768 0.40784 2.07509 130.591 83.7296 18.7098 60.7743 0.00403318 0 -40 10
0.68 1.97059e-08 2.5389e-06 0.0908371 0.0908338 0.012041 8.95724e-06 0.00115405 0.113546 0.000657354 0.114199 0.86805 101.856 0.244991 0.729967 4.14367 0.0550086 0.0390912 0.960909 0.0198492 0.00426208 0.0191119 0.00410006 0.00515081 0.00588807 0.206032 0.235523 57.9813 -87.8951 126.186 15.9756 145.014 0.000141957 0.267112 192.902 0.310648 0.0673811 0.00409525 0.000561666 0.00138279 0.986989 0.991733 -2.97415e-06 -85.667 0.0929923 31193 301.065 0.983519 0.319147 0.736401 0.736397 9.99958 2.98119e-06 1.19246e-05 0.130837 0.980729 0.931055 -0.0132931 4.89889e-06 0.501646 -1.8878e-20 6.95706e-24 -1.8871e-20 0.00139524 0.997818 8.5937e-05 0.152568 2.85181 0.00139524 0.997843 0.694642 0.00104809 0.0018798 0.00085937 0.455627 0.0018798 0.437099 0.000128151 1.02 0.88759 0.534706 0.285928 1.71658e-07 3.05974e-09 2388.72 3132.24 -0.0562981 0.482128 0.27758 0.254301 -0.593189 -0.169505 0.494338 -0.268056 -0.226291 1.582 1 0 296.789 0 2.07503 1.58 0.00029992 0.86022 0.65025 0.418534 0.407869 2.07526 130.6 83.7309 18.7099 60.775 0.00403312 0 -40 10
0.681 1.97349e-08 2.5389e-06 0.0909153 0.090912 0.012041 8.9704e-06 0.00115405 0.113644 0.000657357 0.114297 0.868108 101.856 0.244985 0.730052 4.14382 0.0550155 0.0390927 0.960907 0.019849 0.00426223 0.0191118 0.00410018 0.00515099 0.00588825 0.20604 0.23553 57.9814 -87.8951 126.187 15.9755 145.014 0.000141952 0.267112 192.902 0.310648 0.067381 0.00409525 0.000561666 0.00138279 0.986989 0.991733 -2.97416e-06 -85.667 0.0929924 31193 301.069 0.983519 0.319147 0.736374 0.736369 9.99958 2.98119e-06 1.19247e-05 0.130838 0.980737 0.931059 -0.0132931 4.89891e-06 0.501652 -1.88788e-20 6.9574e-24 -1.88719e-20 0.00139524 0.997818 8.59371e-05 0.152568 2.85181 0.00139524 0.997843 0.694748 0.00104811 0.00187981 0.000859371 0.455627 0.0018798 0.437108 0.000128154 1.02 0.887591 0.534705 0.28593 1.71658e-07 3.05976e-09 2388.7 3132.12 -0.0562904 0.482128 0.27758 0.254294 -0.59319 -0.169505 0.494361 -0.268054 -0.226315 1.583 1 0 296.797 0 2.0752 1.581 0.000299919 0.860169 0.650303 0.418301 0.407897 2.07544 130.609 83.7323 18.71 60.7756 0.00403307 0 -40 10
0.682 1.97638e-08 2.5389e-06 0.0909935 0.0909902 0.012041 8.98355e-06 0.00115405 0.113742 0.000657361 0.114395 0.868166 101.856 0.244978 0.730138 4.14398 0.0550223 0.0390941 0.960906 0.0198488 0.00426238 0.0191116 0.0041003 0.00515117 0.00588843 0.206047 0.235537 57.9814 -87.8951 126.187 15.9755 145.014 0.000141946 0.267112 192.902 0.310647 0.067381 0.00409526 0.000561667 0.00138279 0.986989 0.991733 -2.97418e-06 -85.667 0.0929925 31192.9 301.073 0.983519 0.319147 0.736346 0.736342 9.99958 2.9812e-06 1.19247e-05 0.13084 0.980746 0.931063 -0.0132931 4.89894e-06 0.501659 -1.88796e-20 6.95774e-24 -1.88727e-20 0.00139524 0.997818 8.59371e-05 0.152569 2.85181 0.00139524 0.997843 0.694855 0.00104813 0.00187981 0.000859371 0.455627 0.00187981 0.437116 0.000128157 1.02 0.887592 0.534705 0.285931 1.71658e-07 3.05978e-09 2388.68 3132 -0.0562827 0.482128 0.27758 0.254286 -0.593191 -0.169505 0.494383 -0.268052 -0.22634 1.584 1 0 296.805 0 2.07537 1.582 0.000299919 0.860117 0.650356 0.418068 0.407926 2.07561 130.618 83.7336 18.7101 60.7763 0.00403301 0 -40 10
0.683 1.97928e-08 2.5389e-06 0.0910717 0.0910684 0.012041 8.99671e-06 0.00115405 0.11384 0.000657364 0.114492 0.868225 101.856 0.244971 0.730224 4.14413 0.0550291 0.0390956 0.960904 0.0198486 0.00426253 0.0191114 0.00410043 0.00515135 0.00588861 0.206054 0.235544 57.9815 -87.8951 126.188 15.9755 145.014 0.000141941 0.267112 192.902 0.310647 0.0673809 0.00409526 0.000561667 0.00138279 0.986989 0.991733 -2.97419e-06 -85.667 0.0929926 31192.9 301.077 0.983519 0.319147 0.736319 0.736314 9.99958 2.9812e-06 1.19247e-05 0.130841 0.980755 0.931067 -0.0132931 4.89897e-06 0.501665 -1.88804e-20 6.95808e-24 -1.88735e-20 0.00139524 0.997818 8.59372e-05 0.152569 2.85181 0.00139524 0.997843 0.694961 0.00104815 0.00187981 0.000859372 0.455627 0.00187981 0.437125 0.000128161 1.02 0.887593 0.534705 0.285933 1.71658e-07 3.0598e-09 2388.67 3131.89 -0.0562751 0.482128 0.277579 0.254279 -0.593193 -0.169505 0.494404 -0.26805 -0.226364 1.585 1 0 296.812 0 2.07554 1.583 0.000299919 0.860066 0.65041 0.417836 0.407955 2.07578 130.627 83.735 18.7101 60.7769 0.00403296 0 -40 10
0.684 1.98217e-08 2.5389e-06 0.0911498 0.0911465 0.0120409 9.00987e-06 0.00115405 0.113937 0.000657367 0.11459 0.868283 101.856 0.244964 0.73031 4.14429 0.055036 0.0390971 0.960903 0.0198485 0.00426268 0.0191112 0.00410055 0.00515154 0.00588879 0.206062 0.235552 57.9816 -87.8951 126.188 15.9754 145.014 0.000141936 0.267112 192.902 0.310647 0.0673809 0.00409526 0.000561668 0.00138279 0.986989 0.991733 -2.9742e-06 -85.667 0.0929927 31192.9 301.081 0.983519 0.319147 0.736292 0.736287 9.99958 2.9812e-06 1.19247e-05 0.130843 0.980763 0.931071 -0.0132931 4.899e-06 0.501671 -1.88812e-20 6.95842e-24 -1.88743e-20 0.00139524 0.997818 8.59373e-05 0.152569 2.85181 0.00139524 0.997843 0.695067 0.00104817 0.00187981 0.000859373 0.455627 0.00187981 0.437134 0.000128164 1.02 0.887594 0.534705 0.285934 1.71659e-07 3.05982e-09 2388.65 3131.77 -0.0562675 0.482128 0.277579 0.254272 -0.593194 -0.169505 0.494426 -0.268048 -0.226387 1.586 1 0 296.82 0 2.07571 1.584 0.000299918 0.860016 0.650463 0.417604 0.407983 2.07595 130.636 83.7363 18.7102 60.7776 0.0040329 0 -40 10
0.685 1.98507e-08 2.5389e-06 0.0912278 0.0912245 0.0120409 9.02303e-06 0.00115405 0.114035 0.00065737 0.114687 0.868341 101.856 0.244957 0.730396 4.14444 0.0550428 0.0390985 0.960901 0.0198483 0.00426283 0.019111 0.00410068 0.00515172 0.00588897 0.206069 0.235559 57.9816 -87.8951 126.189 15.9754 145.014 0.00014193 0.267113 192.901 0.310646 0.0673808 0.00409526 0.000561669 0.0013828 0.986989 0.991733 -2.97422e-06 -85.667 0.0929927 31192.9 301.085 0.983519 0.319147 0.736264 0.73626 9.99958 2.98121e-06 1.19247e-05 0.130844 0.980772 0.931074 -0.0132931 4.89903e-06 0.501677 -1.88821e-20 6.95876e-24 -1.88751e-20 0.00139524 0.997818 8.59374e-05 0.152569 2.85181 0.00139524 0.997843 0.695173 0.00104819 0.00187981 0.000859374 0.455626 0.00187981 0.437143 0.000128168 1.02 0.887595 0.534704 0.285936 1.71659e-07 3.05985e-09 2388.63 3131.65 -0.05626 0.482128 0.277579 0.254264 -0.593195 -0.169505 0.494448 -0.268046 -0.226411 1.587 1 0 296.828 0 2.07588 1.585 0.000299918 0.859965 0.650517 0.417373 0.408012 2.07612 130.645 83.7377 18.7103 60.7782 0.00403285 0 -40 10
0.686 1.98796e-08 2.5389e-06 0.0913057 0.0913025 0.0120409 9.03618e-06 0.00115405 0.114132 0.000657374 0.114785 0.8684 101.855 0.24495 0.730483 4.1446 0.0550497 0.0391 0.9609 0.0198481 0.00426298 0.0191108 0.0041008 0.00515191 0.00588916 0.206076 0.235566 57.9817 -87.8951 126.189 15.9753 145.014 0.000141925 0.267113 192.901 0.310646 0.0673808 0.00409527 0.000561669 0.0013828 0.986989 0.991733 -2.97423e-06 -85.667 0.0929928 31192.8 301.089 0.983519 0.319147 0.736237 0.736233 9.99958 2.98121e-06 1.19247e-05 0.130846 0.980781 0.931078 -0.0132931 4.89906e-06 0.501683 -1.88829e-20 6.9591e-24 -1.88759e-20 0.00139524 0.997818 8.59374e-05 0.152569 2.85181 0.00139524 0.997843 0.695279 0.00104821 0.00187981 0.000859374 0.455626 0.00187981 0.437152 0.000128171 1.02 0.887597 0.534704 0.285937 1.71659e-07 3.05987e-09 2388.62 3131.54 -0.0562525 0.482128 0.277578 0.254257 -0.593197 -0.169505 0.494469 -0.268044 -0.226435 1.588 1 0 296.836 0 2.07605 1.586 0.000299918 0.859915 0.65057 0.417143 0.408041 2.07629 130.655 83.739 18.7104 60.7789 0.00403279 0 -40 10
0.687 1.99086e-08 2.5389e-06 0.0913836 0.0913804 0.0120409 9.04934e-06 0.00115405 0.11423 0.000657377 0.114882 0.868458 101.855 0.244943 0.730569 4.14476 0.0550565 0.0391015 0.960899 0.0198479 0.00426313 0.0191107 0.00410093 0.00515209 0.00588934 0.206084 0.235574 57.9818 -87.8951 126.19 15.9753 145.014 0.00014192 0.267113 192.901 0.310645 0.0673807 0.00409527 0.00056167 0.0013828 0.986989 0.991733 -2.97425e-06 -85.667 0.0929929 31192.8 301.093 0.983519 0.319147 0.73621 0.736206 9.99958 2.98122e-06 1.19248e-05 0.130847 0.980789 0.931082 -0.0132931 4.89908e-06 0.50169 -1.88837e-20 6.95944e-24 -1.88767e-20 0.00139524 0.997818 8.59375e-05 0.152569 2.85181 0.00139524 0.997842 0.695385 0.00104823 0.00187981 0.000859375 0.455626 0.00187981 0.43716 0.000128174 1.02 0.887598 0.534704 0.285938 1.71659e-07 3.05989e-09 2388.6 3131.42 -0.0562451 0.482128 0.277578 0.25425 -0.593198 -0.169505 0.494491 -0.268042 -0.226458 1.589 1 0 296.843 0 2.07622 1.587 0.000299918 0.859865 0.650623 0.416913 0.408069 2.07646 130.664 83.7403 18.7105 60.7795 0.00403274 0 -40 10
0.688 1.99375e-08 2.5389e-06 0.0914614 0.0914582 0.0120409 9.0625e-06 0.00115405 0.114327 0.00065738 0.11498 0.868517 101.855 0.244937 0.730655 4.14491 0.0550634 0.039103 0.960897 0.0198477 0.00426328 0.0191105 0.00410105 0.00515228 0.00588952 0.206091 0.235581 57.9818 -87.8951 126.19 15.9753 145.014 0.000141915 0.267113 192.901 0.310645 0.0673807 0.00409527 0.000561671 0.0013828 0.986988 0.991733 -2.97426e-06 -85.667 0.092993 31192.8 301.097 0.983519 0.319147 0.736184 0.736179 9.99958 2.98122e-06 1.19248e-05 0.130849 0.980798 0.931085 -0.0132931 4.89911e-06 0.501696 -1.88845e-20 6.95978e-24 -1.88775e-20 0.00139525 0.997818 8.59376e-05 0.152569 2.85181 0.00139525 0.997842 0.695491 0.00104825 0.00187982 0.000859376 0.455626 0.00187981 0.437169 0.000128178 1.02 0.887599 0.534703 0.28594 1.7166e-07 3.05991e-09 2388.58 3131.31 -0.0562376 0.482128 0.277578 0.254243 -0.5932 -0.169506 0.494512 -0.268039 -0.226482 1.59 1 0 296.851 0 2.07639 1.588 0.000299917 0.859815 0.650676 0.416683 0.408098 2.07663 130.673 83.7417 18.7105 60.7801 0.00403268 0 -40 10
0.689 1.99664e-08 2.5389e-06 0.0915392 0.091536 0.0120409 9.07566e-06 0.00115405 0.114424 0.000657383 0.115077 0.868575 101.855 0.24493 0.730742 4.14507 0.0550703 0.0391045 0.960896 0.0198475 0.00426343 0.0191103 0.00410118 0.00515246 0.00588971 0.206098 0.235588 57.9819 -87.8951 126.191 15.9752 145.014 0.00014191 0.267113 192.901 0.310645 0.0673806 0.00409528 0.000561671 0.0013828 0.986988 0.991733 -2.97427e-06 -85.6669 0.0929931 31192.8 301.102 0.983519 0.319147 0.736157 0.736153 9.99958 2.98123e-06 1.19248e-05 0.13085 0.980806 0.931089 -0.0132931 4.89914e-06 0.501702 -1.88853e-20 6.96013e-24 -1.88784e-20 0.00139525 0.997818 8.59377e-05 0.15257 2.85182 0.00139525 0.997842 0.695597 0.00104827 0.00187982 0.000859377 0.455626 0.00187982 0.437178 0.000128181 1.02 0.8876 0.534703 0.285941 1.7166e-07 3.05993e-09 2388.57 3131.19 -0.0562303 0.482128 0.277578 0.254235 -0.593201 -0.169506 0.494533 -0.268037 -0.226505 1.591 1 0 296.859 0 2.07656 1.589 0.000299917 0.859766 0.65073 0.416455 0.408126 2.0768 130.682 83.743 18.7106 60.7808 0.00403263 0 -40 10
0.69 1.99954e-08 2.5389e-06 0.0916169 0.0916137 0.0120409 9.08881e-06 0.00115405 0.114521 0.000657387 0.115174 0.868634 101.855 0.244923 0.730828 4.14523 0.0550772 0.0391059 0.960894 0.0198474 0.00426358 0.0191101 0.0041013 0.00515265 0.00588989 0.206106 0.235596 57.9819 -87.8951 126.191 15.9752 145.014 0.000141905 0.267113 192.901 0.310644 0.0673806 0.00409528 0.000561672 0.00138281 0.986988 0.991733 -2.97429e-06 -85.6669 0.0929932 31192.8 301.106 0.983519 0.319147 0.73613 0.736126 9.99958 2.98123e-06 1.19248e-05 0.130852 0.980815 0.931093 -0.0132931 4.89917e-06 0.501709 -1.88861e-20 6.96047e-24 -1.88792e-20 0.00139525 0.997818 8.59377e-05 0.15257 2.85182 0.00139525 0.997842 0.695703 0.00104829 0.00187982 0.000859377 0.455625 0.00187982 0.437187 0.000128185 1.02 0.887601 0.534703 0.285943 1.7166e-07 3.05995e-09 2388.55 3131.08 -0.0562229 0.482128 0.277577 0.254228 -0.593202 -0.169506 0.494555 -0.268035 -0.226528 1.592 1 0 296.866 0 2.07673 1.59 0.000299917 0.859717 0.650783 0.416226 0.408155 2.07697 130.691 83.7443 18.7107 60.7814 0.00403257 0 -40 10
0.691 2.00243e-08 2.5389e-06 0.0916946 0.0916913 0.0120409 9.10197e-06 0.00115405 0.114618 0.00065739 0.115271 0.868693 101.855 0.244916 0.730915 4.14539 0.0550841 0.0391074 0.960893 0.0198472 0.00426373 0.0191099 0.00410143 0.00515283 0.00589008 0.206113 0.235603 57.982 -87.8952 126.191 15.9752 145.014 0.0001419 0.267114 192.9 0.310644 0.0673805 0.00409528 0.000561672 0.00138281 0.986988 0.991733 -2.9743e-06 -85.6669 0.0929932 31192.7 301.11 0.983519 0.319147 0.736104 0.7361 9.99958 2.98124e-06 1.19248e-05 0.130853 0.980823 0.931096 -0.0132931 4.8992e-06 0.501715 -1.88869e-20 6.96081e-24 -1.888e-20 0.00139525 0.997818 8.59378e-05 0.15257 2.85182 0.00139525 0.997842 0.695809 0.00104831 0.00187982 0.000859378 0.455625 0.00187982 0.437196 0.000128188 1.02 0.887602 0.534702 0.285944 1.7166e-07 3.05998e-09 2388.53 3130.97 -0.0562156 0.482128 0.277577 0.254221 -0.593204 -0.169506 0.494576 -0.268033 -0.226551 1.593 1 0 296.874 0 2.0769 1.591 0.000299916 0.859668 0.650836 0.415998 0.408183 2.07714 130.7 83.7456 18.7108 60.782 0.00403252 0 -40 10
0.692 2.00533e-08 2.5389e-06 0.0917721 0.0917689 0.0120408 9.11513e-06 0.00115405 0.114715 0.000657393 0.115368 0.868751 101.854 0.244909 0.731002 4.14555 0.055091 0.0391089 0.960891 0.019847 0.00426389 0.0191097 0.00410156 0.00515302 0.00589026 0.206121 0.23561 57.9821 -87.8952 126.192 15.9751 145.014 0.000141894 0.267114 192.9 0.310643 0.0673805 0.00409528 0.000561673 0.00138281 0.986988 0.991733 -2.97432e-06 -85.6669 0.0929933 31192.7 301.114 0.983519 0.319147 0.736078 0.736073 9.99958 2.98124e-06 1.19249e-05 0.130855 0.980832 0.9311 -0.0132931 4.89923e-06 0.501721 -1.88878e-20 6.96115e-24 -1.88808e-20 0.00139525 0.997818 8.59379e-05 0.15257 2.85182 0.00139525 0.997842 0.695915 0.00104833 0.00187982 0.000859379 0.455625 0.00187982 0.437204 0.000128191 1.02 0.887603 0.534702 0.285946 1.71661e-07 3.06e-09 2388.52 3130.86 -0.0562084 0.482128 0.277577 0.254214 -0.593205 -0.169506 0.494596 -0.268031 -0.226574 1.594 1 0 296.881 0 2.07707 1.592 0.000299916 0.859619 0.650889 0.415771 0.408212 2.07731 130.709 83.7469 18.7108 60.7826 0.00403247 0 -40 10
0.693 2.00822e-08 2.5389e-06 0.0918497 0.0918465 0.0120408 9.12829e-06 0.00115405 0.114812 0.000657396 0.115465 0.86881 101.854 0.244902 0.731089 4.14571 0.0550979 0.0391104 0.96089 0.0198468 0.00426404 0.0191096 0.00410168 0.00515321 0.00589045 0.206128 0.235618 57.9821 -87.8952 126.192 15.9751 145.014 0.000141889 0.267114 192.9 0.310643 0.0673804 0.00409529 0.000561674 0.00138281 0.986988 0.991733 -2.97433e-06 -85.6669 0.0929934 31192.7 301.118 0.983519 0.319147 0.736051 0.736047 9.99958 2.98125e-06 1.19249e-05 0.130857 0.98084 0.931104 -0.0132931 4.89925e-06 0.501728 -1.88886e-20 6.96149e-24 -1.88816e-20 0.00139525 0.997818 8.5938e-05 0.15257 2.85182 0.00139525 0.997841 0.696021 0.00104835 0.00187982 0.00085938 0.455625 0.00187982 0.437213 0.000128195 1.02 0.887604 0.534702 0.285947 1.71661e-07 3.06002e-09 2388.5 3130.74 -0.0562011 0.482128 0.277576 0.254207 -0.593206 -0.169506 0.494617 -0.268029 -0.226597 1.595 1 0 296.889 0 2.07724 1.593 0.000299916 0.85957 0.650942 0.415545 0.40824 2.07748 130.718 83.7482 18.7109 60.7833 0.00403241 0 -40 10
0.694 2.01112e-08 2.5389e-06 0.0919271 0.0919239 0.0120408 9.14144e-06 0.00115405 0.114909 0.000657399 0.115562 0.868869 101.854 0.244895 0.731176 4.14587 0.0551048 0.0391119 0.960888 0.0198466 0.00426419 0.0191094 0.00410181 0.00515339 0.00589063 0.206136 0.235625 57.9822 -87.8952 126.193 15.975 145.014 0.000141884 0.267114 192.9 0.310643 0.0673804 0.00409529 0.000561674 0.00138281 0.986988 0.991733 -2.97434e-06 -85.6669 0.0929935 31192.7 301.122 0.983519 0.319147 0.736025 0.736021 9.99958 2.98125e-06 1.19249e-05 0.130858 0.980848 0.931107 -0.0132931 4.89928e-06 0.501734 -1.88894e-20 6.96183e-24 -1.88824e-20 0.00139525 0.997818 8.59381e-05 0.15257 2.85182 0.00139525 0.997841 0.696127 0.00104837 0.00187982 0.000859381 0.455624 0.00187982 0.437222 0.000128198 1.02 0.887605 0.534702 0.285949 1.71661e-07 3.06004e-09 2388.48 3130.63 -0.056194 0.482129 0.277576 0.2542 -0.593207 -0.169506 0.494638 -0.268027 -0.226619 1.596 1 0 296.896 0 2.07741 1.594 0.000299915 0.859522 0.650995 0.415319 0.408269 2.07764 130.727 83.7495 18.711 60.7839 0.00403236 0 -40 10
0.695 2.01401e-08 2.53891e-06 0.0920045 0.0920013 0.0120408 9.1546e-06 0.00115405 0.115006 0.000657403 0.115658 0.868928 101.854 0.244888 0.731263 4.14603 0.0551117 0.0391135 0.960887 0.0198464 0.00426434 0.0191092 0.00410194 0.00515358 0.00589082 0.206143 0.235633 57.9823 -87.8952 126.193 15.975 145.014 0.000141879 0.267114 192.9 0.310642 0.0673803 0.00409529 0.000561675 0.00138282 0.986988 0.991733 -2.97436e-06 -85.6669 0.0929936 31192.7 301.126 0.983519 0.319147 0.735999 0.735995 9.99958 2.98126e-06 1.19249e-05 0.13086 0.980857 0.931111 -0.0132931 4.89931e-06 0.50174 -1.88902e-20 6.96217e-24 -1.88832e-20 0.00139525 0.997818 8.59381e-05 0.15257 2.85182 0.00139525 0.997841 0.696233 0.00104839 0.00187982 0.000859381 0.455624 0.00187982 0.437231 0.000128202 1.02 0.887606 0.534701 0.28595 1.71661e-07 3.06006e-09 2388.47 3130.52 -0.0561868 0.482129 0.277576 0.254193 -0.593209 -0.169506 0.494658 -0.268025 -0.226642 1.597 1 0 296.904 0 2.07758 1.595 0.000299915 0.859474 0.651048 0.415093 0.408297 2.07781 130.736 83.7507 18.7111 60.7845 0.00403231 0 -40 10
0.696 2.01691e-08 2.53891e-06 0.0920818 0.0920787 0.0120408 9.16776e-06 0.00115405 0.115102 0.000657406 0.115755 0.868987 101.854 0.244881 0.73135 4.14619 0.0551186 0.039115 0.960885 0.0198462 0.0042645 0.019109 0.00410206 0.00515377 0.00589101 0.206151 0.23564 57.9823 -87.8952 126.194 15.975 145.014 0.000141874 0.267115 192.9 0.310642 0.0673803 0.0040953 0.000561676 0.00138282 0.986988 0.991733 -2.97437e-06 -85.6669 0.0929936 31192.6 301.13 0.983519 0.319147 0.735974 0.735969 9.99958 2.98126e-06 1.19249e-05 0.130861 0.980865 0.931114 -0.0132931 4.89934e-06 0.501747 -1.8891e-20 6.96251e-24 -1.88841e-20 0.00139525 0.997818 8.59382e-05 0.152571 2.85182 0.00139525 0.997841 0.696338 0.00104841 0.00187983 0.000859382 0.455624 0.00187983 0.437239 0.000128205 1.02 0.887607 0.534701 0.285952 1.71662e-07 3.06009e-09 2388.45 3130.41 -0.0561797 0.482129 0.277576 0.254186 -0.59321 -0.169506 0.494679 -0.268023 -0.226664 1.598 1 0 296.911 0 2.07775 1.596 0.000299915 0.859426 0.651101 0.414868 0.408326 2.07798 130.745 83.752 18.7111 60.7851 0.00403225 0 -40 10
0.697 2.0198e-08 2.53891e-06 0.0921591 0.0921559 0.0120408 9.18091e-06 0.00115405 0.115199 0.000657409 0.115852 0.869046 101.854 0.244874 0.731437 4.14635 0.0551255 0.0391165 0.960884 0.019846 0.00426465 0.0191088 0.00410219 0.00515396 0.00589119 0.206158 0.235648 57.9824 -87.8952 126.194 15.9749 145.014 0.000141869 0.267115 192.9 0.310641 0.0673802 0.0040953 0.000561676 0.00138282 0.986988 0.991733 -2.97439e-06 -85.6669 0.0929937 31192.6 301.135 0.983519 0.319147 0.735948 0.735943 9.99958 2.98126e-06 1.1925e-05 0.130863 0.980873 0.931118 -0.0132931 4.89937e-06 0.501753 -1.88918e-20 6.96286e-24 -1.88849e-20 0.00139526 0.997818 8.59383e-05 0.152571 2.85182 0.00139526 0.997841 0.696444 0.00104843 0.00187983 0.000859383 0.455624 0.00187983 0.437248 0.000128208 1.02 0.887608 0.534701 0.285953 1.71662e-07 3.06011e-09 2388.43 3130.3 -0.0561727 0.482129 0.277575 0.254179 -0.593211 -0.169506 0.494699 -0.268021 -0.226687 1.599 1 0 296.918 0 2.07792 1.597 0.000299914 0.859378 0.651154 0.414644 0.408354 2.07815 130.754 83.7533 18.7112 60.7857 0.0040322 0 -40 10
0.698 2.0227e-08 2.53891e-06 0.0922363 0.0922332 0.0120408 9.19407e-06 0.00115405 0.115295 0.000657412 0.115948 0.869105 101.853 0.244868 0.731524 4.14651 0.0551325 0.039118 0.960882 0.0198459 0.0042648 0.0191086 0.00410232 0.00515415 0.00589138 0.206166 0.235655 57.9825 -87.8952 126.195 15.9749 145.014 0.000141865 0.267115 192.899 0.310641 0.0673802 0.0040953 0.000561677 0.00138282 0.986988 0.991733 -2.9744e-06 -85.6669 0.0929938 31192.6 301.139 0.983519 0.319147 0.735922 0.735918 9.99958 2.98127e-06 1.1925e-05 0.130864 0.980882 0.931121 -0.0132931 4.8994e-06 0.50176 -1.88927e-20 6.9632e-24 -1.88857e-20 0.00139526 0.997818 8.59384e-05 0.152571 2.85182 0.00139526 0.997841 0.69655 0.00104845 0.00187983 0.000859384 0.455624 0.00187983 0.437257 0.000128212 1.02 0.887609 0.5347 0.285954 1.71662e-07 3.06013e-09 2388.42 3130.19 -0.0561656 0.482129 0.277575 0.254172 -0.593213 -0.169506 0.494719 -0.268019 -0.226709 1.6 1 0 296.926 0 2.07809 1.598 0.000299914 0.859331 0.651207 0.41442 0.408383 2.07832 130.764 83.7546 18.7113 60.7863 0.00403215 0 -40 10
0.699 2.02559e-08 2.53891e-06 0.0923135 0.0923103 0.0120407 9.20723e-06 0.00115405 0.115392 0.000657415 0.116045 0.869164 101.853 0.244861 0.731611 4.14667 0.0551394 0.0391195 0.96088 0.0198457 0.00426496 0.0191084 0.00410245 0.00515434 0.00589157 0.206173 0.235663 57.9825 -87.8952 126.195 15.9749 145.014 0.00014186 0.267115 192.899 0.310641 0.0673801 0.0040953 0.000561677 0.00138282 0.986988 0.991733 -2.97442e-06 -85.6669 0.0929939 31192.6 301.143 0.983519 0.319147 0.735897 0.735892 9.99958 2.98127e-06 1.1925e-05 0.130866 0.98089 0.931125 -0.0132931 4.89942e-06 0.501766 -1.88935e-20 6.96354e-24 -1.88865e-20 0.00139526 0.997818 8.59384e-05 0.152571 2.85182 0.00139526 0.99784 0.696655 0.00104847 0.00187983 0.000859384 0.455623 0.00187983 0.437266 0.000128215 1.02 0.88761 0.5347 0.285956 1.71662e-07 3.06015e-09 2388.4 3130.08 -0.0561586 0.482129 0.277575 0.254165 -0.593214 -0.169506 0.494739 -0.268017 -0.226731 1.601 1 0 296.933 0 2.07825 1.599 0.000299914 0.859284 0.65126 0.414196 0.408411 2.07849 130.773 83.7558 18.7114 60.7869 0.0040321 0 -40 10
0.7 2.02848e-08 2.53891e-06 0.0923905 0.0923874 0.0120407 9.22038e-06 0.00115405 0.115488 0.000657418 0.116141 0.869223 101.853 0.244854 0.731699 4.14683 0.0551464 0.039121 0.960879 0.0198455 0.00426511 0.0191082 0.00410258 0.00515453 0.00589176 0.206181 0.23567 57.9826 -87.8952 126.196 15.9748 145.014 0.000141855 0.267115 192.899 0.31064 0.0673801 0.00409531 0.000561678 0.00138283 0.986988 0.991733 -2.97443e-06 -85.6669 0.092994 31192.6 301.147 0.983519 0.319147 0.735871 0.735867 9.99958 2.98128e-06 1.1925e-05 0.130868 0.980898 0.931128 -0.0132931 4.89945e-06 0.501773 -1.88943e-20 6.96388e-24 -1.88873e-20 0.00139526 0.997818 8.59385e-05 0.152571 2.85182 0.00139526 0.99784 0.696761 0.00104849 0.00187983 0.000859385 0.455623 0.00187983 0.437274 0.000128219 1.02 0.887611 0.5347 0.285957 1.71663e-07 3.06017e-09 2388.38 3129.97 -0.0561517 0.482129 0.277574 0.254159 -0.593215 -0.169506 0.494759 -0.268015 -0.226753 1.602 1 0 296.94 0 2.07842 1.6 0.000299914 0.859237 0.651313 0.413974 0.408439 2.07866 130.782 83.7571 18.7114 60.7876 0.00403205 0 -40 10
0.701 2.03138e-08 2.53891e-06 0.0924676 0.0924644 0.0120407 9.23354e-06 0.00115405 0.115584 0.000657422 0.116237 0.869283 101.853 0.244847 0.731786 4.14699 0.0551533 0.0391226 0.960877 0.0198453 0.00426527 0.0191081 0.00410271 0.00515472 0.00589195 0.206189 0.235678 57.9826 -87.8952 126.196 15.9748 145.014 0.00014185 0.267115 192.899 0.31064 0.06738 0.00409531 0.000561679 0.00138283 0.986988 0.991733 -2.97444e-06 -85.6668 0.0929941 31192.5 301.151 0.983519 0.319147 0.735846 0.735842 9.99958 2.98128e-06 1.1925e-05 0.130869 0.980906 0.931132 -0.0132931 4.89948e-06 0.501779 -1.88951e-20 6.96423e-24 -1.88881e-20 0.00139526 0.997818 8.59386e-05 0.152571 2.85183 0.00139526 0.99784 0.696866 0.0010485 0.00187983 0.000859386 0.455623 0.00187983 0.437283 0.000128222 1.02 0.887612 0.5347 0.285959 1.71663e-07 3.06019e-09 2388.37 3129.86 -0.0561448 0.482129 0.277574 0.254152 -0.593216 -0.169506 0.494779 -0.268013 -0.226775 1.603 1 0 296.947 0 2.07859 1.601 0.000299913 0.85919 0.651366 0.413751 0.408468 2.07883 130.791 83.7583 18.7115 60.7882 0.00403199 0 -40 10
0.702 2.03427e-08 2.53891e-06 0.0925445 0.0925414 0.0120407 9.2467e-06 0.00115405 0.115681 0.000657425 0.116333 0.869342 101.853 0.24484 0.731874 4.14716 0.0551603 0.0391241 0.960876 0.0198451 0.00426542 0.0191079 0.00410283 0.00515491 0.00589214 0.206196 0.235685 57.9827 -87.8952 126.197 15.9747 145.014 0.000141845 0.267116 192.899 0.310639 0.06738 0.00409531 0.000561679 0.00138283 0.986988 0.991733 -2.97446e-06 -85.6668 0.0929941 31192.5 301.155 0.983519 0.319147 0.735821 0.735817 9.99958 2.98129e-06 1.1925e-05 0.130871 0.980914 0.931135 -0.0132931 4.89951e-06 0.501785 -1.88959e-20 6.96457e-24 -1.8889e-20 0.00139526 0.997818 8.59387e-05 0.152571 2.85183 0.00139526 0.99784 0.696972 0.00104852 0.00187983 0.000859387 0.455623 0.00187983 0.437292 0.000128225 1.02 0.887613 0.534699 0.28596 1.71663e-07 3.06022e-09 2388.35 3129.76 -0.0561379 0.482129 0.277574 0.254145 -0.593218 -0.169506 0.494799 -0.268011 -0.226797 1.604 1 0 296.955 0 2.07876 1.602 0.000299913 0.859144 0.651419 0.41353 0.408496 2.079 130.8 83.7596 18.7116 60.7887 0.00403194 0 -40 10
0.703 2.03717e-08 2.53891e-06 0.0926214 0.0926183 0.0120407 9.25985e-06 0.00115405 0.115777 0.000657428 0.11643 0.869401 101.853 0.244833 0.731962 4.14732 0.0551673 0.0391256 0.960874 0.0198449 0.00426558 0.0191077 0.00410296 0.0051551 0.00589232 0.206204 0.235693 57.9828 -87.8952 126.197 15.9747 145.014 0.00014184 0.267116 192.899 0.310639 0.0673799 0.00409532 0.00056168 0.00138283 0.986988 0.991733 -2.97447e-06 -85.6668 0.0929942 31192.5 301.16 0.983519 0.319147 0.735796 0.735792 9.99958 2.98129e-06 1.19251e-05 0.130872 0.980923 0.931139 -0.0132931 4.89954e-06 0.501792 -1.88967e-20 6.96491e-24 -1.88898e-20 0.00139526 0.997818 8.59387e-05 0.152572 2.85183 0.00139526 0.99784 0.697077 0.00104854 0.00187984 0.000859387 0.455623 0.00187983 0.437301 0.000128229 1.02 0.887614 0.534699 0.285962 1.71663e-07 3.06024e-09 2388.33 3129.65 -0.056131 0.482129 0.277574 0.254138 -0.593219 -0.169507 0.494818 -0.268009 -0.226818 1.605 1 0 296.962 0 2.07893 1.603 0.000299913 0.859097 0.651472 0.413309 0.408524 2.07917 130.809 83.7608 18.7116 60.7893 0.00403189 0 -40 10
0.704 2.04006e-08 2.53891e-06 0.0926982 0.0926951 0.0120407 9.27301e-06 0.00115405 0.115873 0.000657431 0.116526 0.869461 101.853 0.244826 0.732049 4.14748 0.0551743 0.0391272 0.960873 0.0198447 0.00426573 0.0191075 0.00410309 0.00515529 0.00589251 0.206212 0.235701 57.9828 -87.8952 126.198 15.9747 145.014 0.000141835 0.267116 192.898 0.310639 0.0673799 0.00409532 0.000561681 0.00138283 0.986988 0.991733 -2.97449e-06 -85.6668 0.0929943 31192.5 301.164 0.983519 0.319147 0.735771 0.735767 9.99958 2.9813e-06 1.19251e-05 0.130874 0.980931 0.931142 -0.0132931 4.89957e-06 0.501798 -1.88976e-20 6.96525e-24 -1.88906e-20 0.00139526 0.997818 8.59388e-05 0.152572 2.85183 0.00139526 0.99784 0.697183 0.00104856 0.00187984 0.000859388 0.455622 0.00187984 0.437309 0.000128232 1.02 0.887615 0.534699 0.285963 1.71664e-07 3.06026e-09 2388.32 3129.54 -0.0561242 0.482129 0.277573 0.254132 -0.59322 -0.169507 0.494838 -0.268007 -0.22684 1.606 1 0 296.969 0 2.0791 1.604 0.000299912 0.859051 0.651525 0.413088 0.408553 2.07934 130.818 83.762 18.7117 60.7899 0.00403184 0 -40 10
0.705 2.04296e-08 2.53891e-06 0.092775 0.0927719 0.0120407 9.28617e-06 0.00115405 0.115969 0.000657434 0.116622 0.86952 101.852 0.244819 0.732137 4.14765 0.0551813 0.0391287 0.960871 0.0198445 0.00426589 0.0191073 0.00410322 0.00515548 0.00589271 0.206219 0.235708 57.9829 -87.8952 126.198 15.9746 145.014 0.000141831 0.267116 192.898 0.310638 0.0673798 0.00409532 0.000561681 0.00138284 0.986988 0.991733 -2.9745e-06 -85.6668 0.0929944 31192.4 301.168 0.983519 0.319147 0.735746 0.735742 9.99958 2.9813e-06 1.19251e-05 0.130876 0.980939 0.931146 -0.0132931 4.8996e-06 0.501805 -1.88984e-20 6.9656e-24 -1.88914e-20 0.00139526 0.997818 8.59389e-05 0.152572 2.85183 0.00139526 0.99784 0.697288 0.00104858 0.00187984 0.000859389 0.455622 0.00187984 0.437318 0.000128235 1.02 0.887617 0.534698 0.285965 1.71664e-07 3.06028e-09 2388.3 3129.44 -0.0561175 0.482129 0.277573 0.254125 -0.593221 -0.169507 0.494857 -0.268005 -0.226861 1.607 1 0 296.976 0 2.07927 1.605 0.000299912 0.859005 0.651578 0.412868 0.408581 2.0795 130.827 83.7632 18.7118 60.7905 0.00403179 0 -40 10
0.706 2.04585e-08 2.53891e-06 0.0928517 0.0928486 0.0120407 9.29932e-06 0.00115405 0.116065 0.000657437 0.116718 0.869579 101.852 0.244812 0.732225 4.14781 0.0551883 0.0391303 0.96087 0.0198443 0.00426604 0.0191071 0.00410335 0.00515567 0.0058929 0.206227 0.235716 57.983 -87.8952 126.198 15.9746 145.014 0.000141826 0.267116 192.898 0.310638 0.0673798 0.00409532 0.000561682 0.00138284 0.986988 0.991733 -2.97451e-06 -85.6668 0.0929945 31192.4 301.172 0.983519 0.319147 0.735722 0.735717 9.99958 2.98131e-06 1.19251e-05 0.130877 0.980947 0.931149 -0.0132931 4.89962e-06 0.501811 -1.88992e-20 6.96594e-24 -1.88922e-20 0.00139526 0.997818 8.5939e-05 0.152572 2.85183 0.00139526 0.997839 0.697394 0.0010486 0.00187984 0.00085939 0.455622 0.00187984 0.437327 0.000128239 1.02 0.887618 0.534698 0.285966 1.71664e-07 3.0603e-09 2388.28 3129.33 -0.0561107 0.482129 0.277573 0.254118 -0.593223 -0.169507 0.494876 -0.268002 -0.226883 1.608 1 0 296.983 0 2.07944 1.606 0.000299912 0.85896 0.651631 0.412648 0.408609 2.07967 130.836 83.7645 18.7119 60.7911 0.00403174 0 -40 10
0.707 2.04875e-08 2.53891e-06 0.0929284 0.0929253 0.0120406 9.31248e-06 0.00115405 0.11616 0.00065744 0.116813 0.869639 101.852 0.244805 0.732313 4.14797 0.0551953 0.0391318 0.960868 0.0198441 0.0042662 0.0191069 0.00410348 0.00515587 0.00589309 0.206235 0.235723 57.983 -87.8952 126.199 15.9745 145.015 0.000141821 0.267117 192.898 0.310637 0.0673797 0.00409533 0.000561682 0.00138284 0.986988 0.991733 -2.97453e-06 -85.6668 0.0929945 31192.4 301.177 0.983519 0.319147 0.735697 0.735693 9.99958 2.98131e-06 1.19251e-05 0.130879 0.980955 0.931153 -0.0132931 4.89965e-06 0.501818 -1.89e-20 6.96628e-24 -1.8893e-20 0.00139527 0.997818 8.5939e-05 0.152572 2.85183 0.00139527 0.997839 0.697499 0.00104862 0.00187984 0.00085939 0.455622 0.00187984 0.437335 0.000128242 1.02 0.887619 0.534698 0.285968 1.71664e-07 3.06033e-09 2388.27 3129.23 -0.0561041 0.482129 0.277572 0.254112 -0.593224 -0.169507 0.494896 -0.268 -0.226904 1.609 1 0 296.99 0 2.07961 1.607 0.000299911 0.858915 0.651683 0.412429 0.408638 2.07984 130.845 83.7657 18.7119 60.7917 0.00403169 0 -40 10
0.708 2.05164e-08 2.53891e-06 0.093005 0.0930019 0.0120406 9.32564e-06 0.00115405 0.116256 0.000657443 0.116909 0.869699 101.852 0.244798 0.732401 4.14814 0.0552023 0.0391334 0.960867 0.0198439 0.00426636 0.0191067 0.00410362 0.00515606 0.00589328 0.206242 0.235731 57.9831 -87.8952 126.199 15.9745 145.015 0.000141816 0.267117 192.898 0.310637 0.0673797 0.00409533 0.000561683 0.00138284 0.986988 0.991733 -2.97454e-06 -85.6668 0.0929946 31192.4 301.181 0.983519 0.319147 0.735673 0.735668 9.99958 2.98132e-06 1.19252e-05 0.13088 0.980963 0.931156 -0.0132931 4.89968e-06 0.501825 -1.89008e-20 6.96662e-24 -1.88939e-20 0.00139527 0.997818 8.59391e-05 0.152572 2.85183 0.00139527 0.997839 0.697604 0.00104864 0.00187984 0.000859391 0.455621 0.00187984 0.437344 0.000128246 1.02 0.88762 0.534697 0.285969 1.71665e-07 3.06035e-09 2388.25 3129.12 -0.0560974 0.48213 0.277572 0.254105 -0.593225 -0.169507 0.494915 -0.267998 -0.226925 1.61 1 0 296.997 0 2.07977 1.608 0.000299911 0.858869 0.651736 0.412211 0.408666 2.08001 130.854 83.7669 18.712 60.7923 0.00403164 0 -40 10
0.709 2.05453e-08 2.53891e-06 0.0930815 0.0930784 0.0120406 9.33879e-06 0.00115405 0.116352 0.000657446 0.117005 0.869758 101.852 0.244791 0.73249 4.1483 0.0552093 0.0391349 0.960865 0.0198437 0.00426652 0.0191065 0.00410375 0.00515625 0.00589347 0.20625 0.235739 57.9832 -87.8952 126.2 15.9745 145.015 0.000141812 0.267117 192.898 0.310637 0.0673796 0.00409533 0.000561684 0.00138284 0.986988 0.991733 -2.97456e-06 -85.6668 0.0929947 31192.4 301.185 0.983519 0.319147 0.735648 0.735644 9.99958 2.98132e-06 1.19252e-05 0.130882 0.980971 0.931159 -0.0132931 4.89971e-06 0.501831 -1.89016e-20 6.96697e-24 -1.88947e-20 0.00139527 0.997818 8.59392e-05 0.152572 2.85183 0.00139527 0.997839 0.69771 0.00104866 0.00187984 0.000859392 0.455621 0.00187984 0.437353 0.000128249 1.02 0.887621 0.534697 0.285971 1.71665e-07 3.06037e-09 2388.23 3129.02 -0.0560908 0.48213 0.277572 0.254099 -0.593226 -0.169507 0.494933 -0.267996 -0.226946 1.611 1 0 297.004 0 2.07994 1.609 0.000299911 0.858824 0.651789 0.411993 0.408694 2.08018 130.863 83.7681 18.7121 60.7929 0.00403159 0 -40 10
0.71 2.05743e-08 2.53891e-06 0.093158 0.0931549 0.0120406 9.35195e-06 0.00115405 0.116447 0.000657449 0.1171 0.869818 101.852 0.244784 0.732578 4.14847 0.0552163 0.0391365 0.960863 0.0198436 0.00426667 0.0191063 0.00410388 0.00515645 0.00589366 0.206258 0.235747 57.9832 -87.8952 126.2 15.9744 145.015 0.000141807 0.267117 192.897 0.310636 0.0673796 0.00409534 0.000561684 0.00138285 0.986988 0.991733 -2.97457e-06 -85.6668 0.0929948 31192.3 301.189 0.983519 0.319147 0.735624 0.73562 9.99958 2.98133e-06 1.19252e-05 0.130884 0.980979 0.931163 -0.0132931 4.89974e-06 0.501838 -1.89025e-20 6.96731e-24 -1.88955e-20 0.00139527 0.997818 8.59393e-05 0.152573 2.85183 0.00139527 0.997839 0.697815 0.00104868 0.00187985 0.000859393 0.455621 0.00187984 0.437361 0.000128252 1.02 0.887622 0.534697 0.285972 1.71665e-07 3.06039e-09 2388.22 3128.91 -0.0560842 0.48213 0.277572 0.254092 -0.593227 -0.169507 0.494952 -0.267994 -0.226967 1.612 1 0 297.01 0 2.08011 1.61 0.00029991 0.85878 0.651842 0.411775 0.408722 2.08035 130.872 83.7693 18.7121 60.7934 0.00403154 0 -40 10
0.711 2.06032e-08 2.53891e-06 0.0932344 0.0932313 0.0120406 9.36511e-06 0.00115405 0.116543 0.000657452 0.117196 0.869878 101.851 0.244777 0.732666 4.14864 0.0552233 0.0391381 0.960862 0.0198434 0.00426683 0.0191061 0.00410401 0.00515664 0.00589386 0.206266 0.235754 57.9833 -87.8952 126.201 15.9744 145.015 0.000141802 0.267117 192.897 0.310636 0.0673795 0.00409534 0.000561685 0.00138285 0.986988 0.991733 -2.97459e-06 -85.6668 0.0929949 31192.3 301.194 0.983519 0.319147 0.7356 0.735596 9.99958 2.98133e-06 1.19252e-05 0.130885 0.980987 0.931166 -0.0132931 4.89977e-06 0.501844 -1.89033e-20 6.96766e-24 -1.88963e-20 0.00139527 0.997818 8.59393e-05 0.152573 2.85183 0.00139527 0.997839 0.69792 0.0010487 0.00187985 0.000859393 0.455621 0.00187985 0.43737 0.000128256 1.02 0.887623 0.534697 0.285974 1.71665e-07 3.06041e-09 2388.2 3128.81 -0.0560777 0.48213 0.277571 0.254086 -0.593229 -0.169507 0.494971 -0.267992 -0.226988 1.613 1 0 297.017 0 2.08028 1.611 0.00029991 0.858735 0.651894 0.411558 0.408751 2.08051 130.881 83.7705 18.7122 60.794 0.00403149 0 -40 10
0.712 2.06322e-08 2.53891e-06 0.0933107 0.0933077 0.0120406 9.37826e-06 0.00115405 0.116638 0.000657455 0.117291 0.869937 101.851 0.24477 0.732755 4.1488 0.0552304 0.0391396 0.96086 0.0198432 0.00426699 0.019106 0.00410414 0.00515684 0.00589405 0.206273 0.235762 57.9833 -87.8952 126.201 15.9744 145.015 0.000141798 0.267117 192.897 0.310635 0.0673795 0.00409534 0.000561686 0.00138285 0.986988 0.991733 -2.9746e-06 -85.6667 0.092995 31192.3 301.198 0.983519 0.319147 0.735576 0.735572 9.99958 2.98133e-06 1.19252e-05 0.130887 0.980995 0.931169 -0.0132931 4.8998e-06 0.501851 -1.89041e-20 6.968e-24 -1.88971e-20 0.00139527 0.997818 8.59394e-05 0.152573 2.85184 0.00139527 0.997839 0.698025 0.00104872 0.00187985 0.000859394 0.455621 0.00187985 0.437379 0.000128259 1.02 0.887624 0.534696 0.285975 1.71666e-07 3.06044e-09 2388.18 3128.71 -0.0560711 0.48213 0.277571 0.254079 -0.59323 -0.169507 0.49499 -0.26799 -0.227008 1.614 1 0 297.024 0 2.08045 1.612 0.00029991 0.858691 0.651947 0.411342 0.408779 2.08068 130.89 83.7716 18.7123 60.7946 0.00403144 0 -40 10
0.713 2.06611e-08 2.53891e-06 0.093387 0.093384 0.0120406 9.39142e-06 0.00115405 0.116734 0.000657459 0.117387 0.869997 101.851 0.244763 0.732843 4.14897 0.0552374 0.0391412 0.960859 0.019843 0.00426715 0.0191058 0.00410427 0.00515703 0.00589424 0.206281 0.23577 57.9834 -87.8952 126.201 15.9743 145.015 0.000141793 0.267118 192.897 0.310635 0.0673794 0.00409534 0.000561686 0.00138285 0.986988 0.991733 -2.97461e-06 -85.6667 0.092995 31192.3 301.202 0.983519 0.319147 0.735552 0.735548 9.99958 2.98134e-06 1.19253e-05 0.130888 0.981003 0.931173 -0.0132931 4.89982e-06 0.501858 -1.89049e-20 6.96834e-24 -1.8898e-20 0.00139527 0.997818 8.59395e-05 0.152573 2.85184 0.00139527 0.997839 0.69813 0.00104874 0.00187985 0.000859395 0.45562 0.00187985 0.437388 0.000128262 1.02 0.887625 0.534696 0.285976 1.71666e-07 3.06046e-09 2388.17 3128.61 -0.0560647 0.48213 0.277571 0.254073 -0.593231 -0.169507 0.495008 -0.267988 -0.227029 1.615 1 0 297.031 0 2.08062 1.613 0.000299909 0.858647 0.652 0.411126 0.408807 2.08085 130.899 83.7728 18.7123 60.7951 0.00403139 0 -40 10
0.714 2.06901e-08 2.53891e-06 0.0934632 0.0934602 0.0120405 9.40457e-06 0.00115405 0.116829 0.000657462 0.117482 0.870057 101.851 0.244756 0.732932 4.14914 0.0552445 0.0391428 0.960857 0.0198428 0.00426731 0.0191056 0.00410441 0.00515723 0.00589444 0.206289 0.235777 57.9835 -87.8952 126.202 15.9743 145.015 0.000141789 0.267118 192.897 0.310635 0.0673794 0.00409535 0.000561687 0.00138286 0.986988 0.991733 -2.97463e-06 -85.6667 0.0929951 31192.3 301.207 0.983518 0.319147 0.735528 0.735524 9.99958 2.98134e-06 1.19253e-05 0.13089 0.981011 0.931176 -0.0132931 4.89985e-06 0.501864 -1.89057e-20 6.96869e-24 -1.88988e-20 0.00139527 0.997818 8.59396e-05 0.152573 2.85184 0.00139527 0.997838 0.698235 0.00104876 0.00187985 0.000859396 0.45562 0.00187985 0.437396 0.000128266 1.02 0.887626 0.534696 0.285978 1.71666e-07 3.06048e-09 2388.15 3128.5 -0.0560582 0.48213 0.27757 0.254066 -0.593232 -0.169507 0.495027 -0.267986 -0.227049 1.616 1 0 297.038 0 2.08078 1.614 0.000299909 0.858603 0.652052 0.41091 0.408835 2.08102 130.908 83.774 18.7124 60.7957 0.00403135 0 -40 10
0.715 2.0719e-08 2.53891e-06 0.0935394 0.0935364 0.0120405 9.41773e-06 0.00115405 0.116924 0.000657465 0.117577 0.870117 101.851 0.244748 0.733021 4.1493 0.0552515 0.0391444 0.960856 0.0198426 0.00426747 0.0191054 0.00410454 0.00515742 0.00589463 0.206297 0.235785 57.9835 -87.8952 126.202 15.9742 145.015 0.000141784 0.267118 192.897 0.310634 0.0673793 0.00409535 0.000561688 0.00138286 0.986988 0.991733 -2.97464e-06 -85.6667 0.0929952 31192.2 301.211 0.983518 0.319147 0.735505 0.7355 9.99958 2.98135e-06 1.19253e-05 0.130892 0.981018 0.931179 -0.0132931 4.89988e-06 0.501871 -1.89066e-20 6.96903e-24 -1.88996e-20 0.00139527 0.997818 8.59396e-05 0.152573 2.85184 0.00139527 0.997838 0.69834 0.00104878 0.00187985 0.000859396 0.45562 0.00187985 0.437405 0.000128269 1.02 0.887627 0.534695 0.285979 1.71666e-07 3.0605e-09 2388.13 3128.4 -0.0560518 0.48213 0.27757 0.25406 -0.593233 -0.169507 0.495045 -0.267984 -0.22707 1.617 1 0 297.044 0 2.08095 1.615 0.000299909 0.858559 0.652105 0.410696 0.408864 2.08119 130.917 83.7752 18.7125 60.7963 0.0040313 0 -40 10
0.716 2.07479e-08 2.53891e-06 0.0936155 0.0936125 0.0120405 9.43089e-06 0.00115405 0.117019 0.000657468 0.117672 0.870177 101.851 0.244741 0.733109 4.14947 0.0552586 0.039146 0.960854 0.0198424 0.00426763 0.0191052 0.00410467 0.00515762 0.00589483 0.206305 0.235793 57.9836 -87.8952 126.203 15.9742 145.015 0.000141779 0.267118 192.897 0.310634 0.0673793 0.00409535 0.000561688 0.00138286 0.986988 0.991733 -2.97466e-06 -85.6667 0.0929953 31192.2 301.215 0.983518 0.319147 0.735481 0.735477 9.99958 2.98135e-06 1.19253e-05 0.130893 0.981026 0.931183 -0.0132931 4.89991e-06 0.501878 -1.89074e-20 6.96938e-24 -1.89004e-20 0.00139528 0.997818 8.59397e-05 0.152573 2.85184 0.00139528 0.997838 0.698445 0.0010488 0.00187985 0.000859397 0.45562 0.00187985 0.437414 0.000128273 1.02 0.887628 0.534695 0.285981 1.71667e-07 3.06052e-09 2388.11 3128.3 -0.0560455 0.48213 0.27757 0.254054 -0.593235 -0.169507 0.495063 -0.267982 -0.22709 1.618 1 0 297.051 0 2.08112 1.616 0.000299908 0.858516 0.652157 0.410481 0.408892 2.08135 130.926 83.7763 18.7125 60.7968 0.00403125 0 -40 10
0.717 2.07769e-08 2.53891e-06 0.0936915 0.0936885 0.0120405 9.44404e-06 0.00115405 0.117114 0.000657471 0.117767 0.870237 101.85 0.244734 0.733198 4.14964 0.0552656 0.0391475 0.960852 0.0198422 0.00426779 0.019105 0.0041048 0.00515781 0.00589502 0.206313 0.235801 57.9837 -87.8952 126.203 15.9742 145.015 0.000141775 0.267118 192.896 0.310633 0.0673792 0.00409536 0.000561689 0.00138286 0.986988 0.991733 -2.97467e-06 -85.6667 0.0929954 31192.2 301.22 0.983518 0.319147 0.735458 0.735453 9.99958 2.98136e-06 1.19253e-05 0.130895 0.981034 0.931186 -0.0132931 4.89994e-06 0.501884 -1.89082e-20 6.96972e-24 -1.89012e-20 0.00139528 0.997818 8.59398e-05 0.152574 2.85184 0.00139528 0.997838 0.69855 0.00104882 0.00187986 0.000859398 0.45562 0.00187985 0.437422 0.000128276 1.02 0.887629 0.534695 0.285982 1.71667e-07 3.06054e-09 2388.1 3128.2 -0.0560391 0.48213 0.27757 0.254047 -0.593236 -0.169507 0.495081 -0.26798 -0.22711 1.619 1 0 297.057 0 2.08129 1.617 0.000299908 0.858473 0.65221 0.410267 0.40892 2.08152 130.935 83.7775 18.7126 60.7974 0.0040312 0 -40 10
0.718 2.08058e-08 2.53891e-06 0.0937675 0.0937645 0.0120405 9.4572e-06 0.00115405 0.117209 0.000657474 0.117862 0.870297 101.85 0.244727 0.733287 4.14981 0.0552727 0.0391491 0.960851 0.019842 0.00426795 0.0191048 0.00410494 0.00515801 0.00589522 0.20632 0.235809 57.9837 -87.8953 126.204 15.9741 145.015 0.00014177 0.267119 192.896 0.310633 0.0673792 0.00409536 0.000561689 0.00138286 0.986988 0.991733 -2.97469e-06 -85.6667 0.0929955 31192.2 301.224 0.983518 0.319147 0.735434 0.73543 9.99958 2.98136e-06 1.19253e-05 0.130897 0.981042 0.931189 -0.0132931 4.89997e-06 0.501891 -1.8909e-20 6.97006e-24 -1.89021e-20 0.00139528 0.997818 8.59399e-05 0.152574 2.85184 0.00139528 0.997838 0.698655 0.00104884 0.00187986 0.000859399 0.455619 0.00187986 0.437431 0.000128279 1.02 0.88763 0.534694 0.285984 1.71667e-07 3.06057e-09 2388.08 3128.1 -0.0560329 0.48213 0.277569 0.254041 -0.593237 -0.169507 0.495099 -0.267978 -0.22713 1.62 1 0 297.064 0 2.08145 1.618 0.000299908 0.85843 0.652262 0.410054 0.408948 2.08169 130.944 83.7786 18.7127 60.7979 0.00403115 0 -40 10
0.719 2.08348e-08 2.53891e-06 0.0938434 0.0938404 0.0120405 9.47035e-06 0.00115405 0.117304 0.000657477 0.117957 0.870357 101.85 0.24472 0.733376 4.14998 0.0552798 0.0391507 0.960849 0.0198418 0.00426811 0.0191046 0.00410507 0.00515821 0.00589541 0.206328 0.235816 57.9838 -87.8953 126.204 15.9741 145.015 0.000141766 0.267119 192.896 0.310632 0.0673791 0.00409536 0.00056169 0.00138287 0.986988 0.991733 -2.9747e-06 -85.6667 0.0929955 31192.1 301.228 0.983518 0.319147 0.735411 0.735407 9.99958 2.98137e-06 1.19254e-05 0.130898 0.981049 0.931192 -0.0132931 4.9e-06 0.501898 -1.89099e-20 6.97041e-24 -1.89029e-20 0.00139528 0.997818 8.594e-05 0.152574 2.85184 0.00139528 0.997838 0.69876 0.00104886 0.00187986 0.0008594 0.455619 0.00187986 0.43744 0.000128283 1.02 0.887631 0.534694 0.285985 1.71668e-07 3.06059e-09 2388.06 3128 -0.0560266 0.48213 0.277569 0.254035 -0.593238 -0.169508 0.495117 -0.267976 -0.22715 1.621 1 0 297.071 0 2.08162 1.619 0.000299907 0.858387 0.652315 0.409841 0.408976 2.08186 130.953 83.7798 18.7127 60.7985 0.00403111 0 -40 10
0.72 2.08637e-08 2.53891e-06 0.0939193 0.0939163 0.0120405 9.48351e-06 0.00115405 0.117399 0.00065748 0.118052 0.870418 101.85 0.244713 0.733465 4.15015 0.0552869 0.0391523 0.960848 0.0198416 0.00426827 0.0191044 0.00410521 0.00515841 0.00589561 0.206336 0.235824 57.9838 -87.8953 126.204 15.9741 145.015 0.000141762 0.267119 192.896 0.310632 0.0673791 0.00409536 0.000561691 0.00138287 0.986988 0.991733 -2.97471e-06 -85.6667 0.0929956 31192.1 301.233 0.983518 0.319147 0.735388 0.735384 9.99958 2.98137e-06 1.19254e-05 0.1309 0.981057 0.931196 -0.0132931 4.90002e-06 0.501904 -1.89107e-20 6.97075e-24 -1.89037e-20 0.00139528 0.997818 8.594e-05 0.152574 2.85184 0.00139528 0.997838 0.698865 0.00104888 0.00187986 0.0008594 0.455619 0.00187986 0.437448 0.000128286 1.02 0.887632 0.534694 0.285987 1.71668e-07 3.06061e-09 2388.05 3127.9 -0.0560204 0.48213 0.277569 0.254029 -0.593239 -0.169508 0.495135 -0.267974 -0.22717 1.622 1 0 297.077 0 2.08179 1.62 0.000299907 0.858345 0.652367 0.409629 0.409004 2.08202 130.962 83.7809 18.7128 60.799 0.00403106 0 -40 10
0.721 2.08927e-08 2.53892e-06 0.0939951 0.0939921 0.0120405 9.49667e-06 0.00115405 0.117494 0.000657483 0.118147 0.870478 101.85 0.244706 0.733555 4.15032 0.055294 0.0391539 0.960846 0.0198414 0.00426843 0.0191042 0.00410534 0.00515861 0.00589581 0.206344 0.235832 57.9839 -87.8953 126.205 15.974 145.015 0.000141757 0.267119 192.896 0.310632 0.067379 0.00409537 0.000561691 0.00138287 0.986988 0.991733 -2.97473e-06 -85.6667 0.0929957 31192.1 301.237 0.983518 0.319147 0.735365 0.735361 9.99958 2.98138e-06 1.19254e-05 0.130901 0.981065 0.931199 -0.0132931 4.90005e-06 0.501911 -1.89115e-20 6.9711e-24 -1.89045e-20 0.00139528 0.997818 8.59401e-05 0.152574 2.85184 0.00139528 0.997837 0.69897 0.0010489 0.00187986 0.000859401 0.455619 0.00187986 0.437457 0.000128289 1.02 0.887633 0.534694 0.285988 1.71668e-07 3.06063e-09 2388.03 3127.8 -0.0560142 0.48213 0.277568 0.254022 -0.59324 -0.169508 0.495152 -0.267972 -0.22719 1.623 1 0 297.084 0 2.08196 1.621 0.000299907 0.858302 0.65242 0.409417 0.409032 2.08219 130.971 83.782 18.7129 60.7996 0.00403101 0 -40 10
0.722 2.09216e-08 2.53892e-06 0.0940708 0.0940678 0.0120404 9.50982e-06 0.00115405 0.117589 0.000657486 0.118241 0.870538 101.85 0.244699 0.733644 4.15049 0.0553011 0.0391555 0.960844 0.0198412 0.00426859 0.019104 0.00410548 0.0051588 0.005896 0.206352 0.23584 57.984 -87.8953 126.205 15.974 145.015 0.000141753 0.267119 192.896 0.310631 0.067379 0.00409537 0.000561692 0.00138287 0.986988 0.991733 -2.97474e-06 -85.6667 0.0929958 31192.1 301.241 0.983518 0.319147 0.735342 0.735338 9.99958 2.98138e-06 1.19254e-05 0.130903 0.981073 0.931202 -0.0132931 4.90008e-06 0.501918 -1.89123e-20 6.97144e-24 -1.89054e-20 0.00139528 0.997818 8.59402e-05 0.152574 2.85184 0.00139528 0.997837 0.699074 0.00104892 0.00187986 0.000859402 0.455618 0.00187986 0.437466 0.000128293 1.02 0.887635 0.534693 0.28599 1.71668e-07 3.06065e-09 2388.01 3127.71 -0.056008 0.482131 0.277568 0.254016 -0.593241 -0.169508 0.49517 -0.26797 -0.227209 1.624 1 0 297.09 0 2.08212 1.622 0.000299906 0.85826 0.652472 0.409206 0.40906 2.08236 130.98 83.7832 18.7129 60.8001 0.00403097 0 -40 10
0.723 2.09506e-08 2.53892e-06 0.0941465 0.0941435 0.0120404 9.52298e-06 0.00115405 0.117683 0.000657489 0.118336 0.870598 101.849 0.244692 0.733733 4.15066 0.0553082 0.0391571 0.960843 0.019841 0.00426875 0.0191038 0.00410561 0.005159 0.0058962 0.20636 0.235848 57.984 -87.8953 126.206 15.9739 145.015 0.000141748 0.267119 192.895 0.310631 0.0673789 0.00409537 0.000561693 0.00138287 0.986988 0.991733 -2.97476e-06 -85.6666 0.0929959 31192.1 301.246 0.983518 0.319147 0.735319 0.735315 9.99958 2.98139e-06 1.19254e-05 0.130905 0.98108 0.931205 -0.0132931 4.90011e-06 0.501925 -1.89132e-20 6.97179e-24 -1.89062e-20 0.00139528 0.997818 8.59403e-05 0.152574 2.85184 0.00139528 0.997837 0.699179 0.00104894 0.00187986 0.000859403 0.455618 0.00187986 0.437474 0.000128296 1.02 0.887636 0.534693 0.285991 1.71669e-07 3.06068e-09 2388 3127.61 -0.0560019 0.482131 0.277568 0.25401 -0.593243 -0.169508 0.495187 -0.267967 -0.227229 1.625 1 0 297.096 0 2.08229 1.623 0.000299906 0.858218 0.652525 0.408995 0.409088 2.08253 130.989 83.7843 18.713 60.8007 0.00403092 0 -40 10
0.724 2.09795e-08 2.53892e-06 0.0942221 0.0942191 0.0120404 9.53613e-06 0.00115405 0.117778 0.000657492 0.118431 0.870659 101.849 0.244685 0.733823 4.15083 0.0553153 0.0391588 0.960841 0.0198408 0.00426891 0.0191036 0.00410575 0.0051592 0.0058964 0.206368 0.235856 57.9841 -87.8953 126.206 15.9739 145.015 0.000141744 0.26712 192.895 0.31063 0.0673789 0.00409538 0.000561693 0.00138288 0.986988 0.991733 -2.97477e-06 -85.6666 0.092996 31192 301.25 0.983518 0.319147 0.735297 0.735292 9.99958 2.98139e-06 1.19255e-05 0.130906 0.981088 0.931208 -0.0132931 4.90014e-06 0.501931 -1.8914e-20 6.97213e-24 -1.8907e-20 0.00139528 0.997818 8.59403e-05 0.152575 2.85185 0.00139528 0.997837 0.699284 0.00104896 0.00187987 0.000859403 0.455618 0.00187986 0.437483 0.000128299 1.02 0.887637 0.534693 0.285993 1.71669e-07 3.0607e-09 2387.98 3127.51 -0.0559959 0.482131 0.277568 0.254004 -0.593244 -0.169508 0.495204 -0.267965 -0.227248 1.626 1 0 297.103 0 2.08246 1.624 0.000299906 0.858177 0.652577 0.408785 0.409117 2.08269 130.998 83.7854 18.7131 60.8012 0.00403087 0 -40 10
0.725 2.10084e-08 2.53892e-06 0.0942977 0.0942947 0.0120404 9.54929e-06 0.00115405 0.117872 0.000657494 0.118525 0.870719 101.849 0.244678 0.733912 4.151 0.0553224 0.0391604 0.96084 0.0198406 0.00426908 0.0191034 0.00410588 0.0051594 0.0058966 0.206376 0.235864 57.9842 -87.8953 126.207 15.9739 145.015 0.00014174 0.26712 192.895 0.31063 0.0673788 0.00409538 0.000561694 0.00138288 0.986988 0.991733 -2.97479e-06 -85.6666 0.092996 31192 301.255 0.983518 0.319147 0.735274 0.73527 9.99958 2.9814e-06 1.19255e-05 0.130908 0.981095 0.931212 -0.0132931 4.90017e-06 0.501938 -1.89148e-20 6.97248e-24 -1.89078e-20 0.00139529 0.997818 8.59404e-05 0.152575 2.85185 0.00139529 0.997837 0.699389 0.00104898 0.00187987 0.000859404 0.455618 0.00187987 0.437491 0.000128303 1.02 0.887638 0.534692 0.285994 1.71669e-07 3.06072e-09 2387.96 3127.42 -0.0559898 0.482131 0.277567 0.253998 -0.593245 -0.169508 0.495222 -0.267963 -0.227267 1.627 1 0 297.109 0 2.08263 1.625 0.000299905 0.858135 0.652629 0.408575 0.409145 2.08286 131.007 83.7865 18.7131 60.8017 0.00403083 0 -40 10
0.726 2.10374e-08 2.53892e-06 0.0943731 0.0943702 0.0120404 9.56244e-06 0.00115405 0.117966 0.000657497 0.118619 0.87078 101.849 0.24467 0.734002 4.15117 0.0553296 0.039162 0.960838 0.0198404 0.00426924 0.0191032 0.00410602 0.0051596 0.0058968 0.206384 0.235872 57.9842 -87.8953 126.207 15.9738 145.015 0.000141735 0.26712 192.895 0.31063 0.0673788 0.00409538 0.000561695 0.00138288 0.986988 0.991733 -2.9748e-06 -85.6666 0.0929961 31192 301.259 0.983518 0.319147 0.735252 0.735247 9.99958 2.9814e-06 1.19255e-05 0.13091 0.981103 0.931215 -0.0132931 4.9002e-06 0.501945 -1.89156e-20 6.97283e-24 -1.89087e-20 0.00139529 0.997818 8.59405e-05 0.152575 2.85185 0.00139529 0.997837 0.699493 0.001049 0.00187987 0.000859405 0.455618 0.00187987 0.4375 0.000128306 1.02 0.887639 0.534692 0.285996 1.71669e-07 3.06074e-09 2387.95 3127.32 -0.0559838 0.482131 0.277567 0.253992 -0.593246 -0.169508 0.495239 -0.267961 -0.227286 1.628 1 0 297.115 0 2.08279 1.626 0.000299905 0.858094 0.652682 0.408366 0.409173 2.08303 131.016 83.7876 18.7132 60.8023 0.00403078 0 -40 10
0.727 2.10663e-08 2.53892e-06 0.0944486 0.0944456 0.0120404 9.5756e-06 0.00115405 0.118061 0.0006575 0.118714 0.87084 101.849 0.244663 0.734092 4.15134 0.0553367 0.0391636 0.960836 0.0198402 0.0042694 0.019103 0.00410615 0.0051598 0.00589699 0.206392 0.23588 57.9843 -87.8953 126.207 15.9738 145.015 0.000141731 0.26712 192.895 0.310629 0.0673787 0.00409538 0.000561695 0.00138288 0.986987 0.991733 -2.97481e-06 -85.6666 0.0929962 31192 301.263 0.983518 0.319147 0.735229 0.735225 9.99958 2.98141e-06 1.19255e-05 0.130911 0.981111 0.931218 -0.0132931 4.90022e-06 0.501952 -1.89165e-20 6.97317e-24 -1.89095e-20 0.00139529 0.997818 8.59406e-05 0.152575 2.85185 0.00139529 0.997837 0.699598 0.00104902 0.00187987 0.000859406 0.455617 0.00187987 0.437509 0.00012831 1.02 0.88764 0.534692 0.285997 1.7167e-07 3.06076e-09 2387.93 3127.22 -0.0559778 0.482131 0.277567 0.253986 -0.593247 -0.169508 0.495256 -0.267959 -0.227306 1.629 1 0 297.122 0 2.08296 1.627 0.000299905 0.858053 0.652734 0.408157 0.409201 2.08319 131.025 83.7887 18.7133 60.8028 0.00403074 0 -40 10
0.728 2.10953e-08 2.53892e-06 0.0945239 0.094521 0.0120404 9.58876e-06 0.00115405 0.118155 0.000657503 0.118808 0.870901 101.848 0.244656 0.734182 4.15152 0.0553439 0.0391652 0.960835 0.01984 0.00426957 0.0191028 0.00410629 0.00516 0.00589719 0.2064 0.235888 57.9844 -87.8953 126.208 15.9738 145.015 0.000141727 0.26712 192.895 0.310629 0.0673787 0.00409539 0.000561696 0.00138288 0.986987 0.991733 -2.97483e-06 -85.6666 0.0929963 31192 301.268 0.983518 0.319147 0.735207 0.735203 9.99958 2.98141e-06 1.19255e-05 0.130913 0.981118 0.931221 -0.0132931 4.90025e-06 0.501959 -1.89173e-20 6.97352e-24 -1.89103e-20 0.00139529 0.997818 8.59406e-05 0.152575 2.85185 0.00139529 0.997837 0.699702 0.00104904 0.00187987 0.000859406 0.455617 0.00187987 0.437517 0.000128313 1.02 0.887641 0.534692 0.285998 1.7167e-07 3.06079e-09 2387.91 3127.13 -0.0559719 0.482131 0.277566 0.25398 -0.593248 -0.169508 0.495273 -0.267957 -0.227324 1.63 1 0 297.128 0 2.08313 1.628 0.000299904 0.858012 0.652786 0.407949 0.409229 2.08336 131.033 83.7898 18.7133 60.8033 0.00403069 0 -40 10
0.729 2.11242e-08 2.53892e-06 0.0945993 0.0945963 0.0120403 9.60191e-06 0.00115405 0.118249 0.000657506 0.118902 0.870962 101.848 0.244649 0.734271 4.15169 0.055351 0.0391669 0.960833 0.0198398 0.00426973 0.0191026 0.00410643 0.0051602 0.00589739 0.206408 0.235896 57.9844 -87.8953 126.208 15.9737 145.015 0.000141722 0.267121 192.895 0.310628 0.0673786 0.00409539 0.000561696 0.00138289 0.986987 0.991733 -2.97484e-06 -85.6666 0.0929964 31191.9 301.272 0.983518 0.319147 0.735185 0.735181 9.99958 2.98141e-06 1.19256e-05 0.130915 0.981126 0.931224 -0.0132931 4.90028e-06 0.501966 -1.89181e-20 6.97386e-24 -1.89111e-20 0.00139529 0.997818 8.59407e-05 0.152575 2.85185 0.00139529 0.997836 0.699807 0.00104906 0.00187987 0.000859407 0.455617 0.00187987 0.437526 0.000128316 1.02 0.887642 0.534691 0.286 1.7167e-07 3.06081e-09 2387.9 3127.03 -0.055966 0.482131 0.277566 0.253974 -0.593249 -0.169508 0.495289 -0.267955 -0.227343 1.631 1 0 297.134 0 2.08329 1.629 0.000299904 0.857971 0.652839 0.407741 0.409257 2.08353 131.042 83.7909 18.7134 60.8039 0.00403065 0 -40 10
0.73 2.11531e-08 2.53892e-06 0.0946745 0.0946716 0.0120403 9.61507e-06 0.00115405 0.118343 0.000657509 0.118996 0.871022 101.848 0.244642 0.734361 4.15186 0.0553582 0.0391685 0.960831 0.0198396 0.00426989 0.0191024 0.00410656 0.00516041 0.00589759 0.206416 0.235904 57.9845 -87.8953 126.209 15.9737 145.015 0.000141718 0.267121 192.894 0.310628 0.0673786 0.00409539 0.000561697 0.00138289 0.986987 0.991733 -2.97486e-06 -85.6666 0.0929965 31191.9 301.277 0.983518 0.319147 0.735163 0.735159 9.99958 2.98142e-06 1.19256e-05 0.130916 0.981133 0.931227 -0.0132931 4.90031e-06 0.501972 -1.89189e-20 6.97421e-24 -1.8912e-20 0.00139529 0.997818 8.59408e-05 0.152575 2.85185 0.00139529 0.997836 0.699911 0.00104908 0.00187987 0.000859408 0.455617 0.00187987 0.437535 0.00012832 1.02 0.887643 0.534691 0.286001 1.7167e-07 3.06083e-09 2387.88 3126.94 -0.0559601 0.482131 0.277566 0.253968 -0.59325 -0.169508 0.495306 -0.267953 -0.227362 1.632 1 0 297.14 0 2.08346 1.63 0.000299904 0.857931 0.652891 0.407534 0.409285 2.08369 131.051 83.792 18.7134 60.8044 0.0040306 0 -40 10
0.731 2.11821e-08 2.53892e-06 0.0947497 0.0947468 0.0120403 9.62822e-06 0.00115405 0.118437 0.000657512 0.11909 0.871083 101.848 0.244635 0.734451 4.15203 0.0553653 0.0391701 0.96083 0.0198394 0.00427006 0.0191022 0.0041067 0.00516061 0.0058978 0.206424 0.235912 57.9845 -87.8953 126.209 15.9736 145.015 0.000141714 0.267121 192.894 0.310628 0.0673785 0.0040954 0.000561698 0.00138289 0.986987 0.991733 -2.97487e-06 -85.6666 0.0929965 31191.9 301.281 0.983518 0.319147 0.735141 0.735137 9.99958 2.98142e-06 1.19256e-05 0.130918 0.981141 0.93123 -0.0132931 4.90034e-06 0.501979 -1.89198e-20 6.97456e-24 -1.89128e-20 0.00139529 0.997818 8.59409e-05 0.152576 2.85185 0.00139529 0.997836 0.700016 0.00104909 0.00187988 0.000859409 0.455617 0.00187987 0.437543 0.000128323 1.02 0.887644 0.534691 0.286003 1.71671e-07 3.06085e-09 2387.86 3126.85 -0.0559543 0.482131 0.277566 0.253962 -0.593251 -0.169508 0.495323 -0.267951 -0.227381 1.633 1 0 297.146 0 2.08363 1.631 0.000299903 0.857891 0.652943 0.407327 0.409313 2.08386 131.06 83.7931 18.7135 60.8049 0.00403056 0 -40 10
0.732 2.1211e-08 2.53892e-06 0.0948248 0.0948219 0.0120403 9.64138e-06 0.00115405 0.118531 0.000657515 0.119184 0.871144 101.848 0.244628 0.734542 4.15221 0.0553725 0.0391718 0.960828 0.0198392 0.00427022 0.019102 0.00410684 0.00516081 0.005898 0.206432 0.23592 57.9846 -87.8953 126.209 15.9736 145.015 0.00014171 0.267121 192.894 0.310627 0.0673785 0.0040954 0.000561698 0.00138289 0.986987 0.991733 -2.97489e-06 -85.6666 0.0929966 31191.9 301.286 0.983518 0.319147 0.735119 0.735115 9.99958 2.98143e-06 1.19256e-05 0.13092 0.981148 0.931233 -0.0132931 4.90037e-06 0.501986 -1.89206e-20 6.9749e-24 -1.89136e-20 0.00139529 0.997818 8.59409e-05 0.152576 2.85185 0.00139529 0.997836 0.70012 0.00104911 0.00187988 0.000859409 0.455616 0.00187988 0.437552 0.000128326 1.02 0.887645 0.53469 0.286004 1.71671e-07 3.06088e-09 2387.85 3126.75 -0.0559485 0.482131 0.277565 0.253956 -0.593253 -0.169508 0.495339 -0.267949 -0.227399 1.634 1 0 297.152 0 2.0838 1.632 0.000299903 0.857851 0.652995 0.407121 0.409341 2.08403 131.069 83.7942 18.7136 60.8054 0.00403051 0 -40 10
0.733 2.124e-08 2.53892e-06 0.0948999 0.094897 0.0120403 9.65453e-06 0.00115405 0.118625 0.000657518 0.119278 0.871205 101.848 0.24462 0.734632 4.15238 0.0553797 0.0391734 0.960827 0.019839 0.00427039 0.0191018 0.00410697 0.00516101 0.0058982 0.206441 0.235928 57.9847 -87.8953 126.21 15.9736 145.015 0.000141706 0.267121 192.894 0.310627 0.0673784 0.0040954 0.000561699 0.00138289 0.986987 0.991733 -2.9749e-06 -85.6666 0.0929967 31191.8 301.29 0.983518 0.319147 0.735098 0.735093 9.99958 2.98143e-06 1.19256e-05 0.130922 0.981155 0.931237 -0.0132931 4.9004e-06 0.501993 -1.89214e-20 6.97525e-24 -1.89144e-20 0.00139529 0.997818 8.5941e-05 0.152576 2.85185 0.00139529 0.997836 0.700225 0.00104913 0.00187988 0.00085941 0.455616 0.00187988 0.43756 0.00012833 1.02 0.887646 0.53469 0.286006 1.71671e-07 3.0609e-09 2387.83 3126.66 -0.0559427 0.482131 0.277565 0.25395 -0.593254 -0.169508 0.495356 -0.267947 -0.227418 1.635 1 0 297.159 0 2.08396 1.633 0.000299903 0.857811 0.653047 0.406915 0.409368 2.08419 131.078 83.7952 18.7136 60.8059 0.00403047 0 -40 10
0.734 2.12689e-08 2.53892e-06 0.0949749 0.094972 0.0120403 9.66769e-06 0.00115405 0.118719 0.000657521 0.119372 0.871266 101.847 0.244613 0.734722 4.15256 0.0553869 0.0391751 0.960825 0.0198388 0.00427055 0.0191016 0.00410711 0.00516122 0.0058984 0.206449 0.235936 57.9847 -87.8953 126.21 15.9735 145.015 0.000141701 0.267121 192.894 0.310626 0.0673784 0.00409541 0.0005617 0.0013829 0.986987 0.991733 -2.97491e-06 -85.6665 0.0929968 31191.8 301.295 0.983518 0.319147 0.735076 0.735072 9.99958 2.98144e-06 1.19256e-05 0.130923 0.981163 0.93124 -0.0132931 4.90043e-06 0.502 -1.89222e-20 6.9756e-24 -1.89153e-20 0.0013953 0.997818 8.59411e-05 0.152576 2.85185 0.0013953 0.997836 0.700329 0.00104915 0.00187988 0.000859411 0.455616 0.00187988 0.437569 0.000128333 1.02 0.887647 0.53469 0.286007 1.71671e-07 3.06092e-09 2387.81 3126.57 -0.055937 0.482131 0.277565 0.253945 -0.593255 -0.169509 0.495372 -0.267945 -0.227436 1.636 1 0 297.165 0 2.08413 1.634 0.000299902 0.857771 0.653099 0.406709 0.409396 2.08436 131.087 83.7963 18.7137 60.8065 0.00403043 0 -40 10
0.735 2.12979e-08 2.53892e-06 0.0950499 0.095047 0.0120403 9.68084e-06 0.00115405 0.118812 0.000657524 0.119465 0.871326 101.847 0.244606 0.734812 4.15273 0.0553941 0.0391767 0.960823 0.0198386 0.00427072 0.0191014 0.00410725 0.00516142 0.0058986 0.206457 0.235944 57.9848 -87.8953 126.211 15.9735 145.015 0.000141697 0.267122 192.894 0.310626 0.0673783 0.00409541 0.0005617 0.0013829 0.986987 0.991733 -2.97493e-06 -85.6665 0.0929969 31191.8 301.299 0.983518 0.319147 0.735055 0.73505 9.99958 2.98144e-06 1.19257e-05 0.130925 0.98117 0.931243 -0.0132931 4.90045e-06 0.502007 -1.89231e-20 6.97594e-24 -1.89161e-20 0.0013953 0.997818 8.59412e-05 0.152576 2.85186 0.0013953 0.997836 0.700433 0.00104917 0.00187988 0.000859412 0.455616 0.00187988 0.437578 0.000128336 1.02 0.887648 0.534689 0.286009 1.71672e-07 3.06094e-09 2387.8 3126.47 -0.0559313 0.482131 0.277564 0.253939 -0.593256 -0.169509 0.495388 -0.267943 -0.227454 1.637 1 0 297.171 0 2.08429 1.635 0.000299902 0.857732 0.653152 0.406505 0.409424 2.08453 131.096 83.7974 18.7138 60.807 0.00403038 0 -40 10
0.736 2.13268e-08 2.53892e-06 0.0951247 0.0951219 0.0120403 9.694e-06 0.00115406 0.118906 0.000657526 0.119559 0.871387 101.847 0.244599 0.734903 4.15291 0.0554012 0.0391784 0.960822 0.0198384 0.00427089 0.0191012 0.00410739 0.00516163 0.00589881 0.206465 0.235952 57.9849 -87.8953 126.211 15.9734 145.015 0.000141693 0.267122 192.893 0.310626 0.0673783 0.00409541 0.000561701 0.0013829 0.986987 0.991733 -2.97494e-06 -85.6665 0.092997 31191.8 301.304 0.983518 0.319147 0.735033 0.735029 9.99958 2.98145e-06 1.19257e-05 0.130927 0.981178 0.931246 -0.0132931 4.90048e-06 0.502014 -1.89239e-20 6.97629e-24 -1.89169e-20 0.0013953 0.997818 8.59413e-05 0.152576 2.85186 0.0013953 0.997836 0.700537 0.00104919 0.00187988 0.000859413 0.455615 0.00187988 0.437586 0.00012834 1.02 0.887649 0.534689 0.28601 1.71672e-07 3.06096e-09 2387.78 3126.38 -0.0559256 0.482132 0.277564 0.253933 -0.593257 -0.169509 0.495404 -0.267941 -0.227472 1.638 1 0 297.176 0 2.08446 1.636 0.000299902 0.857693 0.653204 0.4063 0.409452 2.08469 131.105 83.7984 18.7138 60.8075 0.00403034 0 -40 10
0.737 2.13557e-08 2.53892e-06 0.0951996 0.0951967 0.0120402 9.70715e-06 0.00115406 0.118999 0.000657529 0.119652 0.871448 101.847 0.244592 0.734993 4.15308 0.0554085 0.03918 0.96082 0.0198382 0.00427105 0.019101 0.00410753 0.00516183 0.00589901 0.206473 0.23596 57.9849 -87.8953 126.211 15.9734 145.015 0.000141689 0.267122 192.893 0.310625 0.0673782 0.00409541 0.000561702 0.0013829 0.986987 0.991733 -2.97496e-06 -85.6665 0.092997 31191.8 301.308 0.983518 0.319147 0.735012 0.735008 9.99958 2.98145e-06 1.19257e-05 0.130928 0.981185 0.931249 -0.0132931 4.90051e-06 0.502021 -1.89247e-20 6.97664e-24 -1.89177e-20 0.0013953 0.997818 8.59413e-05 0.152576 2.85186 0.0013953 0.997835 0.700642 0.00104921 0.00187988 0.000859413 0.455615 0.00187988 0.437595 0.000128343 1.02 0.88765 0.534689 0.286012 1.71672e-07 3.06099e-09 2387.76 3126.29 -0.05592 0.482132 0.277564 0.253927 -0.593258 -0.169509 0.49542 -0.267939 -0.227491 1.639 1 0 297.182 0 2.08463 1.637 0.000299901 0.857654 0.653256 0.406096 0.40948 2.08486 131.114 83.7995 18.7139 60.808 0.00403029 0 -40 10
0.738 2.13847e-08 2.53892e-06 0.0952743 0.0952715 0.0120402 9.72031e-06 0.00115406 0.119093 0.000657532 0.119746 0.87151 101.847 0.244584 0.735084 4.15326 0.0554157 0.0391817 0.960818 0.019838 0.00427122 0.0191008 0.00410767 0.00516204 0.00589921 0.206481 0.235969 57.985 -87.8953 126.212 15.9734 145.015 0.000141685 0.267122 192.893 0.310625 0.0673782 0.00409542 0.000561702 0.0013829 0.986987 0.991733 -2.97497e-06 -85.6665 0.0929971 31191.7 301.313 0.983518 0.319147 0.734991 0.734986 9.99958 2.98146e-06 1.19257e-05 0.13093 0.981192 0.931252 -0.0132931 4.90054e-06 0.502028 -1.89256e-20 6.97698e-24 -1.89186e-20 0.0013953 0.997818 8.59414e-05 0.152577 2.85186 0.0013953 0.997835 0.700746 0.00104923 0.00187989 0.000859414 0.455615 0.00187988 0.437603 0.000128346 1.02 0.887652 0.534689 0.286013 1.71672e-07 3.06101e-09 2387.75 3126.2 -0.0559144 0.482132 0.277564 0.253922 -0.593259 -0.169509 0.495436 -0.267936 -0.227508 1.64 1 0 297.188 0 2.08479 1.638 0.000299901 0.857615 0.653308 0.405893 0.409508 2.08503 131.123 83.8005 18.7139 60.8085 0.00403025 0 -40 10
0.739 2.14136e-08 2.53892e-06 0.095349 0.0953462 0.0120402 9.73346e-06 0.00115406 0.119186 0.000657535 0.119839 0.871571 101.847 0.244577 0.735175 4.15344 0.0554229 0.0391834 0.960817 0.0198378 0.00427139 0.0191006 0.00410781 0.00516224 0.00589942 0.20649 0.235977 57.985 -87.8953 126.212 15.9733 145.015 0.000141681 0.267122 192.893 0.310624 0.0673781 0.00409542 0.000561703 0.00138291 0.986987 0.991733 -2.97499e-06 -85.6665 0.0929972 31191.7 301.317 0.983518 0.319147 0.73497 0.734965 9.99958 2.98146e-06 1.19257e-05 0.130932 0.981199 0.931255 -0.0132931 4.90057e-06 0.502035 -1.89264e-20 6.97733e-24 -1.89194e-20 0.0013953 0.997818 8.59415e-05 0.152577 2.85186 0.0013953 0.997835 0.70085 0.00104925 0.00187989 0.000859415 0.455615 0.00187989 0.437612 0.00012835 1.02 0.887653 0.534688 0.286015 1.71673e-07 3.06103e-09 2387.73 3126.11 -0.0559088 0.482132 0.277563 0.253916 -0.59326 -0.169509 0.495452 -0.267934 -0.227526 1.641 1 0 297.194 0 2.08496 1.639 0.000299901 0.857576 0.65336 0.40569 0.409536 2.08519 131.132 83.8016 18.714 60.809 0.00403021 0 -40 10
0.74 2.14426e-08 2.53892e-06 0.0954237 0.0954209 0.0120402 9.74662e-06 0.00115406 0.11928 0.000657538 0.119933 0.871632 101.846 0.24457 0.735266 4.15361 0.0554301 0.039185 0.960815 0.0198376 0.00427155 0.0191004 0.00410795 0.00516245 0.00589962 0.206498 0.235985 57.9851 -87.8953 126.212 15.9733 145.015 0.000141677 0.267123 192.893 0.310624 0.0673781 0.00409542 0.000561703 0.00138291 0.986987 0.991733 -2.975e-06 -85.6665 0.0929973 31191.7 301.322 0.983518 0.319147 0.734949 0.734944 9.99958 2.98147e-06 1.19258e-05 0.130933 0.981207 0.931258 -0.0132931 4.9006e-06 0.502042 -1.89272e-20 6.97768e-24 -1.89202e-20 0.0013953 0.997818 8.59416e-05 0.152577 2.85186 0.0013953 0.997835 0.700954 0.00104927 0.00187989 0.000859416 0.455615 0.00187989 0.43762 0.000128353 1.02 0.887654 0.534688 0.286016 1.71673e-07 3.06105e-09 2387.71 3126.02 -0.0559033 0.482132 0.277563 0.25391 -0.593261 -0.169509 0.495467 -0.267932 -0.227544 1.642 1 0 297.2 0 2.08513 1.64 0.0002999 0.857538 0.653412 0.405488 0.409564 2.08536 131.14 83.8026 18.7141 60.8095 0.00403017 0 -40 10
0.741 2.14715e-08 2.53892e-06 0.0954983 0.0954954 0.0120402 9.75977e-06 0.00115406 0.119373 0.000657541 0.120026 0.871693 101.846 0.244563 0.735356 4.15379 0.0554373 0.0391867 0.960813 0.0198373 0.00427172 0.0191002 0.00410809 0.00516265 0.00589983 0.206506 0.235993 57.9852 -87.8953 126.213 15.9733 145.015 0.000141673 0.267123 192.893 0.310623 0.067378 0.00409543 0.000561704 0.00138291 0.986987 0.991733 -2.97501e-06 -85.6665 0.0929974 31191.7 301.326 0.983518 0.319147 0.734928 0.734924 9.99958 2.98147e-06 1.19258e-05 0.130935 0.981214 0.931261 -0.0132931 4.90063e-06 0.502049 -1.8928e-20 6.97803e-24 -1.89211e-20 0.0013953 0.997818 8.59416e-05 0.152577 2.85186 0.0013953 0.997835 0.701058 0.00104929 0.00187989 0.000859416 0.455614 0.00187989 0.437629 0.000128356 1.02 0.887655 0.534688 0.286018 1.71673e-07 3.06107e-09 2387.7 3125.93 -0.0558978 0.482132 0.277563 0.253905 -0.593262 -0.169509 0.495483 -0.26793 -0.227562 1.643 1 0 297.206 0 2.08529 1.641 0.0002999 0.8575 0.653464 0.405286 0.409591 2.08552 131.149 83.8036 18.7141 60.81 0.00403012 0 -40 10
0.742 2.15004e-08 2.53892e-06 0.0955728 0.09557 0.0120402 9.77293e-06 0.00115406 0.119466 0.000657544 0.120119 0.871754 101.846 0.244555 0.735447 4.15397 0.0554446 0.0391884 0.960812 0.0198371 0.00427189 0.0191 0.00410823 0.00516286 0.00590003 0.206514 0.236001 57.9852 -87.8953 126.213 15.9732 145.015 0.000141669 0.267123 192.892 0.310623 0.067378 0.00409543 0.000561705 0.00138291 0.986987 0.991733 -2.97503e-06 -85.6665 0.0929975 31191.7 301.331 0.983518 0.319147 0.734907 0.734903 9.99958 2.98148e-06 1.19258e-05 0.130937 0.981221 0.931264 -0.0132931 4.90066e-06 0.502056 -1.89289e-20 6.97838e-24 -1.89219e-20 0.0013953 0.997818 8.59417e-05 0.152577 2.85186 0.0013953 0.997835 0.701162 0.00104931 0.00187989 0.000859417 0.455614 0.00187989 0.437638 0.00012836 1.02 0.887656 0.534687 0.286019 1.71673e-07 3.0611e-09 2387.68 3125.84 -0.0558923 0.482132 0.277562 0.253899 -0.593263 -0.169509 0.495498 -0.267928 -0.227579 1.644 1 0 297.212 0 2.08546 1.642 0.0002999 0.857462 0.653516 0.405084 0.409619 2.08569 131.158 83.8046 18.7142 60.8105 0.00403008 0 -40 10
0.743 2.15294e-08 2.53892e-06 0.0956473 0.0956445 0.0120402 9.78608e-06 0.00115406 0.119559 0.000657546 0.120212 0.871816 101.846 0.244548 0.735538 4.15415 0.0554518 0.0391901 0.96081 0.0198369 0.00427206 0.0190998 0.00410837 0.00516307 0.00590024 0.206523 0.236009 57.9853 -87.8953 126.214 15.9732 145.015 0.000141665 0.267123 192.892 0.310623 0.0673779 0.00409543 0.000561705 0.00138291 0.986987 0.991733 -2.97504e-06 -85.6665 0.0929975 31191.6 301.335 0.983518 0.319147 0.734887 0.734882 9.99958 2.98148e-06 1.19258e-05 0.130939 0.981228 0.931266 -0.0132931 4.90068e-06 0.502063 -1.89297e-20 6.97872e-24 -1.89227e-20 0.00139531 0.997818 8.59418e-05 0.152577 2.85186 0.00139531 0.997835 0.701266 0.00104933 0.00187989 0.000859418 0.455614 0.00187989 0.437646 0.000128363 1.02 0.887657 0.534687 0.286021 1.71674e-07 3.06112e-09 2387.66 3125.75 -0.0558869 0.482132 0.277562 0.253894 -0.593264 -0.169509 0.495514 -0.267926 -0.227597 1.645 1 0 297.217 0 2.08562 1.643 0.000299899 0.857424 0.653568 0.404883 0.409647 2.08585 131.167 83.8057 18.7142 60.811 0.00403004 0 -40 10
0.744 2.15583e-08 2.53892e-06 0.0957217 0.0957189 0.0120401 9.79924e-06 0.00115406 0.119652 0.000657549 0.120305 0.871877 101.846 0.244541 0.73563 4.15433 0.0554591 0.0391918 0.960808 0.0198367 0.00427223 0.0190996 0.00410851 0.00516327 0.00590044 0.206531 0.236018 57.9854 -87.8954 126.214 15.9731 145.015 0.000141661 0.267123 192.892 0.310622 0.0673779 0.00409543 0.000561706 0.00138292 0.986987 0.991732 -2.97506e-06 -85.6665 0.0929976 31191.6 301.34 0.983518 0.319147 0.734866 0.734862 9.99958 2.98149e-06 1.19258e-05 0.13094 0.981235 0.931269 -0.013293 4.90071e-06 0.50207 -1.89305e-20 6.97907e-24 -1.89236e-20 0.00139531 0.997818 8.59419e-05 0.152578 2.85186 0.00139531 0.997835 0.70137 0.00104935 0.00187989 0.000859419 0.455614 0.00187989 0.437655 0.000128366 1.02 0.887658 0.534687 0.286022 1.71674e-07 3.06114e-09 2387.65 3125.67 -0.0558815 0.482132 0.277562 0.253888 -0.593265 -0.169509 0.495529 -0.267924 -0.227614 1.646 1 0 297.223 0 2.08579 1.644 0.000299899 0.857387 0.65362 0.404683 0.409675 2.08602 131.176 83.8067 18.7143 60.8115 0.00403 0 -40 10
0.745 2.15873e-08 2.53893e-06 0.095796 0.0957932 0.0120401 9.81239e-06 0.00115406 0.119745 0.000657552 0.120398 0.871939 101.845 0.244534 0.735721 4.15451 0.0554663 0.0391935 0.960807 0.0198365 0.0042724 0.0190994 0.00410865 0.00516348 0.00590065 0.206539 0.236026 57.9854 -87.8954 126.214 15.9731 145.015 0.000141657 0.267123 192.892 0.310622 0.0673778 0.00409544 0.000561707 0.00138292 0.986987 0.991732 -2.97507e-06 -85.6665 0.0929977 31191.6 301.345 0.983518 0.319147 0.734846 0.734841 9.99958 2.98149e-06 1.19259e-05 0.130942 0.981243 0.931272 -0.013293 4.90074e-06 0.502077 -1.89314e-20 6.97942e-24 -1.89244e-20 0.00139531 0.997818 8.59419e-05 0.152578 2.85186 0.00139531 0.997835 0.701474 0.00104937 0.0018799 0.000859419 0.455614 0.00187989 0.437663 0.00012837 1.02 0.887659 0.534686 0.286024 1.71674e-07 3.06116e-09 2387.63 3125.58 -0.0558762 0.482132 0.277562 0.253883 -0.593266 -0.169509 0.495544 -0.267922 -0.227631 1.647 1 0 297.229 0 2.08596 1.645 0.000299899 0.857349 0.653672 0.404483 0.409703 2.08619 131.185 83.8077 18.7144 60.8119 0.00402996 0 -40 10
0.746 2.16162e-08 2.53893e-06 0.0958703 0.0958675 0.0120401 9.82555e-06 0.00115406 0.119838 0.000657555 0.120491 0.872 101.845 0.244526 0.735812 4.15469 0.0554736 0.0391951 0.960805 0.0198363 0.00427256 0.0190991 0.00410879 0.00516369 0.00590086 0.206548 0.236034 57.9855 -87.8954 126.215 15.9731 145.015 0.000141653 0.267124 192.892 0.310621 0.0673778 0.00409544 0.000561707 0.00138292 0.986987 0.991732 -2.97509e-06 -85.6664 0.0929978 31191.6 301.349 0.983518 0.319147 0.734825 0.734821 9.99958 2.9815e-06 1.19259e-05 0.130944 0.98125 0.931275 -0.013293 4.90077e-06 0.502084 -1.89322e-20 6.97977e-24 -1.89252e-20 0.00139531 0.997818 8.5942e-05 0.152578 2.85187 0.00139531 0.997834 0.701578 0.00104939 0.0018799 0.00085942 0.455613 0.0018799 0.437672 0.000128373 1.02 0.88766 0.534686 0.286025 1.71674e-07 3.06118e-09 2387.61 3125.49 -0.0558708 0.482132 0.277561 0.253877 -0.593267 -0.169509 0.495559 -0.26792 -0.227648 1.648 1 0 297.234 0 2.08612 1.646 0.000299898 0.857312 0.653723 0.404283 0.40973 2.08635 131.194 83.8087 18.7144 60.8124 0.00402991 0 -40 10
0.747 2.16451e-08 2.53893e-06 0.0959446 0.0959418 0.0120401 9.8387e-06 0.00115406 0.119931 0.000657558 0.120584 0.872062 101.845 0.244519 0.735903 4.15487 0.0554808 0.0391968 0.960803 0.0198361 0.00427273 0.0190989 0.00410893 0.0051639 0.00590106 0.206556 0.236043 57.9856 -87.8954 126.215 15.973 145.015 0.000141649 0.267124 192.892 0.310621 0.0673777 0.00409544 0.000561708 0.00138292 0.986987 0.991732 -2.9751e-06 -85.6664 0.0929979 31191.5 301.354 0.983518 0.319147 0.734805 0.734801 9.99958 2.9815e-06 1.19259e-05 0.130946 0.981257 0.931278 -0.013293 4.9008e-06 0.502091 -1.8933e-20 6.98012e-24 -1.89261e-20 0.00139531 0.997818 8.59421e-05 0.152578 2.85187 0.00139531 0.997834 0.701682 0.00104941 0.0018799 0.000859421 0.455613 0.0018799 0.43768 0.000128376 1.02 0.887661 0.534686 0.286027 1.71675e-07 3.06121e-09 2387.6 3125.41 -0.0558655 0.482132 0.277561 0.253872 -0.593268 -0.169509 0.495574 -0.267918 -0.227665 1.649 1 0 297.24 0 2.08629 1.647 0.000299898 0.857275 0.653775 0.404084 0.409758 2.08652 131.203 83.8097 18.7145 60.8129 0.00402987 0 -40 10
0.748 2.16741e-08 2.53893e-06 0.0960187 0.0960159 0.0120401 9.85186e-06 0.00115406 0.120023 0.00065756 0.120676 0.872123 101.845 0.244512 0.735995 4.15505 0.0554881 0.0391985 0.960801 0.0198359 0.0042729 0.0190987 0.00410907 0.00516411 0.00590127 0.206564 0.236051 57.9856 -87.8954 126.215 15.973 145.015 0.000141645 0.267124 192.892 0.310621 0.0673777 0.00409545 0.000561709 0.00138293 0.986987 0.991732 -2.97512e-06 -85.6664 0.092998 31191.5 301.358 0.983518 0.319147 0.734785 0.734781 9.99958 2.9815e-06 1.19259e-05 0.130947 0.981264 0.931281 -0.013293 4.90083e-06 0.502098 -1.89339e-20 6.98047e-24 -1.89269e-20 0.00139531 0.997818 8.59422e-05 0.152578 2.85187 0.00139531 0.997834 0.701786 0.00104943 0.0018799 0.000859422 0.455613 0.0018799 0.437689 0.00012838 1.02 0.887662 0.534686 0.286028 1.71675e-07 3.06123e-09 2387.58 3125.32 -0.0558603 0.482132 0.277561 0.253866 -0.593269 -0.169509 0.495589 -0.267916 -0.227682 1.65 1 0 297.245 0 2.08645 1.648 0.000299898 0.857238 0.653827 0.403886 0.409786 2.08668 131.211 83.8107 18.7145 60.8134 0.00402983 0 -40 10
0.749 2.1703e-08 2.53893e-06 0.0960928 0.0960901 0.0120401 9.86501e-06 0.00115406 0.120116 0.000657563 0.120769 0.872185 101.845 0.244505 0.736086 4.15523 0.0554954 0.0392002 0.9608 0.0198357 0.00427307 0.0190985 0.00410922 0.00516432 0.00590148 0.206573 0.236059 57.9857 -87.8954 126.216 15.973 145.015 0.000141641 0.267124 192.891 0.31062 0.0673776 0.00409545 0.000561709 0.00138293 0.986987 0.991732 -2.97513e-06 -85.6664 0.092998 31191.5 301.363 0.983518 0.319147 0.734765 0.734761 9.99958 2.98151e-06 1.19259e-05 0.130949 0.981271 0.931284 -0.013293 4.90086e-06 0.502105 -1.89347e-20 6.98082e-24 -1.89277e-20 0.00139531 0.997818 8.59423e-05 0.152578 2.85187 0.00139531 0.997834 0.701889 0.00104945 0.0018799 0.000859423 0.455613 0.0018799 0.437697 0.000128383 1.02 0.887663 0.534685 0.286029 1.71675e-07 3.06125e-09 2387.56 3125.23 -0.055855 0.482132 0.27756 0.253861 -0.59327 -0.169509 0.495604 -0.267914 -0.227699 1.651 1 0 297.251 0 2.08662 1.649 0.000299897 0.857202 0.653879 0.403688 0.409814 2.08685 131.22 83.8117 18.7146 60.8139 0.00402979 0 -40 10
0.75 2.1732e-08 2.53893e-06 0.0961669 0.0961641 0.0120401 9.87817e-06 0.00115406 0.120209 0.000657566 0.120862 0.872247 101.845 0.244497 0.736178 4.15541 0.0555027 0.039202 0.960798 0.0198355 0.00427325 0.0190983 0.00410936 0.00516453 0.00590169 0.206581 0.236068 57.9857 -87.8954 126.216 15.9729 145.015 0.000141638 0.267124 192.891 0.31062 0.0673776 0.00409545 0.00056171 0.00138293 0.986987 0.991732 -2.97514e-06 -85.6664 0.0929981 31191.5 301.368 0.983518 0.319147 0.734745 0.734741 9.99958 2.98151e-06 1.19259e-05 0.130951 0.981278 0.931287 -0.013293 4.90089e-06 0.502113 -1.89355e-20 6.98117e-24 -1.89286e-20 0.00139531 0.997818 8.59423e-05 0.152578 2.85187 0.00139531 0.997834 0.701993 0.00104947 0.0018799 0.000859423 0.455612 0.0018799 0.437706 0.000128386 1.02 0.887664 0.534685 0.286031 1.71675e-07 3.06127e-09 2387.55 3125.15 -0.0558498 0.482133 0.27756 0.253855 -0.593271 -0.16951 0.495619 -0.267912 -0.227716 1.652 1 0 297.257 0 2.08678 1.65 0.000299897 0.857165 0.653931 0.40349 0.409841 2.08701 131.229 83.8127 18.7146 60.8143 0.00402975 0 -40 10
0.751 2.17609e-08 2.53893e-06 0.0962409 0.0962381 0.0120401 9.89132e-06 0.00115406 0.120301 0.000657569 0.120954 0.872308 101.844 0.24449 0.73627 4.15559 0.05551 0.0392037 0.960796 0.0198353 0.00427342 0.0190981 0.0041095 0.00516474 0.0059019 0.206589 0.236076 57.9858 -87.8954 126.217 15.9729 145.015 0.000141634 0.267125 192.891 0.310619 0.0673775 0.00409545 0.000561711 0.00138293 0.986987 0.991732 -2.97516e-06 -85.6664 0.0929982 31191.5 301.372 0.983518 0.319147 0.734725 0.734721 9.99958 2.98152e-06 1.1926e-05 0.130952 0.981285 0.93129 -0.013293 4.90092e-06 0.50212 -1.89364e-20 6.98151e-24 -1.89294e-20 0.00139531 0.997818 8.59424e-05 0.152579 2.85187 0.00139531 0.997834 0.702097 0.00104949 0.0018799 0.000859424 0.455612 0.0018799 0.437714 0.00012839 1.02 0.887665 0.534685 0.286032 1.71676e-07 3.0613e-09 2387.53 3125.06 -0.0558447 0.482133 0.27756 0.25385 -0.593272 -0.16951 0.495633 -0.26791 -0.227733 1.653 1 0 297.262 0 2.08695 1.651 0.000299897 0.857129 0.653983 0.403293 0.409869 2.08718 131.238 83.8136 18.7147 60.8148 0.00402971 0 -40 10
0.752 2.17898e-08 2.53893e-06 0.0963148 0.0963121 0.01204 9.90448e-06 0.00115406 0.120394 0.000657572 0.121047 0.87237 101.844 0.244483 0.736361 4.15577 0.0555173 0.0392054 0.960795 0.0198351 0.00427359 0.0190979 0.00410964 0.00516495 0.00590211 0.206598 0.236084 57.9859 -87.8954 126.217 15.9728 145.015 0.00014163 0.267125 192.891 0.310619 0.0673775 0.00409546 0.000561711 0.00138293 0.986987 0.991732 -2.97517e-06 -85.6664 0.0929983 31191.4 301.377 0.983518 0.319147 0.734705 0.734701 9.99958 2.98152e-06 1.1926e-05 0.130954 0.981292 0.931292 -0.013293 4.90094e-06 0.502127 -1.89372e-20 6.98186e-24 -1.89302e-20 0.00139531 0.997818 8.59425e-05 0.152579 2.85187 0.00139531 0.997834 0.702201 0.00104951 0.00187991 0.000859425 0.455612 0.0018799 0.437723 0.000128393 1.02 0.887666 0.534684 0.286034 1.71676e-07 3.06132e-09 2387.51 3124.98 -0.0558395 0.482133 0.27756 0.253845 -0.593273 -0.16951 0.495648 -0.267907 -0.227749 1.654 1 0 297.267 0 2.08711 1.652 0.000299896 0.857093 0.654034 0.403096 0.409897 2.08734 131.247 83.8146 18.7148 60.8153 0.00402967 0 -40 10
0.753 2.18188e-08 2.53893e-06 0.0963887 0.0963859 0.01204 9.91763e-06 0.00115406 0.120486 0.000657574 0.121139 0.872432 101.844 0.244475 0.736453 4.15595 0.0555246 0.0392071 0.960793 0.0198348 0.00427376 0.0190977 0.00410979 0.00516516 0.00590232 0.206606 0.236093 57.9859 -87.8954 126.217 15.9728 145.015 0.000141626 0.267125 192.891 0.310619 0.0673774 0.00409546 0.000561712 0.00138294 0.986987 0.991732 -2.97519e-06 -85.6664 0.0929984 31191.4 301.381 0.983518 0.319147 0.734686 0.734681 9.99958 2.98153e-06 1.1926e-05 0.130956 0.981299 0.931295 -0.013293 4.90097e-06 0.502134 -1.8938e-20 6.98221e-24 -1.89311e-20 0.00139532 0.997818 8.59426e-05 0.152579 2.85187 0.00139532 0.997834 0.702304 0.00104953 0.00187991 0.000859426 0.455612 0.00187991 0.437731 0.000128396 1.02 0.887668 0.534684 0.286035 1.71676e-07 3.06134e-09 2387.5 3124.89 -0.0558344 0.482133 0.277559 0.25384 -0.593274 -0.16951 0.495662 -0.267905 -0.227766 1.655 1 0 297.273 0 2.08728 1.653 0.000299896 0.857058 0.654086 0.4029 0.409924 2.08751 131.256 83.8156 18.7148 60.8157 0.00402963 0 -40 10
0.754 2.18477e-08 2.53893e-06 0.0964625 0.0964598 0.01204 9.93078e-06 0.00115406 0.120578 0.000657577 0.121231 0.872494 101.844 0.244468 0.736545 4.15613 0.0555319 0.0392088 0.960791 0.0198346 0.00427393 0.0190975 0.00410993 0.00516537 0.00590253 0.206615 0.236101 57.986 -87.8954 126.218 15.9728 145.015 0.000141622 0.267125 192.891 0.310618 0.0673774 0.00409546 0.000561712 0.00138294 0.986987 0.991732 -2.9752e-06 -85.6664 0.0929985 31191.4 301.386 0.983518 0.319147 0.734666 0.734662 9.99958 2.98153e-06 1.1926e-05 0.130958 0.981306 0.931298 -0.013293 4.901e-06 0.502141 -1.89389e-20 6.98256e-24 -1.89319e-20 0.00139532 0.997818 8.59426e-05 0.152579 2.85187 0.00139532 0.997834 0.702408 0.00104955 0.00187991 0.000859426 0.455612 0.00187991 0.43774 0.0001284 1.02 0.887669 0.534684 0.286037 1.71677e-07 3.06136e-09 2387.48 3124.81 -0.0558294 0.482133 0.277559 0.253834 -0.593275 -0.16951 0.495676 -0.267903 -0.227782 1.656 1 0 297.278 0 2.08744 1.654 0.000299896 0.857022 0.654138 0.402704 0.409952 2.08767 131.265 83.8165 18.7149 60.8162 0.00402959 0 -40 10
0.755 2.18767e-08 2.53893e-06 0.0965363 0.0965335 0.01204 9.94394e-06 0.00115406 0.12067 0.00065758 0.121323 0.872556 101.844 0.244461 0.736637 4.15632 0.0555392 0.0392105 0.960789 0.0198344 0.0042741 0.0190973 0.00411007 0.00516558 0.00590274 0.206623 0.236109 57.9861 -87.8954 126.218 15.9727 145.015 0.000141619 0.267125 192.89 0.310618 0.0673773 0.00409547 0.000561713 0.00138294 0.986987 0.991732 -2.97522e-06 -85.6664 0.0929985 31191.4 301.391 0.983518 0.319147 0.734647 0.734643 9.99958 2.98154e-06 1.1926e-05 0.13096 0.981313 0.931301 -0.013293 4.90103e-06 0.502149 -1.89397e-20 6.98291e-24 -1.89327e-20 0.00139532 0.997818 8.59427e-05 0.152579 2.85187 0.00139532 0.997834 0.702511 0.00104957 0.00187991 0.000859427 0.455611 0.00187991 0.437748 0.000128403 1.02 0.88767 0.534683 0.286038 1.71677e-07 3.06138e-09 2387.46 3124.73 -0.0558243 0.482133 0.277559 0.253829 -0.593276 -0.16951 0.49569 -0.267901 -0.227798 1.657 1 0 297.284 0 2.08761 1.655 0.000299895 0.856987 0.654189 0.402509 0.40998 2.08784 131.273 83.8175 18.7149 60.8167 0.00402955 0 -40 10
0.756 2.19056e-08 2.53893e-06 0.09661 0.0966072 0.01204 9.95709e-06 0.00115406 0.120762 0.000657583 0.121415 0.872618 101.843 0.244453 0.736729 4.1565 0.0555466 0.0392123 0.960788 0.0198342 0.00427428 0.0190971 0.00411022 0.00516579 0.00590295 0.206632 0.236118 57.9861 -87.8954 126.218 15.9727 145.016 0.000141615 0.267125 192.89 0.310617 0.0673773 0.00409547 0.000561714 0.00138294 0.986987 0.991732 -2.97523e-06 -85.6664 0.0929986 31191.4 301.395 0.983518 0.319147 0.734628 0.734623 9.99958 2.98154e-06 1.19261e-05 0.130961 0.98132 0.931304 -0.013293 4.90106e-06 0.502156 -1.89405e-20 6.98326e-24 -1.89336e-20 0.00139532 0.997818 8.59428e-05 0.152579 2.85187 0.00139532 0.997833 0.702615 0.00104959 0.00187991 0.000859428 0.455611 0.00187991 0.437757 0.000128406 1.02 0.887671 0.534683 0.28604 1.71677e-07 3.06141e-09 2387.45 3124.64 -0.0558193 0.482133 0.277558 0.253824 -0.593277 -0.16951 0.495705 -0.267899 -0.227814 1.658 1 0 297.289 0 2.08777 1.656 0.000299895 0.856951 0.654241 0.402314 0.410007 2.088 131.282 83.8185 18.715 60.8171 0.00402951 0 -40 10
0.757 2.19345e-08 2.53893e-06 0.0966836 0.0966809 0.01204 9.97025e-06 0.00115406 0.120855 0.000657585 0.121507 0.87268 101.843 0.244446 0.736821 4.15668 0.0555539 0.039214 0.960786 0.019834 0.00427445 0.0190968 0.00411036 0.00516601 0.00590316 0.20664 0.236126 57.9862 -87.8954 126.219 15.9727 145.016 0.000141611 0.267126 192.89 0.310617 0.0673772 0.00409547 0.000561714 0.00138294 0.986987 0.991732 -2.97525e-06 -85.6663 0.0929987 31191.3 301.4 0.983518 0.319147 0.734608 0.734604 9.99958 2.98155e-06 1.19261e-05 0.130963 0.981327 0.931306 -0.013293 4.90109e-06 0.502163 -1.89414e-20 6.98361e-24 -1.89344e-20 0.00139532 0.997818 8.59429e-05 0.152579 2.85187 0.00139532 0.997833 0.702718 0.00104961 0.00187991 0.000859429 0.455611 0.00187991 0.437765 0.00012841 1.02 0.887672 0.534683 0.286041 1.71677e-07 3.06143e-09 2387.43 3124.56 -0.0558144 0.482133 0.277558 0.253819 -0.593278 -0.16951 0.495719 -0.267897 -0.227831 1.659 1 0 297.294 0 2.08794 1.657 0.000299894 0.856916 0.654293 0.402119 0.410035 2.08817 131.291 83.8194 18.715 60.8176 0.00402947 0 -40 10
0.758 2.19635e-08 2.53893e-06 0.0967572 0.0967545 0.01204 9.9834e-06 0.00115406 0.120946 0.000657588 0.121599 0.872742 101.843 0.244439 0.736913 4.15687 0.0555612 0.0392157 0.960784 0.0198338 0.00427462 0.0190966 0.00411051 0.00516622 0.00590337 0.206649 0.236135 57.9863 -87.8954 126.219 15.9726 145.016 0.000141608 0.267126 192.89 0.310617 0.0673772 0.00409548 0.000561715 0.00138295 0.986987 0.991732 -2.97526e-06 -85.6663 0.0929988 31191.3 301.405 0.983518 0.319147 0.734589 0.734585 9.99958 2.98155e-06 1.19261e-05 0.130965 0.981333 0.931309 -0.013293 4.90112e-06 0.50217 -1.89422e-20 6.98396e-24 -1.89352e-20 0.00139532 0.997818 8.5943e-05 0.15258 2.85188 0.00139532 0.997833 0.702822 0.00104962 0.00187991 0.00085943 0.455611 0.00187991 0.437774 0.000128413 1.02 0.887673 0.534683 0.286043 1.71678e-07 3.06145e-09 2387.41 3124.48 -0.0558094 0.482133 0.277558 0.253814 -0.593279 -0.16951 0.495732 -0.267895 -0.227846 1.66 1 0 297.299 0 2.0881 1.658 0.000299894 0.856881 0.654344 0.401925 0.410063 2.08833 131.3 83.8203 18.7151 60.818 0.00402943 0 -40 10
0.759 2.19924e-08 2.53893e-06 0.0968307 0.096828 0.0120399 9.99656e-06 0.00115406 0.121038 0.000657591 0.121691 0.872804 101.843 0.244431 0.737006 4.15705 0.0555686 0.0392175 0.960783 0.0198336 0.0042748 0.0190964 0.00411065 0.00516643 0.00590358 0.206657 0.236143 57.9863 -87.8954 126.219 15.9726 145.016 0.000141604 0.267126 192.89 0.310616 0.0673771 0.00409548 0.000561716 0.00138295 0.986987 0.991732 -2.97527e-06 -85.6663 0.0929989 31191.3 301.41 0.983518 0.319147 0.73457 0.734566 9.99958 2.98156e-06 1.19261e-05 0.130967 0.98134 0.931312 -0.013293 4.90115e-06 0.502178 -1.89431e-20 6.98432e-24 -1.89361e-20 0.00139532 0.997818 8.5943e-05 0.15258 2.85188 0.00139532 0.997833 0.702925 0.00104964 0.00187992 0.00085943 0.45561 0.00187991 0.437782 0.000128416 1.02 0.887674 0.534682 0.286044 1.71678e-07 3.06147e-09 2387.4 3124.4 -0.0558045 0.482133 0.277558 0.253808 -0.59328 -0.16951 0.495746 -0.267893 -0.227862 1.661 1 0 297.305 0 2.08827 1.659 0.000299894 0.856847 0.654396 0.401732 0.41009 2.0885 131.309 83.8213 18.7151 60.8185 0.0040294 0 -40 10
0.76 2.20214e-08 2.53893e-06 0.0969042 0.0969015 0.0120399 1.00097e-05 0.00115406 0.12113 0.000657594 0.121783 0.872866 101.843 0.244424 0.737098 4.15724 0.0555759 0.0392192 0.960781 0.0198334 0.00427497 0.0190962 0.0041108 0.00516665 0.0059038 0.206666 0.236152 57.9864 -87.8954 126.22 15.9725 145.016 0.0001416 0.267126 192.89 0.310616 0.0673771 0.00409548 0.000561716 0.00138295 0.986987 0.991732 -2.97529e-06 -85.6663 0.092999 31191.3 301.414 0.983518 0.319147 0.734551 0.734547 9.99958 2.98156e-06 1.19261e-05 0.130968 0.981347 0.931315 -0.013293 4.90117e-06 0.502185 -1.89439e-20 6.98467e-24 -1.89369e-20 0.00139532 0.997818 8.59431e-05 0.15258 2.85188 0.00139532 0.997833 0.703029 0.00104966 0.00187992 0.000859431 0.45561 0.00187992 0.437791 0.00012842 1.02 0.887675 0.534682 0.286046 1.71678e-07 3.06149e-09 2387.38 3124.32 -0.0557996 0.482133 0.277557 0.253803 -0.593281 -0.16951 0.49576 -0.267891 -0.227878 1.662 1 0 297.31 0 2.08843 1.66 0.000299893 0.856812 0.654448 0.401539 0.410118 2.08866 131.318 83.8222 18.7152 60.8189 0.00402936 0 -40 10
0.761 2.20503e-08 2.53893e-06 0.0969776 0.0969749 0.0120399 1.00229e-05 0.00115406 0.121222 0.000657596 0.121875 0.872928 101.843 0.244417 0.737191 4.15742 0.0555833 0.039221 0.960779 0.0198331 0.00427514 0.019096 0.00411094 0.00516686 0.00590401 0.206674 0.23616 57.9864 -87.8954 126.22 15.9725 145.016 0.000141597 0.267126 192.889 0.310615 0.067377 0.00409548 0.000561717 0.00138295 0.986987 0.991732 -2.9753e-06 -85.6663 0.092999 31191.2 301.419 0.983518 0.319147 0.734532 0.734528 9.99958 2.98157e-06 1.19262e-05 0.13097 0.981354 0.931317 -0.013293 4.9012e-06 0.502192 -1.89447e-20 6.98502e-24 -1.89378e-20 0.00139532 0.997818 8.59432e-05 0.15258 2.85188 0.00139532 0.997833 0.703132 0.00104968 0.00187992 0.000859432 0.45561 0.00187992 0.437799 0.000128423 1.02 0.887676 0.534682 0.286047 1.71678e-07 3.06152e-09 2387.36 3124.24 -0.0557948 0.482133 0.277557 0.253798 -0.593282 -0.16951 0.495774 -0.267889 -0.227894 1.663 1 0 297.315 0 2.0886 1.661 0.000299893 0.856778 0.654499 0.401346 0.410145 2.08883 131.326 83.8231 18.7153 60.8194 0.00402932 0 -40 10
0.762 2.20792e-08 2.53893e-06 0.0970509 0.0970482 0.0120399 1.0036e-05 0.00115406 0.121314 0.000657599 0.121967 0.87299 101.842 0.244409 0.737283 4.15761 0.0555907 0.0392227 0.960777 0.0198329 0.00427532 0.0190958 0.00411109 0.00516707 0.00590422 0.206683 0.236169 57.9865 -87.8954 126.22 15.9725 145.016 0.000141593 0.267127 192.889 0.310615 0.067377 0.00409549 0.000561718 0.00138295 0.986987 0.991732 -2.97532e-06 -85.6663 0.0929991 31191.2 301.424 0.983518 0.319147 0.734514 0.734509 9.99958 2.98157e-06 1.19262e-05 0.130972 0.981361 0.93132 -0.013293 4.90123e-06 0.502199 -1.89456e-20 6.98537e-24 -1.89386e-20 0.00139533 0.997818 8.59433e-05 0.15258 2.85188 0.00139533 0.997833 0.703235 0.0010497 0.00187992 0.000859433 0.45561 0.00187992 0.437808 0.000128426 1.02 0.887677 0.534681 0.286049 1.71679e-07 3.06154e-09 2387.35 3124.16 -0.05579 0.482133 0.277557 0.253793 -0.593283 -0.16951 0.495787 -0.267887 -0.227909 1.664 1 0 297.32 0 2.08876 1.662 0.000299893 0.856744 0.654551 0.401154 0.410173 2.08899 131.335 83.8241 18.7153 60.8198 0.00402928 0 -40 10
0.763 2.21082e-08 2.53893e-06 0.0971242 0.0971215 0.0120399 1.00492e-05 0.00115406 0.121405 0.000657602 0.122058 0.873053 101.842 0.244402 0.737376 4.1578 0.055598 0.0392245 0.960776 0.0198327 0.00427549 0.0190956 0.00411123 0.00516729 0.00590444 0.206692 0.236177 57.9866 -87.8954 126.221 15.9724 145.016 0.000141589 0.267127 192.889 0.310614 0.0673769 0.00409549 0.000561718 0.00138296 0.986987 0.991732 -2.97533e-06 -85.6663 0.0929992 31191.2 301.428 0.983518 0.319147 0.734495 0.734491 9.99958 2.98158e-06 1.19262e-05 0.130974 0.981367 0.931323 -0.013293 4.90126e-06 0.502207 -1.89464e-20 6.98572e-24 -1.89394e-20 0.00139533 0.997818 8.59433e-05 0.15258 2.85188 0.00139533 0.997833 0.703339 0.00104972 0.00187992 0.000859433 0.45561 0.00187992 0.437816 0.00012843 1.02 0.887678 0.534681 0.28605 1.71679e-07 3.06156e-09 2387.33 3124.08 -0.0557852 0.482133 0.277556 0.253788 -0.593284 -0.16951 0.495801 -0.267885 -0.227925 1.665 1 0 297.325 0 2.08893 1.663 0.000299892 0.85671 0.654602 0.400962 0.410201 2.08916 131.344 83.825 18.7154 60.8203 0.00402924 0 -40 10
0.764 2.21371e-08 2.53893e-06 0.0971974 0.0971947 0.0120399 1.00623e-05 0.00115406 0.121497 0.000657604 0.12215 0.873115 101.842 0.244395 0.737468 4.15798 0.0556054 0.0392262 0.960774 0.0198325 0.00427567 0.0190953 0.00411138 0.0051675 0.00590465 0.2067 0.236186 57.9866 -87.8954 126.221 15.9724 145.016 0.000141586 0.267127 192.889 0.310614 0.0673769 0.00409549 0.000561719 0.00138296 0.986987 0.991732 -2.97535e-06 -85.6663 0.0929993 31191.2 301.433 0.983518 0.319147 0.734477 0.734472 9.99958 2.98158e-06 1.19262e-05 0.130976 0.981374 0.931325 -0.013293 4.90129e-06 0.502214 -1.89473e-20 6.98607e-24 -1.89403e-20 0.00139533 0.997818 8.59434e-05 0.15258 2.85188 0.00139533 0.997833 0.703442 0.00104974 0.00187992 0.000859434 0.455609 0.00187992 0.437825 0.000128433 1.02 0.887679 0.534681 0.286052 1.71679e-07 3.06158e-09 2387.31 3124 -0.0557804 0.482134 0.277556 0.253783 -0.593284 -0.16951 0.495814 -0.267883 -0.22794 1.666 1 0 297.33 0 2.08909 1.664 0.000299892 0.856677 0.654654 0.400771 0.410228 2.08932 131.353 83.8259 18.7154 60.8207 0.0040292 0 -40 10
0.765 2.21661e-08 2.53893e-06 0.0972706 0.0972679 0.0120399 1.00755e-05 0.00115406 0.121588 0.000657607 0.122241 0.873178 101.842 0.244387 0.737561 4.15817 0.0556128 0.039228 0.960772 0.0198323 0.00427584 0.0190951 0.00411153 0.00516772 0.00590487 0.206709 0.236195 57.9867 -87.8954 126.221 15.9724 145.016 0.000141582 0.267127 192.889 0.310614 0.0673768 0.0040955 0.00056172 0.00138296 0.986986 0.991732 -2.97536e-06 -85.6663 0.0929994 31191.2 301.438 0.983517 0.319147 0.734458 0.734454 9.99958 2.98159e-06 1.19262e-05 0.130977 0.981381 0.931328 -0.013293 4.90132e-06 0.502221 -1.89481e-20 6.98642e-24 -1.89411e-20 0.00139533 0.997818 8.59435e-05 0.152581 2.85188 0.00139533 0.997833 0.703545 0.00104976 0.00187992 0.000859435 0.455609 0.00187992 0.437833 0.000128436 1.02 0.88768 0.53468 0.286053 1.71679e-07 3.06161e-09 2387.3 3123.92 -0.0557757 0.482134 0.277556 0.253778 -0.593285 -0.169511 0.495827 -0.26788 -0.227956 1.667 1 0 297.335 0 2.08926 1.665 0.000299892 0.856643 0.654705 0.40058 0.410256 2.08948 131.362 83.8268 18.7155 60.8212 0.00402917 0 -40 10
0.766 2.2195e-08 2.53893e-06 0.0973437 0.097341 0.0120399 1.00886e-05 0.00115406 0.12168 0.00065761 0.122333 0.87324 101.842 0.24438 0.737654 4.15836 0.0556202 0.0392298 0.96077 0.0198321 0.00427602 0.0190949 0.00411167 0.00516794 0.00590508 0.206717 0.236203 57.9868 -87.8954 126.222 15.9723 145.016 0.000141579 0.267127 192.889 0.310613 0.0673768 0.0040955 0.00056172 0.00138296 0.986986 0.991732 -2.97538e-06 -85.6663 0.0929995 31191.1 301.443 0.983517 0.319147 0.73444 0.734435 9.99958 2.98159e-06 1.19263e-05 0.130979 0.981388 0.931331 -0.013293 4.90135e-06 0.502229 -1.89489e-20 6.98678e-24 -1.89419e-20 0.00139533 0.997818 8.59436e-05 0.152581 2.85188 0.00139533 0.997832 0.703648 0.00104978 0.00187993 0.000859436 0.455609 0.00187992 0.437842 0.00012844 1.02 0.887681 0.53468 0.286055 1.7168e-07 3.06163e-09 2387.28 3123.84 -0.055771 0.482134 0.277556 0.253773 -0.593286 -0.169511 0.49584 -0.267878 -0.227971 1.668 1 0 297.34 0 2.08942 1.666 0.000299891 0.85661 0.654757 0.40039 0.410283 2.08965 131.37 83.8277 18.7155 60.8216 0.00402913 0 -40 10
0.767 2.22239e-08 2.53893e-06 0.0974167 0.0974141 0.0120398 1.01018e-05 0.00115406 0.121771 0.000657612 0.122424 0.873302 101.841 0.244372 0.737747 4.15854 0.0556276 0.0392315 0.960768 0.0198318 0.0042762 0.0190947 0.00411182 0.00516815 0.0059053 0.206726 0.236212 57.9868 -87.8954 126.222 15.9723 145.016 0.000141575 0.267127 192.889 0.310613 0.0673767 0.0040955 0.000561721 0.00138296 0.986986 0.991732 -2.97539e-06 -85.6663 0.0929995 31191.1 301.448 0.983517 0.319147 0.734422 0.734417 9.99958 2.98159e-06 1.19263e-05 0.130981 0.981394 0.931333 -0.013293 4.90138e-06 0.502236 -1.89498e-20 6.98713e-24 -1.89428e-20 0.00139533 0.997818 8.59437e-05 0.152581 2.85188 0.00139533 0.997832 0.703751 0.0010498 0.00187993 0.000859437 0.455609 0.00187993 0.43785 0.000128443 1.02 0.887682 0.53468 0.286056 1.7168e-07 3.06165e-09 2387.26 3123.76 -0.0557664 0.482134 0.277555 0.253768 -0.593287 -0.169511 0.495853 -0.267876 -0.227986 1.669 1 0 297.345 0 2.08958 1.667 0.000299891 0.856577 0.654808 0.4002 0.410311 2.08981 131.379 83.8286 18.7156 60.822 0.00402909 0 -40 10
0.768 2.22529e-08 2.53894e-06 0.0974897 0.0974871 0.0120398 1.01149e-05 0.00115406 0.121862 0.000657615 0.122515 0.873365 101.841 0.244365 0.73784 4.15873 0.055635 0.0392333 0.960767 0.0198316 0.00427637 0.0190945 0.00411197 0.00516837 0.00590551 0.206735 0.23622 57.9869 -87.8954 126.222 15.9722 145.016 0.000141572 0.267128 192.888 0.310612 0.0673767 0.0040955 0.000561721 0.00138297 0.986986 0.991732 -2.9754e-06 -85.6662 0.0929996 31191.1 301.452 0.983517 0.319147 0.734403 0.734399 9.99958 2.9816e-06 1.19263e-05 0.130983 0.981401 0.931336 -0.013293 4.90141e-06 0.502244 -1.89506e-20 6.98748e-24 -1.89436e-20 0.00139533 0.997818 8.59437e-05 0.152581 2.85188 0.00139533 0.997832 0.703854 0.00104982 0.00187993 0.000859437 0.455609 0.00187993 0.437859 0.000128446 1.02 0.887684 0.53468 0.286058 1.7168e-07 3.06167e-09 2387.25 3123.68 -0.0557617 0.482134 0.277555 0.253764 -0.593288 -0.169511 0.495866 -0.267874 -0.228001 1.67 1 0 297.35 0 2.08975 1.668 0.000299891 0.856544 0.654859 0.40001 0.410338 2.08998 131.388 83.8295 18.7156 60.8225 0.00402906 0 -40 10
0.769 2.22818e-08 2.53894e-06 0.0975627 0.09756 0.0120398 1.01281e-05 0.00115406 0.121953 0.000657618 0.122606 0.873428 101.841 0.244358 0.737933 4.15892 0.0556424 0.0392351 0.960765 0.0198314 0.00427655 0.0190943 0.00411212 0.00516859 0.00590573 0.206744 0.236229 57.987 -87.8954 126.223 15.9722 145.016 0.000141568 0.267128 192.888 0.310612 0.0673766 0.00409551 0.000561722 0.00138297 0.986986 0.991732 -2.97542e-06 -85.6662 0.0929997 31191.1 301.457 0.983517 0.319147 0.734385 0.734381 9.99958 2.9816e-06 1.19263e-05 0.130985 0.981407 0.931339 -0.013293 4.90144e-06 0.502251 -1.89515e-20 6.98783e-24 -1.89445e-20 0.00139533 0.997818 8.59438e-05 0.152581 2.85189 0.00139533 0.997832 0.703958 0.00104984 0.00187993 0.000859438 0.455608 0.00187993 0.437867 0.00012845 1.02 0.887685 0.534679 0.286059 1.7168e-07 3.06169e-09 2387.23 3123.6 -0.0557571 0.482134 0.277555 0.253759 -0.593289 -0.169511 0.495879 -0.267872 -0.228016 1.671 1 0 297.355 0 2.08991 1.669 0.00029989 0.856511 0.654911 0.399821 0.410366 2.09014 131.397 83.8304 18.7157 60.8229 0.00402902 0 -40 10
0.77 2.23107e-08 2.53894e-06 0.0976355 0.0976329 0.0120398 1.01412e-05 0.00115406 0.122044 0.00065762 0.122697 0.87349 101.841 0.24435 0.738026 4.15911 0.0556498 0.0392369 0.960763 0.0198312 0.00427673 0.0190941 0.00411226 0.00516881 0.00590594 0.206752 0.236238 57.987 -87.8954 126.223 15.9722 145.016 0.000141565 0.267128 192.888 0.310612 0.0673766 0.00409551 0.000561723 0.00138297 0.986986 0.991732 -2.97543e-06 -85.6662 0.0929998 31191 301.462 0.983517 0.319147 0.734367 0.734363 9.99958 2.98161e-06 1.19263e-05 0.130986 0.981414 0.931341 -0.013293 4.90146e-06 0.502258 -1.89523e-20 6.98818e-24 -1.89453e-20 0.00139533 0.997818 8.59439e-05 0.152581 2.85189 0.00139533 0.997832 0.704061 0.00104986 0.00187993 0.000859439 0.455608 0.00187993 0.437876 0.000128453 1.02 0.887686 0.534679 0.286061 1.71681e-07 3.06172e-09 2387.21 3123.53 -0.0557526 0.482134 0.277554 0.253754 -0.59329 -0.169511 0.495892 -0.26787 -0.228031 1.672 1 0 297.36 0 2.09008 1.67 0.00029989 0.856478 0.654962 0.399633 0.410393 2.0903 131.406 83.8313 18.7157 60.8233 0.00402898 0 -40 10
0.771 2.23397e-08 2.53894e-06 0.0977084 0.0977057 0.0120398 1.01544e-05 0.00115406 0.122135 0.000657623 0.122788 0.873553 101.841 0.244343 0.73812 4.1593 0.0556572 0.0392387 0.960761 0.019831 0.0042769 0.0190938 0.00411241 0.00516902 0.00590616 0.206761 0.236246 57.9871 -87.8955 126.223 15.9721 145.016 0.000141561 0.267128 192.888 0.310611 0.0673765 0.00409551 0.000561723 0.00138297 0.986986 0.991732 -2.97545e-06 -85.6662 0.0929999 31191 301.467 0.983517 0.319147 0.734349 0.734345 9.99958 2.98161e-06 1.19263e-05 0.130988 0.981421 0.931344 -0.013293 4.90149e-06 0.502266 -1.89531e-20 6.98854e-24 -1.89462e-20 0.00139534 0.997818 8.5944e-05 0.152582 2.85189 0.00139534 0.997832 0.704164 0.00104988 0.00187993 0.00085944 0.455608 0.00187993 0.437884 0.000128456 1.02 0.887687 0.534679 0.286062 1.71681e-07 3.06174e-09 2387.2 3123.45 -0.055748 0.482134 0.277554 0.253749 -0.593291 -0.169511 0.495905 -0.267868 -0.228046 1.673 1 0 297.365 0 2.09024 1.671 0.000299889 0.856446 0.655013 0.399445 0.410421 2.09047 131.414 83.8322 18.7158 60.8237 0.00402895 0 -40 10
0.772 2.23686e-08 2.53894e-06 0.0977811 0.0977785 0.0120398 1.01676e-05 0.00115406 0.122226 0.000657626 0.122879 0.873616 101.841 0.244335 0.738213 4.15949 0.0556647 0.0392405 0.96076 0.0198308 0.00427708 0.0190936 0.00411256 0.00516924 0.00590638 0.20677 0.236255 57.9871 -87.8955 126.224 15.9721 145.016 0.000141558 0.267128 192.888 0.310611 0.0673765 0.00409552 0.000561724 0.00138298 0.986986 0.991732 -2.97546e-06 -85.6662 0.093 31191 301.472 0.983517 0.319147 0.734332 0.734327 9.99958 2.98162e-06 1.19264e-05 0.13099 0.981427 0.931347 -0.013293 4.90152e-06 0.502273 -1.8954e-20 6.98889e-24 -1.8947e-20 0.00139534 0.997818 8.5944e-05 0.152582 2.85189 0.00139534 0.997832 0.704266 0.0010499 0.00187993 0.00085944 0.455608 0.00187993 0.437893 0.00012846 1.02 0.887688 0.534678 0.286064 1.71681e-07 3.06176e-09 2387.18 3123.37 -0.0557435 0.482134 0.277554 0.253744 -0.593292 -0.169511 0.495917 -0.267866 -0.22806 1.674 1 0 297.37 0 2.0904 1.672 0.000299889 0.856414 0.655065 0.399257 0.410448 2.09063 131.423 83.8331 18.7158 60.8242 0.00402891 0 -40 10
0.773 2.23976e-08 2.53894e-06 0.0978538 0.0978512 0.0120398 1.01807e-05 0.00115406 0.122317 0.000657628 0.12297 0.873678 101.84 0.244328 0.738306 4.15968 0.0556721 0.0392422 0.960758 0.0198305 0.00427726 0.0190934 0.00411271 0.00516946 0.0059066 0.206778 0.236264 57.9872 -87.8955 126.224 15.972 145.016 0.000141555 0.267129 192.888 0.31061 0.0673764 0.00409552 0.000561725 0.00138298 0.986986 0.991732 -2.97548e-06 -85.6662 0.0930001 31191 301.476 0.983517 0.319147 0.734314 0.73431 9.99958 2.98162e-06 1.19264e-05 0.130992 0.981434 0.931349 -0.013293 4.90155e-06 0.502281 -1.89548e-20 6.98924e-24 -1.89478e-20 0.00139534 0.997818 8.59441e-05 0.152582 2.85189 0.00139534 0.997832 0.704369 0.00104992 0.00187994 0.000859441 0.455607 0.00187993 0.437901 0.000128463 1.02 0.887689 0.534678 0.286065 1.71681e-07 3.06178e-09 2387.16 3123.3 -0.0557391 0.482134 0.277554 0.253739 -0.593292 -0.169511 0.49593 -0.267864 -0.228075 1.675 1 0 297.375 0 2.09057 1.673 0.000299889 0.856382 0.655116 0.39907 0.410475 2.0908 131.432 83.8339 18.7159 60.8246 0.00402887 0 -40 10
0.774 2.24265e-08 2.53894e-06 0.0979265 0.0979238 0.0120397 1.01939e-05 0.00115406 0.122408 0.000657631 0.123061 0.873741 101.84 0.24432 0.7384 4.15987 0.0556795 0.039244 0.960756 0.0198303 0.00427744 0.0190932 0.00411286 0.00516968 0.00590682 0.206787 0.236273 57.9873 -87.8955 126.224 15.972 145.016 0.000141551 0.267129 192.887 0.31061 0.0673763 0.00409552 0.000561725 0.00138298 0.986986 0.991732 -2.97549e-06 -85.6662 0.0930001 31191 301.481 0.983517 0.319147 0.734296 0.734292 9.99958 2.98163e-06 1.19264e-05 0.130994 0.98144 0.931352 -0.013293 4.90158e-06 0.502288 -1.89557e-20 6.9896e-24 -1.89487e-20 0.00139534 0.997818 8.59442e-05 0.152582 2.85189 0.00139534 0.997832 0.704472 0.00104994 0.00187994 0.000859442 0.455607 0.00187994 0.437909 0.000128466 1.02 0.88769 0.534678 0.286067 1.71682e-07 3.06181e-09 2387.15 3123.22 -0.0557346 0.482134 0.277553 0.253735 -0.593293 -0.169511 0.495942 -0.267862 -0.228089 1.676 1 0 297.379 0 2.09073 1.674 0.000299888 0.85635 0.655167 0.398883 0.410503 2.09096 131.441 83.8348 18.7159 60.825 0.00402884 0 -40 10
0.775 2.24554e-08 2.53894e-06 0.097999 0.0979964 0.0120397 1.0207e-05 0.00115406 0.122499 0.000657634 0.123152 0.873804 101.84 0.244313 0.738493 4.16006 0.055687 0.0392458 0.960754 0.0198301 0.00427762 0.019093 0.00411301 0.0051699 0.00590703 0.206796 0.236281 57.9873 -87.8955 126.225 15.972 145.016 0.000141548 0.267129 192.887 0.310609 0.0673763 0.00409552 0.000561726 0.00138298 0.986986 0.991732 -2.97551e-06 -85.6662 0.0930002 31190.9 301.486 0.983517 0.319147 0.734279 0.734275 9.99958 2.98163e-06 1.19264e-05 0.130995 0.981447 0.931354 -0.013293 4.90161e-06 0.502296 -1.89565e-20 6.98995e-24 -1.89495e-20 0.00139534 0.997818 8.59443e-05 0.152582 2.85189 0.00139534 0.997832 0.704575 0.00104996 0.00187994 0.000859443 0.455607 0.00187994 0.437918 0.00012847 1.02 0.887691 0.534677 0.286068 1.71682e-07 3.06183e-09 2387.13 3123.15 -0.0557302 0.482134 0.277553 0.25373 -0.593294 -0.169511 0.495954 -0.26786 -0.228104 1.677 1 0 297.384 0 2.0909 1.675 0.000299888 0.856319 0.655219 0.398696 0.41053 2.09112 131.449 83.8357 18.716 60.8254 0.0040288 0 -40 10
0.776 2.24844e-08 2.53894e-06 0.0980716 0.0980689 0.0120397 1.02202e-05 0.00115406 0.122589 0.000657636 0.123242 0.873867 101.84 0.244306 0.738587 4.16025 0.0556944 0.0392476 0.960752 0.0198299 0.0042778 0.0190927 0.00411316 0.00517012 0.00590725 0.206805 0.23629 57.9874 -87.8955 126.225 15.9719 145.016 0.000141544 0.267129 192.887 0.310609 0.0673762 0.00409553 0.000561727 0.00138298 0.986986 0.991732 -2.97552e-06 -85.6662 0.0930003 31190.9 301.491 0.983517 0.319147 0.734262 0.734257 9.99958 2.98164e-06 1.19264e-05 0.130997 0.981453 0.931357 -0.013293 4.90164e-06 0.502303 -1.89574e-20 6.9903e-24 -1.89504e-20 0.00139534 0.997818 8.59444e-05 0.152582 2.85189 0.00139534 0.997831 0.704678 0.00104998 0.00187994 0.000859444 0.455607 0.00187994 0.437926 0.000128473 1.02 0.887692 0.534677 0.286069 1.71682e-07 3.06185e-09 2387.11 3123.07 -0.0557258 0.482134 0.277553 0.253725 -0.593295 -0.169511 0.495967 -0.267858 -0.228118 1.678 1 0 297.389 0 2.09106 1.676 0.000299888 0.856287 0.65527 0.39851 0.410558 2.09129 131.458 83.8365 18.716 60.8258 0.00402877 0 -40 10
0.777 2.25133e-08 2.53894e-06 0.098144 0.0981414 0.0120397 1.02333e-05 0.00115406 0.12268 0.000657639 0.123333 0.87393 101.84 0.244298 0.738681 4.16044 0.0557019 0.0392495 0.960751 0.0198297 0.00427798 0.0190925 0.00411331 0.00517034 0.00590747 0.206814 0.236299 57.9875 -87.8955 126.225 15.9719 145.016 0.000141541 0.267129 192.887 0.310609 0.0673762 0.00409553 0.000561727 0.00138299 0.986986 0.991732 -2.97553e-06 -85.6662 0.0930004 31190.9 301.496 0.983517 0.319147 0.734244 0.73424 9.99958 2.98164e-06 1.19265e-05 0.130999 0.98146 0.931359 -0.013293 4.90167e-06 0.502311 -1.89582e-20 6.99066e-24 -1.89512e-20 0.00139534 0.997818 8.59444e-05 0.152582 2.85189 0.00139534 0.997831 0.704781 0.00105 0.00187994 0.000859444 0.455607 0.00187994 0.437935 0.000128476 1.02 0.887693 0.534677 0.286071 1.71682e-07 3.06187e-09 2387.1 3123 -0.0557215 0.482134 0.277552 0.253721 -0.593296 -0.169511 0.495979 -0.267855 -0.228132 1.679 1 0 297.393 0 2.09122 1.677 0.000299887 0.856256 0.655321 0.398325 0.410585 2.09145 131.467 83.8374 18.7161 60.8262 0.00402873 0 -40 10
0.778 2.25423e-08 2.53894e-06 0.0982164 0.0982138 0.0120397 1.02465e-05 0.00115406 0.122771 0.000657641 0.123424 0.873993 101.839 0.244291 0.738775 4.16063 0.0557094 0.0392513 0.960749 0.0198294 0.00427816 0.0190923 0.00411346 0.00517056 0.00590769 0.206822 0.236308 57.9875 -87.8955 126.226 15.9719 145.016 0.000141538 0.267129 192.887 0.310608 0.0673761 0.00409553 0.000561728 0.00138299 0.986986 0.991732 -2.97555e-06 -85.6662 0.0930005 31190.9 301.501 0.983517 0.319147 0.734227 0.734223 9.99958 2.98165e-06 1.19265e-05 0.131001 0.981466 0.931362 -0.013293 4.9017e-06 0.502318 -1.89591e-20 6.99101e-24 -1.89521e-20 0.00139534 0.997818 8.59445e-05 0.152583 2.85189 0.00139534 0.997831 0.704883 0.00105002 0.00187994 0.000859445 0.455606 0.00187994 0.437943 0.000128479 1.02 0.887694 0.534677 0.286072 1.71683e-07 3.0619e-09 2387.08 3122.93 -0.0557172 0.482135 0.277552 0.253716 -0.593297 -0.169511 0.495991 -0.267853 -0.228146 1.68 1 0 297.398 0 2.09139 1.678 0.000299887 0.856225 0.655372 0.39814 0.410612 2.09161 131.476 83.8382 18.7161 60.8267 0.0040287 0 -40 10
0.779 2.25712e-08 2.53894e-06 0.0982888 0.0982862 0.0120397 1.02596e-05 0.00115406 0.122861 0.000657644 0.123514 0.874056 101.839 0.244283 0.738868 4.16083 0.0557168 0.0392531 0.960747 0.0198292 0.00427834 0.0190921 0.00411361 0.00517078 0.00590791 0.206831 0.236317 57.9876 -87.8955 126.226 15.9718 145.016 0.000141534 0.26713 192.887 0.310608 0.0673761 0.00409554 0.000561729 0.00138299 0.986986 0.991732 -2.97556e-06 -85.6661 0.0930006 31190.9 301.506 0.983517 0.319147 0.73421 0.734206 9.99958 2.98165e-06 1.19265e-05 0.131003 0.981473 0.931364 -0.013293 4.90172e-06 0.502326 -1.89599e-20 6.99137e-24 -1.89529e-20 0.00139534 0.997818 8.59446e-05 0.152583 2.85189 0.00139534 0.997831 0.704986 0.00105004 0.00187994 0.000859446 0.455606 0.00187994 0.437951 0.000128483 1.02 0.887695 0.534676 0.286074 1.71683e-07 3.06192e-09 2387.06 3122.85 -0.0557129 0.482135 0.277552 0.253711 -0.593298 -0.169511 0.496003 -0.267851 -0.228161 1.681 1 0 297.403 0 2.09155 1.679 0.000299886 0.856194 0.655423 0.397955 0.41064 2.09178 131.484 83.8391 18.7162 60.8271 0.00402866 0 -40 10
0.78 2.26001e-08 2.53894e-06 0.0983611 0.0983585 0.0120397 1.02728e-05 0.00115406 0.122951 0.000657647 0.123604 0.874119 101.839 0.244276 0.738962 4.16102 0.0557243 0.0392549 0.960745 0.019829 0.00427852 0.0190919 0.00411376 0.00517101 0.00590813 0.20684 0.236325 57.9876 -87.8955 126.226 15.9718 145.016 0.000141531 0.26713 192.886 0.310607 0.067376 0.00409554 0.000561729 0.00138299 0.986986 0.991732 -2.97558e-06 -85.6661 0.0930006 31190.8 301.51 0.983517 0.319147 0.734193 0.734189 9.99958 2.98166e-06 1.19265e-05 0.131005 0.981479 0.931367 -0.013293 4.90175e-06 0.502333 -1.89608e-20 6.99172e-24 -1.89538e-20 0.00139535 0.997818 8.59447e-05 0.152583 2.8519 0.00139535 0.997831 0.705089 0.00105006 0.00187995 0.000859447 0.455606 0.00187994 0.43796 0.000128486 1.02 0.887696 0.534676 0.286075 1.71683e-07 3.06194e-09 2387.05 3122.78 -0.0557086 0.482135 0.277552 0.253707 -0.593298 -0.169511 0.496015 -0.267849 -0.228174 1.682 1 0 297.407 0 2.09171 1.68 0.000299886 0.856163 0.655475 0.397771 0.410667 2.09194 131.493 83.8399 18.7162 60.8275 0.00402863 0 -40 10
0.781 2.26291e-08 2.53894e-06 0.0984333 0.0984307 0.0120396 1.02859e-05 0.00115406 0.123042 0.000657649 0.123695 0.874182 101.839 0.244268 0.739056 4.16121 0.0557318 0.0392567 0.960743 0.0198288 0.0042787 0.0190916 0.00411391 0.00517123 0.00590836 0.206849 0.236334 57.9877 -87.8955 126.226 15.9717 145.016 0.000141528 0.26713 192.886 0.310607 0.067376 0.00409554 0.00056173 0.00138299 0.986986 0.991732 -2.97559e-06 -85.6661 0.0930007 31190.8 301.515 0.983517 0.319147 0.734176 0.734172 9.99958 2.98166e-06 1.19265e-05 0.131006 0.981485 0.931369 -0.013293 4.90178e-06 0.502341 -1.89616e-20 6.99207e-24 -1.89546e-20 0.00139535 0.997818 8.59447e-05 0.152583 2.8519 0.00139535 0.997831 0.705191 0.00105007 0.00187995 0.000859447 0.455606 0.00187995 0.437968 0.000128489 1.02 0.887697 0.534676 0.286077 1.71684e-07 3.06196e-09 2387.03 3122.71 -0.0557044 0.482135 0.277551 0.253702 -0.593299 -0.169512 0.496026 -0.267847 -0.228188 1.683 1 0 297.412 0 2.09188 1.681 0.000299886 0.856133 0.655526 0.397587 0.410694 2.0921 131.502 83.8408 18.7163 60.8279 0.00402859 0 -40 10
0.782 2.2658e-08 2.53894e-06 0.0985055 0.0985029 0.0120396 1.02991e-05 0.00115406 0.123132 0.000657652 0.123785 0.874246 101.839 0.244261 0.73915 4.16141 0.0557393 0.0392585 0.960741 0.0198285 0.00427888 0.0190914 0.00411406 0.00517145 0.00590858 0.206858 0.236343 57.9878 -87.8955 126.227 15.9717 145.016 0.000141525 0.26713 192.886 0.310607 0.0673759 0.00409555 0.000561731 0.001383 0.986986 0.991732 -2.97561e-06 -85.6661 0.0930008 31190.8 301.52 0.983517 0.319147 0.734159 0.734155 9.99958 2.98167e-06 1.19266e-05 0.131008 0.981492 0.931372 -0.013293 4.90181e-06 0.502349 -1.89624e-20 6.99243e-24 -1.89555e-20 0.00139535 0.997818 8.59448e-05 0.152583 2.8519 0.00139535 0.997831 0.705294 0.00105009 0.00187995 0.000859448 0.455605 0.00187995 0.437977 0.000128493 1.02 0.887699 0.534675 0.286078 1.71684e-07 3.06198e-09 2387.01 3122.63 -0.0557002 0.482135 0.277551 0.253698 -0.5933 -0.169512 0.496038 -0.267845 -0.228202 1.684 1 0 297.416 0 2.09204 1.682 0.000299885 0.856102 0.655577 0.397404 0.410722 2.09227 131.511 83.8416 18.7163 60.8283 0.00402856 0 -40 10
0.783 2.26869e-08 2.53894e-06 0.0985776 0.098575 0.0120396 1.03122e-05 0.00115406 0.123222 0.000657654 0.123875 0.874309 101.838 0.244253 0.739245 4.1616 0.0557468 0.0392604 0.96074 0.0198283 0.00427906 0.0190912 0.00411421 0.00517167 0.0059088 0.206867 0.236352 57.9878 -87.8955 126.227 15.9717 145.016 0.000141521 0.26713 192.886 0.310606 0.0673759 0.00409555 0.000561731 0.001383 0.986986 0.991732 -2.97562e-06 -85.6661 0.0930009 31190.8 301.525 0.983517 0.319147 0.734142 0.734138 9.99958 2.98167e-06 1.19266e-05 0.13101 0.981498 0.931374 -0.013293 4.90184e-06 0.502356 -1.89633e-20 6.99278e-24 -1.89563e-20 0.00139535 0.997818 8.59449e-05 0.152583 2.8519 0.00139535 0.997831 0.705397 0.00105011 0.00187995 0.000859449 0.455605 0.00187995 0.437985 0.000128496 1.02 0.8877 0.534675 0.28608 1.71684e-07 3.06201e-09 2387 3122.56 -0.055696 0.482135 0.277551 0.253693 -0.593301 -0.169512 0.49605 -0.267843 -0.228216 1.685 1 0 297.421 0 2.0922 1.683 0.000299885 0.856072 0.655628 0.397221 0.410749 2.09243 131.519 83.8424 18.7164 60.8287 0.00402852 0 -40 10
0.784 2.27159e-08 2.53894e-06 0.0986497 0.0986471 0.0120396 1.03254e-05 0.00115406 0.123312 0.000657657 0.123965 0.874372 101.838 0.244246 0.739339 4.16179 0.0557543 0.0392622 0.960738 0.0198281 0.00427924 0.019091 0.00411437 0.0051719 0.00590902 0.206876 0.236361 57.9879 -87.8955 126.227 15.9716 145.016 0.000141518 0.267131 192.886 0.310606 0.0673758 0.00409555 0.000561732 0.001383 0.986986 0.991732 -2.97564e-06 -85.6661 0.093001 31190.7 301.53 0.983517 0.319147 0.734126 0.734121 9.99958 2.98168e-06 1.19266e-05 0.131012 0.981504 0.931377 -0.013293 4.90187e-06 0.502364 -1.89641e-20 6.99314e-24 -1.89572e-20 0.00139535 0.997818 8.5945e-05 0.152583 2.8519 0.00139535 0.997831 0.705499 0.00105013 0.00187995 0.00085945 0.455605 0.00187995 0.437993 0.000128499 1.02 0.887701 0.534675 0.286081 1.71684e-07 3.06203e-09 2386.98 3122.49 -0.0556918 0.482135 0.27755 0.253689 -0.593302 -0.169512 0.496061 -0.267841 -0.228229 1.686 1 0 297.425 0 2.09237 1.684 0.000299885 0.856042 0.655679 0.397038 0.410776 2.09259 131.528 83.8432 18.7164 60.8291 0.00402849 0 -40 10
0.785 2.27448e-08 2.53894e-06 0.0987217 0.0987191 0.0120396 1.03386e-05 0.00115406 0.123402 0.000657659 0.124055 0.874436 101.838 0.244238 0.739433 4.16199 0.0557618 0.039264 0.960736 0.0198279 0.00427942 0.0190908 0.00411452 0.00517212 0.00590924 0.206885 0.23637 57.988 -87.8955 126.228 15.9716 145.016 0.000141515 0.267131 192.886 0.310605 0.0673758 0.00409555 0.000561732 0.001383 0.986986 0.991732 -2.97565e-06 -85.6661 0.0930011 31190.7 301.535 0.983517 0.319147 0.734109 0.734105 9.99958 2.98168e-06 1.19266e-05 0.131014 0.981511 0.931379 -0.013293 4.9019e-06 0.502371 -1.8965e-20 6.99349e-24 -1.8958e-20 0.00139535 0.997818 8.59451e-05 0.152584 2.8519 0.00139535 0.997831 0.705602 0.00105015 0.00187995 0.000859451 0.455605 0.00187995 0.438002 0.000128503 1.02 0.887702 0.534674 0.286083 1.71685e-07 3.06205e-09 2386.96 3122.42 -0.0556877 0.482135 0.27755 0.253684 -0.593303 -0.169512 0.496073 -0.267839 -0.228243 1.687 1 0 297.43 0 2.09253 1.685 0.000299884 0.856012 0.65573 0.396856 0.410804 2.09276 131.537 83.8441 18.7165 60.8295 0.00402846 0 -40 10
0.786 2.27737e-08 2.53894e-06 0.0987936 0.098791 0.0120396 1.03517e-05 0.00115407 0.123492 0.000657662 0.124145 0.874499 101.838 0.244231 0.739528 4.16218 0.0557693 0.0392659 0.960734 0.0198277 0.0042796 0.0190905 0.00411467 0.00517234 0.00590947 0.206894 0.236379 57.988 -87.8955 126.228 15.9716 145.016 0.000141512 0.267131 192.886 0.310605 0.0673757 0.00409556 0.000561733 0.001383 0.986986 0.991732 -2.97567e-06 -85.6661 0.0930012 31190.7 301.54 0.983517 0.319147 0.734093 0.734088 9.99958 2.98169e-06 1.19266e-05 0.131016 0.981517 0.931382 -0.013293 4.90193e-06 0.502379 -1.89658e-20 6.99385e-24 -1.89588e-20 0.00139535 0.997818 8.59451e-05 0.152584 2.8519 0.00139535 0.997831 0.705704 0.00105017 0.00187995 0.000859451 0.455605 0.00187995 0.43801 0.000128506 1.02 0.887703 0.534674 0.286084 1.71685e-07 3.06207e-09 2386.95 3122.35 -0.0556836 0.482135 0.27755 0.25368 -0.593303 -0.169512 0.496084 -0.267837 -0.228256 1.688 1 0 297.434 0 2.09269 1.686 0.000299884 0.855983 0.655781 0.396674 0.410831 2.09292 131.546 83.8449 18.7165 60.8299 0.00402842 0 -40 10
0.787 2.28027e-08 2.53894e-06 0.0988655 0.0988629 0.0120396 1.03649e-05 0.00115407 0.123582 0.000657665 0.124235 0.874562 101.838 0.244223 0.739622 4.16238 0.0557768 0.0392677 0.960732 0.0198274 0.00427979 0.0190903 0.00411482 0.00517257 0.00590969 0.206903 0.236388 57.9881 -87.8955 126.228 15.9715 145.016 0.000141509 0.267131 192.885 0.310605 0.0673757 0.00409556 0.000561734 0.00138301 0.986986 0.991732 -2.97568e-06 -85.6661 0.0930012 31190.7 301.545 0.983517 0.319147 0.734076 0.734072 9.99958 2.98169e-06 1.19267e-05 0.131018 0.981523 0.931384 -0.013293 4.90196e-06 0.502387 -1.89667e-20 6.99421e-24 -1.89597e-20 0.00139535 0.997818 8.59452e-05 0.152584 2.8519 0.00139535 0.997831 0.705806 0.00105019 0.00187996 0.000859452 0.455604 0.00187995 0.438019 0.000128509 1.02 0.887704 0.534674 0.286086 1.71685e-07 3.0621e-09 2386.93 3122.28 -0.0556796 0.482135 0.27755 0.253675 -0.593304 -0.169512 0.496095 -0.267835 -0.22827 1.689 1 0 297.439 0 2.09286 1.687 0.000299883 0.855953 0.655832 0.396493 0.410858 2.09308 131.554 83.8457 18.7166 60.8302 0.00402839 0 -40 10
0.788 2.28316e-08 2.53894e-06 0.0989373 0.0989348 0.0120396 1.0378e-05 0.00115407 0.123672 0.000657667 0.124325 0.874626 101.837 0.244216 0.739717 4.16258 0.0557844 0.0392696 0.96073 0.0198272 0.00427997 0.0190901 0.00411498 0.00517279 0.00590991 0.206912 0.236397 57.9882 -87.8955 126.229 15.9715 145.016 0.000141506 0.267131 192.885 0.310604 0.0673756 0.00409556 0.000561734 0.00138301 0.986986 0.991732 -2.97569e-06 -85.6661 0.0930013 31190.7 301.55 0.983517 0.319147 0.73406 0.734056 9.99958 2.9817e-06 1.19267e-05 0.13102 0.981529 0.931387 -0.013293 4.90199e-06 0.502394 -1.89675e-20 6.99456e-24 -1.89605e-20 0.00139535 0.997818 8.59453e-05 0.152584 2.8519 0.00139535 0.99783 0.705909 0.00105021 0.00187996 0.000859453 0.455604 0.00187996 0.438027 0.000128512 1.02 0.887705 0.534674 0.286087 1.71685e-07 3.06212e-09 2386.91 3122.21 -0.0556756 0.482135 0.277549 0.253671 -0.593305 -0.169512 0.496106 -0.267833 -0.228283 1.69 1 0 297.443 0 2.09302 1.688 0.000299883 0.855924 0.655883 0.396312 0.410886 2.09324 131.563 83.8465 18.7166 60.8306 0.00402836 0 -40 10
0.789 2.28606e-08 2.53894e-06 0.0990091 0.0990066 0.0120395 1.03912e-05 0.00115407 0.123761 0.00065767 0.124414 0.874689 101.837 0.244208 0.739811 4.16277 0.0557919 0.0392714 0.960729 0.019827 0.00428015 0.0190899 0.00411513 0.00517302 0.00591014 0.206921 0.236406 57.9882 -87.8955 126.229 15.9714 145.016 0.000141502 0.267132 192.885 0.310604 0.0673756 0.00409557 0.000561735 0.00138301 0.986986 0.991732 -2.97571e-06 -85.6661 0.0930014 31190.6 301.555 0.983517 0.319147 0.734044 0.734039 9.99958 2.9817e-06 1.19267e-05 0.131021 0.981536 0.931389 -0.013293 4.90201e-06 0.502402 -1.89684e-20 6.99492e-24 -1.89614e-20 0.00139536 0.997818 8.59454e-05 0.152584 2.8519 0.00139536 0.99783 0.706011 0.00105023 0.00187996 0.000859454 0.455604 0.00187996 0.438035 0.000128516 1.02 0.887706 0.534673 0.286089 1.71686e-07 3.06214e-09 2386.9 3122.14 -0.0556716 0.482135 0.277549 0.253667 -0.593306 -0.169512 0.496117 -0.267831 -0.228296 1.691 1 0 297.447 0 2.09318 1.689 0.000299883 0.855895 0.655934 0.396132 0.410913 2.09341 131.572 83.8473 18.7167 60.831 0.00402832 0 -40 10
0.79 2.28895e-08 2.53895e-06 0.0990808 0.0990783 0.0120395 1.04043e-05 0.00115407 0.123851 0.000657672 0.124504 0.874753 101.837 0.244201 0.739906 4.16297 0.0557995 0.0392733 0.960727 0.0198268 0.00428034 0.0190896 0.00411528 0.00517325 0.00591036 0.20693 0.236415 57.9883 -87.8955 126.229 15.9714 145.016 0.000141499 0.267132 192.885 0.310603 0.0673755 0.00409557 0.000561736 0.00138301 0.986986 0.991732 -2.97572e-06 -85.666 0.0930015 31190.6 301.56 0.983517 0.319147 0.734028 0.734023 9.99958 2.98171e-06 1.19267e-05 0.131023 0.981542 0.931391 -0.013293 4.90204e-06 0.50241 -1.89692e-20 6.99527e-24 -1.89622e-20 0.00139536 0.997818 8.59454e-05 0.152584 2.8519 0.00139536 0.99783 0.706113 0.00105025 0.00187996 0.000859454 0.455604 0.00187996 0.438044 0.000128519 1.02 0.887707 0.534673 0.28609 1.71686e-07 3.06216e-09 2386.88 3122.07 -0.0556676 0.482135 0.277549 0.253662 -0.593307 -0.169512 0.496128 -0.267828 -0.228309 1.692 1 0 297.452 0 2.09334 1.69 0.000299882 0.855866 0.655985 0.395952 0.41094 2.09357 131.58 83.8481 18.7167 60.8314 0.00402829 0 -40 10
0.791 2.29184e-08 2.53895e-06 0.0991525 0.0991499 0.0120395 1.04175e-05 0.00115407 0.123941 0.000657675 0.124594 0.874817 101.837 0.244193 0.740001 4.16317 0.055807 0.0392751 0.960725 0.0198265 0.00428052 0.0190894 0.00411544 0.00517347 0.00591059 0.206939 0.236424 57.9883 -87.8955 126.229 15.9714 145.016 0.000141496 0.267132 192.885 0.310603 0.0673755 0.00409557 0.000561736 0.00138302 0.986986 0.991732 -2.97574e-06 -85.666 0.0930016 31190.6 301.565 0.983517 0.319147 0.734012 0.734007 9.99958 2.98171e-06 1.19267e-05 0.131025 0.981548 0.931394 -0.013293 4.90207e-06 0.502417 -1.89701e-20 6.99563e-24 -1.89631e-20 0.00139536 0.997818 8.59455e-05 0.152584 2.85191 0.00139536 0.99783 0.706216 0.00105027 0.00187996 0.000859455 0.455603 0.00187996 0.438052 0.000128522 1.02 0.887708 0.534673 0.286092 1.71686e-07 3.06219e-09 2386.86 3122 -0.0556637 0.482136 0.277548 0.253658 -0.593307 -0.169512 0.496139 -0.267826 -0.228322 1.693 1 0 297.456 0 2.09351 1.691 0.000299882 0.855837 0.656036 0.395772 0.410967 2.09373 131.589 83.8489 18.7167 60.8318 0.00402826 0 -40 10
0.792 2.29474e-08 2.53895e-06 0.0992241 0.0992215 0.0120395 1.04306e-05 0.00115407 0.12403 0.000657677 0.124683 0.87488 101.837 0.244185 0.740096 4.16336 0.0558146 0.039277 0.960723 0.0198263 0.00428071 0.0190892 0.00411559 0.0051737 0.00591081 0.206948 0.236433 57.9884 -87.8955 126.23 15.9713 145.016 0.000141493 0.267132 192.885 0.310602 0.0673754 0.00409557 0.000561737 0.00138302 0.986986 0.991732 -2.97575e-06 -85.666 0.0930017 31190.6 301.57 0.983517 0.319147 0.733996 0.733991 9.99958 2.98171e-06 1.19268e-05 0.131027 0.981554 0.931396 -0.013293 4.9021e-06 0.502425 -1.89709e-20 6.99599e-24 -1.8964e-20 0.00139536 0.997818 8.59456e-05 0.152585 2.85191 0.00139536 0.99783 0.706318 0.00105029 0.00187996 0.000859456 0.455603 0.00187996 0.43806 0.000128526 1.02 0.887709 0.534672 0.286093 1.71686e-07 3.06221e-09 2386.85 3121.93 -0.0556597 0.482136 0.277548 0.253654 -0.593308 -0.169512 0.49615 -0.267824 -0.228335 1.694 1 0 297.46 0 2.09367 1.692 0.000299882 0.855808 0.656087 0.395593 0.410994 2.09389 131.598 83.8497 18.7168 60.8322 0.00402823 0 -40 10
0.793 2.29763e-08 2.53895e-06 0.0992956 0.0992931 0.0120395 1.04438e-05 0.00115407 0.124119 0.00065768 0.124773 0.874944 101.836 0.244178 0.740191 4.16356 0.0558221 0.0392789 0.960721 0.0198261 0.00428089 0.019089 0.00411574 0.00517393 0.00591104 0.206957 0.236442 57.9885 -87.8955 126.23 15.9713 145.016 0.00014149 0.267132 192.884 0.310602 0.0673754 0.00409558 0.000561738 0.00138302 0.986986 0.991732 -2.97577e-06 -85.666 0.0930017 31190.5 301.575 0.983517 0.319147 0.73398 0.733976 9.99958 2.98172e-06 1.19268e-05 0.131029 0.98156 0.931399 -0.013293 4.90213e-06 0.502433 -1.89718e-20 6.99634e-24 -1.89648e-20 0.00139536 0.997818 8.59457e-05 0.152585 2.85191 0.00139536 0.99783 0.70642 0.00105031 0.00187996 0.000859457 0.455603 0.00187996 0.438069 0.000128529 1.02 0.88771 0.534672 0.286095 1.71687e-07 3.06223e-09 2386.83 3121.86 -0.0556559 0.482136 0.277548 0.253649 -0.593309 -0.169512 0.496161 -0.267822 -0.228348 1.695 1 0 297.464 0 2.09383 1.693 0.000299881 0.85578 0.656138 0.395414 0.411022 2.09406 131.607 83.8504 18.7168 60.8325 0.00402819 0 -40 10
0.794 2.30052e-08 2.53895e-06 0.0993671 0.0993646 0.0120395 1.04569e-05 0.00115407 0.124209 0.000657682 0.124862 0.875008 101.836 0.24417 0.740286 4.16376 0.0558297 0.0392808 0.960719 0.0198258 0.00428108 0.0190887 0.0041159 0.00517415 0.00591127 0.206966 0.236451 57.9885 -87.8955 126.23 15.9713 145.016 0.000141487 0.267132 192.884 0.310602 0.0673753 0.00409558 0.000561738 0.00138302 0.986986 0.991732 -2.97578e-06 -85.666 0.0930018 31190.5 301.58 0.983517 0.319147 0.733964 0.73396 9.99958 2.98172e-06 1.19268e-05 0.131031 0.981566 0.931401 -0.013293 4.90216e-06 0.502441 -1.89727e-20 6.9967e-24 -1.89657e-20 0.00139536 0.997818 8.59458e-05 0.152585 2.85191 0.00139536 0.99783 0.706522 0.00105033 0.00187997 0.000859458 0.455603 0.00187996 0.438077 0.000128532 1.02 0.887711 0.534672 0.286096 1.71687e-07 3.06225e-09 2386.81 3121.8 -0.055652 0.482136 0.277548 0.253645 -0.59331 -0.169512 0.496172 -0.26782 -0.228361 1.696 1 0 297.468 0 2.09399 1.694 0.000299881 0.855752 0.656189 0.395235 0.411049 2.09422 131.615 83.8512 18.7169 60.8329 0.00402816 0 -40 10
0.795 2.30342e-08 2.53895e-06 0.0994385 0.099436 0.0120395 1.04701e-05 0.00115407 0.124298 0.000657685 0.124951 0.875072 101.836 0.244163 0.740381 4.16396 0.0558372 0.0392826 0.960717 0.0198256 0.00428126 0.0190885 0.00411605 0.00517438 0.00591149 0.206975 0.23646 57.9886 -87.8955 126.231 15.9712 145.016 0.000141484 0.267133 192.884 0.310601 0.0673753 0.00409558 0.000561739 0.00138302 0.986986 0.991732 -2.9758e-06 -85.666 0.0930019 31190.5 301.585 0.983517 0.319147 0.733949 0.733944 9.99958 2.98173e-06 1.19268e-05 0.131033 0.981573 0.931403 -0.013293 4.90219e-06 0.502448 -1.89735e-20 6.99706e-24 -1.89665e-20 0.00139536 0.997818 8.59458e-05 0.152585 2.85191 0.00139536 0.99783 0.706624 0.00105035 0.00187997 0.000859458 0.455603 0.00187997 0.438085 0.000128536 1.02 0.887713 0.534671 0.286098 1.71687e-07 3.06227e-09 2386.8 3121.73 -0.0556482 0.482136 0.277547 0.253641 -0.593311 -0.169512 0.496182 -0.267818 -0.228373 1.697 1 0 297.473 0 2.09416 1.695 0.00029988 0.855724 0.65624 0.395058 0.411076 2.09438 131.624 83.852 18.7169 60.8333 0.00402813 0 -40 10
0.796 2.30631e-08 2.53895e-06 0.0995099 0.0995074 0.0120394 1.04832e-05 0.00115407 0.124387 0.000657687 0.12504 0.875135 101.836 0.244155 0.740476 4.16416 0.0558448 0.0392845 0.960715 0.0198254 0.00428145 0.0190883 0.00411621 0.00517461 0.00591172 0.206984 0.236469 57.9887 -87.8955 126.231 15.9712 145.016 0.000141481 0.267133 192.884 0.310601 0.0673752 0.00409559 0.00056174 0.00138303 0.986986 0.991732 -2.97581e-06 -85.666 0.093002 31190.5 301.59 0.983517 0.319147 0.733933 0.733929 9.99958 2.98173e-06 1.19268e-05 0.131035 0.981579 0.931406 -0.013293 4.90222e-06 0.502456 -1.89744e-20 6.99741e-24 -1.89674e-20 0.00139536 0.997818 8.59459e-05 0.152585 2.85191 0.00139536 0.99783 0.706726 0.00105037 0.00187997 0.000859459 0.455602 0.00187997 0.438094 0.000128539 1.02 0.887714 0.534671 0.286099 1.71687e-07 3.0623e-09 2386.78 3121.66 -0.0556444 0.482136 0.277547 0.253637 -0.593311 -0.169512 0.496193 -0.267816 -0.228386 1.698 1 0 297.477 0 2.09432 1.696 0.00029988 0.855696 0.65629 0.39488 0.411103 2.09454 131.633 83.8528 18.717 60.8337 0.0040281 0 -40 10
0.797 2.3092e-08 2.53895e-06 0.0995812 0.0995787 0.0120394 1.04964e-05 0.00115407 0.124476 0.00065769 0.12513 0.875199 101.836 0.244148 0.740571 4.16436 0.0558524 0.0392864 0.960714 0.0198252 0.00428163 0.0190881 0.00411636 0.00517484 0.00591195 0.206994 0.236478 57.9887 -87.8956 126.231 15.9711 145.016 0.000141478 0.267133 192.884 0.3106 0.0673752 0.00409559 0.00056174 0.00138303 0.986986 0.991732 -2.97583e-06 -85.666 0.0930021 31190.5 301.595 0.983517 0.319147 0.733917 0.733913 9.99958 2.98174e-06 1.19268e-05 0.131037 0.981585 0.931408 -0.013293 4.90225e-06 0.502464 -1.89752e-20 6.99777e-24 -1.89682e-20 0.00139536 0.997818 8.5946e-05 0.152585 2.85191 0.00139536 0.99783 0.706829 0.00105039 0.00187997 0.00085946 0.455602 0.00187997 0.438102 0.000128542 1.02 0.887715 0.534671 0.286101 1.71688e-07 3.06232e-09 2386.76 3121.6 -0.0556406 0.482136 0.277547 0.253633 -0.593312 -0.169513 0.496203 -0.267814 -0.228398 1.699 1 0 297.481 0 2.09448 1.697 0.00029988 0.855668 0.656341 0.394703 0.41113 2.09471 131.641 83.8535 18.717 60.834 0.00402807 0 -40 10
0.798 2.3121e-08 2.53895e-06 0.0996524 0.09965 0.0120394 1.05095e-05 0.00115407 0.124566 0.000657692 0.125219 0.875263 101.835 0.24414 0.740666 4.16456 0.05586 0.0392883 0.960712 0.0198249 0.00428182 0.0190878 0.00411652 0.00517507 0.00591218 0.207003 0.236487 57.9888 -87.8956 126.231 15.9711 145.016 0.000141475 0.267133 192.884 0.3106 0.0673751 0.00409559 0.000561741 0.00138303 0.986986 0.991732 -2.97584e-06 -85.666 0.0930022 31190.4 301.6 0.983517 0.319147 0.733902 0.733898 9.99958 2.98174e-06 1.19269e-05 0.131038 0.981591 0.93141 -0.013293 4.90228e-06 0.502472 -1.89761e-20 6.99813e-24 -1.89691e-20 0.00139537 0.997818 8.59461e-05 0.152586 2.85191 0.00139537 0.99783 0.706931 0.00105041 0.00187997 0.000859461 0.455602 0.00187997 0.43811 0.000128545 1.02 0.887716 0.534671 0.286102 1.71688e-07 3.06234e-09 2386.74 3121.53 -0.0556369 0.482136 0.277546 0.253628 -0.593313 -0.169513 0.496213 -0.267812 -0.228411 1.7 1 0 297.485 0 2.09464 1.698 0.000299879 0.85564 0.656392 0.394526 0.411157 2.09487 131.65 83.8543 18.7171 60.8344 0.00402803 0 -40 10
0.799 2.31499e-08 2.53895e-06 0.0997236 0.0997212 0.0120394 1.05227e-05 0.00115407 0.124655 0.000657695 0.125308 0.875327 101.835 0.244132 0.740762 4.16476 0.0558676 0.0392902 0.96071 0.0198247 0.00428201 0.0190876 0.00411668 0.0051753 0.00591241 0.207012 0.236496 57.9889 -87.8956 126.232 15.9711 145.016 0.000141472 0.267133 192.883 0.3106 0.0673751 0.0040956 0.000561742 0.00138303 0.986986 0.991732 -2.97585e-06 -85.666 0.0930023 31190.4 301.605 0.983517 0.319147 0.733887 0.733882 9.99958 2.98175e-06 1.19269e-05 0.13104 0.981597 0.931413 -0.013293 4.90231e-06 0.50248 -1.89769e-20 6.99849e-24 -1.89699e-20 0.00139537 0.997818 8.59461e-05 0.152586 2.85191 0.00139537 0.99783 0.707033 0.00105043 0.00187997 0.000859461 0.455602 0.00187997 0.438119 0.000128549 1.02 0.887717 0.53467 0.286104 1.71688e-07 3.06236e-09 2386.73 3121.46 -0.0556332 0.482136 0.277546 0.253624 -0.593314 -0.169513 0.496223 -0.26781 -0.228423 1.701 1 0 297.489 0 2.09481 1.699 0.000299879 0.855613 0.656443 0.39435 0.411185 2.09503 131.659 83.855 18.7171 60.8348 0.004028 0 -40 10
0.8 2.31789e-08 2.53895e-06 0.0997948 0.0997923 0.0120394 1.05358e-05 0.00115407 0.124743 0.000657697 0.125397 0.875391 101.835 0.244125 0.740857 4.16496 0.0558752 0.0392921 0.960708 0.0198245 0.00428219 0.0190874 0.00411683 0.00517553 0.00591263 0.207021 0.236505 57.9889 -87.8956 126.232 15.971 145.016 0.000141469 0.267134 192.883 0.310599 0.067375 0.0040956 0.000561742 0.00138303 0.986986 0.991732 -2.97587e-06 -85.666 0.0930023 31190.4 301.61 0.983517 0.319147 0.733872 0.733867 9.99958 2.98175e-06 1.19269e-05 0.131042 0.981603 0.931415 -0.013293 4.90233e-06 0.502487 -1.89778e-20 6.99885e-24 -1.89708e-20 0.00139537 0.997818 8.59462e-05 0.152586 2.85191 0.00139537 0.997829 0.707134 0.00105045 0.00187997 0.000859462 0.455602 0.00187997 0.438127 0.000128552 1.02 0.887718 0.53467 0.286105 1.71688e-07 3.06239e-09 2386.71 3121.4 -0.0556295 0.482136 0.277546 0.25362 -0.593314 -0.169513 0.496234 -0.267808 -0.228435 1.702 1 0 297.493 0 2.09497 1.7 0.000299878 0.855586 0.656494 0.394174 0.411212 2.09519 131.667 83.8558 18.7171 60.8351 0.00402797 0 -40 10
0.801 2.32078e-08 2.53895e-06 0.0998659 0.0998634 0.0120394 1.0549e-05 0.00115407 0.124832 0.0006577 0.125485 0.875455 101.835 0.244117 0.740953 4.16516 0.0558828 0.039294 0.960706 0.0198242 0.00428238 0.0190871 0.00411699 0.00517576 0.00591286 0.20703 0.236515 57.989 -87.8956 126.232 15.971 145.016 0.000141466 0.267134 192.883 0.310599 0.067375 0.0040956 0.000561743 0.00138304 0.986986 0.991732 -2.97588e-06 -85.6659 0.0930024 31190.4 301.615 0.983517 0.319147 0.733856 0.733852 9.99958 2.98176e-06 1.19269e-05 0.131044 0.981609 0.931417 -0.013293 4.90236e-06 0.502495 -1.89786e-20 6.9992e-24 -1.89716e-20 0.00139537 0.997818 8.59463e-05 0.152586 2.85191 0.00139537 0.997829 0.707236 0.00105046 0.00187998 0.000859463 0.455601 0.00187997 0.438135 0.000128555 1.02 0.887719 0.53467 0.286107 1.71689e-07 3.06241e-09 2386.69 3121.33 -0.0556258 0.482136 0.277546 0.253616 -0.593315 -0.169513 0.496244 -0.267805 -0.228447 1.703 1 0 297.497 0 2.09513 1.701 0.000299878 0.855559 0.656544 0.393998 0.411239 2.09535 131.676 83.8565 18.7172 60.8355 0.00402794 0 -40 10
0.802 2.32367e-08 2.53895e-06 0.0999369 0.0999344 0.0120394 1.05621e-05 0.00115407 0.124921 0.000657702 0.125574 0.87552 101.835 0.24411 0.741048 4.16536 0.0558904 0.0392959 0.960704 0.019824 0.00428257 0.0190869 0.00411715 0.00517599 0.00591309 0.207039 0.236524 57.989 -87.8956 126.233 15.9709 145.016 0.000141463 0.267134 192.883 0.310598 0.0673749 0.0040956 0.000561744 0.00138304 0.986986 0.991732 -2.9759e-06 -85.6659 0.0930025 31190.4 301.62 0.983517 0.319147 0.733841 0.733837 9.99958 2.98176e-06 1.19269e-05 0.131046 0.981615 0.931419 -0.013293 4.90239e-06 0.502503 -1.89795e-20 6.99956e-24 -1.89725e-20 0.00139537 0.997818 8.59464e-05 0.152586 2.85191 0.00139537 0.997829 0.707338 0.00105048 0.00187998 0.000859464 0.455601 0.00187998 0.438144 0.000128559 1.02 0.88772 0.534669 0.286108 1.71689e-07 3.06243e-09 2386.68 3121.27 -0.0556222 0.482136 0.277545 0.253612 -0.593316 -0.169513 0.496254 -0.267803 -0.228459 1.704 1 0 297.501 0 2.09529 1.702 0.000299878 0.855532 0.656595 0.393823 0.411266 2.09552 131.685 83.8573 18.7172 60.8358 0.00402791 0 -40 10
0.803 2.32657e-08 2.53895e-06 0.100008 0.100005 0.0120394 1.05753e-05 0.00115407 0.12501 0.000657705 0.125663 0.875584 101.834 0.244102 0.741144 4.16556 0.055898 0.0392978 0.960702 0.0198238 0.00428276 0.0190867 0.0041173 0.00517622 0.00591332 0.207049 0.236533 57.9891 -87.8956 126.233 15.9709 145.016 0.000141461 0.267134 192.883 0.310598 0.0673749 0.00409561 0.000561744 0.00138304 0.986985 0.991732 -2.97591e-06 -85.6659 0.0930026 31190.3 301.625 0.983517 0.319147 0.733826 0.733822 9.99958 2.98177e-06 1.1927e-05 0.131048 0.981621 0.931422 -0.013293 4.90242e-06 0.502511 -1.89804e-20 6.99992e-24 -1.89734e-20 0.00139537 0.997818 8.59465e-05 0.152586 2.85192 0.00139537 0.997829 0.70744 0.0010505 0.00187998 0.000859465 0.455601 0.00187998 0.438152 0.000128562 1.02 0.887721 0.534669 0.28611 1.71689e-07 3.06245e-09 2386.66 3121.2 -0.0556186 0.482136 0.277545 0.253608 -0.593317 -0.169513 0.496263 -0.267801 -0.228471 1.705 1 0 297.505 0 2.09545 1.703 0.000299877 0.855505 0.656646 0.393648 0.411293 2.09568 131.693 83.858 18.7173 60.8362 0.00402788 0 -40 10
0.804 2.32946e-08 2.53895e-06 0.100079 0.100076 0.0120393 1.05885e-05 0.00115407 0.125098 0.000657707 0.125752 0.875648 101.834 0.244094 0.74124 4.16577 0.0559057 0.0392997 0.9607 0.0198236 0.00428294 0.0190864 0.00411746 0.00517645 0.00591355 0.207058 0.236542 57.9892 -87.8956 126.233 15.9709 145.016 0.000141458 0.267134 192.883 0.310597 0.0673748 0.00409561 0.000561745 0.00138304 0.986985 0.991732 -2.97593e-06 -85.6659 0.0930027 31190.3 301.63 0.983517 0.319147 0.733812 0.733807 9.99958 2.98177e-06 1.1927e-05 0.13105 0.981627 0.931424 -0.013293 4.90245e-06 0.502519 -1.89812e-20 7.00028e-24 -1.89742e-20 0.00139537 0.997818 8.59465e-05 0.152586 2.85192 0.00139537 0.997829 0.707542 0.00105052 0.00187998 0.000859465 0.455601 0.00187998 0.43816 0.000128565 1.02 0.887722 0.534669 0.286111 1.7169e-07 3.06248e-09 2386.64 3121.14 -0.055615 0.482136 0.277545 0.253604 -0.593317 -0.169513 0.496273 -0.267799 -0.228483 1.706 1 0 297.509 0 2.09562 1.704 0.000299877 0.855479 0.656697 0.393474 0.41132 2.09584 131.702 83.8588 18.7173 60.8365 0.00402785 0 -40 10
0.805 2.33235e-08 2.53895e-06 0.10015 0.100147 0.0120393 1.06016e-05 0.00115407 0.125187 0.00065771 0.12584 0.875712 101.834 0.244087 0.741336 4.16597 0.0559133 0.0393016 0.960698 0.0198233 0.00428313 0.0190862 0.00411762 0.00517668 0.00591379 0.207067 0.236551 57.9892 -87.8956 126.233 15.9708 145.017 0.000141455 0.267135 192.882 0.310597 0.0673748 0.00409561 0.000561745 0.00138304 0.986985 0.991732 -2.97594e-06 -85.6659 0.0930028 31190.3 301.636 0.983517 0.319147 0.733797 0.733792 9.99958 2.98178e-06 1.1927e-05 0.131052 0.981632 0.931426 -0.013293 4.90248e-06 0.502527 -1.89821e-20 7.00064e-24 -1.89751e-20 0.00139537 0.997818 8.59466e-05 0.152587 2.85192 0.00139537 0.997829 0.707644 0.00105054 0.00187998 0.000859466 0.4556 0.00187998 0.438169 0.000128568 1.02 0.887723 0.534668 0.286113 1.7169e-07 3.0625e-09 2386.63 3121.08 -0.0556115 0.482137 0.277544 0.2536 -0.593318 -0.169513 0.496283 -0.267797 -0.228495 1.707 1 0 297.513 0 2.09578 1.705 0.000299876 0.855452 0.656747 0.3933 0.411347 2.096 131.711 83.8595 18.7174 60.8369 0.00402782 0 -40 10
0.806 2.33525e-08 2.53895e-06 0.10022 0.100218 0.0120393 1.06148e-05 0.00115407 0.125276 0.000657712 0.125929 0.875777 101.834 0.244079 0.741432 4.16617 0.0559209 0.0393035 0.960696 0.0198231 0.00428332 0.019086 0.00411778 0.00517691 0.00591402 0.207077 0.236561 57.9893 -87.8956 126.234 15.9708 145.017 0.000141452 0.267135 192.882 0.310597 0.0673747 0.00409562 0.000561746 0.00138305 0.986985 0.991732 -2.97596e-06 -85.6659 0.0930028 31190.3 301.641 0.983517 0.319147 0.733782 0.733778 9.99958 2.98178e-06 1.1927e-05 0.131054 0.981638 0.931428 -0.013293 4.90251e-06 0.502535 -1.89829e-20 7.001e-24 -1.89759e-20 0.00139537 0.997818 8.59467e-05 0.152587 2.85192 0.00139537 0.997829 0.707745 0.00105056 0.00187998 0.000859467 0.4556 0.00187998 0.438177 0.000128572 1.02 0.887724 0.534668 0.286114 1.7169e-07 3.06252e-09 2386.61 3121.01 -0.055608 0.482137 0.277544 0.253596 -0.593319 -0.169513 0.496293 -0.267795 -0.228507 1.708 1 0 297.516 0 2.09594 1.706 0.000299876 0.855426 0.656798 0.393127 0.411374 2.09616 131.719 83.8602 18.7174 60.8372 0.00402779 0 -40 10
0.807 2.33814e-08 2.53895e-06 0.100291 0.100289 0.0120393 1.06279e-05 0.00115407 0.125364 0.000657714 0.126017 0.875841 101.834 0.244071 0.741527 4.16637 0.0559286 0.0393054 0.960695 0.0198229 0.00428351 0.0190858 0.00411794 0.00517715 0.00591425 0.207086 0.23657 57.9894 -87.8956 126.234 15.9708 145.017 0.000141449 0.267135 192.882 0.310596 0.0673747 0.00409562 0.000561747 0.00138305 0.986985 0.991732 -2.97597e-06 -85.6659 0.0930029 31190.2 301.646 0.983517 0.319147 0.733767 0.733763 9.99958 2.98179e-06 1.1927e-05 0.131056 0.981644 0.931431 -0.013293 4.90254e-06 0.502543 -1.89838e-20 7.00136e-24 -1.89768e-20 0.00139538 0.997818 8.59468e-05 0.152587 2.85192 0.00139538 0.997829 0.707847 0.00105058 0.00187998 0.000859468 0.4556 0.00187998 0.438185 0.000128575 1.02 0.887725 0.534668 0.286116 1.7169e-07 3.06254e-09 2386.59 3120.95 -0.0556045 0.482137 0.277544 0.253592 -0.593319 -0.169513 0.496302 -0.267793 -0.228518 1.709 1 0 297.52 0 2.0961 1.707 0.000299876 0.8554 0.656848 0.392953 0.411401 2.09632 131.728 83.8609 18.7174 60.8376 0.00402776 0 -40 10
0.808 2.34103e-08 2.53895e-06 0.100362 0.100359 0.0120393 1.06411e-05 0.00115407 0.125452 0.000657717 0.126105 0.875905 101.833 0.244064 0.741624 4.16658 0.0559362 0.0393073 0.960693 0.0198226 0.0042837 0.0190855 0.00411809 0.00517738 0.00591448 0.207095 0.236579 57.9894 -87.8956 126.234 15.9707 145.017 0.000141446 0.267135 192.882 0.310596 0.0673746 0.00409562 0.000561747 0.00138305 0.986985 0.991732 -2.97599e-06 -85.6659 0.093003 31190.2 301.651 0.983517 0.319147 0.733753 0.733749 9.99958 2.98179e-06 1.19271e-05 0.131058 0.98165 0.931433 -0.013293 4.90257e-06 0.502551 -1.89847e-20 7.00172e-24 -1.89777e-20 0.00139538 0.997818 8.59469e-05 0.152587 2.85192 0.00139538 0.997829 0.707949 0.0010506 0.00187999 0.000859469 0.4556 0.00187999 0.438194 0.000128578 1.02 0.887727 0.534668 0.286117 1.71691e-07 3.06257e-09 2386.58 3120.89 -0.055601 0.482137 0.277544 0.253588 -0.59332 -0.169513 0.496312 -0.267791 -0.22853 1.71 1 0 297.524 0 2.09626 1.708 0.000299875 0.855374 0.656899 0.392781 0.411428 2.09649 131.737 83.8617 18.7175 60.8379 0.00402773 0 -40 10
0.809 2.34393e-08 2.53895e-06 0.100432 0.10043 0.0120393 1.06542e-05 0.00115407 0.125541 0.000657719 0.126194 0.87597 101.833 0.244056 0.74172 4.16678 0.0559439 0.0393093 0.960691 0.0198224 0.00428389 0.0190853 0.00411825 0.00517761 0.00591471 0.207105 0.236589 57.9895 -87.8956 126.234 15.9707 145.017 0.000141444 0.267135 192.882 0.310595 0.0673746 0.00409562 0.000561748 0.00138305 0.986985 0.991731 -2.976e-06 -85.6659 0.0930031 31190.2 301.656 0.983517 0.319147 0.733738 0.733734 9.99958 2.9818e-06 1.19271e-05 0.13106 0.981656 0.931435 -0.013293 4.9026e-06 0.502559 -1.89855e-20 7.00208e-24 -1.89785e-20 0.00139538 0.997818 8.59469e-05 0.152587 2.85192 0.00139538 0.997829 0.70805 0.00105062 0.00187999 0.000859469 0.4556 0.00187999 0.438202 0.000128581 1.02 0.887728 0.534667 0.286119 1.71691e-07 3.06259e-09 2386.56 3120.83 -0.0555976 0.482137 0.277543 0.253584 -0.593321 -0.169513 0.496321 -0.267789 -0.228541 1.711 1 0 297.528 0 2.09642 1.709 0.000299875 0.855348 0.65695 0.392608 0.411455 2.09665 131.745 83.8624 18.7175 60.8383 0.0040277 0 -40 10
0.81 2.34682e-08 2.53895e-06 0.100503 0.100501 0.0120393 1.06674e-05 0.00115407 0.125629 0.000657722 0.126282 0.876034 101.833 0.244048 0.741816 4.16699 0.0559515 0.0393112 0.960689 0.0198222 0.00428408 0.0190851 0.00411841 0.00517785 0.00591495 0.207114 0.236598 57.9896 -87.8956 126.235 15.9706 145.017 0.000141441 0.267135 192.882 0.310595 0.0673745 0.00409563 0.000561749 0.00138306 0.986985 0.991731 -2.97602e-06 -85.6659 0.0930032 31190.2 301.661 0.983517 0.319147 0.733724 0.73372 9.99958 2.9818e-06 1.19271e-05 0.131062 0.981662 0.931437 -0.013293 4.90263e-06 0.502567 -1.89864e-20 7.00244e-24 -1.89794e-20 0.00139538 0.997818 8.5947e-05 0.152587 2.85192 0.00139538 0.997829 0.708152 0.00105064 0.00187999 0.00085947 0.455599 0.00187999 0.43821 0.000128585 1.02 0.887729 0.534667 0.28612 1.71691e-07 3.06261e-09 2386.54 3120.76 -0.0555942 0.482137 0.277543 0.253581 -0.593322 -0.169513 0.49633 -0.267787 -0.228553 1.712 1 0 297.532 0 2.09659 1.71 0.000299875 0.855323 0.657 0.392436 0.411482 2.09681 131.754 83.8631 18.7176 60.8386 0.00402767 0 -40 10
0.811 2.34971e-08 2.53896e-06 0.100574 0.100571 0.0120392 1.06805e-05 0.00115407 0.125717 0.000657724 0.12637 0.876099 101.833 0.244041 0.741912 4.16719 0.0559592 0.0393131 0.960687 0.0198219 0.00428427 0.0190848 0.00411857 0.00517808 0.00591518 0.207123 0.236607 57.9896 -87.8956 126.235 15.9706 145.017 0.000141438 0.267136 192.882 0.310595 0.0673745 0.00409563 0.000561749 0.00138306 0.986985 0.991731 -2.97603e-06 -85.6659 0.0930033 31190.2 301.666 0.983517 0.319147 0.73371 0.733705 9.99958 2.98181e-06 1.19271e-05 0.131064 0.981668 0.931439 -0.013293 4.90265e-06 0.502575 -1.89872e-20 7.0028e-24 -1.89802e-20 0.00139538 0.997818 8.59471e-05 0.152587 2.85192 0.00139538 0.997829 0.708253 0.00105066 0.00187999 0.000859471 0.455599 0.00187999 0.438218 0.000128588 1.02 0.88773 0.534667 0.286122 1.71691e-07 3.06263e-09 2386.53 3120.7 -0.0555908 0.482137 0.277543 0.253577 -0.593322 -0.169513 0.496339 -0.267785 -0.228564 1.713 1 0 297.535 0 2.09675 1.711 0.000299874 0.855297 0.657051 0.392265 0.411509 2.09697 131.763 83.8638 18.7176 60.839 0.00402764 0 -40 10
0.812 2.35261e-08 2.53896e-06 0.100644 0.100642 0.0120392 1.06937e-05 0.00115407 0.125805 0.000657727 0.126458 0.876163 101.833 0.244033 0.742008 4.1674 0.0559669 0.0393151 0.960685 0.0198217 0.00428446 0.0190846 0.00411873 0.00517832 0.00591541 0.207133 0.236617 57.9897 -87.8956 126.235 15.9706 145.017 0.000141435 0.267136 192.881 0.310594 0.0673744 0.00409563 0.00056175 0.00138306 0.986985 0.991731 -2.97604e-06 -85.6658 0.0930034 31190.1 301.672 0.983517 0.319147 0.733696 0.733691 9.99958 2.98181e-06 1.19271e-05 0.131065 0.981673 0.931442 -0.013293 4.90268e-06 0.502583 -1.89881e-20 7.00316e-24 -1.89811e-20 0.00139538 0.997818 8.59472e-05 0.152588 2.85192 0.00139538 0.997829 0.708355 0.00105068 0.00187999 0.000859472 0.455599 0.00187999 0.438227 0.000128591 1.02 0.887731 0.534666 0.286123 1.71692e-07 3.06266e-09 2386.51 3120.64 -0.0555874 0.482137 0.277542 0.253573 -0.593323 -0.169514 0.496349 -0.267783 -0.228575 1.714 1 0 297.539 0 2.09691 1.712 0.000299874 0.855272 0.657101 0.392094 0.411536 2.09713 131.771 83.8645 18.7176 60.8393 0.00402761 0 -40 10
0.813 2.3555e-08 2.53896e-06 0.100714 0.100712 0.0120392 1.07068e-05 0.00115407 0.125893 0.000657729 0.126546 0.876228 101.832 0.244025 0.742105 4.1676 0.0559746 0.039317 0.960683 0.0198214 0.00428465 0.0190844 0.00411889 0.00517855 0.00591565 0.207142 0.236626 57.9897 -87.8956 126.235 15.9705 145.017 0.000141433 0.267136 192.881 0.310594 0.0673744 0.00409564 0.000561751 0.00138306 0.986985 0.991731 -2.97606e-06 -85.6658 0.0930034 31190.1 301.677 0.983517 0.319147 0.733681 0.733677 9.99958 2.98182e-06 1.19272e-05 0.131067 0.981679 0.931444 -0.013293 4.90271e-06 0.502591 -1.8989e-20 7.00352e-24 -1.8982e-20 0.00139538 0.997818 8.59472e-05 0.152588 2.85192 0.00139538 0.997828 0.708456 0.0010507 0.00187999 0.000859472 0.455599 0.00187999 0.438235 0.000128595 1.02 0.887732 0.534666 0.286125 1.71692e-07 3.06268e-09 2386.49 3120.58 -0.0555841 0.482137 0.277542 0.253569 -0.593324 -0.169514 0.496358 -0.26778 -0.228586 1.715 1 0 297.543 0 2.09707 1.713 0.000299873 0.855247 0.657152 0.391923 0.411563 2.09729 131.78 83.8652 18.7177 60.8396 0.00402759 0 -40 10
0.814 2.35839e-08 2.53896e-06 0.100785 0.100782 0.0120392 1.072e-05 0.00115407 0.125981 0.000657731 0.126634 0.876293 101.832 0.244018 0.742201 4.16781 0.0559823 0.039319 0.960681 0.0198212 0.00428484 0.0190841 0.00411905 0.00517879 0.00591588 0.207151 0.236635 57.9898 -87.8956 126.236 15.9705 145.017 0.00014143 0.267136 192.881 0.310593 0.0673743 0.00409564 0.000561751 0.00138306 0.986985 0.991731 -2.97607e-06 -85.6658 0.0930035 31190.1 301.682 0.983517 0.319147 0.733667 0.733663 9.99958 2.98182e-06 1.19272e-05 0.131069 0.981685 0.931446 -0.013293 4.90274e-06 0.502599 -1.89898e-20 7.00388e-24 -1.89828e-20 0.00139538 0.997818 8.59473e-05 0.152588 2.85193 0.00139538 0.997828 0.708558 0.00105072 0.00187999 0.000859473 0.455598 0.00187999 0.438243 0.000128598 1.02 0.887733 0.534666 0.286126 1.71692e-07 3.0627e-09 2386.48 3120.52 -0.0555808 0.482137 0.277542 0.253565 -0.593324 -0.169514 0.496367 -0.267778 -0.228597 1.716 1 0 297.546 0 2.09723 1.714 0.000299873 0.855222 0.657202 0.391752 0.41159 2.09745 131.789 83.8659 18.7177 60.84 0.00402756 0 -40 10
0.815 2.36129e-08 2.53896e-06 0.100855 0.100853 0.0120392 1.07331e-05 0.00115407 0.126069 0.000657734 0.126722 0.876357 101.832 0.24401 0.742298 4.16802 0.0559899 0.0393209 0.960679 0.019821 0.00428504 0.0190839 0.00411921 0.00517902 0.00591612 0.207161 0.236645 57.9899 -87.8956 126.236 15.9705 145.017 0.000141427 0.267136 192.881 0.310593 0.0673743 0.00409564 0.000561752 0.00138307 0.986985 0.991731 -2.97609e-06 -85.6658 0.0930036 31190.1 301.687 0.983517 0.319147 0.733654 0.733649 9.99958 2.98183e-06 1.19272e-05 0.131071 0.981691 0.931448 -0.013293 4.90277e-06 0.502607 -1.89907e-20 7.00424e-24 -1.89837e-20 0.00139538 0.997818 8.59474e-05 0.152588 2.85193 0.00139538 0.997828 0.708659 0.00105074 0.00188 0.000859474 0.455598 0.00188 0.438251 0.000128601 1.02 0.887734 0.534665 0.286128 1.71692e-07 3.06272e-09 2386.46 3120.46 -0.0555775 0.482137 0.277542 0.253562 -0.593325 -0.169514 0.496376 -0.267776 -0.228608 1.717 1 0 297.55 0 2.09739 1.715 0.000299873 0.855198 0.657253 0.391582 0.411617 2.09762 131.797 83.8666 18.7178 60.8403 0.00402753 0 -40 10
0.816 2.36418e-08 2.53896e-06 0.100925 0.100923 0.0120392 1.07463e-05 0.00115407 0.126157 0.000657736 0.12681 0.876422 101.832 0.244002 0.742395 4.16822 0.0559976 0.0393229 0.960677 0.0198207 0.00428523 0.0190836 0.00411937 0.00517926 0.00591635 0.20717 0.236654 57.9899 -87.8956 126.236 15.9704 145.017 0.000141425 0.267137 192.881 0.310592 0.0673742 0.00409565 0.000561753 0.00138307 0.986985 0.991731 -2.9761e-06 -85.6658 0.0930037 31190 301.692 0.983516 0.319147 0.73364 0.733635 9.99958 2.98183e-06 1.19272e-05 0.131073 0.981696 0.93145 -0.0132929 4.9028e-06 0.502615 -1.89916e-20 7.0046e-24 -1.89845e-20 0.00139539 0.997818 8.59475e-05 0.152588 2.85193 0.00139539 0.997828 0.708761 0.00105076 0.00188 0.000859475 0.455598 0.00188 0.43826 0.000128604 1.02 0.887735 0.534665 0.286129 1.71693e-07 3.06274e-09 2386.44 3120.4 -0.0555743 0.482137 0.277541 0.253558 -0.593326 -0.169514 0.496384 -0.267774 -0.228619 1.718 1 0 297.554 0 2.09755 1.716 0.000299872 0.855173 0.657303 0.391413 0.411644 2.09778 131.806 83.8673 18.7178 60.8406 0.0040275 0 -40 10
0.817 2.36707e-08 2.53896e-06 0.100995 0.100993 0.0120392 1.07594e-05 0.00115407 0.126244 0.000657739 0.126897 0.876487 101.832 0.243995 0.742491 4.16843 0.0560053 0.0393248 0.960675 0.0198205 0.00428542 0.0190834 0.00411953 0.00517949 0.00591659 0.20718 0.236664 57.99 -87.8956 126.237 15.9704 145.017 0.000141422 0.267137 192.881 0.310592 0.0673742 0.00409565 0.000561753 0.00138307 0.986985 0.991731 -2.97612e-06 -85.6658 0.0930038 31190 301.698 0.983516 0.319147 0.733626 0.733622 9.99958 2.98183e-06 1.19272e-05 0.131075 0.981702 0.931452 -0.0132929 4.90283e-06 0.502623 -1.89924e-20 7.00496e-24 -1.89854e-20 0.00139539 0.997818 8.59476e-05 0.152588 2.85193 0.00139539 0.997828 0.708862 0.00105078 0.00188 0.000859476 0.455598 0.00188 0.438268 0.000128608 1.02 0.887736 0.534665 0.286131 1.71693e-07 3.06277e-09 2386.43 3120.34 -0.0555711 0.482137 0.277541 0.253554 -0.593326 -0.169514 0.496393 -0.267772 -0.22863 1.719 1 0 297.557 0 2.09771 1.717 0.000299872 0.855149 0.657354 0.391244 0.411671 2.09794 131.814 83.8679 18.7178 60.841 0.00402747 0 -40 10
0.818 2.36997e-08 2.53896e-06 0.101066 0.101063 0.0120392 1.07726e-05 0.00115407 0.126332 0.000657741 0.126985 0.876552 101.831 0.243987 0.742588 4.16864 0.0560131 0.0393268 0.960673 0.0198203 0.00428561 0.0190832 0.00411969 0.00517973 0.00591683 0.207189 0.236673 57.9901 -87.8956 126.237 15.9703 145.017 0.000141419 0.267137 192.88 0.310592 0.0673741 0.00409565 0.000561754 0.00138307 0.986985 0.991731 -2.97613e-06 -85.6658 0.0930039 31190 301.703 0.983516 0.319147 0.733612 0.733608 9.99958 2.98184e-06 1.19273e-05 0.131077 0.981708 0.931454 -0.0132929 4.90286e-06 0.502631 -1.89933e-20 7.00532e-24 -1.89863e-20 0.00139539 0.997817 8.59476e-05 0.152589 2.85193 0.00139539 0.997828 0.708963 0.0010508 0.00188 0.000859476 0.455598 0.00188 0.438276 0.000128611 1.02 0.887737 0.534664 0.286132 1.71693e-07 3.06279e-09 2386.41 3120.28 -0.0555679 0.482137 0.277541 0.25355 -0.593327 -0.169514 0.496402 -0.26777 -0.228641 1.72 1 0 297.561 0 2.09788 1.718 0.000299871 0.855124 0.657404 0.391075 0.411698 2.0981 131.823 83.8686 18.7179 60.8413 0.00402744 0 -40 10
0.819 2.37286e-08 2.53896e-06 0.101136 0.101133 0.0120391 1.07857e-05 0.00115407 0.12642 0.000657743 0.127073 0.876617 101.831 0.243979 0.742685 4.16885 0.0560208 0.0393288 0.960671 0.01982 0.00428581 0.0190829 0.00411986 0.00517997 0.00591706 0.207199 0.236683 57.9901 -87.8956 126.237 15.9703 145.017 0.000141417 0.267137 192.88 0.310591 0.067374 0.00409565 0.000561755 0.00138307 0.986985 0.991731 -2.97615e-06 -85.6658 0.093004 31190 301.708 0.983516 0.319147 0.733599 0.733594 9.99958 2.98184e-06 1.19273e-05 0.131079 0.981713 0.931456 -0.0132929 4.90289e-06 0.502639 -1.89942e-20 7.00569e-24 -1.89871e-20 0.00139539 0.997817 8.59477e-05 0.152589 2.85193 0.00139539 0.997828 0.709065 0.00105082 0.00188 0.000859477 0.455597 0.00188 0.438284 0.000128614 1.02 0.887738 0.534664 0.286134 1.71693e-07 3.06281e-09 2386.39 3120.22 -0.0555647 0.482138 0.27754 0.253547 -0.593328 -0.169514 0.49641 -0.267768 -0.228652 1.721 1 0 297.564 0 2.09804 1.719 0.000299871 0.8551 0.657455 0.390906 0.411725 2.09826 131.832 83.8693 18.7179 60.8416 0.00402742 0 -40 10
0.82 2.37575e-08 2.53896e-06 0.101206 0.101203 0.0120391 1.07989e-05 0.00115407 0.126507 0.000657746 0.12716 0.876682 101.831 0.243972 0.742782 4.16906 0.0560285 0.0393307 0.960669 0.0198198 0.004286 0.0190827 0.00412002 0.00518021 0.0059173 0.207208 0.236692 57.9902 -87.8956 126.237 15.9703 145.017 0.000141414 0.267137 192.88 0.310591 0.067374 0.00409566 0.000561755 0.00138308 0.986985 0.991731 -2.97616e-06 -85.6658 0.093004 31190 301.713 0.983516 0.319147 0.733585 0.733581 9.99958 2.98185e-06 1.19273e-05 0.131081 0.981719 0.931459 -0.0132929 4.90292e-06 0.502647 -1.8995e-20 7.00605e-24 -1.8988e-20 0.00139539 0.997817 8.59478e-05 0.152589 2.85193 0.00139539 0.997828 0.709166 0.00105083 0.00188 0.000859478 0.455597 0.00188 0.438293 0.000128617 1.02 0.887739 0.534664 0.286135 1.71694e-07 3.06283e-09 2386.38 3120.17 -0.0555616 0.482138 0.27754 0.253543 -0.593328 -0.169514 0.496419 -0.267766 -0.228662 1.722 1 0 297.568 0 2.0982 1.72 0.000299871 0.855076 0.657505 0.390738 0.411752 2.09842 131.84 83.87 18.718 60.8419 0.00402739 0 -40 10
0.821 2.37865e-08 2.53896e-06 0.101276 0.101273 0.0120391 1.0812e-05 0.00115407 0.126595 0.000657748 0.127248 0.876747 101.831 0.243964 0.742879 4.16927 0.0560362 0.0393327 0.960667 0.0198196 0.00428619 0.0190825 0.00412018 0.00518045 0.00591754 0.207218 0.236701 57.9902 -87.8956 126.237 15.9702 145.017 0.000141411 0.267137 192.88 0.31059 0.0673739 0.00409566 0.000561756 0.00138308 0.986985 0.991731 -2.97618e-06 -85.6658 0.0930041 31189.9 301.719 0.983516 0.319147 0.733572 0.733567 9.99958 2.98185e-06 1.19273e-05 0.131083 0.981725 0.931461 -0.0132929 4.90295e-06 0.502655 -1.89959e-20 7.00641e-24 -1.89889e-20 0.00139539 0.997817 8.59479e-05 0.152589 2.85193 0.00139539 0.997828 0.709267 0.00105085 0.00188001 0.000859479 0.455597 0.00188 0.438301 0.000128621 1.02 0.887741 0.534664 0.286137 1.71694e-07 3.06286e-09 2386.36 3120.11 -0.0555585 0.482138 0.27754 0.253539 -0.593329 -0.169514 0.496427 -0.267764 -0.228673 1.723 1 0 297.571 0 2.09836 1.721 0.00029987 0.855053 0.657555 0.39057 0.411779 2.09858 131.849 83.8706 18.718 60.8423 0.00402736 0 -40 10
0.822 2.38154e-08 2.53896e-06 0.101346 0.101343 0.0120391 1.08252e-05 0.00115407 0.126682 0.00065775 0.127335 0.876812 101.831 0.243956 0.742976 4.16948 0.0560439 0.0393347 0.960665 0.0198193 0.00428639 0.0190822 0.00412034 0.00518068 0.00591778 0.207227 0.236711 57.9903 -87.8956 126.238 15.9702 145.017 0.000141409 0.267138 192.88 0.31059 0.0673739 0.00409566 0.000561757 0.00138308 0.986985 0.991731 -2.97619e-06 -85.6658 0.0930042 31189.9 301.724 0.983516 0.319147 0.733558 0.733554 9.99958 2.98186e-06 1.19273e-05 0.131085 0.98173 0.931463 -0.0132929 4.90298e-06 0.502664 -1.89968e-20 7.00677e-24 -1.89897e-20 0.00139539 0.997817 8.59479e-05 0.152589 2.85193 0.00139539 0.997828 0.709368 0.00105087 0.00188001 0.000859479 0.455597 0.00188001 0.438309 0.000128624 1.02 0.887742 0.534663 0.286138 1.71694e-07 3.06288e-09 2386.34 3120.05 -0.0555554 0.482138 0.27754 0.253536 -0.59333 -0.169514 0.496436 -0.267762 -0.228683 1.724 1 0 297.575 0 2.09852 1.722 0.00029987 0.855029 0.657606 0.390403 0.411805 2.09874 131.858 83.8713 18.718 60.8426 0.00402733 0 -40 10
0.823 2.38443e-08 2.53896e-06 0.101415 0.101413 0.0120391 1.08383e-05 0.00115407 0.126769 0.000657753 0.127422 0.876877 101.83 0.243948 0.743073 4.16969 0.0560517 0.0393367 0.960663 0.0198191 0.00428658 0.019082 0.00412051 0.00518092 0.00591801 0.207237 0.236721 57.9904 -87.8956 126.238 15.9702 145.017 0.000141406 0.267138 192.88 0.310589 0.0673738 0.00409567 0.000561757 0.00138308 0.986985 0.991731 -2.97621e-06 -85.6657 0.0930043 31189.9 301.729 0.983516 0.319147 0.733545 0.733541 9.99958 2.98186e-06 1.19273e-05 0.131087 0.981736 0.931465 -0.0132929 4.903e-06 0.502672 -1.89976e-20 7.00713e-24 -1.89906e-20 0.00139539 0.997817 8.5948e-05 0.152589 2.85193 0.00139539 0.997828 0.709469 0.00105089 0.00188001 0.00085948 0.455596 0.00188001 0.438317 0.000128627 1.02 0.887743 0.534663 0.28614 1.71695e-07 3.0629e-09 2386.33 3119.99 -0.0555523 0.482138 0.277539 0.253532 -0.59333 -0.169514 0.496444 -0.26776 -0.228693 1.725 1 0 297.578 0 2.09868 1.723 0.000299869 0.855006 0.657656 0.390236 0.411832 2.0989 131.866 83.8719 18.7181 60.8429 0.00402731 0 -40 10
0.824 2.38733e-08 2.53896e-06 0.101485 0.101483 0.0120391 1.08515e-05 0.00115407 0.126856 0.000657755 0.12751 0.876942 101.83 0.243941 0.74317 4.1699 0.0560594 0.0393386 0.960661 0.0198188 0.00428678 0.0190817 0.00412067 0.00518116 0.00591825 0.207247 0.23673 57.9904 -87.8957 126.238 15.9701 145.017 0.000141404 0.267138 192.879 0.310589 0.0673738 0.00409567 0.000561758 0.00138308 0.986985 0.991731 -2.97622e-06 -85.6657 0.0930044 31189.9 301.734 0.983516 0.319147 0.733532 0.733527 9.99958 2.98187e-06 1.19274e-05 0.131089 0.981741 0.931467 -0.0132929 4.90303e-06 0.50268 -1.89985e-20 7.0075e-24 -1.89915e-20 0.00139539 0.997817 8.59481e-05 0.152589 2.85193 0.00139539 0.997828 0.70957 0.00105091 0.00188001 0.000859481 0.455596 0.00188001 0.438326 0.00012863 1.02 0.887744 0.534663 0.286141 1.71695e-07 3.06292e-09 2386.31 3119.94 -0.0555493 0.482138 0.277539 0.253529 -0.593331 -0.169514 0.496452 -0.267757 -0.228704 1.726 1 0 297.581 0 2.09884 1.724 0.000299869 0.854982 0.657706 0.39007 0.411859 2.09906 131.875 83.8726 18.7181 60.8432 0.00402728 0 -40 10
0.825 2.39022e-08 2.53896e-06 0.101555 0.101553 0.0120391 1.08646e-05 0.00115407 0.126944 0.000657757 0.127597 0.877007 101.83 0.243933 0.743268 4.17011 0.0560672 0.0393406 0.960659 0.0198186 0.00428697 0.0190815 0.00412083 0.0051814 0.00591849 0.207256 0.23674 57.9905 -87.8957 126.238 15.9701 145.017 0.000141401 0.267138 192.879 0.310589 0.0673737 0.00409567 0.000561759 0.00138309 0.986985 0.991731 -2.97623e-06 -85.6657 0.0930045 31189.8 301.74 0.983516 0.319147 0.733519 0.733514 9.99958 2.98187e-06 1.19274e-05 0.131091 0.981747 0.931469 -0.0132929 4.90306e-06 0.502688 -1.89994e-20 7.00786e-24 -1.89923e-20 0.0013954 0.997817 8.59482e-05 0.15259 2.85194 0.0013954 0.997828 0.709671 0.00105093 0.00188001 0.000859482 0.455596 0.00188001 0.438334 0.000128634 1.02 0.887745 0.534662 0.286143 1.71695e-07 3.06295e-09 2386.29 3119.88 -0.0555463 0.482138 0.277539 0.253525 -0.593332 -0.169514 0.49646 -0.267755 -0.228714 1.727 1 0 297.585 0 2.099 1.725 0.000299868 0.854959 0.657757 0.389903 0.411886 2.09922 131.883 83.8732 18.7182 60.8435 0.00402725 0 -40 10
0.826 2.39311e-08 2.53896e-06 0.101625 0.101622 0.012039 1.08778e-05 0.00115407 0.127031 0.00065776 0.127684 0.877072 101.83 0.243925 0.743365 4.17032 0.0560749 0.0393426 0.960657 0.0198184 0.00428717 0.0190813 0.004121 0.00518164 0.00591873 0.207266 0.236749 57.9906 -87.8957 126.239 15.97 145.017 0.000141399 0.267138 192.879 0.310588 0.0673737 0.00409568 0.000561759 0.00138309 0.986985 0.991731 -2.97625e-06 -85.6657 0.0930045 31189.8 301.745 0.983516 0.319147 0.733506 0.733501 9.99958 2.98188e-06 1.19274e-05 0.131093 0.981752 0.931471 -0.0132929 4.90309e-06 0.502696 -1.90002e-20 7.00822e-24 -1.89932e-20 0.0013954 0.997817 8.59483e-05 0.15259 2.85194 0.0013954 0.997828 0.709772 0.00105095 0.00188001 0.000859483 0.455596 0.00188001 0.438342 0.000128637 1.02 0.887746 0.534662 0.286144 1.71695e-07 3.06297e-09 2386.28 3119.82 -0.0555433 0.482138 0.277538 0.253522 -0.593332 -0.169514 0.496468 -0.267753 -0.228724 1.728 1 0 297.588 0 2.09916 1.726 0.000299868 0.854936 0.657807 0.389738 0.411913 2.09938 131.892 83.8739 18.7182 60.8438 0.00402723 0 -40 10
0.827 2.39601e-08 2.53896e-06 0.101694 0.101692 0.012039 1.08909e-05 0.00115407 0.127118 0.000657762 0.127771 0.877138 101.829 0.243917 0.743462 4.17053 0.0560827 0.0393446 0.960655 0.0198181 0.00428736 0.019081 0.00412116 0.00518188 0.00591897 0.207275 0.236759 57.9906 -87.8957 126.239 15.97 145.017 0.000141396 0.267139 192.879 0.310588 0.0673736 0.00409568 0.00056176 0.00138309 0.986985 0.991731 -2.97626e-06 -85.6657 0.0930046 31189.8 301.75 0.983516 0.319147 0.733493 0.733488 9.99958 2.98188e-06 1.19274e-05 0.131095 0.981758 0.931473 -0.0132929 4.90312e-06 0.502704 -1.90011e-20 7.00859e-24 -1.89941e-20 0.0013954 0.997817 8.59483e-05 0.15259 2.85194 0.0013954 0.997828 0.709873 0.00105097 0.00188001 0.000859483 0.455596 0.00188001 0.43835 0.00012864 1.02 0.887747 0.534662 0.286146 1.71696e-07 3.06299e-09 2386.26 3119.77 -0.0555404 0.482138 0.277538 0.253518 -0.593333 -0.169514 0.496476 -0.267751 -0.228734 1.729 1 0 297.591 0 2.09932 1.727 0.000299868 0.854913 0.657857 0.389572 0.41194 2.09954 131.901 83.8745 18.7182 60.8441 0.0040272 0 -40 10
0.828 2.3989e-08 2.53896e-06 0.101764 0.101761 0.012039 1.09041e-05 0.00115407 0.127205 0.000657764 0.127858 0.877203 101.829 0.24391 0.74356 4.17074 0.0560905 0.0393466 0.960653 0.0198179 0.00428756 0.0190808 0.00412132 0.00518212 0.00591921 0.207285 0.236768 57.9907 -87.8957 126.239 15.97 145.017 0.000141394 0.267139 192.879 0.310587 0.0673736 0.00409568 0.000561761 0.00138309 0.986985 0.991731 -2.97628e-06 -85.6657 0.0930047 31189.8 301.756 0.983516 0.319147 0.73348 0.733475 9.99958 2.98189e-06 1.19274e-05 0.131097 0.981763 0.931475 -0.0132929 4.90315e-06 0.502713 -1.9002e-20 7.00895e-24 -1.8995e-20 0.0013954 0.997817 8.59484e-05 0.15259 2.85194 0.0013954 0.997827 0.709974 0.00105099 0.00188002 0.000859484 0.455595 0.00188001 0.438359 0.000128643 1.02 0.887748 0.534661 0.286147 1.71696e-07 3.06301e-09 2386.24 3119.71 -0.0555374 0.482138 0.277538 0.253515 -0.593334 -0.169515 0.496484 -0.267749 -0.228744 1.73 1 0 297.595 0 2.09948 1.728 0.000299867 0.854891 0.657907 0.389407 0.411966 2.0997 131.909 83.8752 18.7183 60.8444 0.00402717 0 -40 10
0.829 2.40179e-08 2.53896e-06 0.101833 0.101831 0.012039 1.09172e-05 0.00115407 0.127292 0.000657767 0.127945 0.877268 101.829 0.243902 0.743658 4.17095 0.0560982 0.0393486 0.960651 0.0198176 0.00428776 0.0190805 0.00412149 0.00518237 0.00591945 0.207295 0.236778 57.9908 -87.8957 126.239 15.9699 145.017 0.000141391 0.267139 192.879 0.310587 0.0673735 0.00409568 0.000561761 0.0013831 0.986985 0.991731 -2.97629e-06 -85.6657 0.0930048 31189.8 301.761 0.983516 0.319147 0.733467 0.733463 9.99958 2.98189e-06 1.19275e-05 0.131099 0.981769 0.931477 -0.0132929 4.90318e-06 0.502721 -1.90028e-20 7.00931e-24 -1.89958e-20 0.0013954 0.997817 8.59485e-05 0.15259 2.85194 0.0013954 0.997827 0.710075 0.00105101 0.00188002 0.000859485 0.455595 0.00188002 0.438367 0.000128647 1.02 0.887749 0.534661 0.286149 1.71696e-07 3.06304e-09 2386.23 3119.66 -0.0555345 0.482138 0.277538 0.253511 -0.593334 -0.169515 0.496492 -0.267747 -0.228754 1.731 1 0 297.598 0 2.09964 1.729 0.000299867 0.854868 0.657958 0.389242 0.411993 2.09987 131.918 83.8758 18.7183 60.8447 0.00402715 0 -40 10
0.83 2.40469e-08 2.53896e-06 0.101903 0.1019 0.012039 1.09304e-05 0.00115407 0.127378 0.000657769 0.128032 0.877334 101.829 0.243894 0.743755 4.17117 0.056106 0.0393506 0.960649 0.0198174 0.00428795 0.0190803 0.00412165 0.00518261 0.00591969 0.207304 0.236788 57.9908 -87.8957 126.24 15.9699 145.017 0.000141389 0.267139 192.878 0.310587 0.0673735 0.00409569 0.000561762 0.0013831 0.986985 0.991731 -2.97631e-06 -85.6657 0.0930049 31189.7 301.766 0.983516 0.319147 0.733454 0.73345 9.99958 2.9819e-06 1.19275e-05 0.131101 0.981774 0.931479 -0.0132929 4.90321e-06 0.502729 -1.90037e-20 7.00968e-24 -1.89967e-20 0.0013954 0.997817 8.59486e-05 0.15259 2.85194 0.0013954 0.997827 0.710176 0.00105103 0.00188002 0.000859486 0.455595 0.00188002 0.438375 0.00012865 1.02 0.88775 0.534661 0.28615 1.71696e-07 3.06306e-09 2386.21 3119.6 -0.0555317 0.482138 0.277537 0.253508 -0.593335 -0.169515 0.496499 -0.267745 -0.228764 1.732 1 0 297.601 0 2.0998 1.73 0.000299866 0.854846 0.658008 0.389078 0.41202 2.10003 131.926 83.8764 18.7183 60.8451 0.00402712 0 -40 10
0.831 2.40758e-08 2.53897e-06 0.101972 0.10197 0.012039 1.09435e-05 0.00115408 0.127465 0.000657771 0.128118 0.877399 101.829 0.243886 0.743853 4.17138 0.0561138 0.0393527 0.960647 0.0198171 0.00428815 0.0190801 0.00412182 0.00518285 0.00591994 0.207314 0.236797 57.9909 -87.8957 126.24 15.9698 145.017 0.000141386 0.267139 192.878 0.310586 0.0673734 0.00409569 0.000561762 0.0013831 0.986985 0.991731 -2.97632e-06 -85.6657 0.093005 31189.7 301.772 0.983516 0.319147 0.733442 0.733437 9.99958 2.9819e-06 1.19275e-05 0.131103 0.98178 0.931481 -0.0132929 4.90324e-06 0.502738 -1.90046e-20 7.01004e-24 -1.89976e-20 0.0013954 0.997817 8.59487e-05 0.15259 2.85194 0.0013954 0.997827 0.710277 0.00105105 0.00188002 0.000859487 0.455595 0.00188002 0.438383 0.000128653 1.02 0.887751 0.534661 0.286152 1.71697e-07 3.06308e-09 2386.19 3119.55 -0.0555288 0.482138 0.277537 0.253504 -0.593335 -0.169515 0.496507 -0.267743 -0.228773 1.733 1 0 297.604 0 2.09996 1.731 0.000299866 0.854824 0.658058 0.388914 0.412047 2.10019 131.935 83.877 18.7184 60.8454 0.0040271 0 -40 10
0.832 2.41047e-08 2.53897e-06 0.102041 0.102039 0.012039 1.09567e-05 0.00115408 0.127552 0.000657774 0.128205 0.877464 101.828 0.243878 0.743951 4.17159 0.0561216 0.0393547 0.960645 0.0198169 0.00428835 0.0190798 0.00412198 0.00518309 0.00592018 0.207324 0.236807 57.9909 -87.8957 126.24 15.9698 145.017 0.000141384 0.26714 192.878 0.310586 0.0673734 0.00409569 0.000561763 0.0013831 0.986985 0.991731 -2.97634e-06 -85.6657 0.0930051 31189.7 301.777 0.983516 0.319147 0.733429 0.733425 9.99958 2.98191e-06 1.19275e-05 0.131105 0.981785 0.931483 -0.0132929 4.90327e-06 0.502746 -1.90055e-20 7.01041e-24 -1.89984e-20 0.0013954 0.997817 8.59487e-05 0.152591 2.85194 0.0013954 0.997827 0.710378 0.00105107 0.00188002 0.000859487 0.455594 0.00188002 0.438391 0.000128657 1.02 0.887752 0.53466 0.286153 1.71697e-07 3.0631e-09 2386.18 3119.49 -0.055526 0.482139 0.277537 0.253501 -0.593336 -0.169515 0.496515 -0.267741 -0.228783 1.734 1 0 297.607 0 2.10012 1.732 0.000299866 0.854802 0.658108 0.38875 0.412074 2.10035 131.944 83.8777 18.7184 60.8457 0.00402707 0 -40 10
0.833 2.41337e-08 2.53897e-06 0.102111 0.102108 0.012039 1.09698e-05 0.00115408 0.127638 0.000657776 0.128292 0.87753 101.828 0.243871 0.744049 4.17181 0.0561294 0.0393567 0.960643 0.0198167 0.00428854 0.0190796 0.00412215 0.00518334 0.00592042 0.207333 0.236817 57.991 -87.8957 126.24 15.9698 145.017 0.000141382 0.26714 192.878 0.310585 0.0673733 0.0040957 0.000561764 0.0013831 0.986985 0.991731 -2.97635e-06 -85.6657 0.0930051 31189.7 301.782 0.983516 0.319147 0.733417 0.733412 9.99958 2.98191e-06 1.19275e-05 0.131107 0.981791 0.931485 -0.0132929 4.9033e-06 0.502754 -1.90063e-20 7.01077e-24 -1.89993e-20 0.0013954 0.997817 8.59488e-05 0.152591 2.85194 0.0013954 0.997827 0.710479 0.00105109 0.00188002 0.000859488 0.455594 0.00188002 0.438399 0.00012866 1.02 0.887754 0.53466 0.286155 1.71697e-07 3.06313e-09 2386.16 3119.44 -0.0555232 0.482139 0.277536 0.253498 -0.593337 -0.169515 0.496522 -0.267739 -0.228793 1.735 1 0 297.611 0 2.10028 1.733 0.000299865 0.85478 0.658158 0.388587 0.4121 2.10051 131.952 83.8783 18.7184 60.8459 0.00402705 0 -40 10
0.834 2.41626e-08 2.53897e-06 0.10218 0.102178 0.0120389 1.0983e-05 0.00115408 0.127725 0.000657778 0.128378 0.877596 101.828 0.243863 0.744146 4.17202 0.0561372 0.0393587 0.960641 0.0198164 0.00428874 0.0190793 0.00412231 0.00518358 0.00592066 0.207343 0.236827 57.9911 -87.8957 126.241 15.9697 145.017 0.000141379 0.26714 192.878 0.310585 0.0673733 0.0040957 0.000561764 0.00138311 0.986985 0.991731 -2.97637e-06 -85.6656 0.0930052 31189.6 301.788 0.983516 0.319147 0.733404 0.7334 9.99958 2.98192e-06 1.19276e-05 0.131109 0.981796 0.931487 -0.0132929 4.90333e-06 0.502762 -1.90072e-20 7.01114e-24 -1.90002e-20 0.00139541 0.997817 8.59489e-05 0.152591 2.85194 0.00139541 0.997827 0.710579 0.00105111 0.00188002 0.000859489 0.455594 0.00188002 0.438408 0.000128663 1.02 0.887755 0.53466 0.286156 1.71697e-07 3.06315e-09 2386.14 3119.39 -0.0555204 0.482139 0.277536 0.253494 -0.593337 -0.169515 0.496529 -0.267737 -0.228802 1.736 1 0 297.614 0 2.10044 1.734 0.000299865 0.854758 0.658209 0.388424 0.412127 2.10067 131.961 83.8789 18.7185 60.8462 0.00402702 0 -40 10
0.835 2.41915e-08 2.53897e-06 0.102249 0.102247 0.0120389 1.09961e-05 0.00115408 0.127811 0.000657781 0.128465 0.877661 101.828 0.243855 0.744244 4.17224 0.056145 0.0393607 0.960639 0.0198162 0.00428894 0.0190791 0.00412248 0.00518382 0.00592091 0.207353 0.236836 57.9911 -87.8957 126.241 15.9697 145.017 0.000141377 0.26714 192.878 0.310584 0.0673732 0.0040957 0.000561765 0.00138311 0.986985 0.991731 -2.97638e-06 -85.6656 0.0930053 31189.6 301.793 0.983516 0.319147 0.733392 0.733387 9.99958 2.98192e-06 1.19276e-05 0.131111 0.981802 0.931489 -0.0132929 4.90336e-06 0.502771 -1.90081e-20 7.0115e-24 -1.90011e-20 0.00139541 0.997817 8.5949e-05 0.152591 2.85194 0.00139541 0.997827 0.71068 0.00105113 0.00188003 0.00085949 0.455594 0.00188002 0.438416 0.000128666 1.02 0.887756 0.534659 0.286158 1.71698e-07 3.06317e-09 2386.13 3119.33 -0.0555177 0.482139 0.277536 0.253491 -0.593338 -0.169515 0.496537 -0.267734 -0.228812 1.737 1 0 297.617 0 2.1006 1.735 0.000299864 0.854737 0.658259 0.388262 0.412154 2.10083 131.969 83.8795 18.7185 60.8465 0.004027 0 -40 10
0.836 2.42205e-08 2.53897e-06 0.102318 0.102316 0.0120389 1.10093e-05 0.00115408 0.127898 0.000657783 0.128551 0.877727 101.828 0.243847 0.744343 4.17245 0.0561528 0.0393628 0.960637 0.0198159 0.00428914 0.0190789 0.00412265 0.00518407 0.00592115 0.207363 0.236846 57.9912 -87.8957 126.241 15.9697 145.017 0.000141374 0.26714 192.877 0.310584 0.0673732 0.0040957 0.000561766 0.00138311 0.986985 0.991731 -2.9764e-06 -85.6656 0.0930054 31189.6 301.798 0.983516 0.319147 0.73338 0.733375 9.99958 2.98193e-06 1.19276e-05 0.131113 0.981807 0.931491 -0.0132929 4.90338e-06 0.502779 -1.9009e-20 7.01187e-24 -1.90019e-20 0.00139541 0.997817 8.59491e-05 0.152591 2.85195 0.00139541 0.997827 0.710781 0.00105115 0.00188003 0.000859491 0.455594 0.00188003 0.438424 0.000128669 1.02 0.887757 0.534659 0.286159 1.71698e-07 3.06319e-09 2386.11 3119.28 -0.0555149 0.482139 0.277536 0.253488 -0.593339 -0.169515 0.496544 -0.267732 -0.228821 1.738 1 0 297.62 0 2.10076 1.736 0.000299864 0.854715 0.658309 0.3881 0.412181 2.10099 131.978 83.8801 18.7186 60.8468 0.00402697 0 -40 10
0.837 2.42494e-08 2.53897e-06 0.102387 0.102385 0.0120389 1.10225e-05 0.00115408 0.127984 0.000657785 0.128637 0.877793 101.827 0.243839 0.744441 4.17267 0.0561606 0.0393648 0.960635 0.0198157 0.00428934 0.0190786 0.00412281 0.00518431 0.00592139 0.207373 0.236856 57.9913 -87.8957 126.241 15.9696 145.017 0.000141372 0.26714 192.877 0.310584 0.0673731 0.00409571 0.000561766 0.00138311 0.986985 0.991731 -2.97641e-06 -85.6656 0.0930055 31189.6 301.804 0.983516 0.319147 0.733367 0.733363 9.99958 2.98193e-06 1.19276e-05 0.131115 0.981812 0.931493 -0.0132929 4.90341e-06 0.502787 -1.90098e-20 7.01223e-24 -1.90028e-20 0.00139541 0.997817 8.59491e-05 0.152591 2.85195 0.00139541 0.997827 0.710881 0.00105116 0.00188003 0.000859491 0.455593 0.00188003 0.438432 0.000128673 1.02 0.887758 0.534659 0.286161 1.71698e-07 3.06322e-09 2386.09 3119.23 -0.0555122 0.482139 0.277535 0.253484 -0.593339 -0.169515 0.496551 -0.26773 -0.22883 1.739 1 0 297.623 0 2.10092 1.737 0.000299864 0.854694 0.658359 0.387938 0.412207 2.10115 131.986 83.8807 18.7186 60.8471 0.00402695 0 -40 10
0.838 2.42783e-08 2.53897e-06 0.102456 0.102454 0.0120389 1.10356e-05 0.00115408 0.12807 0.000657787 0.128724 0.877858 101.827 0.243832 0.744539 4.17289 0.0561685 0.0393668 0.960633 0.0198154 0.00428954 0.0190784 0.00412298 0.00518456 0.00592164 0.207382 0.236866 57.9913 -87.8957 126.241 15.9696 145.017 0.00014137 0.267141 192.877 0.310583 0.0673731 0.00409571 0.000561767 0.00138311 0.986985 0.991731 -2.97643e-06 -85.6656 0.0930056 31189.6 301.809 0.983516 0.319147 0.733355 0.733351 9.99958 2.98194e-06 1.19276e-05 0.131117 0.981818 0.931495 -0.0132929 4.90344e-06 0.502796 -1.90107e-20 7.0126e-24 -1.90037e-20 0.00139541 0.997817 8.59492e-05 0.152592 2.85195 0.00139541 0.997827 0.710982 0.00105118 0.00188003 0.000859492 0.455593 0.00188003 0.43844 0.000128676 1.02 0.887759 0.534658 0.286162 1.71698e-07 3.06324e-09 2386.08 3119.18 -0.0555096 0.482139 0.277535 0.253481 -0.59334 -0.169515 0.496558 -0.267728 -0.228839 1.74 1 0 297.626 0 2.10108 1.738 0.000299863 0.854673 0.658409 0.387777 0.412234 2.10131 131.995 83.8813 18.7186 60.8474 0.00402692 0 -40 10
0.839 2.43073e-08 2.53897e-06 0.102525 0.102523 0.0120389 1.10488e-05 0.00115408 0.128157 0.00065779 0.12881 0.877924 101.827 0.243824 0.744637 4.1731 0.0561763 0.0393689 0.960631 0.0198152 0.00428974 0.0190781 0.00412315 0.0051848 0.00592188 0.207392 0.236875 57.9914 -87.8957 126.242 15.9695 145.017 0.000141367 0.267141 192.877 0.310583 0.067373 0.00409571 0.000561768 0.00138312 0.986985 0.991731 -2.97644e-06 -85.6656 0.0930057 31189.5 301.815 0.983516 0.319147 0.733343 0.733339 9.99958 2.98194e-06 1.19277e-05 0.131119 0.981823 0.931496 -0.0132929 4.90347e-06 0.502804 -1.90116e-20 7.01296e-24 -1.90046e-20 0.00139541 0.997817 8.59493e-05 0.152592 2.85195 0.00139541 0.997827 0.711082 0.0010512 0.00188003 0.000859493 0.455593 0.00188003 0.438449 0.000128679 1.02 0.88776 0.534658 0.286164 1.71699e-07 3.06326e-09 2386.06 3119.12 -0.0555069 0.482139 0.277535 0.253478 -0.59334 -0.169515 0.496565 -0.267726 -0.228848 1.741 1 0 297.629 0 2.10124 1.739 0.000299863 0.854652 0.658459 0.387615 0.412261 2.10146 132.004 83.8819 18.7187 60.8477 0.0040269 0 -40 10
0.84 2.43362e-08 2.53897e-06 0.102594 0.102592 0.0120389 1.10619e-05 0.00115408 0.128243 0.000657792 0.128896 0.87799 101.827 0.243816 0.744736 4.17332 0.0561841 0.0393709 0.960629 0.019815 0.00428994 0.0190779 0.00412332 0.00518505 0.00592213 0.207402 0.236885 57.9915 -87.8957 126.242 15.9695 145.017 0.000141365 0.267141 192.877 0.310582 0.067373 0.00409572 0.000561768 0.00138312 0.986985 0.991731 -2.97645e-06 -85.6656 0.0930057 31189.5 301.82 0.983516 0.319147 0.733331 0.733327 9.99958 2.98195e-06 1.19277e-05 0.131121 0.981828 0.931498 -0.0132929 4.9035e-06 0.502813 -1.90125e-20 7.01333e-24 -1.90054e-20 0.00139541 0.997817 8.59494e-05 0.152592 2.85195 0.00139541 0.997827 0.711183 0.00105122 0.00188003 0.000859494 0.455593 0.00188003 0.438457 0.000128682 1.02 0.887761 0.534658 0.286165 1.71699e-07 3.06328e-09 2386.04 3119.07 -0.0555043 0.482139 0.277534 0.253475 -0.593341 -0.169515 0.496572 -0.267724 -0.228858 1.742 1 0 297.632 0 2.1014 1.74 0.000299862 0.854631 0.658509 0.387455 0.412287 2.10162 132.012 83.8825 18.7187 60.848 0.00402687 0 -40 10
0.841 2.43651e-08 2.53897e-06 0.102663 0.102661 0.0120388 1.10751e-05 0.00115408 0.128329 0.000657794 0.128982 0.878056 101.826 0.243808 0.744834 4.17354 0.056192 0.039373 0.960627 0.0198147 0.00429014 0.0190776 0.00412348 0.0051853 0.00592237 0.207412 0.236895 57.9915 -87.8957 126.242 15.9695 145.017 0.000141363 0.267141 192.877 0.310582 0.0673729 0.00409572 0.000561769 0.00138312 0.986984 0.991731 -2.97647e-06 -85.6656 0.0930058 31189.5 301.825 0.983516 0.319147 0.73332 0.733315 9.99958 2.98195e-06 1.19277e-05 0.131124 0.981833 0.9315 -0.0132929 4.90353e-06 0.502821 -1.90133e-20 7.0137e-24 -1.90063e-20 0.00139541 0.997817 8.59494e-05 0.152592 2.85195 0.00139541 0.997827 0.711283 0.00105124 0.00188003 0.000859494 0.455592 0.00188003 0.438465 0.000128686 1.02 0.887762 0.534658 0.286167 1.71699e-07 3.06331e-09 2386.03 3119.02 -0.0555017 0.482139 0.277534 0.253472 -0.593341 -0.169515 0.496579 -0.267722 -0.228866 1.743 1 0 297.635 0 2.10156 1.741 0.000299862 0.854611 0.658559 0.387294 0.412314 2.10178 132.021 83.8831 18.7187 60.8483 0.00402685 0 -40 10
0.842 2.4394e-08 2.53897e-06 0.102732 0.102729 0.0120388 1.10882e-05 0.00115408 0.128415 0.000657797 0.129068 0.878122 101.826 0.2438 0.744933 4.17375 0.0561998 0.039375 0.960625 0.0198145 0.00429034 0.0190774 0.00412365 0.00518554 0.00592262 0.207422 0.236905 57.9916 -87.8957 126.242 15.9694 145.017 0.000141361 0.267141 192.877 0.310582 0.0673729 0.00409572 0.00056177 0.00138312 0.986984 0.991731 -2.97648e-06 -85.6656 0.0930059 31189.5 301.831 0.983516 0.319147 0.733308 0.733303 9.99958 2.98196e-06 1.19277e-05 0.131126 0.981839 0.931502 -0.0132929 4.90356e-06 0.502829 -1.90142e-20 7.01406e-24 -1.90072e-20 0.00139541 0.997817 8.59495e-05 0.152592 2.85195 0.00139541 0.997827 0.711384 0.00105126 0.00188004 0.000859495 0.455592 0.00188003 0.438473 0.000128689 1.02 0.887763 0.534657 0.286168 1.717e-07 3.06333e-09 2386.01 3118.97 -0.0554991 0.482139 0.277534 0.253468 -0.593342 -0.169515 0.496586 -0.26772 -0.228875 1.744 1 0 297.638 0 2.10172 1.742 0.000299861 0.85459 0.658609 0.387135 0.412341 2.10194 132.029 83.8837 18.7188 60.8485 0.00402682 0 -40 10
0.843 2.4423e-08 2.53897e-06 0.1028 0.102798 0.0120388 1.11014e-05 0.00115408 0.128501 0.000657799 0.129154 0.878188 101.826 0.243792 0.745031 4.17397 0.0562077 0.0393771 0.960623 0.0198142 0.00429054 0.0190771 0.00412382 0.00518579 0.00592287 0.207432 0.236915 57.9916 -87.8957 126.243 15.9694 145.017 0.000141358 0.267142 192.876 0.310581 0.0673728 0.00409573 0.00056177 0.00138312 0.986984 0.991731 -2.9765e-06 -85.6656 0.093006 31189.5 301.836 0.983516 0.319147 0.733296 0.733292 9.99958 2.98196e-06 1.19277e-05 0.131128 0.981844 0.931504 -0.0132929 4.90359e-06 0.502838 -1.90151e-20 7.01443e-24 -1.90081e-20 0.00139542 0.997817 8.59496e-05 0.152592 2.85195 0.00139542 0.997827 0.711484 0.00105128 0.00188004 0.000859496 0.455592 0.00188004 0.438481 0.000128692 1.02 0.887764 0.534657 0.28617 1.717e-07 3.06335e-09 2385.99 3118.92 -0.0554966 0.482139 0.277534 0.253465 -0.593343 -0.169516 0.496593 -0.267718 -0.228884 1.745 1 0 297.641 0 2.10188 1.743 0.000299861 0.85457 0.658659 0.386975 0.412367 2.1021 132.038 83.8842 18.7188 60.8488 0.0040268 0 -40 10
0.844 2.44519e-08 2.53897e-06 0.102869 0.102867 0.0120388 1.11145e-05 0.00115408 0.128586 0.000657801 0.12924 0.878254 101.826 0.243784 0.74513 4.17419 0.0562155 0.0393792 0.960621 0.019814 0.00429074 0.0190769 0.00412399 0.00518604 0.00592311 0.207441 0.236925 57.9917 -87.8957 126.243 15.9694 145.017 0.000141356 0.267142 192.876 0.310581 0.0673728 0.00409573 0.000561771 0.00138313 0.986984 0.991731 -2.97651e-06 -85.6655 0.0930061 31189.4 301.842 0.983516 0.319147 0.733284 0.73328 9.99958 2.98197e-06 1.19278e-05 0.13113 0.981849 0.931506 -0.0132929 4.90362e-06 0.502846 -1.9016e-20 7.0148e-24 -1.9009e-20 0.00139542 0.997817 8.59497e-05 0.152592 2.85195 0.00139542 0.997826 0.711585 0.0010513 0.00188004 0.000859497 0.455592 0.00188004 0.438489 0.000128695 1.02 0.887765 0.534657 0.286171 1.717e-07 3.06337e-09 2385.98 3118.87 -0.0554941 0.482139 0.277533 0.253462 -0.593343 -0.169516 0.496599 -0.267716 -0.228893 1.746 1 0 297.644 0 2.10204 1.744 0.000299861 0.85455 0.658709 0.386816 0.412394 2.10226 132.046 83.8848 18.7188 60.8491 0.00402678 0 -40 10
0.845 2.44808e-08 2.53897e-06 0.102938 0.102935 0.0120388 1.11277e-05 0.00115408 0.128672 0.000657803 0.129325 0.87832 101.826 0.243777 0.745228 4.17441 0.0562234 0.0393812 0.960619 0.0198137 0.00429094 0.0190766 0.00412416 0.00518629 0.00592336 0.207451 0.236934 57.9918 -87.8957 126.243 15.9693 145.017 0.000141354 0.267142 192.876 0.31058 0.0673727 0.00409573 0.000561772 0.00138313 0.986984 0.991731 -2.97653e-06 -85.6655 0.0930062 31189.4 301.847 0.983516 0.319147 0.733273 0.733269 9.99958 2.98197e-06 1.19278e-05 0.131132 0.981854 0.931508 -0.0132929 4.90365e-06 0.502855 -1.90169e-20 7.01516e-24 -1.90098e-20 0.00139542 0.997817 8.59498e-05 0.152593 2.85195 0.00139542 0.997826 0.711685 0.00105132 0.00188004 0.000859498 0.455592 0.00188004 0.438497 0.000128699 1.02 0.887767 0.534656 0.286173 1.717e-07 3.0634e-09 2385.96 3118.82 -0.0554916 0.482139 0.277533 0.253459 -0.593344 -0.169516 0.496606 -0.267713 -0.228902 1.747 1 0 297.646 0 2.1022 1.745 0.00029986 0.85453 0.658759 0.386657 0.412421 2.10242 132.055 83.8854 18.7189 60.8494 0.00402675 0 -40 10
0.846 2.45098e-08 2.53897e-06 0.103006 0.103004 0.0120388 1.11408e-05 0.00115408 0.128758 0.000657806 0.129411 0.878386 101.825 0.243769 0.745327 4.17463 0.0562313 0.0393833 0.960617 0.0198135 0.00429115 0.0190764 0.00412433 0.00518653 0.00592361 0.207461 0.236944 57.9918 -87.8957 126.243 15.9693 145.017 0.000141352 0.267142 192.876 0.31058 0.0673727 0.00409573 0.000561772 0.00138313 0.986984 0.991731 -2.97654e-06 -85.6655 0.0930063 31189.4 301.853 0.983516 0.319147 0.733261 0.733257 9.99958 2.98198e-06 1.19278e-05 0.131134 0.98186 0.93151 -0.0132929 4.90368e-06 0.502863 -1.90177e-20 7.01553e-24 -1.90107e-20 0.00139542 0.997817 8.59498e-05 0.152593 2.85195 0.00139542 0.997826 0.711785 0.00105134 0.00188004 0.000859498 0.455591 0.00188004 0.438506 0.000128702 1.02 0.887768 0.534656 0.286174 1.71701e-07 3.06342e-09 2385.94 3118.77 -0.0554891 0.48214 0.277533 0.253456 -0.593344 -0.169516 0.496612 -0.267711 -0.22891 1.748 1 0 297.649 0 2.10236 1.746 0.00029986 0.85451 0.658809 0.386498 0.412447 2.10258 132.063 83.8859 18.7189 60.8496 0.00402673 0 -40 10
0.847 2.45387e-08 2.53897e-06 0.103075 0.103073 0.0120388 1.1154e-05 0.00115408 0.128844 0.000657808 0.129497 0.878452 101.825 0.243761 0.745426 4.17485 0.0562392 0.0393854 0.960615 0.0198132 0.00429135 0.0190761 0.0041245 0.00518678 0.00592386 0.207471 0.236954 57.9919 -87.8957 126.243 15.9692 145.017 0.000141349 0.267142 192.876 0.310579 0.0673726 0.00409574 0.000561773 0.00138313 0.986984 0.991731 -2.97656e-06 -85.6655 0.0930063 31189.4 301.858 0.983516 0.319147 0.73325 0.733246 9.99958 2.98198e-06 1.19278e-05 0.131136 0.981865 0.931511 -0.0132929 4.90371e-06 0.502872 -1.90186e-20 7.0159e-24 -1.90116e-20 0.00139542 0.997817 8.59499e-05 0.152593 2.85196 0.00139542 0.997826 0.711886 0.00105136 0.00188004 0.000859499 0.455591 0.00188004 0.438514 0.000128705 1.02 0.887769 0.534656 0.286176 1.71701e-07 3.06344e-09 2385.93 3118.72 -0.0554866 0.48214 0.277532 0.253453 -0.593345 -0.169516 0.496619 -0.267709 -0.228919 1.749 1 0 297.652 0 2.10252 1.747 0.000299859 0.85449 0.658859 0.38634 0.412474 2.10274 132.072 83.8865 18.7189 60.8499 0.00402671 0 -40 10
0.848 2.45676e-08 2.53897e-06 0.103143 0.103141 0.0120388 1.11671e-05 0.00115408 0.128929 0.00065781 0.129582 0.878518 101.825 0.243753 0.745525 4.17507 0.056247 0.0393874 0.960613 0.019813 0.00429155 0.0190759 0.00412467 0.00518703 0.00592411 0.207481 0.236964 57.992 -87.8957 126.244 15.9692 145.017 0.000141347 0.267143 192.876 0.310579 0.0673726 0.00409574 0.000561774 0.00138314 0.986984 0.991731 -2.97657e-06 -85.6655 0.0930064 31189.3 301.864 0.983516 0.319147 0.733239 0.733234 9.99958 2.98199e-06 1.19278e-05 0.131138 0.98187 0.931513 -0.0132929 4.90374e-06 0.50288 -1.90195e-20 7.01627e-24 -1.90125e-20 0.00139542 0.997817 8.595e-05 0.152593 2.85196 0.00139542 0.997826 0.711986 0.00105138 0.00188004 0.0008595 0.455591 0.00188004 0.438522 0.000128708 1.02 0.88777 0.534655 0.286177 1.71701e-07 3.06346e-09 2385.91 3118.67 -0.0554842 0.48214 0.277532 0.25345 -0.593345 -0.169516 0.496625 -0.267707 -0.228927 1.75 1 0 297.655 0 2.10268 1.748 0.000299859 0.85447 0.658909 0.386182 0.412501 2.1029 132.08 83.8871 18.719 60.8502 0.00402668 0 -40 10
0.849 2.45966e-08 2.53897e-06 0.103212 0.103209 0.0120387 1.11803e-05 0.00115408 0.129015 0.000657812 0.129668 0.878584 101.825 0.243745 0.745624 4.17529 0.0562549 0.0393895 0.96061 0.0198127 0.00429175 0.0190756 0.00412484 0.00518728 0.00592435 0.207491 0.236974 57.992 -87.8957 126.244 15.9692 145.017 0.000141345 0.267143 192.875 0.310579 0.0673725 0.00409574 0.000561774 0.00138314 0.986984 0.991731 -2.97659e-06 -85.6655 0.0930065 31189.3 301.869 0.983516 0.319147 0.733228 0.733223 9.99958 2.98199e-06 1.19279e-05 0.13114 0.981875 0.931515 -0.0132929 4.90376e-06 0.502889 -1.90204e-20 7.01663e-24 -1.90134e-20 0.00139542 0.997817 8.59501e-05 0.152593 2.85196 0.00139542 0.997826 0.712086 0.0010514 0.00188005 0.000859501 0.455591 0.00188004 0.43853 0.000128712 1.02 0.887771 0.534655 0.286179 1.71701e-07 3.06349e-09 2385.89 3118.62 -0.0554818 0.48214 0.277532 0.253447 -0.593346 -0.169516 0.496631 -0.267705 -0.228936 1.751 1 0 297.658 0 2.10284 1.749 0.000299858 0.854451 0.658959 0.386025 0.412527 2.10306 132.089 83.8876 18.719 60.8505 0.00402666 0 -40 10
0.85 2.46255e-08 2.53897e-06 0.10328 0.103278 0.0120387 1.11934e-05 0.00115408 0.1291 0.000657814 0.129753 0.878651 101.824 0.243737 0.745723 4.17551 0.0562628 0.0393916 0.960608 0.0198125 0.00429196 0.0190754 0.00412501 0.00518753 0.0059246 0.207501 0.236984 57.9921 -87.8958 126.244 15.9691 145.017 0.000141343 0.267143 192.875 0.310578 0.0673725 0.00409575 0.000561775 0.00138314 0.986984 0.991731 -2.9766e-06 -85.6655 0.0930066 31189.3 301.875 0.983516 0.319147 0.733216 0.733212 9.99958 2.98199e-06 1.19279e-05 0.131142 0.98188 0.931517 -0.0132929 4.90379e-06 0.502897 -1.90213e-20 7.017e-24 -1.90142e-20 0.00139542 0.997817 8.59502e-05 0.152593 2.85196 0.00139542 0.997826 0.712186 0.00105142 0.00188005 0.000859502 0.45559 0.00188005 0.438538 0.000128715 1.02 0.887772 0.534655 0.28618 1.71702e-07 3.06351e-09 2385.88 3118.58 -0.0554794 0.48214 0.277532 0.253444 -0.593346 -0.169516 0.496638 -0.267703 -0.228944 1.752 1 0 297.66 0 2.103 1.75 0.000299858 0.854432 0.659008 0.385868 0.412554 2.10322 132.097 83.8882 18.719 60.8507 0.00402664 0 -40 10
0.851 2.46544e-08 2.53898e-06 0.103348 0.103346 0.0120387 1.12066e-05 0.00115408 0.129185 0.000657817 0.129839 0.878717 101.824 0.243729 0.745822 4.17573 0.0562707 0.0393937 0.960606 0.0198122 0.00429216 0.0190751 0.00412518 0.00518778 0.00592485 0.207511 0.236994 57.9922 -87.8958 126.244 15.9691 145.017 0.000141341 0.267143 192.875 0.310578 0.0673724 0.00409575 0.000561776 0.00138314 0.986984 0.991731 -2.97662e-06 -85.6655 0.0930067 31189.3 301.88 0.983516 0.319147 0.733205 0.733201 9.99958 2.982e-06 1.19279e-05 0.131144 0.981885 0.931519 -0.0132929 4.90382e-06 0.502906 -1.90221e-20 7.01737e-24 -1.90151e-20 0.00139543 0.997817 8.59502e-05 0.152593 2.85196 0.00139542 0.997826 0.712286 0.00105144 0.00188005 0.000859502 0.45559 0.00188005 0.438546 0.000128718 1.02 0.887773 0.534654 0.286182 1.71702e-07 3.06353e-09 2385.86 3118.53 -0.0554771 0.48214 0.277531 0.253441 -0.593347 -0.169516 0.496644 -0.267701 -0.228952 1.753 1 0 297.663 0 2.10316 1.751 0.000299858 0.854412 0.659058 0.385711 0.41258 2.10338 132.106 83.8887 18.7191 60.851 0.00402662 0 -40 10
0.852 2.46834e-08 2.53898e-06 0.103417 0.103414 0.0120387 1.12197e-05 0.00115408 0.129271 0.000657819 0.129924 0.878783 101.824 0.243721 0.745921 4.17595 0.0562786 0.0393958 0.960604 0.019812 0.00429236 0.0190749 0.00412535 0.00518803 0.0059251 0.207521 0.237004 57.9922 -87.8958 126.244 15.9691 145.017 0.000141339 0.267143 192.875 0.310577 0.0673723 0.00409575 0.000561776 0.00138314 0.986984 0.991731 -2.97663e-06 -85.6655 0.0930068 31189.3 301.886 0.983516 0.319147 0.733194 0.73319 9.99958 2.982e-06 1.19279e-05 0.131146 0.98189 0.93152 -0.0132929 4.90385e-06 0.502915 -1.9023e-20 7.01774e-24 -1.9016e-20 0.00139543 0.997817 8.59503e-05 0.152594 2.85196 0.00139543 0.997826 0.712387 0.00105145 0.00188005 0.000859503 0.45559 0.00188005 0.438554 0.000128721 1.02 0.887774 0.534654 0.286183 1.71702e-07 3.06355e-09 2385.84 3118.48 -0.0554747 0.48214 0.277531 0.253438 -0.593348 -0.169516 0.49665 -0.267699 -0.22896 1.754 1 0 297.666 0 2.10332 1.752 0.000299857 0.854393 0.659108 0.385554 0.412607 2.10354 132.115 83.8893 18.7191 60.8512 0.00402659 0 -40 10
0.853 2.47123e-08 2.53898e-06 0.103485 0.103483 0.0120387 1.12329e-05 0.00115408 0.129356 0.000657821 0.130009 0.87885 101.824 0.243713 0.746021 4.17618 0.0562865 0.0393979 0.960602 0.0198117 0.00429257 0.0190746 0.00412552 0.00518828 0.00592536 0.207531 0.237014 57.9923 -87.8958 126.245 15.969 145.018 0.000141337 0.267143 192.875 0.310577 0.0673723 0.00409576 0.000561777 0.00138315 0.986984 0.991731 -2.97665e-06 -85.6655 0.0930069 31189.2 301.891 0.983516 0.319147 0.733183 0.733179 9.99958 2.98201e-06 1.19279e-05 0.131148 0.981896 0.931522 -0.0132929 4.90388e-06 0.502923 -1.90239e-20 7.01811e-24 -1.90169e-20 0.00139543 0.997817 8.59504e-05 0.152594 2.85196 0.00139543 0.997826 0.712487 0.00105147 0.00188005 0.000859504 0.45559 0.00188005 0.438562 0.000128725 1.02 0.887775 0.534654 0.286185 1.71702e-07 3.06358e-09 2385.83 3118.43 -0.0554724 0.48214 0.277531 0.253435 -0.593348 -0.169516 0.496656 -0.267697 -0.228968 1.755 1 0 297.668 0 2.10348 1.753 0.000299857 0.854375 0.659158 0.385398 0.412633 2.1037 132.123 83.8898 18.7191 60.8515 0.00402657 0 -40 10
0.854 2.47412e-08 2.53898e-06 0.103553 0.103551 0.0120387 1.1246e-05 0.00115408 0.129441 0.000657823 0.130094 0.878916 101.824 0.243706 0.74612 4.1764 0.0562945 0.0394 0.9606 0.0198115 0.00429277 0.0190744 0.00412569 0.00518853 0.00592561 0.207541 0.237024 57.9923 -87.8958 126.245 15.969 145.018 0.000141334 0.267144 192.875 0.310576 0.0673722 0.00409576 0.000561778 0.00138315 0.986984 0.991731 -2.97666e-06 -85.6655 0.0930069 31189.2 301.897 0.983516 0.319147 0.733172 0.733168 9.99958 2.98201e-06 1.19279e-05 0.13115 0.981901 0.931524 -0.0132929 4.90391e-06 0.502932 -1.90248e-20 7.01848e-24 -1.90178e-20 0.00139543 0.997817 8.59505e-05 0.152594 2.85196 0.00139543 0.997826 0.712587 0.00105149 0.00188005 0.000859505 0.45559 0.00188005 0.438571 0.000128728 1.02 0.887776 0.534654 0.286186 1.71703e-07 3.0636e-09 2385.81 3118.39 -0.0554702 0.48214 0.27753 0.253432 -0.593349 -0.169516 0.496662 -0.267695 -0.228976 1.756 1 0 297.671 0 2.10363 1.754 0.000299856 0.854356 0.659208 0.385242 0.41266 2.10385 132.132 83.8904 18.7191 60.8518 0.00402655 0 -40 10
0.855 2.47701e-08 2.53898e-06 0.103621 0.103619 0.0120387 1.12592e-05 0.00115408 0.129526 0.000657825 0.130179 0.878982 101.823 0.243698 0.746219 4.17662 0.0563024 0.0394021 0.960598 0.0198112 0.00429298 0.0190741 0.00412586 0.00518879 0.00592586 0.207551 0.237034 57.9924 -87.8958 126.245 15.9689 145.018 0.000141332 0.267144 192.874 0.310576 0.0673722 0.00409576 0.000561778 0.00138315 0.986984 0.991731 -2.97668e-06 -85.6654 0.093007 31189.2 301.902 0.983516 0.319147 0.733162 0.733157 9.99958 2.98202e-06 1.1928e-05 0.131153 0.981906 0.931526 -0.0132929 4.90394e-06 0.50294 -1.90257e-20 7.01885e-24 -1.90187e-20 0.00139543 0.997817 8.59506e-05 0.152594 2.85196 0.00139543 0.997826 0.712687 0.00105151 0.00188005 0.000859506 0.455589 0.00188005 0.438579 0.000128731 1.02 0.887777 0.534653 0.286188 1.71703e-07 3.06362e-09 2385.79 3118.34 -0.0554679 0.48214 0.27753 0.253429 -0.593349 -0.169516 0.496668 -0.267693 -0.228984 1.757 1 0 297.674 0 2.10379 1.755 0.000299856 0.854337 0.659257 0.385087 0.412686 2.10401 132.14 83.8909 18.7192 60.852 0.00402653 0 -40 10
0.856 2.47991e-08 2.53898e-06 0.103689 0.103687 0.0120386 1.12723e-05 0.00115408 0.129611 0.000657828 0.130264 0.879049 101.823 0.24369 0.746319 4.17684 0.0563103 0.0394042 0.960596 0.019811 0.00429318 0.0190739 0.00412603 0.00518904 0.00592611 0.207562 0.237044 57.9925 -87.8958 126.245 15.9689 145.018 0.00014133 0.267144 192.874 0.310576 0.0673721 0.00409576 0.000561779 0.00138315 0.986984 0.991731 -2.97669e-06 -85.6654 0.0930071 31189.2 301.908 0.983516 0.319147 0.733151 0.733147 9.99958 2.98202e-06 1.1928e-05 0.131155 0.981911 0.931528 -0.0132929 4.90397e-06 0.502949 -1.90266e-20 7.01922e-24 -1.90195e-20 0.00139543 0.997817 8.59506e-05 0.152594 2.85196 0.00139543 0.997826 0.712787 0.00105153 0.00188006 0.000859506 0.455589 0.00188005 0.438587 0.000128734 1.02 0.887778 0.534653 0.286189 1.71703e-07 3.06364e-09 2385.77 3118.29 -0.0554657 0.48214 0.27753 0.253426 -0.59335 -0.169516 0.496673 -0.26769 -0.228992 1.758 1 0 297.676 0 2.10395 1.756 0.000299855 0.854319 0.659307 0.384932 0.412713 2.10417 132.149 83.8914 18.7192 60.8523 0.00402651 0 -40 10
0.857 2.4828e-08 2.53898e-06 0.103757 0.103755 0.0120386 1.12855e-05 0.00115408 0.129696 0.00065783 0.130349 0.879116 101.823 0.243682 0.746418 4.17707 0.0563182 0.0394063 0.960594 0.0198107 0.00429339 0.0190736 0.00412621 0.00518929 0.00592636 0.207572 0.237054 57.9925 -87.8958 126.245 15.9689 145.018 0.000141328 0.267144 192.874 0.310575 0.0673721 0.00409577 0.00056178 0.00138315 0.986984 0.991731 -2.9767e-06 -85.6654 0.0930072 31189.1 301.914 0.983516 0.319147 0.73314 0.733136 9.99958 2.98203e-06 1.1928e-05 0.131157 0.981916 0.931529 -0.0132929 4.904e-06 0.502958 -1.90275e-20 7.01959e-24 -1.90204e-20 0.00139543 0.997817 8.59507e-05 0.152594 2.85196 0.00139543 0.997826 0.712886 0.00105155 0.00188006 0.000859507 0.455589 0.00188006 0.438595 0.000128737 1.02 0.88778 0.534653 0.286191 1.71703e-07 3.06367e-09 2385.76 3118.25 -0.0554635 0.48214 0.27753 0.253423 -0.59335 -0.169516 0.496679 -0.267688 -0.229 1.759 1 0 297.679 0 2.10411 1.757 0.000299855 0.854301 0.659357 0.384777 0.41274 2.10433 132.157 83.8919 18.7192 60.8525 0.00402648 0 -40 10
0.858 2.48569e-08 2.53898e-06 0.103825 0.103823 0.0120386 1.12986e-05 0.00115408 0.129781 0.000657832 0.130434 0.879182 101.823 0.243674 0.746518 4.17729 0.0563262 0.0394084 0.960592 0.0198105 0.00429359 0.0190734 0.00412638 0.00518954 0.00592661 0.207582 0.237065 57.9926 -87.8958 126.246 15.9688 145.018 0.000141326 0.267144 192.874 0.310575 0.067372 0.00409577 0.00056178 0.00138316 0.986984 0.991731 -2.97672e-06 -85.6654 0.0930073 31189.1 301.919 0.983516 0.319147 0.73313 0.733125 9.99958 2.98203e-06 1.1928e-05 0.131159 0.981921 0.931531 -0.0132929 4.90403e-06 0.502966 -1.90283e-20 7.01996e-24 -1.90213e-20 0.00139543 0.997817 8.59508e-05 0.152595 2.85197 0.00139543 0.997826 0.712986 0.00105157 0.00188006 0.000859508 0.455589 0.00188006 0.438603 0.000128741 1.02 0.887781 0.534652 0.286192 1.71704e-07 3.06369e-09 2385.74 3118.2 -0.0554613 0.48214 0.277529 0.25342 -0.593351 -0.169516 0.496685 -0.267686 -0.229008 1.76 1 0 297.681 0 2.10427 1.758 0.000299855 0.854282 0.659407 0.384623 0.412766 2.10449 132.166 83.8925 18.7193 60.8528 0.00402646 0 -40 10
0.859 2.48859e-08 2.53898e-06 0.103893 0.10389 0.0120386 1.13118e-05 0.00115408 0.129866 0.000657834 0.130519 0.879249 101.822 0.243666 0.746618 4.17752 0.0563341 0.0394105 0.960589 0.0198102 0.0042938 0.0190731 0.00412655 0.0051898 0.00592687 0.207592 0.237075 57.9927 -87.8958 126.246 15.9688 145.018 0.000141324 0.267145 192.874 0.310574 0.067372 0.00409577 0.000561781 0.00138316 0.986984 0.991731 -2.97673e-06 -85.6654 0.0930074 31189.1 301.925 0.983516 0.319147 0.733119 0.733115 9.99958 2.98204e-06 1.1928e-05 0.131161 0.981926 0.931533 -0.0132929 4.90406e-06 0.502975 -1.90292e-20 7.02033e-24 -1.90222e-20 0.00139543 0.997817 8.59509e-05 0.152595 2.85197 0.00139543 0.997826 0.713086 0.00105159 0.00188006 0.000859509 0.455588 0.00188006 0.438611 0.000128744 1.02 0.887782 0.534652 0.286194 1.71704e-07 3.06371e-09 2385.72 3118.16 -0.0554591 0.48214 0.277529 0.253418 -0.593351 -0.169517 0.49669 -0.267684 -0.229015 1.761 1 0 297.684 0 2.10443 1.759 0.000299854 0.854264 0.659456 0.384469 0.412793 2.10465 132.174 83.893 18.7193 60.853 0.00402644 0 -40 10
0.86 2.49148e-08 2.53898e-06 0.10396 0.103958 0.0120386 1.13249e-05 0.00115408 0.129951 0.000657836 0.130604 0.879315 101.822 0.243658 0.746717 4.17774 0.0563421 0.0394127 0.960587 0.0198099 0.00429401 0.0190729 0.00412672 0.00519005 0.00592712 0.207602 0.237085 57.9927 -87.8958 126.246 15.9687 145.018 0.000141322 0.267145 192.874 0.310574 0.0673719 0.00409578 0.000561781 0.00138316 0.986984 0.991731 -2.97675e-06 -85.6654 0.0930075 31189.1 301.93 0.983516 0.319147 0.733109 0.733104 9.99958 2.98204e-06 1.19281e-05 0.131163 0.981931 0.931534 -0.0132929 4.90409e-06 0.502984 -1.90301e-20 7.0207e-24 -1.90231e-20 0.00139544 0.997817 8.59509e-05 0.152595 2.85197 0.00139544 0.997826 0.713186 0.00105161 0.00188006 0.000859509 0.455588 0.00188006 0.438619 0.000128747 1.02 0.887783 0.534652 0.286195 1.71704e-07 3.06373e-09 2385.71 3118.11 -0.055457 0.482141 0.277529 0.253415 -0.593352 -0.169517 0.496696 -0.267682 -0.229023 1.762 1 0 297.686 0 2.10459 1.76 0.000299854 0.854247 0.659506 0.384315 0.412819 2.10481 132.183 83.8935 18.7193 60.8533 0.00402642 0 -40 10
0.861 2.49437e-08 2.53898e-06 0.104028 0.104026 0.0120386 1.13381e-05 0.00115408 0.130035 0.000657839 0.130688 0.879382 101.822 0.24365 0.746817 4.17797 0.05635 0.0394148 0.960585 0.0198097 0.00429421 0.0190726 0.0041269 0.00519031 0.00592738 0.207612 0.237095 57.9928 -87.8958 126.246 15.9687 145.018 0.00014132 0.267145 192.873 0.310574 0.0673719 0.00409578 0.000561782 0.00138316 0.986984 0.991731 -2.97676e-06 -85.6654 0.0930075 31189.1 301.936 0.983516 0.319147 0.733098 0.733094 9.99958 2.98205e-06 1.19281e-05 0.131165 0.981936 0.931536 -0.0132929 4.90412e-06 0.502992 -1.9031e-20 7.02107e-24 -1.9024e-20 0.00139544 0.997817 8.5951e-05 0.152595 2.85197 0.00139544 0.997825 0.713286 0.00105163 0.00188006 0.00085951 0.455588 0.00188006 0.438627 0.00012875 1.02 0.887784 0.534651 0.286197 1.71705e-07 3.06376e-09 2385.69 3118.07 -0.0554549 0.482141 0.277528 0.253412 -0.593352 -0.169517 0.496701 -0.26768 -0.22903 1.763 1 0 297.689 0 2.10475 1.761 0.000299853 0.854229 0.659556 0.384162 0.412845 2.10497 132.191 83.894 18.7194 60.8535 0.0040264 0 -40 10
0.862 2.49727e-08 2.53898e-06 0.104096 0.104094 0.0120386 1.13512e-05 0.00115408 0.13012 0.000657841 0.130773 0.879449 101.822 0.243642 0.746917 4.17819 0.056358 0.0394169 0.960583 0.0198094 0.00429442 0.0190724 0.00412707 0.00519056 0.00592763 0.207622 0.237105 57.9929 -87.8958 126.246 15.9687 145.018 0.000141318 0.267145 192.873 0.310573 0.0673718 0.00409578 0.000561783 0.00138317 0.986984 0.991731 -2.97678e-06 -85.6654 0.0930076 31189 301.942 0.983516 0.319147 0.733088 0.733084 9.99958 2.98205e-06 1.19281e-05 0.131167 0.981941 0.931538 -0.0132929 4.90415e-06 0.503001 -1.90319e-20 7.02144e-24 -1.90249e-20 0.00139544 0.997817 8.59511e-05 0.152595 2.85197 0.00139544 0.997825 0.713386 0.00105165 0.00188006 0.000859511 0.455588 0.00188006 0.438635 0.000128754 1.02 0.887785 0.534651 0.286198 1.71705e-07 3.06378e-09 2385.67 3118.02 -0.0554528 0.482141 0.277528 0.253409 -0.593353 -0.169517 0.496707 -0.267678 -0.229038 1.764 1 0 297.691 0 2.1049 1.762 0.000299853 0.854211 0.659605 0.384009 0.412872 2.10512 132.2 83.8945 18.7194 60.8538 0.00402638 0 -40 10
0.863 2.50016e-08 2.53898e-06 0.104163 0.104161 0.0120386 1.13644e-05 0.00115408 0.130204 0.000657843 0.130858 0.879516 101.822 0.243634 0.747017 4.17842 0.056366 0.0394191 0.960581 0.0198092 0.00429463 0.0190721 0.00412725 0.00519082 0.00592788 0.207633 0.237115 57.9929 -87.8958 126.246 15.9686 145.018 0.000141316 0.267145 192.873 0.310573 0.0673718 0.00409579 0.000561783 0.00138317 0.986984 0.991731 -2.97679e-06 -85.6654 0.0930077 31189 301.947 0.983516 0.319147 0.733078 0.733074 9.99958 2.98206e-06 1.19281e-05 0.131169 0.981945 0.93154 -0.0132929 4.90417e-06 0.50301 -1.90328e-20 7.02181e-24 -1.90258e-20 0.00139544 0.997817 8.59512e-05 0.152595 2.85197 0.00139544 0.997825 0.713485 0.00105167 0.00188007 0.000859512 0.455588 0.00188007 0.438643 0.000128757 1.02 0.887786 0.534651 0.2862 1.71705e-07 3.0638e-09 2385.66 3117.98 -0.0554507 0.482141 0.277528 0.253406 -0.593353 -0.169517 0.496712 -0.267676 -0.229045 1.765 1 0 297.694 0 2.10506 1.763 0.000299852 0.854194 0.659655 0.383856 0.412898 2.10528 132.208 83.895 18.7194 60.854 0.00402636 0 -40 10
0.864 2.50305e-08 2.53898e-06 0.104231 0.104229 0.0120385 1.13775e-05 0.00115408 0.130289 0.000657845 0.130942 0.879583 101.821 0.243626 0.747117 4.17865 0.0563739 0.0394212 0.960579 0.0198089 0.00429484 0.0190719 0.00412742 0.00519107 0.00592814 0.207643 0.237126 57.993 -87.8958 126.247 15.9686 145.018 0.000141314 0.267146 192.873 0.310572 0.0673717 0.00409579 0.000561784 0.00138317 0.986984 0.991731 -2.97681e-06 -85.6654 0.0930078 31189 301.953 0.983516 0.319147 0.733068 0.733063 9.99958 2.98206e-06 1.19281e-05 0.131172 0.98195 0.931541 -0.0132929 4.9042e-06 0.503018 -1.90337e-20 7.02218e-24 -1.90267e-20 0.00139544 0.997817 8.59513e-05 0.152595 2.85197 0.00139544 0.997825 0.713585 0.00105169 0.00188007 0.000859513 0.455587 0.00188007 0.438651 0.00012876 1.02 0.887787 0.534651 0.286201 1.71705e-07 3.06382e-09 2385.64 3117.93 -0.0554487 0.482141 0.277528 0.253404 -0.593354 -0.169517 0.496717 -0.267674 -0.229053 1.766 1 0 297.696 0 2.10522 1.764 0.000299852 0.854177 0.659705 0.383704 0.412925 2.10544 132.217 83.8955 18.7194 60.8543 0.00402634 0 -40 10
0.865 2.50594e-08 2.53898e-06 0.104299 0.104296 0.0120385 1.13907e-05 0.00115408 0.130373 0.000657847 0.131026 0.87965 101.821 0.243618 0.747217 4.17887 0.0563819 0.0394233 0.960577 0.0198087 0.00429504 0.0190716 0.00412759 0.00519133 0.0059284 0.207653 0.237136 57.993 -87.8958 126.247 15.9686 145.018 0.000141312 0.267146 192.873 0.310572 0.0673717 0.00409579 0.000561785 0.00138317 0.986984 0.991731 -2.97682e-06 -85.6654 0.0930079 31189 301.958 0.983516 0.319147 0.733058 0.733053 9.99958 2.98207e-06 1.19282e-05 0.131174 0.981955 0.931543 -0.0132929 4.90423e-06 0.503027 -1.90346e-20 7.02255e-24 -1.90275e-20 0.00139544 0.997817 8.59513e-05 0.152596 2.85197 0.00139544 0.997825 0.713685 0.00105171 0.00188007 0.000859513 0.455587 0.00188007 0.438659 0.000128763 1.02 0.887788 0.53465 0.286203 1.71706e-07 3.06385e-09 2385.62 3117.89 -0.0554466 0.482141 0.277527 0.253401 -0.593354 -0.169517 0.496722 -0.267672 -0.22906 1.767 1 0 297.699 0 2.10538 1.765 0.000299851 0.85416 0.659754 0.383552 0.412951 2.1056 132.225 83.896 18.7195 60.8545 0.00402632 0 -40 10
0.866 2.50884e-08 2.53898e-06 0.104366 0.104364 0.0120385 1.14038e-05 0.00115408 0.130458 0.000657849 0.131111 0.879716 101.821 0.24361 0.747317 4.1791 0.0563899 0.0394255 0.960575 0.0198084 0.00429525 0.0190713 0.00412777 0.00519158 0.00592865 0.207663 0.237146 57.9931 -87.8958 126.247 15.9685 145.018 0.00014131 0.267146 192.873 0.310571 0.0673716 0.00409579 0.000561785 0.00138317 0.986984 0.991731 -2.97684e-06 -85.6653 0.093008 31188.9 301.964 0.983516 0.319147 0.733048 0.733043 9.99958 2.98207e-06 1.19282e-05 0.131176 0.98196 0.931545 -0.0132929 4.90426e-06 0.503036 -1.90355e-20 7.02293e-24 -1.90284e-20 0.00139544 0.997817 8.59514e-05 0.152596 2.85197 0.00139544 0.997825 0.713784 0.00105173 0.00188007 0.000859514 0.455587 0.00188007 0.438668 0.000128766 1.02 0.887789 0.53465 0.286204 1.71706e-07 3.06387e-09 2385.61 3117.85 -0.0554446 0.482141 0.277527 0.253398 -0.593355 -0.169517 0.496727 -0.267669 -0.229067 1.768 1 0 297.701 0 2.10554 1.766 0.000299851 0.854143 0.659804 0.3834 0.412978 2.10576 132.234 83.8965 18.7195 60.8547 0.0040263 0 -40 10
0.867 2.51173e-08 2.53898e-06 0.104433 0.104431 0.0120385 1.1417e-05 0.00115408 0.130542 0.000657851 0.131195 0.879783 101.821 0.243602 0.747418 4.17933 0.0563979 0.0394276 0.960572 0.0198082 0.00429546 0.0190711 0.00412794 0.00519184 0.00592891 0.207674 0.237156 57.9932 -87.8958 126.247 15.9685 145.018 0.000141309 0.267146 192.872 0.310571 0.0673716 0.0040958 0.000561786 0.00138318 0.986984 0.991731 -2.97685e-06 -85.6653 0.0930081 31188.9 301.97 0.983515 0.319147 0.733038 0.733034 9.99958 2.98208e-06 1.19282e-05 0.131178 0.981965 0.931546 -0.0132929 4.90429e-06 0.503045 -1.90364e-20 7.0233e-24 -1.90293e-20 0.00139544 0.997817 8.59515e-05 0.152596 2.85197 0.00139544 0.997825 0.713884 0.00105174 0.00188007 0.000859515 0.455587 0.00188007 0.438676 0.00012877 1.02 0.88779 0.53465 0.286206 1.71706e-07 3.06389e-09 2385.59 3117.81 -0.0554427 0.482141 0.277527 0.253396 -0.593355 -0.169517 0.496732 -0.267667 -0.229074 1.769 1 0 297.703 0 2.1057 1.767 0.000299851 0.854126 0.659853 0.383249 0.413004 2.10592 132.242 83.897 18.7195 60.855 0.00402628 0 -40 10
0.868 2.51462e-08 2.53898e-06 0.104501 0.104499 0.0120385 1.14301e-05 0.00115408 0.130626 0.000657854 0.131279 0.87985 101.82 0.243594 0.747518 4.17956 0.0564059 0.0394298 0.96057 0.0198079 0.00429567 0.0190708 0.00412812 0.0051921 0.00592916 0.207684 0.237167 57.9932 -87.8958 126.247 15.9684 145.018 0.000141307 0.267146 192.872 0.310571 0.0673715 0.0040958 0.000561787 0.00138318 0.986984 0.991731 -2.97687e-06 -85.6653 0.0930081 31188.9 301.975 0.983515 0.319147 0.733028 0.733024 9.99958 2.98208e-06 1.19282e-05 0.13118 0.98197 0.931548 -0.0132929 4.90432e-06 0.503054 -1.90372e-20 7.02367e-24 -1.90302e-20 0.00139544 0.997817 8.59516e-05 0.152596 2.85197 0.00139544 0.997825 0.713983 0.00105176 0.00188007 0.000859516 0.455586 0.00188007 0.438684 0.000128773 1.02 0.887791 0.534649 0.286207 1.71706e-07 3.06392e-09 2385.57 3117.76 -0.0554407 0.482141 0.277526 0.253393 -0.593356 -0.169517 0.496737 -0.267665 -0.229081 1.77 1 0 297.706 0 2.10586 1.768 0.00029985 0.854109 0.659903 0.383098 0.413031 2.10607 132.25 83.8975 18.7196 60.8552 0.00402626 0 -40 10
0.869 2.51752e-08 2.53899e-06 0.104568 0.104566 0.0120385 1.14433e-05 0.00115408 0.13071 0.000657856 0.131363 0.879918 101.82 0.243586 0.747618 4.17979 0.0564139 0.039432 0.960568 0.0198076 0.00429588 0.0190706 0.00412829 0.00519236 0.00592942 0.207694 0.237177 57.9933 -87.8958 126.248 15.9684 145.018 0.000141305 0.267146 192.872 0.31057 0.0673715 0.0040958 0.000561787 0.00138318 0.986984 0.991731 -2.97688e-06 -85.6653 0.0930082 31188.9 301.981 0.983515 0.319147 0.733018 0.733014 9.99958 2.98209e-06 1.19282e-05 0.131182 0.981975 0.93155 -0.0132929 4.90435e-06 0.503062 -1.90381e-20 7.02404e-24 -1.90311e-20 0.00139545 0.997817 8.59517e-05 0.152596 2.85198 0.00139545 0.997825 0.714083 0.00105178 0.00188008 0.000859517 0.455586 0.00188007 0.438692 0.000128776 1.02 0.887793 0.534649 0.286209 1.71707e-07 3.06394e-09 2385.56 3117.72 -0.0554388 0.482141 0.277526 0.25339 -0.593356 -0.169517 0.496742 -0.267663 -0.229088 1.771 1 0 297.708 0 2.10601 1.769 0.00029985 0.854092 0.659953 0.382947 0.413057 2.10623 132.259 83.898 18.7196 60.8554 0.00402624 0 -40 10
0.87 2.52041e-08 2.53899e-06 0.104635 0.104633 0.0120385 1.14564e-05 0.00115408 0.130794 0.000657858 0.131448 0.879985 101.82 0.243578 0.747719 4.18002 0.0564219 0.0394341 0.960566 0.0198074 0.00429609 0.0190703 0.00412847 0.00519261 0.00592968 0.207705 0.237187 57.9934 -87.8958 126.248 15.9684 145.018 0.000141303 0.267147 192.872 0.31057 0.0673714 0.00409581 0.000561788 0.00138318 0.986984 0.991731 -2.9769e-06 -85.6653 0.0930083 31188.9 301.987 0.983515 0.319147 0.733009 0.733004 9.99958 2.98209e-06 1.19283e-05 0.131184 0.98198 0.931551 -0.0132929 4.90438e-06 0.503071 -1.9039e-20 7.02441e-24 -1.9032e-20 0.00139545 0.997817 8.59517e-05 0.152596 2.85198 0.00139545 0.997825 0.714182 0.0010518 0.00188008 0.000859517 0.455586 0.00188008 0.4387 0.000128779 1.02 0.887794 0.534649 0.28621 1.71707e-07 3.06396e-09 2385.54 3117.68 -0.0554369 0.482141 0.277526 0.253388 -0.593357 -0.169517 0.496747 -0.267661 -0.229095 1.772 1 0 297.71 0 2.10617 1.77 0.000299849 0.854076 0.660002 0.382797 0.413083 2.10639 132.267 83.8985 18.7196 60.8557 0.00402622 0 -40 10
0.871 2.5233e-08 2.53899e-06 0.104703 0.1047 0.0120384 1.14696e-05 0.00115408 0.130878 0.00065786 0.131532 0.880052 101.82 0.24357 0.747819 4.18025 0.0564299 0.0394363 0.960564 0.0198071 0.0042963 0.0190701 0.00412865 0.00519287 0.00592994 0.207715 0.237197 57.9934 -87.8958 126.248 15.9683 145.018 0.000141301 0.267147 192.872 0.310569 0.0673714 0.00409581 0.000561789 0.00138318 0.986984 0.991731 -2.97691e-06 -85.6653 0.0930084 31188.8 301.993 0.983515 0.319147 0.732999 0.732995 9.99958 2.9821e-06 1.19283e-05 0.131187 0.981984 0.931553 -0.0132929 4.90441e-06 0.50308 -1.90399e-20 7.02479e-24 -1.90329e-20 0.00139545 0.997817 8.59518e-05 0.152596 2.85198 0.00139545 0.997825 0.714282 0.00105182 0.00188008 0.000859518 0.455586 0.00188008 0.438708 0.000128782 1.02 0.887795 0.534648 0.286212 1.71707e-07 3.06398e-09 2385.52 3117.64 -0.055435 0.482141 0.277526 0.253385 -0.593357 -0.169517 0.496752 -0.267659 -0.229102 1.773 1 0 297.712 0 2.10633 1.771 0.000299849 0.85406 0.660052 0.382647 0.41311 2.10655 132.276 83.8989 18.7196 60.8559 0.0040262 0 -40 10
0.872 2.52619e-08 2.53899e-06 0.10477 0.104768 0.0120384 1.14827e-05 0.00115408 0.130962 0.000657862 0.131615 0.880119 101.82 0.243562 0.74792 4.18048 0.0564379 0.0394385 0.960562 0.0198069 0.00429651 0.0190698 0.00412882 0.00519313 0.0059302 0.207725 0.237208 57.9935 -87.8958 126.248 15.9683 145.018 0.000141299 0.267147 192.872 0.310569 0.0673713 0.00409581 0.000561789 0.00138319 0.986984 0.99173 -2.97693e-06 -85.6653 0.0930085 31188.8 301.998 0.983515 0.319147 0.732989 0.732985 9.99958 2.9821e-06 1.19283e-05 0.131189 0.981989 0.931554 -0.0132929 4.90444e-06 0.503089 -1.90408e-20 7.02516e-24 -1.90338e-20 0.00139545 0.997817 8.59519e-05 0.152597 2.85198 0.00139545 0.997825 0.714381 0.00105184 0.00188008 0.000859519 0.455586 0.00188008 0.438716 0.000128786 1.02 0.887796 0.534648 0.286213 1.71707e-07 3.06401e-09 2385.51 3117.6 -0.0554331 0.482141 0.277525 0.253383 -0.593357 -0.169517 0.496756 -0.267657 -0.229109 1.774 1 0 297.715 0 2.10649 1.772 0.000299848 0.854044 0.660101 0.382497 0.413136 2.10671 132.284 83.8994 18.7197 60.8561 0.00402618 0 -40 10
0.873 2.52909e-08 2.53899e-06 0.104837 0.104835 0.0120384 1.14959e-05 0.00115409 0.131046 0.000657864 0.131699 0.880186 101.819 0.243554 0.74802 4.18071 0.0564459 0.0394406 0.960559 0.0198066 0.00429672 0.0190695 0.004129 0.00519339 0.00593045 0.207736 0.237218 57.9936 -87.8958 126.248 15.9683 145.018 0.000141297 0.267147 192.872 0.310568 0.0673713 0.00409582 0.00056179 0.00138319 0.986984 0.99173 -2.97694e-06 -85.6653 0.0930086 31188.8 302.004 0.983515 0.319147 0.73298 0.732975 9.99958 2.98211e-06 1.19283e-05 0.131191 0.981994 0.931556 -0.0132929 4.90447e-06 0.503098 -1.90417e-20 7.02553e-24 -1.90347e-20 0.00139545 0.997817 8.5952e-05 0.152597 2.85198 0.00139545 0.997825 0.714481 0.00105186 0.00188008 0.00085952 0.455585 0.00188008 0.438724 0.000128789 1.02 0.887797 0.534648 0.286215 1.71708e-07 3.06403e-09 2385.49 3117.55 -0.0554313 0.482142 0.277525 0.25338 -0.593358 -0.169517 0.496761 -0.267655 -0.229115 1.775 1 0 297.717 0 2.10665 1.773 0.000299848 0.854028 0.660151 0.382348 0.413162 2.10686 132.293 83.8999 18.7197 60.8563 0.00402616 0 -40 10
0.874 2.53198e-08 2.53899e-06 0.104904 0.104902 0.0120384 1.1509e-05 0.00115409 0.13113 0.000657866 0.131783 0.880254 101.819 0.243546 0.748121 4.18094 0.056454 0.0394428 0.960557 0.0198064 0.00429693 0.0190693 0.00412918 0.00519365 0.00593071 0.207746 0.237229 57.9936 -87.8958 126.248 15.9682 145.018 0.000141296 0.267147 192.871 0.310568 0.0673712 0.00409582 0.000561791 0.00138319 0.986984 0.99173 -2.97696e-06 -85.6653 0.0930087 31188.8 302.01 0.983515 0.319147 0.73297 0.732966 9.99958 2.98211e-06 1.19283e-05 0.131193 0.981999 0.931558 -0.0132929 4.9045e-06 0.503107 -1.90426e-20 7.02591e-24 -1.90356e-20 0.00139545 0.997817 8.59521e-05 0.152597 2.85198 0.00139545 0.997825 0.71458 0.00105188 0.00188008 0.000859521 0.455585 0.00188008 0.438732 0.000128792 1.02 0.887798 0.534647 0.286216 1.71708e-07 3.06405e-09 2385.47 3117.51 -0.0554295 0.482142 0.277525 0.253377 -0.593358 -0.169517 0.496765 -0.267653 -0.229122 1.776 1 0 297.719 0 2.1068 1.774 0.000299848 0.854012 0.6602 0.382199 0.413189 2.10702 132.301 83.9003 18.7197 60.8566 0.00402614 0 -40 10
0.875 2.53487e-08 2.53899e-06 0.104971 0.104969 0.0120384 1.15221e-05 0.00115409 0.131214 0.000657868 0.131867 0.880321 101.819 0.243538 0.748222 4.18117 0.056462 0.039445 0.960555 0.0198061 0.00429714 0.019069 0.00412935 0.00519391 0.00593097 0.207756 0.237239 57.9937 -87.8958 126.249 15.9682 145.018 0.000141294 0.267148 192.871 0.310568 0.0673712 0.00409582 0.000561791 0.00138319 0.986984 0.99173 -2.97697e-06 -85.6653 0.0930087 31188.7 302.015 0.983515 0.319147 0.732961 0.732957 9.99958 2.98212e-06 1.19284e-05 0.131195 0.982003 0.931559 -0.0132929 4.90453e-06 0.503116 -1.90435e-20 7.02628e-24 -1.90365e-20 0.00139545 0.997817 8.59521e-05 0.152597 2.85198 0.00139545 0.997825 0.714679 0.0010519 0.00188008 0.000859521 0.455585 0.00188008 0.43874 0.000128795 1.02 0.887799 0.534647 0.286218 1.71708e-07 3.06407e-09 2385.46 3117.47 -0.0554277 0.482142 0.277524 0.253375 -0.593359 -0.169518 0.49677 -0.267651 -0.229128 1.777 1 0 297.721 0 2.10696 1.775 0.000299847 0.853996 0.660249 0.38205 0.413215 2.10718 132.31 83.9008 18.7198 60.8568 0.00402612 0 -40 10
0.876 2.53777e-08 2.53899e-06 0.105038 0.105036 0.0120384 1.15353e-05 0.00115409 0.131297 0.000657871 0.131951 0.880388 101.819 0.24353 0.748323 4.1814 0.05647 0.0394472 0.960553 0.0198058 0.00429736 0.0190688 0.00412953 0.00519417 0.00593123 0.207767 0.237249 57.9937 -87.8958 126.249 15.9681 145.018 0.000141292 0.267148 192.871 0.310567 0.0673711 0.00409582 0.000561792 0.0013832 0.986984 0.99173 -2.97699e-06 -85.6653 0.0930088 31188.7 302.021 0.983515 0.319147 0.732952 0.732947 9.99958 2.98212e-06 1.19284e-05 0.131197 0.982008 0.931561 -0.0132929 4.90456e-06 0.503124 -1.90444e-20 7.02666e-24 -1.90374e-20 0.00139545 0.997817 8.59522e-05 0.152597 2.85198 0.00139545 0.997825 0.714778 0.00105192 0.00188009 0.000859522 0.455585 0.00188008 0.438748 0.000128799 1.02 0.8878 0.534647 0.286219 1.71709e-07 3.0641e-09 2385.44 3117.43 -0.0554259 0.482142 0.277524 0.253372 -0.593359 -0.169518 0.496774 -0.267648 -0.229135 1.778 1 0 297.723 0 2.10712 1.776 0.000299847 0.85398 0.660299 0.381902 0.413241 2.10734 132.318 83.9013 18.7198 60.857 0.0040261 0 -40 10
0.877 2.54066e-08 2.53899e-06 0.105105 0.105103 0.0120384 1.15484e-05 0.00115409 0.131381 0.000657873 0.132034 0.880456 101.818 0.243522 0.748424 4.18163 0.0564781 0.0394494 0.960551 0.0198056 0.00429757 0.0190685 0.00412971 0.00519443 0.00593149 0.207777 0.23726 57.9938 -87.8959 126.249 15.9681 145.018 0.00014129 0.267148 192.871 0.310567 0.0673711 0.00409583 0.000561793 0.0013832 0.986984 0.99173 -2.977e-06 -85.6652 0.0930089 31188.7 302.027 0.983515 0.319147 0.732943 0.732938 9.99958 2.98213e-06 1.19284e-05 0.131199 0.982013 0.931562 -0.0132929 4.90459e-06 0.503133 -1.90453e-20 7.02703e-24 -1.90383e-20 0.00139545 0.997817 8.59523e-05 0.152597 2.85198 0.00139545 0.997825 0.714878 0.00105194 0.00188009 0.000859523 0.455584 0.00188009 0.438756 0.000128802 1.02 0.887801 0.534647 0.286221 1.71709e-07 3.06412e-09 2385.42 3117.39 -0.0554242 0.482142 0.277524 0.25337 -0.59336 -0.169518 0.496779 -0.267646 -0.229141 1.779 1 0 297.725 0 2.10728 1.777 0.000299846 0.853965 0.660348 0.381754 0.413268 2.10749 132.327 83.9017 18.7198 60.8572 0.00402608 0 -40 10
0.878 2.54355e-08 2.53899e-06 0.105172 0.105169 0.0120384 1.15616e-05 0.00115409 0.131464 0.000657875 0.132118 0.880523 101.818 0.243514 0.748525 4.18187 0.0564861 0.0394516 0.960548 0.0198053 0.00429778 0.0190682 0.00412989 0.00519469 0.00593176 0.207788 0.23727 57.9939 -87.8959 126.249 15.9681 145.018 0.000141288 0.267148 192.871 0.310566 0.067371 0.00409583 0.000561793 0.0013832 0.986983 0.99173 -2.97701e-06 -85.6652 0.093009 31188.7 302.033 0.983515 0.319147 0.732933 0.732929 9.99958 2.98213e-06 1.19284e-05 0.131202 0.982018 0.931564 -0.0132929 4.90461e-06 0.503142 -1.90462e-20 7.0274e-24 -1.90392e-20 0.00139546 0.997817 8.59524e-05 0.152598 2.85198 0.00139546 0.997825 0.714977 0.00105196 0.00188009 0.000859524 0.455584 0.00188009 0.438764 0.000128805 1.02 0.887802 0.534646 0.286222 1.71709e-07 3.06414e-09 2385.41 3117.35 -0.0554225 0.482142 0.277524 0.253368 -0.59336 -0.169518 0.496783 -0.267644 -0.229148 1.78 1 0 297.727 0 2.10743 1.778 0.000299846 0.85395 0.660398 0.381606 0.413294 2.10765 132.335 83.9022 18.7198 60.8575 0.00402606 0 -40 10
0.879 2.54644e-08 2.53899e-06 0.105238 0.105236 0.0120383 1.15747e-05 0.00115409 0.131548 0.000657877 0.132201 0.880591 101.818 0.243506 0.748626 4.1821 0.0564942 0.0394538 0.960546 0.019805 0.00429799 0.019068 0.00413007 0.00519495 0.00593202 0.207798 0.237281 57.9939 -87.8959 126.249 15.968 145.018 0.000141287 0.267148 192.871 0.310566 0.067371 0.00409583 0.000561794 0.0013832 0.986983 0.99173 -2.97703e-06 -85.6652 0.0930091 31188.7 302.038 0.983515 0.319147 0.732924 0.73292 9.99958 2.98214e-06 1.19284e-05 0.131204 0.982022 0.931565 -0.0132929 4.90464e-06 0.503151 -1.90471e-20 7.02778e-24 -1.90401e-20 0.00139546 0.997817 8.59525e-05 0.152598 2.85198 0.00139546 0.997825 0.715076 0.00105198 0.00188009 0.000859525 0.455584 0.00188009 0.438772 0.000128808 1.02 0.887803 0.534646 0.286224 1.71709e-07 3.06416e-09 2385.39 3117.31 -0.0554208 0.482142 0.277523 0.253365 -0.593361 -0.169518 0.496787 -0.267642 -0.229154 1.781 1 0 297.73 0 2.10759 1.779 0.000299845 0.853934 0.660447 0.381459 0.41332 2.10781 132.344 83.9026 18.7199 60.8577 0.00402604 0 -40 10
0.88 2.54934e-08 2.53899e-06 0.105305 0.105303 0.0120383 1.15879e-05 0.00115409 0.131631 0.000657879 0.132285 0.880658 101.818 0.243498 0.748727 4.18233 0.0565022 0.039456 0.960544 0.0198048 0.00429821 0.0190677 0.00413024 0.00519522 0.00593228 0.207809 0.237291 57.994 -87.8959 126.249 15.968 145.018 0.000141285 0.267149 192.87 0.310566 0.0673709 0.00409584 0.000561795 0.0013832 0.986983 0.99173 -2.97704e-06 -85.6652 0.0930092 31188.6 302.044 0.983515 0.319147 0.732915 0.732911 9.99958 2.98214e-06 1.19285e-05 0.131206 0.982027 0.931567 -0.0132929 4.90467e-06 0.50316 -1.9048e-20 7.02815e-24 -1.9041e-20 0.00139546 0.997817 8.59525e-05 0.152598 2.85199 0.00139546 0.997825 0.715175 0.001052 0.00188009 0.000859525 0.455584 0.00188009 0.43878 0.000128811 1.02 0.887804 0.534646 0.286225 1.7171e-07 3.06419e-09 2385.37 3117.28 -0.0554191 0.482142 0.277523 0.253363 -0.593361 -0.169518 0.496791 -0.26764 -0.22916 1.782 1 0 297.732 0 2.10775 1.78 0.000299845 0.853919 0.660496 0.381311 0.413347 2.10797 132.352 83.9031 18.7199 60.8579 0.00402603 0 -40 10
0.881 2.55223e-08 2.53899e-06 0.105372 0.10537 0.0120383 1.1601e-05 0.00115409 0.131715 0.000657881 0.132368 0.880726 101.817 0.24349 0.748828 4.18257 0.0565103 0.0394582 0.960542 0.0198045 0.00429842 0.0190675 0.00413042 0.00519548 0.00593254 0.207819 0.237302 57.9941 -87.8959 126.25 15.9679 145.018 0.000141283 0.267149 192.87 0.310565 0.0673708 0.00409584 0.000561795 0.00138321 0.986983 0.99173 -2.97706e-06 -85.6652 0.0930093 31188.6 302.05 0.983515 0.319147 0.732906 0.732902 9.99958 2.98215e-06 1.19285e-05 0.131208 0.982032 0.931569 -0.0132929 4.9047e-06 0.503169 -1.90489e-20 7.02853e-24 -1.90419e-20 0.00139546 0.997817 8.59526e-05 0.152598 2.85199 0.00139546 0.997824 0.715274 0.00105201 0.00188009 0.000859526 0.455584 0.00188009 0.438788 0.000128815 1.02 0.887806 0.534645 0.286227 1.7171e-07 3.06421e-09 2385.36 3117.24 -0.0554174 0.482142 0.277523 0.25336 -0.593361 -0.169518 0.496795 -0.267638 -0.229166 1.783 1 0 297.734 0 2.10791 1.781 0.000299844 0.853904 0.660546 0.381165 0.413373 2.10813 132.36 83.9035 18.7199 60.8581 0.00402601 0 -40 10
0.882 2.55512e-08 2.53899e-06 0.105438 0.105436 0.0120383 1.16142e-05 0.00115409 0.131798 0.000657883 0.132451 0.880793 101.817 0.243482 0.748929 4.1828 0.0565184 0.0394604 0.96054 0.0198043 0.00429863 0.0190672 0.0041306 0.00519574 0.0059328 0.20783 0.237312 57.9941 -87.8959 126.25 15.9679 145.018 0.000141281 0.267149 192.87 0.310565 0.0673708 0.00409584 0.000561796 0.00138321 0.986983 0.99173 -2.97707e-06 -85.6652 0.0930093 31188.6 302.056 0.983515 0.319147 0.732898 0.732893 9.99958 2.98215e-06 1.19285e-05 0.13121 0.982036 0.93157 -0.0132929 4.90473e-06 0.503178 -1.90498e-20 7.02891e-24 -1.90428e-20 0.00139546 0.997817 8.59527e-05 0.152598 2.85199 0.00139546 0.997824 0.715373 0.00105203 0.00188009 0.000859527 0.455583 0.00188009 0.438796 0.000128818 1.02 0.887807 0.534645 0.286228 1.7171e-07 3.06423e-09 2385.34 3117.2 -0.0554158 0.482142 0.277522 0.253358 -0.593362 -0.169518 0.496799 -0.267636 -0.229173 1.784 1 0 297.736 0 2.10807 1.782 0.000299844 0.85389 0.660595 0.381018 0.413399 2.10828 132.369 83.9039 18.7199 60.8583 0.00402599 0 -40 10
0.883 2.55802e-08 2.53899e-06 0.105505 0.105503 0.0120383 1.16273e-05 0.00115409 0.131881 0.000657885 0.132534 0.880861 101.817 0.243474 0.74903 4.18303 0.0565265 0.0394626 0.960537 0.019804 0.00429885 0.0190669 0.00413078 0.005196 0.00593307 0.20784 0.237323 57.9942 -87.8959 126.25 15.9679 145.018 0.00014128 0.267149 192.87 0.310564 0.0673707 0.00409585 0.000561797 0.00138321 0.986983 0.99173 -2.97709e-06 -85.6652 0.0930094 31188.6 302.062 0.983515 0.319147 0.732889 0.732884 9.99958 2.98216e-06 1.19285e-05 0.131213 0.982041 0.931572 -0.0132929 4.90476e-06 0.503187 -1.90507e-20 7.02928e-24 -1.90437e-20 0.00139546 0.997817 8.59528e-05 0.152598 2.85199 0.00139546 0.997824 0.715472 0.00105205 0.0018801 0.000859528 0.455583 0.00188009 0.438804 0.000128821 1.02 0.887808 0.534645 0.28623 1.7171e-07 3.06425e-09 2385.32 3117.16 -0.0554142 0.482142 0.277522 0.253355 -0.593362 -0.169518 0.496803 -0.267634 -0.229179 1.785 1 0 297.738 0 2.10822 1.783 0.000299843 0.853875 0.660645 0.380872 0.413426 2.10844 132.377 83.9044 18.72 60.8585 0.00402597 0 -40 10
0.884 2.56091e-08 2.53899e-06 0.105571 0.105569 0.0120383 1.16405e-05 0.00115409 0.131964 0.000657887 0.132617 0.880929 101.817 0.243465 0.749132 4.18327 0.0565345 0.0394648 0.960535 0.0198037 0.00429906 0.0190667 0.00413096 0.00519627 0.00593333 0.207851 0.237333 57.9942 -87.8959 126.25 15.9678 145.018 0.000141278 0.267149 192.87 0.310564 0.0673707 0.00409585 0.000561797 0.00138321 0.986983 0.99173 -2.9771e-06 -85.6652 0.0930095 31188.5 302.067 0.983515 0.319147 0.73288 0.732876 9.99958 2.98216e-06 1.19285e-05 0.131215 0.982045 0.931573 -0.0132929 4.90479e-06 0.503196 -1.90516e-20 7.02966e-24 -1.90446e-20 0.00139546 0.997817 8.59528e-05 0.152598 2.85199 0.00139546 0.997824 0.715571 0.00105207 0.0018801 0.000859528 0.455583 0.0018801 0.438812 0.000128824 1.02 0.887809 0.534644 0.286231 1.71711e-07 3.06428e-09 2385.31 3117.12 -0.0554126 0.482142 0.277522 0.253353 -0.593363 -0.169518 0.496807 -0.267632 -0.229184 1.786 1 0 297.74 0 2.10838 1.784 0.000299843 0.85386 0.660694 0.380726 0.413452 2.1086 132.386 83.9048 18.72 60.8587 0.00402595 0 -40 10
0.885 2.5638e-08 2.53899e-06 0.105638 0.105636 0.0120383 1.16536e-05 0.00115409 0.132047 0.000657889 0.132701 0.880996 101.816 0.243457 0.749233 4.1835 0.0565426 0.039467 0.960533 0.0198035 0.00429928 0.0190664 0.00413114 0.00519653 0.00593359 0.207861 0.237344 57.9943 -87.8959 126.25 15.9678 145.018 0.000141276 0.267149 192.87 0.310563 0.0673706 0.00409585 0.000561798 0.00138321 0.986983 0.99173 -2.97712e-06 -85.6652 0.0930096 31188.5 302.073 0.983515 0.319147 0.732871 0.732867 9.99958 2.98217e-06 1.19286e-05 0.131217 0.98205 0.931575 -0.0132929 4.90482e-06 0.503205 -1.90525e-20 7.03003e-24 -1.90455e-20 0.00139546 0.997817 8.59529e-05 0.152599 2.85199 0.00139546 0.997824 0.71567 0.00105209 0.0018801 0.000859529 0.455583 0.0018801 0.43882 0.000128827 1.02 0.88781 0.534644 0.286233 1.71711e-07 3.0643e-09 2385.29 3117.08 -0.055411 0.482142 0.277522 0.253351 -0.593363 -0.169518 0.496811 -0.26763 -0.22919 1.787 1 0 297.741 0 2.10854 1.785 0.000299843 0.853846 0.660743 0.380581 0.413478 2.10875 132.394 83.9052 18.72 60.8589 0.00402594 0 -40 10
0.886 2.56669e-08 2.53899e-06 0.105704 0.105702 0.0120382 1.16668e-05 0.00115409 0.13213 0.000657891 0.132784 0.881064 101.816 0.243449 0.749335 4.18374 0.0565507 0.0394693 0.960531 0.0198032 0.00429949 0.0190661 0.00413132 0.0051968 0.00593386 0.207872 0.237354 57.9944 -87.8959 126.25 15.9678 145.018 0.000141275 0.26715 192.869 0.310563 0.0673706 0.00409585 0.000561799 0.00138322 0.986983 0.99173 -2.97713e-06 -85.6652 0.0930097 31188.5 302.079 0.983515 0.319147 0.732863 0.732858 9.99958 2.98217e-06 1.19286e-05 0.131219 0.982055 0.931576 -0.0132929 4.90485e-06 0.503214 -1.90534e-20 7.03041e-24 -1.90464e-20 0.00139546 0.997817 8.5953e-05 0.152599 2.85199 0.00139546 0.997824 0.715769 0.00105211 0.0018801 0.00085953 0.455582 0.0018801 0.438828 0.000128831 1.02 0.887811 0.534644 0.286234 1.71711e-07 3.06432e-09 2385.27 3117.05 -0.0554095 0.482142 0.277521 0.253348 -0.593364 -0.169518 0.496814 -0.267627 -0.229196 1.788 1 0 297.743 0 2.10869 1.786 0.000299842 0.853832 0.660792 0.380436 0.413504 2.10891 132.403 83.9057 18.72 60.8591 0.00402592 0 -40 10
0.887 2.56959e-08 2.53899e-06 0.105771 0.105768 0.0120382 1.16799e-05 0.00115409 0.132213 0.000657893 0.132866 0.881132 101.816 0.243441 0.749436 4.18398 0.0565588 0.0394715 0.960529 0.0198029 0.00429971 0.0190659 0.0041315 0.00519706 0.00593412 0.207882 0.237365 57.9944 -87.8959 126.251 15.9677 145.018 0.000141273 0.26715 192.869 0.310563 0.0673705 0.00409586 0.000561799 0.00138322 0.986983 0.99173 -2.97715e-06 -85.6652 0.0930098 31188.5 302.085 0.983515 0.319147 0.732854 0.73285 9.99958 2.98217e-06 1.19286e-05 0.131221 0.982059 0.931578 -0.0132928 4.90488e-06 0.503223 -1.90543e-20 7.03079e-24 -1.90473e-20 0.00139547 0.997817 8.59531e-05 0.152599 2.85199 0.00139547 0.997824 0.715868 0.00105213 0.0018801 0.000859531 0.455582 0.0018801 0.438836 0.000128834 1.02 0.887812 0.534644 0.286236 1.71711e-07 3.06434e-09 2385.26 3117.01 -0.0554079 0.482143 0.277521 0.253346 -0.593364 -0.169518 0.496818 -0.267625 -0.229202 1.789 1 0 297.745 0 2.10885 1.787 0.000299842 0.853818 0.660842 0.380291 0.41353 2.10907 132.411 83.9061 18.7201 60.8593 0.0040259 0 -40 10
0.888 2.57248e-08 2.539e-06 0.105837 0.105835 0.0120382 1.16931e-05 0.00115409 0.132296 0.000657895 0.132949 0.8812 101.816 0.243433 0.749538 4.18421 0.0565669 0.0394737 0.960526 0.0198027 0.00429992 0.0190656 0.00413168 0.00519733 0.00593439 0.207893 0.237375 57.9945 -87.8959 126.251 15.9677 145.018 0.000141271 0.26715 192.869 0.310562 0.0673705 0.00409586 0.0005618 0.00138322 0.986983 0.99173 -2.97716e-06 -85.6651 0.0930099 31188.5 302.091 0.983515 0.319147 0.732846 0.732841 9.99958 2.98218e-06 1.19286e-05 0.131224 0.982064 0.931579 -0.0132928 4.90491e-06 0.503232 -1.90552e-20 7.03116e-24 -1.90482e-20 0.00139547 0.997817 8.59532e-05 0.152599 2.85199 0.00139547 0.997824 0.715967 0.00105215 0.0018801 0.000859532 0.455582 0.0018801 0.438844 0.000128837 1.02 0.887813 0.534643 0.286237 1.71712e-07 3.06437e-09 2385.24 3116.97 -0.0554064 0.482143 0.277521 0.253344 -0.593364 -0.169518 0.496822 -0.267623 -0.229208 1.79 1 0 297.747 0 2.10901 1.788 0.000299841 0.853804 0.660891 0.380146 0.413557 2.10923 132.419 83.9065 18.7201 60.8595 0.00402588 0 -40 10
0.889 2.57537e-08 2.539e-06 0.105903 0.105901 0.0120382 1.17062e-05 0.00115409 0.132379 0.000657897 0.133032 0.881268 101.816 0.243425 0.74964 4.18445 0.056575 0.0394759 0.960524 0.0198024 0.00430014 0.0190653 0.00413187 0.00519759 0.00593465 0.207904 0.237386 57.9946 -87.8959 126.251 15.9676 145.018 0.00014127 0.26715 192.869 0.310562 0.0673704 0.00409586 0.000561801 0.00138322 0.986983 0.99173 -2.97718e-06 -85.6651 0.0930099 31188.4 302.097 0.983515 0.319147 0.732837 0.732833 9.99958 2.98218e-06 1.19286e-05 0.131226 0.982068 0.931581 -0.0132928 4.90494e-06 0.503242 -1.90561e-20 7.03154e-24 -1.90491e-20 0.00139547 0.997817 8.59532e-05 0.152599 2.85199 0.00139547 0.997824 0.716066 0.00105217 0.0018801 0.000859532 0.455582 0.0018801 0.438852 0.00012884 1.02 0.887814 0.534643 0.286239 1.71712e-07 3.06439e-09 2385.22 3116.94 -0.0554049 0.482143 0.27752 0.253342 -0.593365 -0.169518 0.496825 -0.267621 -0.229213 1.791 1 0 297.749 0 2.10917 1.789 0.000299841 0.85379 0.66094 0.380002 0.413583 2.10938 132.428 83.9069 18.7201 60.8597 0.00402587 0 -40 10
0.89 2.57826e-08 2.539e-06 0.105969 0.105967 0.0120382 1.17194e-05 0.00115409 0.132462 0.0006579 0.133115 0.881336 101.815 0.243417 0.749741 4.18469 0.0565831 0.0394782 0.960522 0.0198021 0.00430035 0.0190651 0.00413205 0.00519786 0.00593492 0.207914 0.237397 57.9946 -87.8959 126.251 15.9676 145.018 0.000141268 0.26715 192.869 0.310561 0.0673704 0.00409587 0.000561801 0.00138322 0.986983 0.99173 -2.97719e-06 -85.6651 0.09301 31188.4 302.102 0.983515 0.319147 0.732829 0.732825 9.99958 2.98219e-06 1.19287e-05 0.131228 0.982073 0.931582 -0.0132928 4.90497e-06 0.503251 -1.9057e-20 7.03192e-24 -1.905e-20 0.00139547 0.997817 8.59533e-05 0.152599 2.85199 0.00139547 0.997824 0.716164 0.00105219 0.00188011 0.000859533 0.455582 0.0018801 0.43886 0.000128843 1.02 0.887815 0.534643 0.28624 1.71712e-07 3.06441e-09 2385.21 3116.9 -0.0554035 0.482143 0.27752 0.253339 -0.593365 -0.169519 0.496829 -0.267619 -0.229219 1.792 1 0 297.751 0 2.10932 1.79 0.00029984 0.853776 0.660989 0.379858 0.413609 2.10954 132.436 83.9073 18.7201 60.8599 0.00402585 0 -40 10
0.891 2.58116e-08 2.539e-06 0.106035 0.106033 0.0120382 1.17325e-05 0.00115409 0.132544 0.000657902 0.133198 0.881404 101.815 0.243409 0.749843 4.18493 0.0565913 0.0394804 0.96052 0.0198019 0.00430057 0.0190648 0.00413223 0.00519812 0.00593518 0.207925 0.237407 57.9947 -87.8959 126.251 15.9676 145.018 0.000141267 0.267151 192.869 0.310561 0.0673703 0.00409587 0.000561802 0.00138323 0.986983 0.99173 -2.97721e-06 -85.6651 0.0930101 31188.4 302.108 0.983515 0.319147 0.732821 0.732816 9.99958 2.98219e-06 1.19287e-05 0.13123 0.982077 0.931584 -0.0132928 4.905e-06 0.50326 -1.9058e-20 7.0323e-24 -1.90509e-20 0.00139547 0.997817 8.59534e-05 0.1526 2.852 0.00139547 0.997824 0.716263 0.00105221 0.00188011 0.000859534 0.455581 0.00188011 0.438868 0.000128846 1.02 0.887816 0.534642 0.286242 1.71713e-07 3.06443e-09 2385.19 3116.87 -0.055402 0.482143 0.27752 0.253337 -0.593366 -0.169519 0.496832 -0.267617 -0.229224 1.793 1 0 297.753 0 2.10948 1.791 0.00029984 0.853762 0.661038 0.379714 0.413635 2.1097 132.445 83.9077 18.7202 60.8601 0.00402583 0 -40 10
0.892 2.58405e-08 2.539e-06 0.106101 0.106099 0.0120382 1.17457e-05 0.00115409 0.132627 0.000657904 0.13328 0.881472 101.815 0.243401 0.749945 4.18516 0.0565994 0.0394827 0.960517 0.0198016 0.00430079 0.0190645 0.00413241 0.00519839 0.00593545 0.207936 0.237418 57.9948 -87.8959 126.251 15.9675 145.018 0.000141265 0.267151 192.868 0.31056 0.0673703 0.00409587 0.000561803 0.00138323 0.986983 0.99173 -2.97722e-06 -85.6651 0.0930102 31188.4 302.114 0.983515 0.319147 0.732813 0.732808 9.99958 2.9822e-06 1.19287e-05 0.131232 0.982082 0.931585 -0.0132928 4.90503e-06 0.503269 -1.90589e-20 7.03267e-24 -1.90518e-20 0.00139547 0.997817 8.59535e-05 0.1526 2.852 0.00139547 0.997824 0.716362 0.00105223 0.00188011 0.000859535 0.455581 0.00188011 0.438876 0.00012885 1.02 0.887818 0.534642 0.286243 1.71713e-07 3.06446e-09 2385.17 3116.83 -0.0554006 0.482143 0.27752 0.253335 -0.593366 -0.169519 0.496835 -0.267615 -0.22923 1.794 1 0 297.754 0 2.10964 1.792 0.000299839 0.853749 0.661088 0.379571 0.413661 2.10985 132.453 83.9081 18.7202 60.8603 0.00402582 0 -40 10
0.893 2.58694e-08 2.539e-06 0.106167 0.106165 0.0120382 1.17588e-05 0.00115409 0.132709 0.000657906 0.133363 0.88154 101.815 0.243392 0.750047 4.1854 0.0566075 0.0394849 0.960515 0.0198013 0.00430101 0.0190643 0.00413259 0.00519866 0.00593572 0.207946 0.237429 57.9948 -87.8959 126.251 15.9675 145.018 0.000141264 0.267151 192.868 0.31056 0.0673702 0.00409587 0.000561803 0.00138323 0.986983 0.99173 -2.97724e-06 -85.6651 0.0930103 31188.3 302.12 0.983515 0.319147 0.732805 0.7328 9.99958 2.9822e-06 1.19287e-05 0.131235 0.982086 0.931586 -0.0132928 4.90505e-06 0.503278 -1.90598e-20 7.03305e-24 -1.90527e-20 0.00139547 0.997817 8.59536e-05 0.1526 2.852 0.00139547 0.997824 0.716461 0.00105224 0.00188011 0.000859536 0.455581 0.00188011 0.438884 0.000128853 1.02 0.887819 0.534642 0.286245 1.71713e-07 3.06448e-09 2385.16 3116.79 -0.0553992 0.482143 0.277519 0.253333 -0.593366 -0.169519 0.496839 -0.267613 -0.229235 1.795 1 0 297.756 0 2.10979 1.793 0.000299839 0.853736 0.661137 0.379428 0.413688 2.11001 132.462 83.9085 18.7202 60.8605 0.0040258 0 -40 10
0.894 2.58983e-08 2.539e-06 0.106233 0.106231 0.0120381 1.1772e-05 0.00115409 0.132792 0.000657908 0.133445 0.881608 101.814 0.243384 0.750149 4.18564 0.0566157 0.0394872 0.960513 0.0198011 0.00430122 0.019064 0.00413278 0.00519893 0.00593599 0.207957 0.237439 57.9949 -87.8959 126.252 15.9675 145.018 0.000141262 0.267151 192.868 0.31056 0.0673702 0.00409588 0.000561804 0.00138323 0.986983 0.99173 -2.97725e-06 -85.6651 0.0930104 31188.3 302.126 0.983515 0.319147 0.732796 0.732792 9.99958 2.98221e-06 1.19287e-05 0.131237 0.982091 0.931588 -0.0132928 4.90508e-06 0.503287 -1.90607e-20 7.03343e-24 -1.90536e-20 0.00139547 0.997817 8.59536e-05 0.1526 2.852 0.00139547 0.997824 0.716559 0.00105226 0.00188011 0.000859536 0.455581 0.00188011 0.438892 0.000128856 1.02 0.88782 0.534641 0.286246 1.71713e-07 3.0645e-09 2385.14 3116.76 -0.0553978 0.482143 0.277519 0.253331 -0.593367 -0.169519 0.496842 -0.267611 -0.22924 1.796 1 0 297.758 0 2.10995 1.794 0.000299838 0.853722 0.661186 0.379286 0.413714 2.11017 132.47 83.9089 18.7202 60.8607 0.00402578 0 -40 10
0.895 2.59273e-08 2.539e-06 0.106299 0.106297 0.0120381 1.17851e-05 0.00115409 0.132874 0.00065791 0.133528 0.881676 101.814 0.243376 0.750251 4.18588 0.0566238 0.0394895 0.960511 0.0198008 0.00430144 0.0190637 0.00413296 0.00519919 0.00593625 0.207968 0.23745 57.9949 -87.8959 126.252 15.9674 145.018 0.00014126 0.267151 192.868 0.310559 0.0673701 0.00409588 0.000561805 0.00138324 0.986983 0.99173 -2.97727e-06 -85.6651 0.0930105 31188.3 302.132 0.983515 0.319147 0.732788 0.732784 9.99958 2.98221e-06 1.19287e-05 0.131239 0.982095 0.931589 -0.0132928 4.90511e-06 0.503296 -1.90616e-20 7.03381e-24 -1.90546e-20 0.00139547 0.997817 8.59537e-05 0.1526 2.852 0.00139547 0.997824 0.716658 0.00105228 0.00188011 0.000859537 0.45558 0.00188011 0.4389 0.000128859 1.02 0.887821 0.534641 0.286248 1.71714e-07 3.06453e-09 2385.12 3116.73 -0.0553965 0.482143 0.277519 0.253328 -0.593367 -0.169519 0.496845 -0.267609 -0.229246 1.797 1 0 297.76 0 2.11011 1.795 0.000299838 0.853709 0.661235 0.379143 0.41374 2.11032 132.478 83.9093 18.7202 60.8609 0.00402577 0 -40 10
0.896 2.59562e-08 2.539e-06 0.106365 0.106363 0.0120381 1.17983e-05 0.00115409 0.132957 0.000657912 0.13361 0.881744 101.814 0.243368 0.750353 4.18612 0.0566319 0.0394917 0.960508 0.0198005 0.00430166 0.0190635 0.00413314 0.00519946 0.00593652 0.207978 0.237461 57.995 -87.8959 126.252 15.9674 145.018 0.000141259 0.267152 192.868 0.310559 0.0673701 0.00409588 0.000561805 0.00138324 0.986983 0.99173 -2.97728e-06 -85.6651 0.0930105 31188.3 302.138 0.983515 0.319147 0.732781 0.732776 9.99958 2.98222e-06 1.19288e-05 0.131241 0.9821 0.931591 -0.0132928 4.90514e-06 0.503306 -1.90625e-20 7.03419e-24 -1.90555e-20 0.00139548 0.997817 8.59538e-05 0.1526 2.852 0.00139548 0.997824 0.716756 0.0010523 0.00188011 0.000859538 0.45558 0.00188011 0.438907 0.000128862 1.02 0.887822 0.534641 0.286249 1.71714e-07 3.06455e-09 2385.11 3116.69 -0.0553952 0.482143 0.277518 0.253326 -0.593368 -0.169519 0.496848 -0.267606 -0.229251 1.798 1 0 297.761 0 2.11027 1.796 0.000299837 0.853696 0.661284 0.379001 0.413766 2.11048 132.487 83.9097 18.7203 60.8611 0.00402575 0 -40 10
0.897 2.59851e-08 2.539e-06 0.106431 0.106429 0.0120381 1.18114e-05 0.00115409 0.133039 0.000657914 0.133692 0.881812 101.814 0.24336 0.750455 4.18636 0.0566401 0.039494 0.960506 0.0198003 0.00430188 0.0190632 0.00413333 0.00519973 0.00593679 0.207989 0.237472 57.9951 -87.8959 126.252 15.9673 145.018 0.000141257 0.267152 192.868 0.310558 0.06737 0.00409589 0.000561806 0.00138324 0.986983 0.99173 -2.9773e-06 -85.6651 0.0930106 31188.3 302.144 0.983515 0.319147 0.732773 0.732768 9.99958 2.98222e-06 1.19288e-05 0.131244 0.982104 0.931592 -0.0132928 4.90517e-06 0.503315 -1.90634e-20 7.03457e-24 -1.90564e-20 0.00139548 0.997817 8.59539e-05 0.1526 2.852 0.00139548 0.997824 0.716855 0.00105232 0.00188012 0.000859539 0.45558 0.00188012 0.438915 0.000128866 1.02 0.887823 0.53464 0.286251 1.71714e-07 3.06457e-09 2385.09 3116.66 -0.0553938 0.482143 0.277518 0.253324 -0.593368 -0.169519 0.496851 -0.267604 -0.229256 1.799 1 0 297.763 0 2.11042 1.797 0.000299837 0.853684 0.661333 0.378859 0.413792 2.11064 132.495 83.9101 18.7203 60.8613 0.00402574 0 -40 10
0.898 2.6014e-08 2.539e-06 0.106497 0.106495 0.0120381 1.18246e-05 0.00115409 0.133121 0.000657916 0.133774 0.881881 101.813 0.243352 0.750558 4.1866 0.0566483 0.0394963 0.960504 0.0198 0.0043021 0.0190629 0.00413351 0.0052 0.00593706 0.208 0.237482 57.9951 -87.8959 126.252 15.9673 145.018 0.000141256 0.267152 192.867 0.310558 0.06737 0.00409589 0.000561807 0.00138324 0.986983 0.99173 -2.97731e-06 -85.6651 0.0930107 31188.2 302.15 0.983515 0.319147 0.732765 0.732761 9.99958 2.98223e-06 1.19288e-05 0.131246 0.982109 0.931594 -0.0132928 4.9052e-06 0.503324 -1.90643e-20 7.03495e-24 -1.90573e-20 0.00139548 0.997817 8.5954e-05 0.152601 2.852 0.00139548 0.997824 0.716953 0.00105234 0.00188012 0.00085954 0.45558 0.00188012 0.438923 0.000128869 1.02 0.887824 0.53464 0.286252 1.71714e-07 3.06459e-09 2385.07 3116.62 -0.0553926 0.482143 0.277518 0.253322 -0.593368 -0.169519 0.496854 -0.267602 -0.229261 1.8 1 0 297.765 0 2.11058 1.798 0.000299837 0.853671 0.661382 0.378718 0.413818 2.1108 132.504 83.9105 18.7203 60.8615 0.00402572 0 -40 10
0.899 2.6043e-08 2.539e-06 0.106563 0.106561 0.0120381 1.18377e-05 0.00115409 0.133203 0.000657918 0.133856 0.881949 101.813 0.243344 0.75066 4.18684 0.0566564 0.0394985 0.960501 0.0197997 0.00430232 0.0190627 0.00413369 0.00520027 0.00593733 0.208011 0.237493 57.9952 -87.8959 126.252 15.9673 145.018 0.000141254 0.267152 192.867 0.310558 0.0673699 0.00409589 0.000561807 0.00138324 0.986983 0.99173 -2.97732e-06 -85.665 0.0930108 31188.2 302.156 0.983515 0.319147 0.732757 0.732753 9.99958 2.98223e-06 1.19288e-05 0.131248 0.982113 0.931595 -0.0132928 4.90523e-06 0.503333 -1.90652e-20 7.03532e-24 -1.90582e-20 0.00139548 0.997817 8.5954e-05 0.152601 2.852 0.00139548 0.997824 0.717052 0.00105236 0.00188012 0.00085954 0.45558 0.00188012 0.438931 0.000128872 1.02 0.887825 0.53464 0.286254 1.71715e-07 3.06462e-09 2385.06 3116.59 -0.0553913 0.482143 0.277518 0.25332 -0.593369 -0.169519 0.496857 -0.2676 -0.229266 1.801 1 0 297.766 0 2.11074 1.799 0.000299836 0.853658 0.661432 0.378577 0.413844 2.11095 132.512 83.9109 18.7203 60.8617 0.0040257 0 -40 10
0.9 2.60719e-08 2.539e-06 0.106628 0.106626 0.0120381 1.18509e-05 0.00115409 0.133285 0.00065792 0.133939 0.882017 101.813 0.243335 0.750762 4.18709 0.0566646 0.0395008 0.960499 0.0197995 0.00430254 0.0190624 0.00413388 0.00520054 0.0059376 0.208022 0.237504 57.9953 -87.8959 126.252 15.9672 145.018 0.000141253 0.267152 192.867 0.310557 0.0673699 0.0040959 0.000561808 0.00138325 0.986983 0.99173 -2.97734e-06 -85.665 0.0930109 31188.2 302.162 0.983515 0.319147 0.73275 0.732745 9.99958 2.98224e-06 1.19288e-05 0.13125 0.982117 0.931596 -0.0132928 4.90526e-06 0.503342 -1.90661e-20 7.0357e-24 -1.90591e-20 0.00139548 0.997817 8.59541e-05 0.152601 2.852 0.00139548 0.997824 0.71715 0.00105238 0.00188012 0.000859541 0.455579 0.00188012 0.438939 0.000128875 1.02 0.887826 0.53464 0.286255 1.71715e-07 3.06464e-09 2385.04 3116.56 -0.05539 0.482144 0.277517 0.253318 -0.593369 -0.169519 0.49686 -0.267598 -0.229271 1.802 1 0 297.768 0 2.11089 1.8 0.000299836 0.853646 0.661481 0.378436 0.413871 2.11111 132.52 83.9113 18.7204 60.8618 0.00402569 0 -40 10
0.901 2.61008e-08 2.539e-06 0.106694 0.106692 0.012038 1.1864e-05 0.00115409 0.133367 0.000657922 0.134021 0.882086 101.813 0.243327 0.750865 4.18733 0.0566728 0.0395031 0.960497 0.0197992 0.00430276 0.0190621 0.00413406 0.00520081 0.00593787 0.208032 0.237515 57.9953 -87.8959 126.253 15.9672 145.018 0.000141251 0.267152 192.867 0.310557 0.0673698 0.0040959 0.000561809 0.00138325 0.986983 0.99173 -2.97735e-06 -85.665 0.093011 31188.2 302.168 0.983515 0.319147 0.732742 0.732738 9.99958 2.98224e-06 1.19289e-05 0.131253 0.982122 0.931598 -0.0132928 4.90529e-06 0.503352 -1.90671e-20 7.03608e-24 -1.906e-20 0.00139548 0.997817 8.59542e-05 0.152601 2.852 0.00139548 0.997824 0.717249 0.0010524 0.00188012 0.000859542 0.455579 0.00188012 0.438947 0.000128878 1.02 0.887827 0.534639 0.286257 1.71715e-07 3.06466e-09 2385.02 3116.52 -0.0553888 0.482144 0.277517 0.253316 -0.593369 -0.169519 0.496863 -0.267596 -0.229276 1.803 1 0 297.77 0 2.11105 1.801 0.000299835 0.853634 0.66153 0.378295 0.413897 2.11126 132.529 83.9116 18.7204 60.862 0.00402567 0 -40 10
0.902 2.61298e-08 2.539e-06 0.106759 0.106757 0.012038 1.18772e-05 0.00115409 0.133449 0.000657924 0.134102 0.882154 101.812 0.243319 0.750967 4.18757 0.0566809 0.0395054 0.960495 0.0197989 0.00430298 0.0190619 0.00413425 0.00520108 0.00593814 0.208043 0.237526 57.9954 -87.8959 126.253 15.9672 145.019 0.00014125 0.267153 192.867 0.310556 0.0673698 0.0040959 0.000561809 0.00138325 0.986983 0.99173 -2.97737e-06 -85.665 0.0930111 31188.1 302.174 0.983515 0.319147 0.732734 0.73273 9.99958 2.98225e-06 1.19289e-05 0.131255 0.982126 0.931599 -0.0132928 4.90532e-06 0.503361 -1.9068e-20 7.03646e-24 -1.90609e-20 0.00139548 0.997817 8.59543e-05 0.152601 2.85201 0.00139548 0.997824 0.717347 0.00105242 0.00188012 0.000859543 0.455579 0.00188012 0.438955 0.000128881 1.02 0.887828 0.534639 0.286258 1.71715e-07 3.06468e-09 2385.01 3116.49 -0.0553876 0.482144 0.277517 0.253314 -0.59337 -0.169519 0.496865 -0.267594 -0.229281 1.804 1 0 297.771 0 2.11121 1.802 0.000299835 0.853621 0.661579 0.378155 0.413923 2.11142 132.537 83.912 18.7204 60.8622 0.00402566 0 -40 10
0.903 2.61587e-08 2.539e-06 0.106825 0.106823 0.012038 1.18903e-05 0.00115409 0.133531 0.000657926 0.134184 0.882223 101.812 0.243311 0.75107 4.18781 0.0566891 0.0395077 0.960492 0.0197986 0.0043032 0.0190616 0.00413443 0.00520135 0.00593841 0.208054 0.237536 57.9955 -87.8959 126.253 15.9671 145.019 0.000141249 0.267153 192.867 0.310556 0.0673697 0.0040959 0.00056181 0.00138325 0.986983 0.99173 -2.97738e-06 -85.665 0.0930111 31188.1 302.179 0.983515 0.319147 0.732727 0.732723 9.99958 2.98225e-06 1.19289e-05 0.131257 0.98213 0.9316 -0.0132928 4.90535e-06 0.50337 -1.90689e-20 7.03684e-24 -1.90619e-20 0.00139548 0.997817 8.59544e-05 0.152601 2.85201 0.00139548 0.997824 0.717445 0.00105244 0.00188013 0.000859544 0.455579 0.00188012 0.438963 0.000128885 1.02 0.88783 0.534639 0.28626 1.71716e-07 3.06471e-09 2384.99 3116.46 -0.0553864 0.482144 0.277517 0.253312 -0.59337 -0.169519 0.496868 -0.267592 -0.229285 1.805 1 0 297.773 0 2.11136 1.803 0.000299834 0.853609 0.661628 0.378015 0.413949 2.11158 132.545 83.9124 18.7204 60.8624 0.00402564 0 -40 10
0.904 2.61876e-08 2.539e-06 0.10689 0.106888 0.012038 1.19035e-05 0.00115409 0.133613 0.000657928 0.134266 0.882291 101.812 0.243303 0.751173 4.18806 0.0566973 0.03951 0.96049 0.0197984 0.00430342 0.0190613 0.00413462 0.00520162 0.00593868 0.208065 0.237547 57.9955 -87.896 126.253 15.9671 145.019 0.000141247 0.267153 192.866 0.310555 0.0673697 0.00409591 0.000561811 0.00138325 0.986983 0.99173 -2.9774e-06 -85.665 0.0930112 31188.1 302.185 0.983515 0.319147 0.732719 0.732715 9.99958 2.98226e-06 1.19289e-05 0.131259 0.982135 0.931602 -0.0132928 4.90538e-06 0.50338 -1.90698e-20 7.03723e-24 -1.90628e-20 0.00139548 0.997817 8.59544e-05 0.152601 2.85201 0.00139548 0.997823 0.717544 0.00105246 0.00188013 0.000859544 0.455578 0.00188013 0.438971 0.000128888 1.02 0.887831 0.534638 0.286261 1.71716e-07 3.06473e-09 2384.97 3116.43 -0.0553852 0.482144 0.277516 0.25331 -0.59337 -0.169519 0.496871 -0.26759 -0.22929 1.806 1 0 297.774 0 2.11152 1.804 0.000299834 0.853597 0.661677 0.377876 0.413975 2.11173 132.554 83.9128 18.7204 60.8625 0.00402563 0 -40 10
0.905 2.62165e-08 2.53901e-06 0.106956 0.106954 0.012038 1.19166e-05 0.00115409 0.133695 0.00065793 0.134348 0.88236 101.812 0.243295 0.751276 4.1883 0.0567055 0.0395123 0.960488 0.0197981 0.00430364 0.019061 0.0041348 0.0052019 0.00593895 0.208076 0.237558 57.9956 -87.896 126.253 15.967 145.019 0.000141246 0.267153 192.866 0.310555 0.0673696 0.00409591 0.000561811 0.00138326 0.986983 0.99173 -2.97741e-06 -85.665 0.0930113 31188.1 302.191 0.983515 0.319147 0.732712 0.732708 9.99958 2.98226e-06 1.19289e-05 0.131262 0.982139 0.931603 -0.0132928 4.90541e-06 0.503389 -1.90707e-20 7.03761e-24 -1.90637e-20 0.00139549 0.997817 8.59545e-05 0.152602 2.85201 0.00139549 0.997823 0.717642 0.00105248 0.00188013 0.000859545 0.455578 0.00188013 0.438979 0.000128891 1.02 0.887832 0.534638 0.286263 1.71716e-07 3.06475e-09 2384.96 3116.39 -0.0553841 0.482144 0.277516 0.253308 -0.593371 -0.169519 0.496873 -0.267588 -0.229295 1.807 1 0 297.776 0 2.11168 1.805 0.000299833 0.853586 0.661726 0.377736 0.414001 2.11189 132.562 83.9131 18.7205 60.8627 0.00402561 0 -40 10
0.906 2.62455e-08 2.53901e-06 0.107021 0.107019 0.012038 1.19298e-05 0.00115409 0.133776 0.000657932 0.13443 0.882428 101.811 0.243286 0.751378 4.18855 0.0567137 0.0395146 0.960485 0.0197978 0.00430386 0.0190608 0.00413499 0.00520217 0.00593923 0.208087 0.237569 57.9956 -87.896 126.253 15.967 145.019 0.000141244 0.267153 192.866 0.310555 0.0673696 0.00409591 0.000561812 0.00138326 0.986983 0.99173 -2.97743e-06 -85.665 0.0930114 31188.1 302.197 0.983515 0.319147 0.732705 0.7327 9.99958 2.98227e-06 1.1929e-05 0.131264 0.982143 0.931604 -0.0132928 4.90544e-06 0.503398 -1.90716e-20 7.03799e-24 -1.90646e-20 0.00139549 0.997817 8.59546e-05 0.152602 2.85201 0.00139549 0.997823 0.71774 0.00105249 0.00188013 0.000859546 0.455578 0.00188013 0.438987 0.000128894 1.02 0.887833 0.534638 0.286264 1.71716e-07 3.06477e-09 2384.94 3116.36 -0.055383 0.482144 0.277516 0.253306 -0.593371 -0.16952 0.496875 -0.267585 -0.229299 1.808 1 0 297.777 0 2.11183 1.806 0.000299833 0.853574 0.661775 0.377597 0.414027 2.11205 132.571 83.9135 18.7205 60.8629 0.0040256 0 -40 10
0.907 2.62744e-08 2.53901e-06 0.107086 0.107084 0.012038 1.19429e-05 0.00115409 0.133858 0.000657934 0.134511 0.882497 101.811 0.243278 0.751481 4.18879 0.0567219 0.0395169 0.960483 0.0197976 0.00430408 0.0190605 0.00413518 0.00520244 0.0059395 0.208098 0.23758 57.9957 -87.896 126.253 15.967 145.019 0.000141243 0.267154 192.866 0.310554 0.0673695 0.00409592 0.000561812 0.00138326 0.986983 0.99173 -2.97744e-06 -85.665 0.0930115 31188 302.203 0.983515 0.319147 0.732698 0.732693 9.99958 2.98227e-06 1.1929e-05 0.131266 0.982148 0.931606 -0.0132928 4.90547e-06 0.503408 -1.90726e-20 7.03837e-24 -1.90655e-20 0.00139549 0.997817 8.59547e-05 0.152602 2.85201 0.00139549 0.997823 0.717838 0.00105251 0.00188013 0.000859547 0.455578 0.00188013 0.438995 0.000128897 1.02 0.887834 0.534637 0.286266 1.71717e-07 3.0648e-09 2384.92 3116.33 -0.0553819 0.482144 0.277515 0.253304 -0.593371 -0.16952 0.496878 -0.267583 -0.229304 1.809 1 0 297.779 0 2.11199 1.807 0.000299832 0.853562 0.661824 0.377458 0.414053 2.1122 132.579 83.9138 18.7205 60.8631 0.00402558 0 -40 10
0.908 2.63033e-08 2.53901e-06 0.107152 0.10715 0.0120379 1.1956e-05 0.00115409 0.133939 0.000657936 0.134593 0.882566 101.811 0.24327 0.751584 4.18903 0.0567301 0.0395192 0.960481 0.0197973 0.0043043 0.0190602 0.00413536 0.00520271 0.00593977 0.208109 0.237591 57.9958 -87.896 126.254 15.9669 145.019 0.000141242 0.267154 192.866 0.310554 0.0673694 0.00409592 0.000561813 0.00138326 0.986983 0.99173 -2.97746e-06 -85.665 0.0930116 31188 302.21 0.983515 0.319147 0.732691 0.732686 9.99958 2.98228e-06 1.1929e-05 0.131268 0.982152 0.931607 -0.0132928 4.9055e-06 0.503417 -1.90735e-20 7.03875e-24 -1.90664e-20 0.00139549 0.997817 8.59548e-05 0.152602 2.85201 0.00139549 0.997823 0.717936 0.00105253 0.00188013 0.000859548 0.455578 0.00188013 0.439002 0.000128901 1.02 0.887835 0.534637 0.286267 1.71717e-07 3.06482e-09 2384.91 3116.3 -0.0553808 0.482144 0.277515 0.253302 -0.593372 -0.16952 0.49688 -0.267581 -0.229308 1.81 1 0 297.78 0 2.11214 1.808 0.000299832 0.853551 0.661872 0.37732 0.414079 2.11236 132.587 83.9142 18.7205 60.8632 0.00402557 0 -40 10
0.909 2.63322e-08 2.53901e-06 0.107217 0.107215 0.0120379 1.19692e-05 0.00115409 0.134021 0.000657938 0.134674 0.882634 101.811 0.243262 0.751687 4.18928 0.0567383 0.0395215 0.960478 0.019797 0.00430453 0.01906 0.00413555 0.00520299 0.00594005 0.208119 0.237602 57.9958 -87.896 126.254 15.9669 145.019 0.00014124 0.267154 192.866 0.310553 0.0673694 0.00409592 0.000561814 0.00138327 0.986983 0.99173 -2.97747e-06 -85.6649 0.0930117 31188 302.216 0.983515 0.319147 0.732683 0.732679 9.99958 2.98228e-06 1.1929e-05 0.131271 0.982156 0.931608 -0.0132928 4.90553e-06 0.503426 -1.90744e-20 7.03913e-24 -1.90674e-20 0.00139549 0.997817 8.59548e-05 0.152602 2.85201 0.00139549 0.997823 0.718035 0.00105255 0.00188013 0.000859548 0.455577 0.00188013 0.43901 0.000128904 1.02 0.887836 0.534637 0.286269 1.71717e-07 3.06484e-09 2384.89 3116.27 -0.0553797 0.482144 0.277515 0.2533 -0.593372 -0.16952 0.496882 -0.267579 -0.229313 1.811 1 0 297.782 0 2.1123 1.809 0.000299831 0.85354 0.661921 0.377182 0.414105 2.11252 132.596 83.9145 18.7205 60.8634 0.00402555 0 -40 10
0.91 2.63612e-08 2.53901e-06 0.107282 0.10728 0.0120379 1.19823e-05 0.00115409 0.134102 0.00065794 0.134756 0.882703 101.81 0.243253 0.75179 4.18953 0.0567465 0.0395238 0.960476 0.0197967 0.00430475 0.0190597 0.00413574 0.00520326 0.00594032 0.20813 0.237613 57.9959 -87.896 126.254 15.9668 145.019 0.000141239 0.267154 192.866 0.310553 0.0673693 0.00409593 0.000561814 0.00138327 0.986983 0.99173 -2.97749e-06 -85.6649 0.0930118 31188 302.222 0.983515 0.319147 0.732676 0.732672 9.99958 2.98229e-06 1.1929e-05 0.131273 0.98216 0.93161 -0.0132928 4.90555e-06 0.503436 -1.90753e-20 7.03951e-24 -1.90683e-20 0.00139549 0.997817 8.59549e-05 0.152602 2.85201 0.00139549 0.997823 0.718133 0.00105257 0.00188014 0.000859549 0.455577 0.00188013 0.439018 0.000128907 1.02 0.887837 0.534637 0.28627 1.71718e-07 3.06486e-09 2384.87 3116.24 -0.0553787 0.482144 0.277515 0.253298 -0.593372 -0.16952 0.496885 -0.267577 -0.229317 1.812 1 0 297.783 0 2.11246 1.81 0.000299831 0.853528 0.66197 0.377044 0.414131 2.11267 132.604 83.9149 18.7206 60.8636 0.00402554 0 -40 10
0.911 2.63901e-08 2.53901e-06 0.107347 0.107345 0.0120379 1.19955e-05 0.00115409 0.134184 0.000657941 0.134837 0.882772 101.81 0.243245 0.751893 4.18977 0.0567548 0.0395262 0.960474 0.0197965 0.00430497 0.0190594 0.00413592 0.00520354 0.0059406 0.208141 0.237624 57.996 -87.896 126.254 15.9668 145.019 0.000141237 0.267154 192.865 0.310552 0.0673693 0.00409593 0.000561815 0.00138327 0.986983 0.99173 -2.9775e-06 -85.6649 0.0930118 31187.9 302.228 0.983515 0.319147 0.732669 0.732665 9.99958 2.98229e-06 1.19291e-05 0.131275 0.982165 0.931611 -0.0132928 4.90558e-06 0.503445 -1.90762e-20 7.0399e-24 -1.90692e-20 0.00139549 0.997817 8.5955e-05 0.152603 2.85201 0.00139549 0.997823 0.718231 0.00105259 0.00188014 0.00085955 0.455577 0.00188014 0.439026 0.00012891 1.02 0.887838 0.534636 0.286272 1.71718e-07 3.06489e-09 2384.85 3116.21 -0.0553777 0.482144 0.277514 0.253296 -0.593373 -0.16952 0.496887 -0.267575 -0.229321 1.813 1 0 297.785 0 2.11261 1.811 0.00029983 0.853517 0.662019 0.376906 0.414157 2.11283 132.612 83.9152 18.7206 60.8637 0.00402553 0 -40 10
0.912 2.6419e-08 2.53901e-06 0.107412 0.10741 0.0120379 1.20086e-05 0.0011541 0.134265 0.000657943 0.134918 0.882841 101.81 0.243237 0.751996 4.19002 0.056763 0.0395285 0.960472 0.0197962 0.0043052 0.0190591 0.00413611 0.00520381 0.00594087 0.208152 0.237635 57.996 -87.896 126.254 15.9668 145.019 0.000141236 0.267155 192.865 0.310552 0.0673692 0.00409593 0.000561816 0.00138327 0.986983 0.99173 -2.97752e-06 -85.6649 0.0930119 31187.9 302.234 0.983515 0.319147 0.732663 0.732658 9.99958 2.9823e-06 1.19291e-05 0.131277 0.982169 0.931612 -0.0132928 4.90561e-06 0.503454 -1.90772e-20 7.04028e-24 -1.90701e-20 0.00139549 0.997817 8.59551e-05 0.152603 2.85201 0.00139549 0.997823 0.718329 0.00105261 0.00188014 0.000859551 0.455577 0.00188014 0.439034 0.000128913 1.02 0.887839 0.534636 0.286273 1.71718e-07 3.06491e-09 2384.84 3116.18 -0.0553767 0.482144 0.277514 0.253294 -0.593373 -0.16952 0.496889 -0.267573 -0.229325 1.814 1 0 297.786 0 2.11277 1.812 0.00029983 0.853506 0.662068 0.376769 0.414183 2.11298 132.621 83.9156 18.7206 60.8639 0.00402551 0 -40 10
0.913 2.64479e-08 2.53901e-06 0.107477 0.107475 0.0120379 1.20218e-05 0.0011541 0.134346 0.000657945 0.134999 0.88291 101.81 0.243229 0.7521 4.19027 0.0567712 0.0395308 0.960469 0.0197959 0.00430542 0.0190589 0.0041363 0.00520409 0.00594115 0.208163 0.237646 57.9961 -87.896 126.254 15.9667 145.019 0.000141235 0.267155 192.865 0.310552 0.0673692 0.00409593 0.000561816 0.00138327 0.986983 0.99173 -2.97753e-06 -85.6649 0.093012 31187.9 302.24 0.983515 0.319147 0.732656 0.732651 9.99958 2.9823e-06 1.19291e-05 0.13128 0.982173 0.931614 -0.0132928 4.90564e-06 0.503464 -1.90781e-20 7.04066e-24 -1.9071e-20 0.00139549 0.997817 8.59552e-05 0.152603 2.85202 0.00139549 0.997823 0.718427 0.00105263 0.00188014 0.000859552 0.455576 0.00188014 0.439042 0.000128916 1.02 0.88784 0.534636 0.286275 1.71718e-07 3.06493e-09 2384.82 3116.15 -0.0553757 0.482144 0.277514 0.253293 -0.593373 -0.16952 0.496891 -0.267571 -0.229329 1.815 1 0 297.787 0 2.11292 1.813 0.000299829 0.853496 0.662117 0.376632 0.414209 2.11314 132.629 83.9159 18.7206 60.8641 0.0040255 0 -40 10
0.914 2.64769e-08 2.53901e-06 0.107542 0.10754 0.0120379 1.20349e-05 0.0011541 0.134427 0.000657947 0.135081 0.882978 101.809 0.243221 0.752203 4.19051 0.0567795 0.0395331 0.960467 0.0197956 0.00430564 0.0190586 0.00413649 0.00520436 0.00594142 0.208174 0.237657 57.9962 -87.896 126.254 15.9667 145.019 0.000141234 0.267155 192.865 0.310551 0.0673691 0.00409594 0.000561817 0.00138328 0.986983 0.99173 -2.97755e-06 -85.6649 0.0930121 31187.9 302.246 0.983515 0.319147 0.732649 0.732645 9.99958 2.98231e-06 1.19291e-05 0.131282 0.982177 0.931615 -0.0132928 4.90567e-06 0.503473 -1.9079e-20 7.04105e-24 -1.9072e-20 0.0013955 0.997817 8.59552e-05 0.152603 2.85202 0.0013955 0.997823 0.718525 0.00105265 0.00188014 0.000859552 0.455576 0.00188014 0.43905 0.00012892 1.02 0.887841 0.534635 0.286276 1.71719e-07 3.06496e-09 2384.8 3116.12 -0.0553747 0.482145 0.277513 0.253291 -0.593374 -0.16952 0.496893 -0.267569 -0.229334 1.816 1 0 297.789 0 2.11308 1.814 0.000299829 0.853485 0.662166 0.376495 0.414235 2.1133 132.638 83.9162 18.7206 60.8642 0.00402548 0 -40 10
0.915 2.65058e-08 2.53901e-06 0.107607 0.107605 0.0120379 1.20481e-05 0.0011541 0.134508 0.000657949 0.135162 0.883047 101.809 0.243212 0.752306 4.19076 0.0567877 0.0395355 0.960465 0.0197954 0.00430587 0.0190583 0.00413668 0.00520464 0.0059417 0.208185 0.237668 57.9962 -87.896 126.254 15.9667 145.019 0.000141232 0.267155 192.865 0.310551 0.0673691 0.00409594 0.000561818 0.00138328 0.986982 0.99173 -2.97756e-06 -85.6649 0.0930122 31187.9 302.252 0.983515 0.319147 0.732642 0.732638 9.99958 2.98231e-06 1.19291e-05 0.131284 0.982181 0.931616 -0.0132928 4.9057e-06 0.503483 -1.90799e-20 7.04143e-24 -1.90729e-20 0.0013955 0.997817 8.59553e-05 0.152603 2.85202 0.0013955 0.997823 0.718623 0.00105267 0.00188014 0.000859553 0.455576 0.00188014 0.439058 0.000128923 1.02 0.887843 0.534635 0.286278 1.71719e-07 3.06498e-09 2384.79 3116.09 -0.0553738 0.482145 0.277513 0.253289 -0.593374 -0.16952 0.496895 -0.267567 -0.229338 1.817 1 0 297.79 0 2.11324 1.815 0.000299828 0.853474 0.662215 0.376359 0.414261 2.11345 132.646 83.9166 18.7207 60.8644 0.00402547 0 -40 10
0.916 2.65347e-08 2.53901e-06 0.107672 0.10767 0.0120378 1.20612e-05 0.0011541 0.134589 0.000657951 0.135243 0.883116 101.809 0.243204 0.75241 4.19101 0.056796 0.0395378 0.960462 0.0197951 0.00430609 0.019058 0.00413686 0.00520491 0.00594197 0.208197 0.237679 57.9963 -87.896 126.255 15.9666 145.019 0.000141231 0.267155 192.865 0.31055 0.067369 0.00409594 0.000561818 0.00138328 0.986982 0.99173 -2.97758e-06 -85.6649 0.0930123 31187.8 302.258 0.983515 0.319147 0.732636 0.732631 9.99958 2.98232e-06 1.19292e-05 0.131287 0.982186 0.931618 -0.0132928 4.90573e-06 0.503492 -1.90808e-20 7.04181e-24 -1.90738e-20 0.0013955 0.997817 8.59554e-05 0.152603 2.85202 0.0013955 0.997823 0.71872 0.00105269 0.00188014 0.000859554 0.455576 0.00188014 0.439065 0.000128926 1.02 0.887844 0.534635 0.28628 1.71719e-07 3.065e-09 2384.77 3116.06 -0.0553728 0.482145 0.277513 0.253287 -0.593374 -0.16952 0.496897 -0.267564 -0.229342 1.818 1 0 297.791 0 2.11339 1.816 0.000299828 0.853464 0.662263 0.376223 0.414287 2.11361 132.654 83.9169 18.7207 60.8645 0.00402546 0 -40 10
0.917 2.65636e-08 2.53901e-06 0.107736 0.107734 0.0120378 1.20744e-05 0.0011541 0.13467 0.000657953 0.135324 0.883185 101.809 0.243196 0.752513 4.19126 0.0568042 0.0395402 0.96046 0.0197948 0.00430632 0.0190577 0.00413705 0.00520519 0.00594225 0.208208 0.23769 57.9963 -87.896 126.255 15.9666 145.019 0.00014123 0.267156 192.864 0.31055 0.067369 0.00409595 0.000561819 0.00138328 0.986982 0.99173 -2.97759e-06 -85.6649 0.0930124 31187.8 302.264 0.983514 0.319147 0.732629 0.732625 9.99958 2.98232e-06 1.19292e-05 0.131289 0.98219 0.931619 -0.0132928 4.90576e-06 0.503502 -1.90818e-20 7.0422e-24 -1.90747e-20 0.0013955 0.997817 8.59555e-05 0.152603 2.85202 0.0013955 0.997823 0.718818 0.0010527 0.00188015 0.000859555 0.455576 0.00188014 0.439073 0.000128929 1.02 0.887845 0.534634 0.286281 1.71719e-07 3.06502e-09 2384.75 3116.03 -0.0553719 0.482145 0.277513 0.253285 -0.593375 -0.16952 0.496898 -0.267562 -0.229345 1.819 1 0 297.793 0 2.11355 1.817 0.000299828 0.853454 0.662312 0.376087 0.414313 2.11376 132.663 83.9172 18.7207 60.8647 0.00402544 0 -40 10
0.918 2.65925e-08 2.53901e-06 0.107801 0.107799 0.0120378 1.20875e-05 0.0011541 0.134751 0.000657955 0.135405 0.883254 101.808 0.243188 0.752617 4.19151 0.0568125 0.0395425 0.960457 0.0197945 0.00430654 0.0190575 0.00413724 0.00520547 0.00594253 0.208219 0.237701 57.9964 -87.896 126.255 15.9665 145.019 0.000141228 0.267156 192.864 0.310549 0.0673689 0.00409595 0.00056182 0.00138328 0.986982 0.99173 -2.97761e-06 -85.6649 0.0930124 31187.8 302.27 0.983514 0.319147 0.732622 0.732618 9.99958 2.98233e-06 1.19292e-05 0.131291 0.982194 0.93162 -0.0132928 4.90579e-06 0.503511 -1.90827e-20 7.04258e-24 -1.90756e-20 0.0013955 0.997817 8.59555e-05 0.152604 2.85202 0.0013955 0.997823 0.718916 0.00105272 0.00188015 0.000859555 0.455575 0.00188015 0.439081 0.000128932 1.02 0.887846 0.534634 0.286283 1.7172e-07 3.06505e-09 2384.74 3116 -0.0553711 0.482145 0.277512 0.253284 -0.593375 -0.16952 0.4969 -0.26756 -0.229349 1.82 1 0 297.794 0 2.1137 1.818 0.000299827 0.853443 0.662361 0.375952 0.414339 2.11392 132.671 83.9176 18.7207 60.8649 0.00402543 0 -40 10
0.919 2.66215e-08 2.53901e-06 0.107866 0.107864 0.0120378 1.21007e-05 0.0011541 0.134832 0.000657957 0.135485 0.883324 101.808 0.243179 0.75272 4.19176 0.0568208 0.0395449 0.960455 0.0197943 0.00430677 0.0190572 0.00413743 0.00520575 0.00594281 0.20823 0.237712 57.9965 -87.896 126.255 15.9665 145.019 0.000141227 0.267156 192.864 0.310549 0.0673689 0.00409595 0.00056182 0.00138329 0.986982 0.99173 -2.97762e-06 -85.6649 0.0930125 31187.8 302.276 0.983514 0.319147 0.732616 0.732612 9.99958 2.98233e-06 1.19292e-05 0.131294 0.982198 0.931621 -0.0132928 4.90582e-06 0.503521 -1.90836e-20 7.04297e-24 -1.90766e-20 0.0013955 0.997817 8.59556e-05 0.152604 2.85202 0.0013955 0.997823 0.719014 0.00105274 0.00188015 0.000859556 0.455575 0.00188015 0.439089 0.000128935 1.02 0.887847 0.534634 0.286284 1.7172e-07 3.06507e-09 2384.72 3115.97 -0.0553702 0.482145 0.277512 0.253282 -0.593375 -0.16952 0.496902 -0.267558 -0.229353 1.821 1 0 297.795 0 2.11386 1.819 0.000299827 0.853433 0.66241 0.375816 0.414365 2.11407 132.679 83.9179 18.7207 60.865 0.00402542 0 -40 10
0.92 2.66504e-08 2.53901e-06 0.10793 0.107928 0.0120378 1.21138e-05 0.0011541 0.134913 0.000657959 0.135566 0.883393 101.808 0.243171 0.752824 4.19201 0.056829 0.0395472 0.960453 0.019794 0.004307 0.0190569 0.00413762 0.00520602 0.00594308 0.208241 0.237723 57.9965 -87.896 126.255 15.9665 145.019 0.000141226 0.267156 192.864 0.310549 0.0673688 0.00409596 0.000561821 0.00138329 0.986982 0.99173 -2.97764e-06 -85.6648 0.0930126 31187.7 302.282 0.983514 0.319147 0.73261 0.732605 9.99958 2.98234e-06 1.19292e-05 0.131296 0.982202 0.931623 -0.0132928 4.90585e-06 0.50353 -1.90845e-20 7.04335e-24 -1.90775e-20 0.0013955 0.997817 8.59557e-05 0.152604 2.85202 0.0013955 0.997823 0.719112 0.00105276 0.00188015 0.000859557 0.455575 0.00188015 0.439097 0.000128939 1.02 0.887848 0.534633 0.286286 1.7172e-07 3.06509e-09 2384.7 3115.95 -0.0553694 0.482145 0.277512 0.25328 -0.593376 -0.16952 0.496903 -0.267556 -0.229357 1.822 1 0 297.796 0 2.11402 1.82 0.000299826 0.853423 0.662459 0.375681 0.414391 2.11423 132.688 83.9182 18.7208 60.8652 0.0040254 0 -40 10
0.921 2.66793e-08 2.53901e-06 0.107995 0.107993 0.0120378 1.2127e-05 0.0011541 0.134994 0.000657961 0.135647 0.883462 101.808 0.243163 0.752928 4.19226 0.0568373 0.0395496 0.96045 0.0197937 0.00430722 0.0190566 0.00413781 0.0052063 0.00594336 0.208252 0.237735 57.9966 -87.896 126.255 15.9664 145.019 0.000141225 0.267156 192.864 0.310548 0.0673688 0.00409596 0.000561822 0.00138329 0.986982 0.99173 -2.97765e-06 -85.6648 0.0930127 31187.7 302.289 0.983514 0.319147 0.732603 0.732599 9.99958 2.98234e-06 1.19293e-05 0.131298 0.982206 0.931624 -0.0132928 4.90588e-06 0.50354 -1.90855e-20 7.04373e-24 -1.90784e-20 0.0013955 0.997817 8.59558e-05 0.152604 2.85202 0.0013955 0.997823 0.719209 0.00105278 0.00188015 0.000859558 0.455575 0.00188015 0.439105 0.000128942 1.02 0.887849 0.534633 0.286287 1.7172e-07 3.06511e-09 2384.69 3115.92 -0.0553685 0.482145 0.277511 0.253278 -0.593376 -0.16952 0.496905 -0.267554 -0.22936 1.823 1 0 297.797 0 2.11417 1.821 0.000299826 0.853414 0.662507 0.375547 0.414417 2.11439 132.696 83.9185 18.7208 60.8653 0.00402539 0 -40 10
0.922 2.67082e-08 2.53902e-06 0.108059 0.108057 0.0120378 1.21401e-05 0.0011541 0.135074 0.000657963 0.135728 0.883531 101.807 0.243154 0.753032 4.19251 0.0568456 0.039552 0.960448 0.0197934 0.00430745 0.0190564 0.004138 0.00520658 0.00594364 0.208263 0.237746 57.9967 -87.896 126.255 15.9664 145.019 0.000141224 0.267156 192.864 0.310548 0.0673687 0.00409596 0.000561822 0.00138329 0.986982 0.99173 -2.97767e-06 -85.6648 0.0930128 31187.7 302.295 0.983514 0.319147 0.732597 0.732593 9.99958 2.98235e-06 1.19293e-05 0.1313 0.98221 0.931625 -0.0132928 4.90591e-06 0.503549 -1.90864e-20 7.04412e-24 -1.90793e-20 0.00139551 0.997817 8.59559e-05 0.152604 2.85202 0.00139551 0.997823 0.719307 0.0010528 0.00188015 0.000859559 0.455574 0.00188015 0.439113 0.000128945 1.02 0.88785 0.534633 0.286289 1.71721e-07 3.06514e-09 2384.67 3115.89 -0.0553677 0.482145 0.277511 0.253277 -0.593376 -0.169521 0.496907 -0.267552 -0.229364 1.824 1 0 297.799 0 2.11433 1.822 0.000299825 0.853404 0.662556 0.375412 0.414443 2.11454 132.704 83.9188 18.7208 60.8655 0.00402538 0 -40 10
0.923 2.67372e-08 2.53902e-06 0.108124 0.108122 0.0120377 1.21533e-05 0.0011541 0.135155 0.000657965 0.135808 0.8836 101.807 0.243146 0.753136 4.19276 0.0568539 0.0395543 0.960446 0.0197931 0.00430768 0.0190561 0.00413819 0.00520686 0.00594392 0.208274 0.237757 57.9967 -87.896 126.255 15.9664 145.019 0.000141222 0.267157 192.863 0.310547 0.0673687 0.00409596 0.000561823 0.0013833 0.986982 0.99173 -2.97768e-06 -85.6648 0.0930129 31187.7 302.301 0.983514 0.319147 0.732591 0.732586 9.99958 2.98235e-06 1.19293e-05 0.131303 0.982214 0.931626 -0.0132928 4.90594e-06 0.503559 -1.90873e-20 7.04451e-24 -1.90803e-20 0.00139551 0.997817 8.59559e-05 0.152604 2.85202 0.00139551 0.997823 0.719405 0.00105282 0.00188015 0.000859559 0.455574 0.00188015 0.43912 0.000128948 1.02 0.887851 0.534633 0.28629 1.71721e-07 3.06516e-09 2384.65 3115.86 -0.0553669 0.482145 0.277511 0.253275 -0.593377 -0.169521 0.496908 -0.26755 -0.229368 1.825 1 0 297.8 0 2.11448 1.823 0.000299825 0.853394 0.662605 0.375278 0.414469 2.1147 132.713 83.9191 18.7208 60.8656 0.00402537 0 -40 10
0.924 2.67661e-08 2.53902e-06 0.108188 0.108186 0.0120377 1.21664e-05 0.0011541 0.135235 0.000657967 0.135889 0.88367 101.807 0.243138 0.753239 4.19301 0.0568622 0.0395567 0.960443 0.0197929 0.0043079 0.0190558 0.00413838 0.00520714 0.0059442 0.208286 0.237768 57.9968 -87.896 126.255 15.9663 145.019 0.000141221 0.267157 192.863 0.310547 0.0673686 0.00409597 0.000561824 0.0013833 0.986982 0.99173 -2.9777e-06 -85.6648 0.093013 31187.7 302.307 0.983514 0.319147 0.732585 0.73258 9.99958 2.98236e-06 1.19293e-05 0.131305 0.982219 0.931627 -0.0132928 4.90597e-06 0.503569 -1.90882e-20 7.04489e-24 -1.90812e-20 0.00139551 0.997817 8.5956e-05 0.152605 2.85203 0.00139551 0.997823 0.719502 0.00105284 0.00188016 0.00085956 0.455574 0.00188015 0.439128 0.000128951 1.02 0.887852 0.534632 0.286292 1.71721e-07 3.06518e-09 2384.64 3115.84 -0.0553662 0.482145 0.277511 0.253273 -0.593377 -0.169521 0.496909 -0.267548 -0.229371 1.826 1 0 297.801 0 2.11464 1.824 0.000299824 0.853385 0.662654 0.375144 0.414495 2.11485 132.721 83.9194 18.7208 60.8658 0.00402535 0 -40 10
0.925 2.6795e-08 2.53902e-06 0.108253 0.108251 0.0120377 1.21796e-05 0.0011541 0.135316 0.000657968 0.135969 0.883739 101.807 0.24313 0.753343 4.19326 0.0568705 0.0395591 0.960441 0.0197926 0.00430813 0.0190555 0.00413858 0.00520742 0.00594448 0.208297 0.237779 57.9969 -87.896 126.256 15.9663 145.019 0.00014122 0.267157 192.863 0.310547 0.0673686 0.00409597 0.000561824 0.0013833 0.986982 0.99173 -2.97771e-06 -85.6648 0.093013 31187.6 302.313 0.983514 0.319147 0.732578 0.732574 9.99958 2.98236e-06 1.19293e-05 0.131307 0.982223 0.931629 -0.0132928 4.906e-06 0.503578 -1.90892e-20 7.04528e-24 -1.90821e-20 0.00139551 0.997817 8.59561e-05 0.152605 2.85203 0.00139551 0.997823 0.7196 0.00105286 0.00188016 0.000859561 0.455574 0.00188016 0.439136 0.000128954 1.02 0.887853 0.534632 0.286293 1.71722e-07 3.06521e-09 2384.62 3115.81 -0.0553654 0.482145 0.27751 0.253272 -0.593377 -0.169521 0.496911 -0.267546 -0.229374 1.827 1 0 297.802 0 2.11479 1.825 0.000299824 0.853375 0.662702 0.375011 0.41452 2.11501 132.729 83.9197 18.7208 60.8659 0.00402534 0 -40 10
0.926 2.68239e-08 2.53902e-06 0.108317 0.108315 0.0120377 1.21927e-05 0.0011541 0.135396 0.00065797 0.136049 0.883808 101.806 0.243121 0.753448 4.19352 0.0568788 0.0395615 0.960439 0.0197923 0.00430836 0.0190552 0.00413877 0.0052077 0.00594476 0.208308 0.23779 57.9969 -87.896 126.256 15.9662 145.019 0.000141219 0.267157 192.863 0.310546 0.0673685 0.00409597 0.000561825 0.0013833 0.986982 0.99173 -2.97772e-06 -85.6648 0.0930131 31187.6 302.319 0.983514 0.319147 0.732572 0.732568 9.99958 2.98237e-06 1.19294e-05 0.13131 0.982227 0.93163 -0.0132928 4.90603e-06 0.503588 -1.90901e-20 7.04566e-24 -1.90831e-20 0.00139551 0.997817 8.59562e-05 0.152605 2.85203 0.00139551 0.997823 0.719697 0.00105288 0.00188016 0.000859562 0.455574 0.00188016 0.439144 0.000128957 1.02 0.887855 0.534632 0.286295 1.71722e-07 3.06523e-09 2384.6 3115.78 -0.0553647 0.482145 0.27751 0.25327 -0.593377 -0.169521 0.496912 -0.267543 -0.229378 1.828 1 0 297.803 0 2.11495 1.826 0.000299823 0.853366 0.662751 0.374878 0.414546 2.11516 132.738 83.92 18.7209 60.8661 0.00402533 0 -40 10
0.927 2.68529e-08 2.53902e-06 0.108381 0.108379 0.0120377 1.22058e-05 0.0011541 0.135476 0.000657972 0.13613 0.883878 101.806 0.243113 0.753552 4.19377 0.0568871 0.0395639 0.960436 0.019792 0.00430859 0.019055 0.00413896 0.00520798 0.00594504 0.208319 0.237802 57.997 -87.896 126.256 15.9662 145.019 0.000141218 0.267157 192.863 0.310546 0.0673685 0.00409598 0.000561826 0.0013833 0.986982 0.99173 -2.97774e-06 -85.6648 0.0930132 31187.6 302.326 0.983514 0.319147 0.732566 0.732562 9.99958 2.98237e-06 1.19294e-05 0.131312 0.982231 0.931631 -0.0132928 4.90606e-06 0.503597 -1.9091e-20 7.04605e-24 -1.9084e-20 0.00139551 0.997817 8.59563e-05 0.152605 2.85203 0.00139551 0.997823 0.719795 0.0010529 0.00188016 0.000859563 0.455573 0.00188016 0.439152 0.000128961 1.02 0.887856 0.534631 0.286296 1.71722e-07 3.06525e-09 2384.59 3115.76 -0.055364 0.482146 0.27751 0.253269 -0.593378 -0.169521 0.496913 -0.267541 -0.229381 1.829 1 0 297.804 0 2.1151 1.827 0.000299823 0.853357 0.6628 0.374745 0.414572 2.11532 132.746 83.9203 18.7209 60.8662 0.00402532 0 -40 10
0.928 2.68818e-08 2.53902e-06 0.108445 0.108443 0.0120377 1.2219e-05 0.0011541 0.135557 0.000657974 0.13621 0.883947 101.806 0.243105 0.753656 4.19402 0.0568954 0.0395663 0.960434 0.0197917 0.00430882 0.0190547 0.00413915 0.00520826 0.00594532 0.20833 0.237813 57.997 -87.896 126.256 15.9662 145.019 0.000141216 0.267158 192.863 0.310545 0.0673684 0.00409598 0.000561826 0.00138331 0.986982 0.99173 -2.97775e-06 -85.6648 0.0930133 31187.6 302.332 0.983514 0.319147 0.732561 0.732556 9.99958 2.98238e-06 1.19294e-05 0.131314 0.982235 0.931632 -0.0132928 4.90608e-06 0.503607 -1.9092e-20 7.04644e-24 -1.90849e-20 0.00139551 0.997817 8.59563e-05 0.152605 2.85203 0.00139551 0.997823 0.719892 0.00105292 0.00188016 0.000859563 0.455573 0.00188016 0.43916 0.000128964 1.02 0.887857 0.534631 0.286298 1.71722e-07 3.06527e-09 2384.57 3115.73 -0.0553633 0.482146 0.277509 0.253267 -0.593378 -0.169521 0.496914 -0.267539 -0.229384 1.83 1 0 297.805 0 2.11526 1.828 0.000299822 0.853348 0.662848 0.374612 0.414598 2.11547 132.754 83.9206 18.7209 60.8663 0.0040253 0 -40 10
0.929 2.69107e-08 2.53902e-06 0.108509 0.108508 0.0120377 1.22321e-05 0.0011541 0.135637 0.000657976 0.13629 0.884017 101.806 0.243096 0.75376 4.19428 0.0569037 0.0395687 0.960431 0.0197915 0.00430904 0.0190544 0.00413934 0.00520854 0.00594561 0.208342 0.237824 57.9971 -87.896 126.256 15.9661 145.019 0.000141215 0.267158 192.862 0.310545 0.0673684 0.00409598 0.000561827 0.00138331 0.986982 0.99173 -2.97777e-06 -85.6648 0.0930134 31187.5 302.338 0.983514 0.319147 0.732555 0.73255 9.99958 2.98238e-06 1.19294e-05 0.131317 0.982239 0.931633 -0.0132928 4.90611e-06 0.503617 -1.90929e-20 7.04682e-24 -1.90858e-20 0.00139551 0.997817 8.59564e-05 0.152605 2.85203 0.00139551 0.997823 0.71999 0.00105293 0.00188016 0.000859564 0.455573 0.00188016 0.439167 0.000128967 1.02 0.887858 0.534631 0.286299 1.71723e-07 3.0653e-09 2384.55 3115.71 -0.0553626 0.482146 0.277509 0.253265 -0.593378 -0.169521 0.496915 -0.267537 -0.229388 1.831 1 0 297.806 0 2.11541 1.829 0.000299822 0.853339 0.662897 0.37448 0.414624 2.11563 132.763 83.9209 18.7209 60.8665 0.00402529 0 -40 10
0.93 2.69396e-08 2.53902e-06 0.108574 0.108572 0.0120377 1.22453e-05 0.0011541 0.135717 0.000657978 0.13637 0.884086 101.805 0.243088 0.753864 4.19453 0.056912 0.0395711 0.960429 0.0197912 0.00430927 0.0190541 0.00413954 0.00520882 0.00594589 0.208353 0.237836 57.9972 -87.8961 126.256 15.9661 145.019 0.000141214 0.267158 192.862 0.310544 0.0673683 0.00409599 0.000561828 0.00138331 0.986982 0.99173 -2.97778e-06 -85.6648 0.0930135 31187.5 302.344 0.983514 0.319147 0.732549 0.732545 9.99958 2.98239e-06 1.19294e-05 0.131319 0.982243 0.931634 -0.0132928 4.90614e-06 0.503626 -1.90938e-20 7.04721e-24 -1.90868e-20 0.00139551 0.997817 8.59565e-05 0.152605 2.85203 0.00139551 0.997823 0.720087 0.00105295 0.00188016 0.000859565 0.455573 0.00188016 0.439175 0.00012897 1.02 0.887859 0.53463 0.286301 1.71723e-07 3.06532e-09 2384.54 3115.68 -0.055362 0.482146 0.277509 0.253264 -0.593378 -0.169521 0.496916 -0.267535 -0.229391 1.832 1 0 297.807 0 2.11557 1.83 0.000299821 0.85333 0.662945 0.374347 0.41465 2.11578 132.771 83.9212 18.7209 60.8666 0.00402528 0 -40 10
0.931 2.69686e-08 2.53902e-06 0.108638 0.108636 0.0120376 1.22584e-05 0.0011541 0.135797 0.00065798 0.13645 0.884156 101.805 0.24308 0.753969 4.19479 0.0569204 0.0395735 0.960427 0.0197909 0.0043095 0.0190538 0.00413973 0.00520911 0.00594617 0.208364 0.237847 57.9972 -87.8961 126.256 15.9661 145.019 0.000141213 0.267158 192.862 0.310544 0.0673683 0.00409599 0.000561828 0.00138331 0.986982 0.99173 -2.9778e-06 -85.6647 0.0930136 31187.5 302.35 0.983514 0.319147 0.732543 0.732539 9.99958 2.98239e-06 1.19295e-05 0.131322 0.982247 0.931636 -0.0132928 4.90617e-06 0.503636 -1.90948e-20 7.0476e-24 -1.90877e-20 0.00139552 0.997817 8.59566e-05 0.152606 2.85203 0.00139552 0.997822 0.720184 0.00105297 0.00188017 0.000859566 0.455572 0.00188017 0.439183 0.000128973 1.02 0.88786 0.53463 0.286302 1.71723e-07 3.06534e-09 2384.52 3115.66 -0.0553614 0.482146 0.277509 0.253262 -0.593379 -0.169521 0.496917 -0.267533 -0.229394 1.833 1 0 297.808 0 2.11573 1.831 0.000299821 0.853322 0.662994 0.374216 0.414676 2.11594 132.779 83.9215 18.7209 60.8667 0.00402527 0 -40 10
0.932 2.69975e-08 2.53902e-06 0.108702 0.1087 0.0120376 1.22716e-05 0.0011541 0.135877 0.000657982 0.13653 0.884226 101.805 0.243071 0.754073 4.19504 0.0569287 0.0395759 0.960424 0.0197906 0.00430973 0.0190535 0.00413992 0.00520939 0.00594645 0.208376 0.237858 57.9973 -87.8961 126.256 15.966 145.019 0.000141212 0.267158 192.862 0.310544 0.0673682 0.00409599 0.000561829 0.00138331 0.986982 0.99173 -2.97781e-06 -85.6647 0.0930137 31187.5 302.357 0.983514 0.319147 0.732537 0.732533 9.99958 2.98239e-06 1.19295e-05 0.131324 0.982251 0.931637 -0.0132928 4.9062e-06 0.503646 -1.90957e-20 7.04798e-24 -1.90886e-20 0.00139552 0.997817 8.59567e-05 0.152606 2.85203 0.00139552 0.997822 0.720282 0.00105299 0.00188017 0.000859567 0.455572 0.00188017 0.439191 0.000128976 1.02 0.887861 0.53463 0.286304 1.71723e-07 3.06536e-09 2384.5 3115.63 -0.0553607 0.482146 0.277508 0.253261 -0.593379 -0.169521 0.496918 -0.267531 -0.229397 1.834 1 0 297.809 0 2.11588 1.832 0.00029982 0.853313 0.663043 0.374084 0.414701 2.11609 132.787 83.9218 18.721 60.8669 0.00402526 0 -40 10
0.933 2.70264e-08 2.53902e-06 0.108765 0.108764 0.0120376 1.22847e-05 0.0011541 0.135957 0.000657984 0.13661 0.884295 101.805 0.243063 0.754178 4.1953 0.056937 0.0395783 0.960422 0.0197903 0.00430996 0.0190533 0.00414012 0.00520967 0.00594674 0.208387 0.237869 57.9974 -87.8961 126.256 15.966 145.019 0.000141211 0.267159 192.862 0.310543 0.0673681 0.00409599 0.00056183 0.00138332 0.986982 0.99173 -2.97783e-06 -85.6647 0.0930137 31187.5 302.363 0.983514 0.319147 0.732532 0.732527 9.99958 2.9824e-06 1.19295e-05 0.131326 0.982255 0.931638 -0.0132928 4.90623e-06 0.503655 -1.90966e-20 7.04837e-24 -1.90896e-20 0.00139552 0.997817 8.59567e-05 0.152606 2.85203 0.00139552 0.997822 0.720379 0.00105301 0.00188017 0.000859567 0.455572 0.00188017 0.439199 0.00012898 1.02 0.887862 0.534629 0.286305 1.71724e-07 3.06539e-09 2384.49 3115.61 -0.0553602 0.482146 0.277508 0.253259 -0.593379 -0.169521 0.496919 -0.267529 -0.2294 1.835 1 0 297.81 0 2.11604 1.833 0.00029982 0.853305 0.663091 0.373953 0.414727 2.11625 132.796 83.922 18.721 60.867 0.00402525 0 -40 10
0.934 2.70553e-08 2.53902e-06 0.108829 0.108827 0.0120376 1.22979e-05 0.0011541 0.136037 0.000657985 0.13669 0.884365 101.804 0.243055 0.754282 4.19555 0.0569454 0.0395807 0.960419 0.01979 0.00431019 0.019053 0.00414031 0.00520996 0.00594702 0.208398 0.237881 57.9974 -87.8961 126.257 15.9659 145.019 0.00014121 0.267159 192.862 0.310543 0.0673681 0.004096 0.00056183 0.00138332 0.986982 0.99173 -2.97784e-06 -85.6647 0.0930138 31187.4 302.369 0.983514 0.319147 0.732526 0.732522 9.99958 2.9824e-06 1.19295e-05 0.131329 0.982259 0.931639 -0.0132928 4.90626e-06 0.503665 -1.90976e-20 7.04876e-24 -1.90905e-20 0.00139552 0.997817 8.59568e-05 0.152606 2.85203 0.00139552 0.997822 0.720476 0.00105303 0.00188017 0.000859568 0.455572 0.00188017 0.439206 0.000128983 1.02 0.887863 0.534629 0.286307 1.71724e-07 3.06541e-09 2384.47 3115.58 -0.0553596 0.482146 0.277508 0.253258 -0.59338 -0.169521 0.49692 -0.267527 -0.229403 1.836 1 0 297.811 0 2.11619 1.834 0.000299819 0.853297 0.66314 0.373822 0.414753 2.1164 132.804 83.9223 18.721 60.8672 0.00402523 0 -40 10
0.935 2.70842e-08 2.53902e-06 0.108893 0.108891 0.0120376 1.2311e-05 0.0011541 0.136116 0.000657987 0.13677 0.884435 101.804 0.243046 0.754387 4.19581 0.0569537 0.0395831 0.960417 0.0197898 0.00431042 0.0190527 0.0041405 0.00521024 0.00594731 0.20841 0.237892 57.9975 -87.8961 126.257 15.9659 145.019 0.000141209 0.267159 192.861 0.310542 0.067368 0.004096 0.000561831 0.00138332 0.986982 0.991729 -2.97786e-06 -85.6647 0.0930139 31187.4 302.375 0.983514 0.319147 0.732521 0.732516 9.99958 2.98241e-06 1.19295e-05 0.131331 0.982262 0.93164 -0.0132928 4.90629e-06 0.503675 -1.90985e-20 7.04915e-24 -1.90915e-20 0.00139552 0.997817 8.59569e-05 0.152606 2.85204 0.00139552 0.997822 0.720574 0.00105305 0.00188017 0.000859569 0.455572 0.00188017 0.439214 0.000128986 1.02 0.887864 0.534629 0.286308 1.71724e-07 3.06543e-09 2384.45 3115.56 -0.055359 0.482146 0.277507 0.253256 -0.59338 -0.169521 0.496921 -0.267524 -0.229405 1.837 1 0 297.812 0 2.11635 1.835 0.000299819 0.853288 0.663188 0.373691 0.414779 2.11656 132.812 83.9226 18.721 60.8673 0.00402522 0 -40 10
0.936 2.71132e-08 2.53902e-06 0.108957 0.108955 0.0120376 1.23242e-05 0.0011541 0.136196 0.000657989 0.13685 0.884505 101.804 0.243038 0.754492 4.19607 0.0569621 0.0395855 0.960414 0.0197895 0.00431066 0.0190524 0.0041407 0.00521052 0.00594759 0.208421 0.237904 57.9976 -87.8961 126.257 15.9659 145.019 0.000141208 0.267159 192.861 0.310542 0.067368 0.004096 0.000561832 0.00138332 0.986982 0.991729 -2.97787e-06 -85.6647 0.093014 31187.4 302.382 0.983514 0.319147 0.732515 0.732511 9.99958 2.98241e-06 1.19296e-05 0.131333 0.982266 0.931641 -0.0132928 4.90632e-06 0.503685 -1.90994e-20 7.04954e-24 -1.90924e-20 0.00139552 0.997817 8.5957e-05 0.152606 2.85204 0.00139552 0.997822 0.720671 0.00105307 0.00188017 0.00085957 0.455571 0.00188017 0.439222 0.000128989 1.02 0.887865 0.534629 0.28631 1.71724e-07 3.06545e-09 2384.44 3115.53 -0.0553585 0.482146 0.277507 0.253255 -0.59338 -0.169521 0.496921 -0.267522 -0.229408 1.838 1 0 297.813 0 2.1165 1.836 0.000299818 0.85328 0.663237 0.373561 0.414805 2.11671 132.821 83.9229 18.721 60.8674 0.00402521 0 -40 10
0.937 2.71421e-08 2.53902e-06 0.109021 0.109019 0.0120376 1.23373e-05 0.0011541 0.136276 0.000657991 0.136929 0.884574 101.804 0.24303 0.754596 4.19632 0.0569704 0.039588 0.960412 0.0197892 0.00431089 0.0190521 0.00414089 0.00521081 0.00594788 0.208432 0.237915 57.9976 -87.8961 126.257 15.9658 145.019 0.000141207 0.267159 192.861 0.310541 0.0673679 0.00409601 0.000561832 0.00138333 0.986982 0.991729 -2.97789e-06 -85.6647 0.0930141 31187.4 302.388 0.983514 0.319147 0.73251 0.732506 9.99958 2.98242e-06 1.19296e-05 0.131336 0.98227 0.931642 -0.0132928 4.90635e-06 0.503694 -1.91004e-20 7.04993e-24 -1.90933e-20 0.00139552 0.997817 8.59571e-05 0.152607 2.85204 0.00139552 0.997822 0.720768 0.00105309 0.00188018 0.000859571 0.455571 0.00188017 0.43923 0.000128992 1.02 0.887867 0.534628 0.286311 1.71725e-07 3.06548e-09 2384.42 3115.51 -0.055358 0.482146 0.277507 0.253253 -0.59338 -0.169522 0.496922 -0.26752 -0.229411 1.839 1 0 297.814 0 2.11666 1.837 0.000299818 0.853272 0.663285 0.37343 0.41483 2.11687 132.829 83.9231 18.721 60.8675 0.0040252 0 -40 10
0.938 2.7171e-08 2.53903e-06 0.109084 0.109083 0.0120375 1.23505e-05 0.0011541 0.136355 0.000657993 0.137009 0.884644 101.803 0.243021 0.754701 4.19658 0.0569788 0.0395904 0.96041 0.0197889 0.00431112 0.0190518 0.00414109 0.00521109 0.00594816 0.208444 0.237926 57.9977 -87.8961 126.257 15.9658 145.019 0.000141206 0.267159 192.861 0.310541 0.0673679 0.00409601 0.000561833 0.00138333 0.986982 0.991729 -2.9779e-06 -85.6647 0.0930142 31187.3 302.394 0.983514 0.319147 0.732505 0.7325 9.99958 2.98242e-06 1.19296e-05 0.131338 0.982274 0.931644 -0.0132928 4.90638e-06 0.503704 -1.91013e-20 7.05032e-24 -1.90943e-20 0.00139552 0.997817 8.59571e-05 0.152607 2.85204 0.00139552 0.997822 0.720865 0.00105311 0.00188018 0.000859571 0.455571 0.00188018 0.439238 0.000128995 1.02 0.887868 0.534628 0.286313 1.71725e-07 3.0655e-09 2384.4 3115.49 -0.0553575 0.482146 0.277507 0.253252 -0.593381 -0.169522 0.496923 -0.267518 -0.229414 1.84 1 0 297.815 0 2.11681 1.838 0.000299817 0.853265 0.663334 0.3733 0.414856 2.11702 132.837 83.9234 18.7211 60.8677 0.00402519 0 -40 10
0.939 2.71999e-08 2.53903e-06 0.109148 0.109146 0.0120375 1.23636e-05 0.0011541 0.136435 0.000657995 0.137088 0.884714 101.803 0.243013 0.754806 4.19684 0.0569872 0.0395928 0.960407 0.0197886 0.00431135 0.0190516 0.00414128 0.00521138 0.00594845 0.208455 0.237938 57.9977 -87.8961 126.257 15.9657 145.019 0.000141205 0.26716 192.861 0.310541 0.0673678 0.00409601 0.000561834 0.00138333 0.986982 0.991729 -2.97792e-06 -85.6647 0.0930143 31187.3 302.401 0.983514 0.319147 0.732499 0.732495 9.99958 2.98243e-06 1.19296e-05 0.13134 0.982278 0.931645 -0.0132928 4.90641e-06 0.503714 -1.91022e-20 7.05071e-24 -1.90952e-20 0.00139552 0.997817 8.59572e-05 0.152607 2.85204 0.00139552 0.997822 0.720962 0.00105312 0.00188018 0.000859572 0.455571 0.00188018 0.439245 0.000128998 1.02 0.887869 0.534628 0.286314 1.71725e-07 3.06552e-09 2384.39 3115.46 -0.055357 0.482146 0.277506 0.25325 -0.593381 -0.169522 0.496923 -0.267516 -0.229416 1.841 1 0 297.816 0 2.11697 1.839 0.000299817 0.853257 0.663382 0.373171 0.414882 2.11718 132.846 83.9236 18.7211 60.8678 0.00402518 0 -40 10
0.94 2.72289e-08 2.53903e-06 0.109212 0.10921 0.0120375 1.23768e-05 0.0011541 0.136515 0.000657997 0.137168 0.884784 101.803 0.243004 0.754911 4.1971 0.0569955 0.0395953 0.960405 0.0197883 0.00431158 0.0190513 0.00414148 0.00521167 0.00594873 0.208467 0.237949 57.9978 -87.8961 126.257 15.9657 145.019 0.000141204 0.26716 192.861 0.31054 0.0673678 0.00409602 0.000561834 0.00138333 0.986982 0.991729 -2.97793e-06 -85.6647 0.0930143 31187.3 302.407 0.983514 0.319147 0.732494 0.73249 9.99958 2.98243e-06 1.19296e-05 0.131343 0.982282 0.931646 -0.0132928 4.90644e-06 0.503724 -1.91032e-20 7.05109e-24 -1.90961e-20 0.00139553 0.997817 8.59573e-05 0.152607 2.85204 0.00139553 0.997822 0.721059 0.00105314 0.00188018 0.000859573 0.45557 0.00188018 0.439253 0.000129001 1.02 0.88787 0.534627 0.286316 1.71726e-07 3.06555e-09 2384.37 3115.44 -0.0553565 0.482146 0.277506 0.253249 -0.593381 -0.169522 0.496924 -0.267514 -0.229419 1.842 1 0 297.817 0 2.11712 1.84 0.000299816 0.853249 0.663431 0.373041 0.414908 2.11733 132.854 83.9239 18.7211 60.8679 0.00402517 0 -40 10
0.941 2.72578e-08 2.53903e-06 0.109275 0.109273 0.0120375 1.23899e-05 0.0011541 0.136594 0.000657998 0.137247 0.884854 101.803 0.242996 0.755016 4.19736 0.0570039 0.0395977 0.960402 0.019788 0.00431182 0.019051 0.00414167 0.00521195 0.00594902 0.208478 0.237961 57.9979 -87.8961 126.257 15.9657 145.019 0.000141203 0.26716 192.86 0.31054 0.0673677 0.00409602 0.000561835 0.00138333 0.986982 0.991729 -2.97795e-06 -85.6647 0.0930144 31187.3 302.413 0.983514 0.319147 0.732489 0.732485 9.99958 2.98244e-06 1.19296e-05 0.131345 0.982286 0.931647 -0.0132928 4.90647e-06 0.503734 -1.91041e-20 7.05148e-24 -1.90971e-20 0.00139553 0.997817 8.59574e-05 0.152607 2.85204 0.00139553 0.997822 0.721156 0.00105316 0.00188018 0.000859574 0.45557 0.00188018 0.439261 0.000129005 1.02 0.887871 0.534627 0.286317 1.71726e-07 3.06557e-09 2384.35 3115.42 -0.0553561 0.482147 0.277506 0.253248 -0.593381 -0.169522 0.496924 -0.267512 -0.229421 1.843 1 0 297.818 0 2.11727 1.841 0.000299816 0.853242 0.663479 0.372912 0.414934 2.11749 132.862 83.9242 18.7211 60.868 0.00402516 0 -40 10
0.942 2.72867e-08 2.53903e-06 0.109339 0.109337 0.0120375 1.2403e-05 0.0011541 0.136673 0.000658 0.137327 0.884924 101.802 0.242988 0.755121 4.19762 0.0570123 0.0396002 0.9604 0.0197878 0.00431205 0.0190507 0.00414187 0.00521224 0.00594931 0.20849 0.237972 57.9979 -87.8961 126.257 15.9656 145.019 0.000141202 0.26716 192.86 0.310539 0.0673677 0.00409602 0.000561836 0.00138334 0.986982 0.991729 -2.97796e-06 -85.6646 0.0930145 31187.3 302.42 0.983514 0.319147 0.732484 0.732479 9.99958 2.98244e-06 1.19297e-05 0.131348 0.98229 0.931648 -0.0132928 4.9065e-06 0.503743 -1.91051e-20 7.05187e-24 -1.9098e-20 0.00139553 0.997817 8.59575e-05 0.152607 2.85204 0.00139553 0.997822 0.721253 0.00105318 0.00188018 0.000859575 0.45557 0.00188018 0.439269 0.000129008 1.02 0.887872 0.534627 0.286319 1.71726e-07 3.06559e-09 2384.34 3115.4 -0.0553557 0.482147 0.277505 0.253246 -0.593381 -0.169522 0.496924 -0.26751 -0.229424 1.844 1 0 297.818 0 2.11743 1.842 0.000299815 0.853234 0.663528 0.372783 0.414959 2.11764 132.87 83.9244 18.7211 60.8682 0.00402515 0 -40 10
0.943 2.73156e-08 2.53903e-06 0.109402 0.1094 0.0120375 1.24162e-05 0.0011541 0.136753 0.000658002 0.137406 0.884994 101.802 0.242979 0.755226 4.19788 0.0570207 0.0396026 0.960397 0.0197875 0.00431228 0.0190504 0.00414207 0.00521253 0.00594959 0.208501 0.237984 57.998 -87.8961 126.257 15.9656 145.019 0.000141201 0.26716 192.86 0.310539 0.0673676 0.00409603 0.000561836 0.00138334 0.986982 0.991729 -2.97798e-06 -85.6646 0.0930146 31187.2 302.426 0.983514 0.319147 0.732479 0.732474 9.99958 2.98245e-06 1.19297e-05 0.13135 0.982293 0.931649 -0.0132928 4.90653e-06 0.503753 -1.9106e-20 7.05227e-24 -1.9099e-20 0.00139553 0.997817 8.59575e-05 0.152607 2.85204 0.00139553 0.997822 0.72135 0.0010532 0.00188018 0.000859575 0.45557 0.00188018 0.439276 0.000129011 1.02 0.887873 0.534626 0.28632 1.71726e-07 3.06561e-09 2384.32 3115.37 -0.0553553 0.482147 0.277505 0.253245 -0.593382 -0.169522 0.496925 -0.267508 -0.229426 1.845 1 0 297.819 0 2.11758 1.843 0.000299815 0.853227 0.663576 0.372655 0.414985 2.1178 132.879 83.9247 18.7211 60.8683 0.00402514 0 -40 10
0.944 2.73445e-08 2.53903e-06 0.109465 0.109464 0.0120375 1.24293e-05 0.0011541 0.136832 0.000658004 0.137485 0.885064 101.802 0.242971 0.755331 4.19814 0.0570291 0.0396051 0.960395 0.0197872 0.00431252 0.0190501 0.00414226 0.00521281 0.00594988 0.208513 0.237995 57.9981 -87.8961 126.257 15.9656 145.019 0.0001412 0.267161 192.86 0.310538 0.0673676 0.00409603 0.000561837 0.00138334 0.986982 0.991729 -2.97799e-06 -85.6646 0.0930147 31187.2 302.432 0.983514 0.319147 0.732474 0.732469 9.99958 2.98245e-06 1.19297e-05 0.131352 0.982297 0.93165 -0.0132928 4.90656e-06 0.503763 -1.91069e-20 7.05266e-24 -1.90999e-20 0.00139553 0.997817 8.59576e-05 0.152608 2.85204 0.00139553 0.997822 0.721447 0.00105322 0.00188019 0.000859576 0.45557 0.00188018 0.439284 0.000129014 1.02 0.887874 0.534626 0.286322 1.71727e-07 3.06564e-09 2384.3 3115.35 -0.0553549 0.482147 0.277505 0.253244 -0.593382 -0.169522 0.496925 -0.267506 -0.229429 1.846 1 0 297.82 0 2.11774 1.844 0.000299814 0.85322 0.663625 0.372527 0.415011 2.11795 132.887 83.9249 18.7211 60.8684 0.00402513 0 -40 10
0.945 2.73735e-08 2.53903e-06 0.109529 0.109527 0.0120375 1.24425e-05 0.0011541 0.136911 0.000658006 0.137564 0.885134 101.802 0.242963 0.755436 4.1984 0.0570375 0.0396075 0.960392 0.0197869 0.00431275 0.0190498 0.00414246 0.0052131 0.00595017 0.208524 0.238007 57.9981 -87.8961 126.258 15.9655 145.019 0.000141199 0.267161 192.86 0.310538 0.0673675 0.00409603 0.000561838 0.00138334 0.986982 0.991729 -2.97801e-06 -85.6646 0.0930148 31187.2 302.439 0.983514 0.319147 0.732469 0.732465 9.99958 2.98246e-06 1.19297e-05 0.131355 0.982301 0.931651 -0.0132928 4.90659e-06 0.503773 -1.91079e-20 7.05305e-24 -1.91008e-20 0.00139553 0.997817 8.59577e-05 0.152608 2.85204 0.00139553 0.997822 0.721544 0.00105324 0.00188019 0.000859577 0.455569 0.00188019 0.439292 0.000129017 1.02 0.887875 0.534626 0.286323 1.71727e-07 3.06566e-09 2384.29 3115.33 -0.0553545 0.482147 0.277505 0.253242 -0.593382 -0.169522 0.496925 -0.267503 -0.229431 1.847 1 0 297.821 0 2.11789 1.845 0.000299814 0.853213 0.663673 0.372399 0.415037 2.11811 132.895 83.9251 18.7212 60.8685 0.00402512 0 -40 10
0.946 2.74024e-08 2.53903e-06 0.109592 0.10959 0.0120374 1.24556e-05 0.0011541 0.13699 0.000658008 0.137643 0.885204 101.801 0.242954 0.755542 4.19866 0.0570459 0.03961 0.96039 0.0197866 0.00431299 0.0190495 0.00414266 0.00521339 0.00595046 0.208536 0.238018 57.9982 -87.8961 126.258 15.9655 145.019 0.000141198 0.267161 192.86 0.310538 0.0673675 0.00409603 0.000561838 0.00138334 0.986982 0.991729 -2.97802e-06 -85.6646 0.0930149 31187.2 302.445 0.983514 0.319147 0.732464 0.73246 9.99958 2.98246e-06 1.19297e-05 0.131357 0.982305 0.931652 -0.0132928 4.90661e-06 0.503783 -1.91088e-20 7.05344e-24 -1.91018e-20 0.00139553 0.997817 8.59578e-05 0.152608 2.85205 0.00139553 0.997822 0.721641 0.00105326 0.00188019 0.000859578 0.455569 0.00188019 0.4393 0.00012902 1.02 0.887876 0.534626 0.286325 1.71727e-07 3.06568e-09 2384.27 3115.31 -0.0553542 0.482147 0.277504 0.253241 -0.593382 -0.169522 0.496925 -0.267501 -0.229433 1.848 1 0 297.821 0 2.11805 1.846 0.000299813 0.853206 0.663721 0.372271 0.415062 2.11826 132.904 83.9254 18.7212 60.8686 0.00402511 0 -40 10
0.947 2.74313e-08 2.53903e-06 0.109655 0.109653 0.0120374 1.24688e-05 0.0011541 0.137069 0.000658009 0.137722 0.885275 101.801 0.242946 0.755647 4.19892 0.0570543 0.0396124 0.960388 0.0197863 0.00431322 0.0190493 0.00414285 0.00521368 0.00595075 0.208547 0.23803 57.9983 -87.8961 126.258 15.9654 145.019 0.000141197 0.267161 192.859 0.310537 0.0673674 0.00409604 0.000561839 0.00138335 0.986982 0.991729 -2.97804e-06 -85.6646 0.0930149 31187.1 302.451 0.983514 0.319147 0.732459 0.732455 9.99958 2.98247e-06 1.19298e-05 0.13136 0.982309 0.931653 -0.0132928 4.90664e-06 0.503793 -1.91098e-20 7.05383e-24 -1.91027e-20 0.00139553 0.997817 8.59579e-05 0.152608 2.85205 0.00139553 0.997822 0.721738 0.00105328 0.00188019 0.000859579 0.455569 0.00188019 0.439307 0.000129023 1.02 0.887877 0.534625 0.286326 1.71727e-07 3.0657e-09 2384.25 3115.29 -0.0553538 0.482147 0.277504 0.25324 -0.593383 -0.169522 0.496925 -0.267499 -0.229435 1.849 1 0 297.822 0 2.1182 1.847 0.000299813 0.853199 0.66377 0.372143 0.415088 2.11841 132.912 83.9256 18.7212 60.8687 0.0040251 0 -40 10
0.948 2.74602e-08 2.53903e-06 0.109718 0.109717 0.0120374 1.24819e-05 0.00115411 0.137148 0.000658011 0.137801 0.885345 101.801 0.242937 0.755752 4.19918 0.0570627 0.0396149 0.960385 0.019786 0.00431346 0.019049 0.00414305 0.00521397 0.00595104 0.208559 0.238042 57.9983 -87.8961 126.258 15.9654 145.019 0.000141196 0.267161 192.859 0.310537 0.0673674 0.00409604 0.00056184 0.00138335 0.986982 0.991729 -2.97805e-06 -85.6646 0.093015 31187.1 302.458 0.983514 0.319147 0.732454 0.73245 9.99958 2.98247e-06 1.19298e-05 0.131362 0.982312 0.931654 -0.0132928 4.90667e-06 0.503803 -1.91107e-20 7.05422e-24 -1.91037e-20 0.00139553 0.997817 8.59579e-05 0.152608 2.85205 0.00139553 0.997822 0.721834 0.0010533 0.00188019 0.000859579 0.455569 0.00188019 0.439315 0.000129027 1.02 0.887879 0.534625 0.286328 1.71728e-07 3.06573e-09 2384.24 3115.27 -0.0553535 0.482147 0.277504 0.253238 -0.593383 -0.169522 0.496925 -0.267497 -0.229437 1.85 1 0 297.823 0 2.11836 1.848 0.000299812 0.853192 0.663818 0.372016 0.415114 2.11857 132.92 83.9259 18.7212 60.8689 0.00402509 0 -40 10
0.949 2.74891e-08 2.53903e-06 0.109782 0.10978 0.0120374 1.24951e-05 0.00115411 0.137227 0.000658013 0.13788 0.885415 101.801 0.242929 0.755858 4.19944 0.0570711 0.0396174 0.960383 0.0197857 0.00431369 0.0190487 0.00414325 0.00521426 0.00595133 0.20857 0.238053 57.9984 -87.8961 126.258 15.9654 145.019 0.000141195 0.267162 192.859 0.310536 0.0673673 0.00409604 0.00056184 0.00138335 0.986982 0.991729 -2.97807e-06 -85.6646 0.0930151 31187.1 302.464 0.983514 0.319147 0.73245 0.732445 9.99958 2.98248e-06 1.19298e-05 0.131364 0.982316 0.931655 -0.0132928 4.9067e-06 0.503813 -1.91117e-20 7.05461e-24 -1.91046e-20 0.00139554 0.997817 8.5958e-05 0.152608 2.85205 0.00139554 0.997822 0.721931 0.00105332 0.00188019 0.00085958 0.455568 0.00188019 0.439323 0.00012903 1.02 0.88788 0.534625 0.286329 1.71728e-07 3.06575e-09 2384.22 3115.25 -0.0553532 0.482147 0.277503 0.253237 -0.593383 -0.169522 0.496925 -0.267495 -0.229439 1.851 1 0 297.823 0 2.11851 1.849 0.000299812 0.853186 0.663867 0.371889 0.415139 2.11872 132.928 83.9261 18.7212 60.869 0.00402508 0 -40 10
0.95 2.75181e-08 2.53903e-06 0.109845 0.109843 0.0120374 1.25082e-05 0.00115411 0.137306 0.000658015 0.137959 0.885485 101.8 0.24292 0.755963 4.19971 0.0570795 0.0396199 0.96038 0.0197855 0.00431393 0.0190484 0.00414345 0.00521455 0.00595162 0.208582 0.238065 57.9984 -87.8961 126.258 15.9653 145.019 0.000141194 0.267162 192.859 0.310536 0.0673673 0.00409605 0.000561841 0.00138335 0.986982 0.991729 -2.97808e-06 -85.6646 0.0930152 31187.1 302.47 0.983514 0.319147 0.732445 0.732441 9.99958 2.98248e-06 1.19298e-05 0.131367 0.98232 0.931656 -0.0132928 4.90673e-06 0.503823 -1.91126e-20 7.05501e-24 -1.91056e-20 0.00139554 0.997817 8.59581e-05 0.152608 2.85205 0.00139554 0.997822 0.722028 0.00105333 0.00188019 0.000859581 0.455568 0.00188019 0.439331 0.000129033 1.02 0.887881 0.534624 0.286331 1.71728e-07 3.06577e-09 2384.2 3115.23 -0.0553529 0.482147 0.277503 0.253236 -0.593383 -0.169522 0.496925 -0.267493 -0.229441 1.852 1 0 297.824 0 2.11867 1.85 0.000299811 0.853179 0.663915 0.371762 0.415165 2.11888 132.937 83.9263 18.7212 60.8691 0.00402507 0 -40 10
0.951 2.7547e-08 2.53903e-06 0.109908 0.109906 0.0120374 1.25214e-05 0.00115411 0.137385 0.000658017 0.138038 0.885556 101.8 0.242912 0.756069 4.19997 0.057088 0.0396224 0.960378 0.0197852 0.00431416 0.0190481 0.00414365 0.00521484 0.00595191 0.208594 0.238076 57.9985 -87.8961 126.258 15.9653 145.02 0.000141193 0.267162 192.859 0.310535 0.0673672 0.00409605 0.000561842 0.00138336 0.986982 0.991729 -2.9781e-06 -85.6646 0.0930153 31187.1 302.477 0.983514 0.319147 0.732441 0.732436 9.99958 2.98249e-06 1.19298e-05 0.131369 0.982324 0.931657 -0.0132928 4.90676e-06 0.503833 -1.91136e-20 7.0554e-24 -1.91065e-20 0.00139554 0.997817 8.59582e-05 0.152609 2.85205 0.00139554 0.997822 0.722125 0.00105335 0.0018802 0.000859582 0.455568 0.00188019 0.439338 0.000129036 1.02 0.887882 0.534624 0.286332 1.71728e-07 3.0658e-09 2384.19 3115.21 -0.0553527 0.482147 0.277503 0.253235 -0.593383 -0.169522 0.496925 -0.267491 -0.229443 1.853 1 0 297.825 0 2.11882 1.851 0.000299811 0.853173 0.663963 0.371636 0.415191 2.11903 132.945 83.9266 18.7212 60.8692 0.00402506 0 -40 10
0.952 2.75759e-08 2.53903e-06 0.109971 0.109969 0.0120374 1.25345e-05 0.00115411 0.137463 0.000658018 0.138117 0.885626 101.8 0.242904 0.756175 4.20023 0.0570964 0.0396248 0.960375 0.0197849 0.0043144 0.0190478 0.00414385 0.00521513 0.0059522 0.208605 0.238088 57.9986 -87.8961 126.258 15.9653 145.02 0.000141192 0.267162 192.859 0.310535 0.0673672 0.00409605 0.000561842 0.00138336 0.986981 0.991729 -2.97811e-06 -85.6645 0.0930154 31187 302.483 0.983514 0.319147 0.732436 0.732432 9.99958 2.98249e-06 1.19299e-05 0.131372 0.982327 0.931658 -0.0132928 4.90679e-06 0.503842 -1.91145e-20 7.05579e-24 -1.91075e-20 0.00139554 0.997817 8.59583e-05 0.152609 2.85205 0.00139554 0.997822 0.722221 0.00105337 0.0018802 0.000859583 0.455568 0.0018802 0.439346 0.000129039 1.02 0.887883 0.534624 0.286334 1.71729e-07 3.06582e-09 2384.17 3115.19 -0.0553524 0.482147 0.277503 0.253233 -0.593384 -0.169522 0.496925 -0.267489 -0.229445 1.854 1 0 297.825 0 2.11897 1.852 0.00029981 0.853167 0.664012 0.37151 0.415216 2.11919 132.953 83.9268 18.7213 60.8693 0.00402505 0 -40 10
0.953 2.76048e-08 2.53903e-06 0.110034 0.110032 0.0120373 1.25476e-05 0.00115411 0.137542 0.00065802 0.138195 0.885697 101.8 0.242895 0.75628 4.2005 0.0571048 0.0396273 0.960373 0.0197846 0.00431464 0.0190475 0.00414404 0.00521542 0.00595249 0.208617 0.2381 57.9986 -87.8961 126.258 15.9652 145.02 0.000141192 0.267162 192.859 0.310535 0.0673671 0.00409606 0.000561843 0.00138336 0.986981 0.991729 -2.97813e-06 -85.6645 0.0930155 31187 302.49 0.983514 0.319147 0.732431 0.732427 9.99958 2.9825e-06 1.19299e-05 0.131374 0.982331 0.931659 -0.0132928 4.90682e-06 0.503852 -1.91155e-20 7.05618e-24 -1.91084e-20 0.00139554 0.997817 8.59583e-05 0.152609 2.85205 0.00139554 0.997822 0.722318 0.00105339 0.0018802 0.000859583 0.455568 0.0018802 0.439354 0.000129042 1.02 0.887884 0.534623 0.286335 1.71729e-07 3.06584e-09 2384.15 3115.17 -0.0553522 0.482147 0.277502 0.253232 -0.593384 -0.169523 0.496925 -0.267487 -0.229447 1.855 1 0 297.826 0 2.11913 1.853 0.00029981 0.85316 0.66406 0.371384 0.415242 2.11934 132.961 83.927 18.7213 60.8694 0.00402504 0 -40 10
0.954 2.76337e-08 2.53904e-06 0.110096 0.110095 0.0120373 1.25608e-05 0.00115411 0.137621 0.000658022 0.138274 0.885767 101.799 0.242887 0.756386 4.20076 0.0571133 0.0396298 0.96037 0.0197843 0.00431487 0.0190472 0.00414424 0.00521571 0.00595278 0.208628 0.238111 57.9987 -87.8961 126.258 15.9652 145.02 0.000141191 0.267163 192.858 0.310534 0.0673671 0.00409606 0.000561844 0.00138336 0.986981 0.991729 -2.97814e-06 -85.6645 0.0930156 31187 302.496 0.983514 0.319147 0.732427 0.732423 9.99958 2.9825e-06 1.19299e-05 0.131376 0.982335 0.93166 -0.0132928 4.90685e-06 0.503862 -1.91164e-20 7.05658e-24 -1.91093e-20 0.00139554 0.997817 8.59584e-05 0.152609 2.85205 0.00139554 0.997822 0.722414 0.00105341 0.0018802 0.000859584 0.455567 0.0018802 0.439361 0.000129045 1.02 0.887885 0.534623 0.286337 1.71729e-07 3.06586e-09 2384.14 3115.15 -0.055352 0.482148 0.277502 0.253231 -0.593384 -0.169523 0.496924 -0.267484 -0.229449 1.856 1 0 297.827 0 2.11928 1.854 0.000299809 0.853154 0.664108 0.371258 0.415268 2.11949 132.97 83.9272 18.7213 60.8695 0.00402503 0 -40 10
0.955 2.76627e-08 2.53904e-06 0.110159 0.110157 0.0120373 1.25739e-05 0.00115411 0.137699 0.000658024 0.138352 0.885838 101.799 0.242878 0.756492 4.20103 0.0571217 0.0396323 0.960368 0.019784 0.00431511 0.0190469 0.00414444 0.005216 0.00595308 0.20864 0.238123 57.9988 -87.8961 126.258 15.9651 145.02 0.00014119 0.267163 192.858 0.310534 0.067367 0.00409606 0.000561844 0.00138336 0.986981 0.991729 -2.97816e-06 -85.6645 0.0930156 31187 302.503 0.983514 0.319147 0.732423 0.732418 9.99958 2.98251e-06 1.19299e-05 0.131379 0.982338 0.931661 -0.0132928 4.90688e-06 0.503872 -1.91174e-20 7.05697e-24 -1.91103e-20 0.00139554 0.997817 8.59585e-05 0.152609 2.85205 0.00139554 0.997822 0.722511 0.00105343 0.0018802 0.000859585 0.455567 0.0018802 0.439369 0.000129048 1.02 0.887886 0.534623 0.286338 1.7173e-07 3.06589e-09 2384.12 3115.13 -0.0553518 0.482148 0.277502 0.25323 -0.593384 -0.169523 0.496924 -0.267482 -0.229451 1.857 1 0 297.827 0 2.11944 1.855 0.000299809 0.853148 0.664156 0.371133 0.415293 2.11965 132.978 83.9274 18.7213 60.8696 0.00402502 0 -40 10
0.956 2.76916e-08 2.53904e-06 0.110222 0.11022 0.0120373 1.25871e-05 0.00115411 0.137777 0.000658026 0.138431 0.885908 101.799 0.24287 0.756598 4.20129 0.0571302 0.0396348 0.960365 0.0197837 0.00431535 0.0190466 0.00414464 0.0052163 0.00595337 0.208652 0.238135 57.9988 -87.8961 126.259 15.9651 145.02 0.000141189 0.267163 192.858 0.310533 0.0673669 0.00409606 0.000561845 0.00138337 0.986981 0.991729 -2.97817e-06 -85.6645 0.0930157 31186.9 302.509 0.983514 0.319147 0.732418 0.732414 9.99958 2.98251e-06 1.19299e-05 0.131381 0.982342 0.931662 -0.0132928 4.90691e-06 0.503883 -1.91183e-20 7.05736e-24 -1.91112e-20 0.00139554 0.997817 8.59586e-05 0.152609 2.85205 0.00139554 0.997822 0.722607 0.00105345 0.0018802 0.000859586 0.455567 0.0018802 0.439377 0.000129052 1.02 0.887887 0.534622 0.28634 1.7173e-07 3.06591e-09 2384.1 3115.11 -0.0553517 0.482148 0.277501 0.253229 -0.593384 -0.169523 0.496923 -0.26748 -0.229452 1.858 1 0 297.828 0 2.11959 1.856 0.000299808 0.853143 0.664205 0.371007 0.415319 2.1198 132.986 83.9276 18.7213 60.8697 0.00402501 0 -40 10
0.957 2.77205e-08 2.53904e-06 0.110285 0.110283 0.0120373 1.26002e-05 0.00115411 0.137856 0.000658027 0.138509 0.885979 101.798 0.242861 0.756704 4.20156 0.0571386 0.0396373 0.960363 0.0197834 0.00431559 0.0190463 0.00414484 0.00521659 0.00595366 0.208664 0.238147 57.9989 -87.8962 126.259 15.9651 145.02 0.000141188 0.267163 192.858 0.310533 0.0673669 0.00409607 0.000561846 0.00138337 0.986981 0.991729 -2.97819e-06 -85.6645 0.0930158 31186.9 302.515 0.983514 0.319147 0.732414 0.73241 9.99958 2.98252e-06 1.193e-05 0.131384 0.982346 0.931663 -0.0132927 4.90694e-06 0.503893 -1.91193e-20 7.05776e-24 -1.91122e-20 0.00139554 0.997817 8.59587e-05 0.15261 2.85206 0.00139554 0.997822 0.722704 0.00105347 0.0018802 0.000859587 0.455567 0.0018802 0.439385 0.000129055 1.02 0.887888 0.534622 0.286341 1.7173e-07 3.06593e-09 2384.09 3115.09 -0.0553515 0.482148 0.277501 0.253228 -0.593385 -0.169523 0.496923 -0.267478 -0.229454 1.859 1 0 297.828 0 2.11974 1.857 0.000299808 0.853137 0.664253 0.370883 0.415345 2.11996 132.995 83.9279 18.7213 60.8698 0.00402501 0 -40 10
0.958 2.77494e-08 2.53904e-06 0.110347 0.110346 0.0120373 1.26134e-05 0.00115411 0.137934 0.000658029 0.138588 0.886049 101.798 0.242853 0.75681 4.20182 0.0571471 0.0396398 0.96036 0.0197831 0.00431582 0.019046 0.00414504 0.00521688 0.00595396 0.208675 0.238158 57.999 -87.8962 126.259 15.965 145.02 0.000141187 0.267163 192.858 0.310533 0.0673668 0.00409607 0.000561846 0.00138337 0.986981 0.991729 -2.9782e-06 -85.6645 0.0930159 31186.9 302.522 0.983514 0.319147 0.73241 0.732406 9.99958 2.98252e-06 1.193e-05 0.131386 0.982349 0.931664 -0.0132927 4.90697e-06 0.503903 -1.91202e-20 7.05815e-24 -1.91131e-20 0.00139555 0.997817 8.59587e-05 0.15261 2.85206 0.00139555 0.997822 0.7228 0.00105349 0.00188021 0.000859587 0.455566 0.0018802 0.439392 0.000129058 1.02 0.887889 0.534622 0.286343 1.7173e-07 3.06595e-09 2384.07 3115.07 -0.0553514 0.482148 0.277501 0.253226 -0.593385 -0.169523 0.496922 -0.267476 -0.229456 1.86 1 0 297.829 0 2.1199 1.858 0.000299807 0.853131 0.664301 0.370758 0.41537 2.12011 133.003 83.9281 18.7213 60.8699 0.004025 0 -40 10
0.959 2.77784e-08 2.53904e-06 0.11041 0.110408 0.0120373 1.26265e-05 0.00115411 0.138012 0.000658031 0.138666 0.88612 101.798 0.242844 0.756916 4.20209 0.0571556 0.0396424 0.960358 0.0197828 0.00431606 0.0190457 0.00414525 0.00521717 0.00595425 0.208687 0.23817 57.999 -87.8962 126.259 15.965 145.02 0.000141187 0.267163 192.858 0.310532 0.0673668 0.00409607 0.000561847 0.00138337 0.986981 0.991729 -2.97822e-06 -85.6645 0.093016 31186.9 302.528 0.983514 0.319147 0.732406 0.732401 9.99958 2.98253e-06 1.193e-05 0.131389 0.982353 0.931665 -0.0132927 4.907e-06 0.503913 -1.91212e-20 7.05855e-24 -1.91141e-20 0.00139555 0.997817 8.59588e-05 0.15261 2.85206 0.00139555 0.997822 0.722897 0.00105351 0.00188021 0.000859588 0.455566 0.00188021 0.4394 0.000129061 1.02 0.887891 0.534622 0.286345 1.71731e-07 3.06598e-09 2384.05 3115.05 -0.0553513 0.482148 0.277501 0.253225 -0.593385 -0.169523 0.496922 -0.267474 -0.229457 1.861 1 0 297.829 0 2.12005 1.859 0.000299807 0.853126 0.664349 0.370634 0.415396 2.12026 133.011 83.9283 18.7213 60.87 0.00402499 0 -40 10
0.96 2.78073e-08 2.53904e-06 0.110473 0.110471 0.0120373 1.26397e-05 0.00115411 0.138091 0.000658033 0.138744 0.886191 101.798 0.242836 0.757022 4.20236 0.057164 0.0396449 0.960355 0.0197825 0.0043163 0.0190455 0.00414545 0.00521747 0.00595455 0.208699 0.238182 57.9991 -87.8962 126.259 15.9649 145.02 0.000141186 0.267164 192.857 0.310532 0.0673667 0.00409608 0.000561848 0.00138337 0.986981 0.991729 -2.97823e-06 -85.6645 0.0930161 31186.9 302.535 0.983514 0.319147 0.732402 0.732397 9.99958 2.98253e-06 1.193e-05 0.131391 0.982357 0.931666 -0.0132927 4.90703e-06 0.503923 -1.91221e-20 7.05894e-24 -1.9115e-20 0.00139555 0.997817 8.59589e-05 0.15261 2.85206 0.00139555 0.997822 0.722993 0.00105352 0.00188021 0.000859589 0.455566 0.00188021 0.439408 0.000129064 1.02 0.887892 0.534621 0.286346 1.71731e-07 3.066e-09 2384.04 3115.03 -0.0553512 0.482148 0.2775 0.253224 -0.593385 -0.169523 0.496921 -0.267472 -0.229459 1.862 1 0 297.83 0 2.12021 1.86 0.000299806 0.85312 0.664398 0.370509 0.415421 2.12042 133.019 83.9285 18.7214 60.8701 0.00402498 0 -40 10
0.961 2.78362e-08 2.53904e-06 0.110535 0.110533 0.0120372 1.26528e-05 0.00115411 0.138169 0.000658034 0.138822 0.886261 101.797 0.242828 0.757128 4.20262 0.0571725 0.0396474 0.960353 0.0197822 0.00431654 0.0190452 0.00414565 0.00521776 0.00595484 0.208711 0.238194 57.9991 -87.8962 126.259 15.9649 145.02 0.000141185 0.267164 192.857 0.310531 0.0673667 0.00409608 0.000561848 0.00138338 0.986981 0.991729 -2.97824e-06 -85.6645 0.0930162 31186.8 302.541 0.983514 0.319147 0.732398 0.732393 9.99958 2.98254e-06 1.193e-05 0.131393 0.98236 0.931667 -0.0132927 4.90706e-06 0.503933 -1.91231e-20 7.05934e-24 -1.9116e-20 0.00139555 0.997817 8.5959e-05 0.15261 2.85206 0.00139555 0.997822 0.723089 0.00105354 0.00188021 0.00085959 0.455566 0.00188021 0.439415 0.000129067 1.02 0.887893 0.534621 0.286348 1.71731e-07 3.06602e-09 2384.02 3115.02 -0.0553511 0.482148 0.2775 0.253223 -0.593385 -0.169523 0.496921 -0.26747 -0.22946 1.863 1 0 297.83 0 2.12036 1.861 0.000299806 0.853115 0.664446 0.370386 0.415447 2.12057 133.028 83.9287 18.7214 60.8702 0.00402497 0 -40 10
0.962 2.78651e-08 2.53904e-06 0.110598 0.110596 0.0120372 1.2666e-05 0.00115411 0.138247 0.000658036 0.1389 0.886332 101.797 0.242819 0.757234 4.20289 0.057181 0.0396499 0.96035 0.0197819 0.00431678 0.0190449 0.00414585 0.00521806 0.00595514 0.208722 0.238205 57.9992 -87.8962 126.259 15.9649 145.02 0.000141184 0.267164 192.857 0.310531 0.0673666 0.00409608 0.000561849 0.00138338 0.986981 0.991729 -2.97826e-06 -85.6645 0.0930162 31186.8 302.548 0.983514 0.319147 0.732394 0.732389 9.99958 2.98254e-06 1.19301e-05 0.131396 0.982364 0.931668 -0.0132927 4.90709e-06 0.503943 -1.9124e-20 7.05973e-24 -1.9117e-20 0.00139555 0.997817 8.59591e-05 0.15261 2.85206 0.00139555 0.997821 0.723186 0.00105356 0.00188021 0.000859591 0.455566 0.00188021 0.439423 0.00012907 1.02 0.887894 0.534621 0.286349 1.71731e-07 3.06605e-09 2384 3115 -0.055351 0.482148 0.2775 0.253222 -0.593386 -0.169523 0.49692 -0.267468 -0.229462 1.864 1 0 297.831 0 2.12051 1.862 0.000299805 0.85311 0.664494 0.370262 0.415473 2.12073 133.036 83.9289 18.7214 60.8703 0.00402496 0 -40 10
0.963 2.7894e-08 2.53904e-06 0.11066 0.110658 0.0120372 1.26791e-05 0.00115411 0.138325 0.000658038 0.138978 0.886403 101.797 0.242811 0.757341 4.20316 0.0571895 0.0396525 0.960348 0.0197816 0.00431702 0.0190446 0.00414605 0.00521835 0.00595543 0.208734 0.238217 57.9993 -87.8962 126.259 15.9648 145.02 0.000141184 0.267164 192.857 0.31053 0.0673666 0.00409609 0.00056185 0.00138338 0.986981 0.991729 -2.97827e-06 -85.6644 0.0930163 31186.8 302.554 0.983514 0.319147 0.73239 0.732385 9.99958 2.98255e-06 1.19301e-05 0.131398 0.982368 0.931669 -0.0132927 4.90712e-06 0.503953 -1.9125e-20 7.06013e-24 -1.91179e-20 0.00139555 0.997817 8.59591e-05 0.15261 2.85206 0.00139555 0.997821 0.723282 0.00105358 0.00188021 0.000859591 0.455565 0.00188021 0.439431 0.000129073 1.02 0.887895 0.53462 0.286351 1.71732e-07 3.06607e-09 2383.99 3114.98 -0.055351 0.482148 0.277499 0.253221 -0.593386 -0.169523 0.496919 -0.267466 -0.229463 1.865 1 0 297.831 0 2.12067 1.863 0.000299804 0.853105 0.664542 0.370139 0.415498 2.12088 133.044 83.9291 18.7214 60.8704 0.00402496 0 -40 10
0.964 2.79229e-08 2.53904e-06 0.110722 0.110721 0.0120372 1.26922e-05 0.00115411 0.138403 0.00065804 0.139056 0.886474 101.797 0.242802 0.757447 4.20343 0.057198 0.039655 0.960345 0.0197814 0.00431726 0.0190443 0.00414625 0.00521865 0.00595573 0.208746 0.238229 57.9993 -87.8962 126.259 15.9648 145.02 0.000141183 0.267164 192.857 0.31053 0.0673665 0.00409609 0.00056185 0.00138338 0.986981 0.991729 -2.97829e-06 -85.6644 0.0930164 31186.8 302.561 0.983514 0.319147 0.732386 0.732381 9.99958 2.98255e-06 1.19301e-05 0.131401 0.982371 0.93167 -0.0132927 4.90715e-06 0.503963 -1.91259e-20 7.06052e-24 -1.91189e-20 0.00139555 0.997817 8.59592e-05 0.152611 2.85206 0.00139555 0.997821 0.723378 0.0010536 0.00188022 0.000859592 0.455565 0.00188021 0.439438 0.000129077 1.02 0.887896 0.53462 0.286352 1.71732e-07 3.06609e-09 2383.97 3114.96 -0.0553509 0.482148 0.277499 0.25322 -0.593386 -0.169523 0.496918 -0.267463 -0.229464 1.866 1 0 297.832 0 2.12082 1.864 0.000299804 0.8531 0.66459 0.370016 0.415524 2.12103 133.052 83.9293 18.7214 60.8705 0.00402495 0 -40 10
0.965 2.79519e-08 2.53904e-06 0.110785 0.110783 0.0120372 1.27054e-05 0.00115411 0.138481 0.000658041 0.139134 0.886545 101.796 0.242794 0.757553 4.2037 0.0572065 0.0396575 0.960342 0.0197811 0.0043175 0.019044 0.00414646 0.00521894 0.00595602 0.208758 0.238241 57.9994 -87.8962 126.259 15.9648 145.02 0.000141182 0.267165 192.857 0.31053 0.0673665 0.00409609 0.000561851 0.00138339 0.986981 0.991729 -2.9783e-06 -85.6644 0.0930165 31186.7 302.567 0.983514 0.319147 0.732382 0.732378 9.99958 2.98256e-06 1.19301e-05 0.131403 0.982375 0.931671 -0.0132927 4.90718e-06 0.503973 -1.91269e-20 7.06092e-24 -1.91198e-20 0.00139555 0.997817 8.59593e-05 0.152611 2.85206 0.00139555 0.997821 0.723475 0.00105362 0.00188022 0.000859593 0.455565 0.00188022 0.439446 0.00012908 1.02 0.887897 0.53462 0.286354 1.71732e-07 3.06611e-09 2383.95 3114.95 -0.0553509 0.482148 0.277499 0.253219 -0.593386 -0.169523 0.496917 -0.267461 -0.229465 1.867 1 0 297.832 0 2.12098 1.865 0.000299803 0.853095 0.664639 0.369893 0.415549 2.12119 133.06 83.9294 18.7214 60.8706 0.00402494 0 -40 10
0.966 2.79808e-08 2.53904e-06 0.110847 0.110845 0.0120372 1.27185e-05 0.00115411 0.138559 0.000658043 0.139212 0.886616 101.796 0.242785 0.75766 4.20397 0.057215 0.0396601 0.96034 0.0197808 0.00431774 0.0190437 0.00414666 0.00521924 0.00595632 0.20877 0.238253 57.9995 -87.8962 126.259 15.9647 145.02 0.000141181 0.267165 192.856 0.310529 0.0673664 0.00409609 0.000561852 0.00138339 0.986981 0.991729 -2.97832e-06 -85.6644 0.0930166 31186.7 302.574 0.983513 0.319147 0.732378 0.732374 9.99958 2.98256e-06 1.19301e-05 0.131406 0.982378 0.931672 -0.0132927 4.9072e-06 0.503984 -1.91278e-20 7.06132e-24 -1.91208e-20 0.00139556 0.997817 8.59594e-05 0.152611 2.85206 0.00139555 0.997821 0.723571 0.00105364 0.00188022 0.000859594 0.455565 0.00188022 0.439454 0.000129083 1.02 0.887898 0.534619 0.286355 1.71732e-07 3.06614e-09 2383.93 3114.93 -0.0553509 0.482148 0.277499 0.253218 -0.593386 -0.169523 0.496916 -0.267459 -0.229467 1.868 1 0 297.832 0 2.12113 1.866 0.000299803 0.85309 0.664687 0.36977 0.415575 2.12134 133.069 83.9296 18.7214 60.8707 0.00402493 0 -40 10
0.967 2.80097e-08 2.53904e-06 0.110909 0.110907 0.0120372 1.27317e-05 0.00115411 0.138636 0.000658045 0.13929 0.886687 101.796 0.242777 0.757766 4.20424 0.0572235 0.0396626 0.960337 0.0197805 0.00431798 0.0190434 0.00414686 0.00521954 0.00595662 0.208781 0.238265 57.9995 -87.8962 126.259 15.9647 145.02 0.000141181 0.267165 192.856 0.310529 0.0673664 0.0040961 0.000561852 0.00138339 0.986981 0.991729 -2.97833e-06 -85.6644 0.0930167 31186.7 302.58 0.983513 0.319147 0.732375 0.73237 9.99958 2.98257e-06 1.19302e-05 0.131408 0.982382 0.931673 -0.0132927 4.90723e-06 0.503994 -1.91288e-20 7.06171e-24 -1.91217e-20 0.00139556 0.997817 8.59595e-05 0.152611 2.85206 0.00139556 0.997821 0.723667 0.00105366 0.00188022 0.000859595 0.455564 0.00188022 0.439461 0.000129086 1.02 0.887899 0.534619 0.286357 1.71733e-07 3.06616e-09 2383.92 3114.91 -0.0553509 0.482149 0.277498 0.253217 -0.593386 -0.169523 0.496915 -0.267457 -0.229468 1.869 1 0 297.833 0 2.12128 1.867 0.000299802 0.853086 0.664735 0.369648 0.4156 2.12149 133.077 83.9298 18.7214 60.8708 0.00402493 0 -40 10
0.968 2.80386e-08 2.53904e-06 0.110971 0.11097 0.0120371 1.27448e-05 0.00115411 0.138714 0.000658047 0.139368 0.886758 101.795 0.242768 0.757873 4.20451 0.057232 0.0396652 0.960335 0.0197802 0.00431823 0.0190431 0.00414706 0.00521983 0.00595692 0.208793 0.238277 57.9996 -87.8962 126.259 15.9646 145.02 0.00014118 0.267165 192.856 0.310528 0.0673663 0.0040961 0.000561853 0.00138339 0.986981 0.991729 -2.97835e-06 -85.6644 0.0930168 31186.7 302.587 0.983513 0.319147 0.732371 0.732367 9.99958 2.98257e-06 1.19302e-05 0.131411 0.982385 0.931674 -0.0132927 4.90726e-06 0.504004 -1.91298e-20 7.06211e-24 -1.91227e-20 0.00139556 0.997817 8.59595e-05 0.152611 2.85207 0.00139556 0.997821 0.723763 0.00105368 0.00188022 0.000859595 0.455564 0.00188022 0.439469 0.000129089 1.02 0.8879 0.534619 0.286358 1.71733e-07 3.06618e-09 2383.9 3114.9 -0.055351 0.482149 0.277498 0.253216 -0.593387 -0.169524 0.496914 -0.267455 -0.229469 1.87 1 0 297.833 0 2.12144 1.868 0.000299802 0.853081 0.664783 0.369526 0.415626 2.12165 133.085 83.93 18.7214 60.8709 0.00402492 0 -40 10
0.969 2.80675e-08 2.53904e-06 0.111033 0.111032 0.0120371 1.2758e-05 0.00115411 0.138792 0.000658048 0.139445 0.886829 101.795 0.24276 0.75798 4.20478 0.0572405 0.0396677 0.960332 0.0197799 0.00431847 0.0190428 0.00414727 0.00522013 0.00595721 0.208805 0.238289 57.9997 -87.8962 126.259 15.9646 145.02 0.000141179 0.267165 192.856 0.310528 0.0673663 0.0040961 0.000561854 0.00138339 0.986981 0.991729 -2.97836e-06 -85.6644 0.0930169 31186.7 302.594 0.983513 0.319147 0.732367 0.732363 9.99958 2.98258e-06 1.19302e-05 0.131413 0.982389 0.931675 -0.0132927 4.90729e-06 0.504014 -1.91307e-20 7.06251e-24 -1.91236e-20 0.00139556 0.997817 8.59596e-05 0.152611 2.85207 0.00139556 0.997821 0.723859 0.00105369 0.00188022 0.000859596 0.455564 0.00188022 0.439477 0.000129092 1.02 0.887902 0.534618 0.28636 1.71733e-07 3.0662e-09 2383.88 3114.88 -0.055351 0.482149 0.277498 0.253215 -0.593387 -0.169524 0.496913 -0.267453 -0.22947 1.871 1 0 297.833 0 2.12159 1.869 0.000299801 0.853077 0.664831 0.369404 0.415651 2.1218 133.093 83.9302 18.7215 60.8709 0.00402491 0 -40 10
0.97 2.80965e-08 2.53905e-06 0.111095 0.111094 0.0120371 1.27711e-05 0.00115411 0.138869 0.00065805 0.139523 0.8869 101.795 0.242751 0.758086 4.20505 0.057249 0.0396703 0.96033 0.0197796 0.00431871 0.0190425 0.00414747 0.00522043 0.00595751 0.208817 0.2383 57.9997 -87.8962 126.259 15.9646 145.02 0.000141179 0.267166 192.856 0.310527 0.0673662 0.00409611 0.000561854 0.0013834 0.986981 0.991729 -2.97838e-06 -85.6644 0.0930169 31186.6 302.6 0.983513 0.319147 0.732364 0.732359 9.99958 2.98258e-06 1.19302e-05 0.131416 0.982392 0.931676 -0.0132927 4.90732e-06 0.504024 -1.91317e-20 7.0629e-24 -1.91246e-20 0.00139556 0.997817 8.59597e-05 0.152612 2.85207 0.00139556 0.997821 0.723955 0.00105371 0.00188022 0.000859597 0.455564 0.00188022 0.439484 0.000129095 1.02 0.887903 0.534618 0.286361 1.71734e-07 3.06623e-09 2383.87 3114.87 -0.0553511 0.482149 0.277497 0.253214 -0.593387 -0.169524 0.496912 -0.267451 -0.229471 1.872 1 0 297.834 0 2.12174 1.87 0.000299801 0.853072 0.664879 0.369282 0.415677 2.12195 133.102 83.9304 18.7215 60.871 0.0040249 0 -40 10
0.971 2.81254e-08 2.53905e-06 0.111158 0.111156 0.0120371 1.27843e-05 0.00115411 0.138947 0.000658052 0.1396 0.886971 101.795 0.242742 0.758193 4.20532 0.0572575 0.0396729 0.960327 0.0197793 0.00431895 0.0190422 0.00414768 0.00522073 0.00595781 0.208829 0.238312 57.9998 -87.8962 126.26 15.9645 145.02 0.000141178 0.267166 192.856 0.310527 0.0673662 0.00409611 0.000561855 0.0013834 0.986981 0.991729 -2.97839e-06 -85.6644 0.093017 31186.6 302.607 0.983513 0.319147 0.73236 0.732356 9.99958 2.98259e-06 1.19302e-05 0.131418 0.982396 0.931676 -0.0132927 4.90735e-06 0.504035 -1.91326e-20 7.0633e-24 -1.91256e-20 0.00139556 0.997817 8.59598e-05 0.152612 2.85207 0.00139556 0.997821 0.724051 0.00105373 0.00188023 0.000859598 0.455563 0.00188022 0.439492 0.000129098 1.02 0.887904 0.534618 0.286363 1.71734e-07 3.06625e-09 2383.85 3114.85 -0.0553512 0.482149 0.277497 0.253213 -0.593387 -0.169524 0.496911 -0.267449 -0.229472 1.873 1 0 297.834 0 2.1219 1.871 0.0002998 0.853068 0.664927 0.369161 0.415703 2.12211 133.11 83.9305 18.7215 60.8711 0.0040249 0 -40 10
0.972 2.81543e-08 2.53905e-06 0.111219 0.111218 0.0120371 1.27974e-05 0.00115411 0.139024 0.000658054 0.139678 0.887042 101.794 0.242734 0.7583 4.20559 0.0572661 0.0396754 0.960325 0.019779 0.00431919 0.0190419 0.00414788 0.00522103 0.00595811 0.208841 0.238324 57.9998 -87.8962 126.26 15.9645 145.02 0.000141177 0.267166 192.855 0.310527 0.0673661 0.00409611 0.000561856 0.0013834 0.986981 0.991729 -2.97841e-06 -85.6644 0.0930171 31186.6 302.613 0.983513 0.319147 0.732357 0.732352 9.99958 2.98259e-06 1.19303e-05 0.131421 0.982399 0.931677 -0.0132927 4.90738e-06 0.504045 -1.91336e-20 7.0637e-24 -1.91265e-20 0.00139556 0.997817 8.59599e-05 0.152612 2.85207 0.00139556 0.997821 0.724147 0.00105375 0.00188023 0.000859599 0.455563 0.00188023 0.4395 0.000129101 1.02 0.887905 0.534618 0.286364 1.71734e-07 3.06627e-09 2383.83 3114.83 -0.0553513 0.482149 0.277497 0.253212 -0.593387 -0.169524 0.49691 -0.267447 -0.229473 1.874 1 0 297.834 0 2.12205 1.872 0.0002998 0.853064 0.664975 0.36904 0.415728 2.12226 133.118 83.9307 18.7215 60.8712 0.00402489 0 -40 10
0.973 2.81832e-08 2.53905e-06 0.111281 0.11128 0.0120371 1.28106e-05 0.00115411 0.139102 0.000658055 0.139755 0.887113 101.794 0.242725 0.758407 4.20587 0.0572746 0.039678 0.960322 0.0197787 0.00431944 0.0190416 0.00414808 0.00522132 0.00595841 0.208853 0.238336 57.9999 -87.8962 126.26 15.9645 145.02 0.000141177 0.267166 192.855 0.310526 0.0673661 0.00409612 0.000561856 0.0013834 0.986981 0.991729 -2.97842e-06 -85.6644 0.0930172 31186.6 302.62 0.983513 0.319147 0.732353 0.732349 9.99958 2.9826e-06 1.19303e-05 0.131423 0.982403 0.931678 -0.0132927 4.90741e-06 0.504055 -1.91346e-20 7.0641e-24 -1.91275e-20 0.00139556 0.997817 8.59599e-05 0.152612 2.85207 0.00139556 0.997821 0.724243 0.00105377 0.00188023 0.000859599 0.455563 0.00188023 0.439507 0.000129104 1.02 0.887906 0.534617 0.286366 1.71734e-07 3.0663e-09 2383.82 3114.82 -0.0553514 0.482149 0.277497 0.253211 -0.593387 -0.169524 0.496908 -0.267444 -0.229473 1.875 1 0 297.835 0 2.1222 1.873 0.000299799 0.85306 0.665023 0.368919 0.415754 2.12241 133.126 83.9309 18.7215 60.8713 0.00402488 0 -40 10
0.974 2.82121e-08 2.53905e-06 0.111343 0.111342 0.0120371 1.28237e-05 0.00115411 0.139179 0.000658057 0.139833 0.887184 101.794 0.242717 0.758514 4.20614 0.0572831 0.0396806 0.960319 0.0197784 0.00431968 0.0190413 0.00414829 0.00522162 0.00595871 0.208865 0.238348 58 -87.8962 126.26 15.9644 145.02 0.000141176 0.267166 192.855 0.310526 0.067366 0.00409612 0.000561857 0.00138341 0.986981 0.991729 -2.97844e-06 -85.6643 0.0930173 31186.5 302.626 0.983513 0.319147 0.73235 0.732346 9.99958 2.9826e-06 1.19303e-05 0.131426 0.982406 0.931679 -0.0132927 4.90744e-06 0.504065 -1.91355e-20 7.0645e-24 -1.91285e-20 0.00139556 0.997817 8.596e-05 0.152612 2.85207 0.00139556 0.997821 0.724339 0.00105379 0.00188023 0.0008596 0.455563 0.00188023 0.439515 0.000129108 1.02 0.887907 0.534617 0.286367 1.71735e-07 3.06632e-09 2383.8 3114.8 -0.0553516 0.482149 0.277496 0.25321 -0.593387 -0.169524 0.496907 -0.267442 -0.229474 1.876 1 0 297.835 0 2.12236 1.874 0.000299799 0.853056 0.665071 0.368798 0.415779 2.12257 133.135 83.931 18.7215 60.8713 0.00402488 0 -40 10
0.975 2.82411e-08 2.53905e-06 0.111405 0.111403 0.0120371 1.28368e-05 0.00115411 0.139256 0.000658059 0.13991 0.887256 101.794 0.242708 0.758621 4.20641 0.0572917 0.0396831 0.960317 0.0197781 0.00431992 0.019041 0.00414849 0.00522192 0.00595901 0.208877 0.23836 58 -87.8962 126.26 15.9644 145.02 0.000141175 0.267166 192.855 0.310525 0.067366 0.00409612 0.000561858 0.00138341 0.986981 0.991729 -2.97845e-06 -85.6643 0.0930174 31186.5 302.633 0.983513 0.319147 0.732347 0.732342 9.99958 2.98261e-06 1.19303e-05 0.131428 0.98241 0.93168 -0.0132927 4.90747e-06 0.504076 -1.91365e-20 7.0649e-24 -1.91294e-20 0.00139557 0.997817 8.59601e-05 0.152612 2.85207 0.00139557 0.997821 0.724435 0.00105381 0.00188023 0.000859601 0.455563 0.00188023 0.439523 0.000129111 1.02 0.887908 0.534617 0.286369 1.71735e-07 3.06634e-09 2383.78 3114.79 -0.0553517 0.482149 0.277496 0.253209 -0.593388 -0.169524 0.496906 -0.26744 -0.229475 1.877 1 0 297.835 0 2.12251 1.875 0.000299798 0.853052 0.665119 0.368678 0.415805 2.12272 133.143 83.9312 18.7215 60.8714 0.00402487 0 -40 10
0.976 2.827e-08 2.53905e-06 0.111467 0.111465 0.012037 1.285e-05 0.00115411 0.139334 0.000658061 0.139987 0.887327 101.793 0.2427 0.758728 4.20669 0.0573002 0.0396857 0.960314 0.0197778 0.00432017 0.0190407 0.0041487 0.00522222 0.00595931 0.208889 0.238372 58.0001 -87.8962 126.26 15.9643 145.02 0.000141175 0.267167 192.855 0.310525 0.0673659 0.00409612 0.000561858 0.00138341 0.986981 0.991729 -2.97847e-06 -85.6643 0.0930175 31186.5 302.64 0.983513 0.319147 0.732343 0.732339 9.99958 2.98261e-06 1.19303e-05 0.131431 0.982413 0.931681 -0.0132927 4.9075e-06 0.504086 -1.91374e-20 7.06529e-24 -1.91304e-20 0.00139557 0.997817 8.59602e-05 0.152612 2.85207 0.00139557 0.997821 0.724531 0.00105383 0.00188023 0.000859602 0.455562 0.00188023 0.43953 0.000129114 1.02 0.887909 0.534616 0.28637 1.71735e-07 3.06636e-09 2383.77 3114.78 -0.0553519 0.482149 0.277496 0.253208 -0.593388 -0.169524 0.496904 -0.267438 -0.229476 1.878 1 0 297.835 0 2.12266 1.876 0.000299798 0.853048 0.665167 0.368558 0.41583 2.12287 133.151 83.9314 18.7215 60.8715 0.00402486 0 -40 10
0.977 2.82989e-08 2.53905e-06 0.111529 0.111527 0.012037 1.28631e-05 0.00115411 0.139411 0.000658062 0.140064 0.887398 101.793 0.242691 0.758835 4.20696 0.0573088 0.0396883 0.960312 0.0197775 0.00432041 0.0190404 0.00414891 0.00522252 0.00595961 0.208901 0.238385 58.0002 -87.8962 126.26 15.9643 145.02 0.000141174 0.267167 192.855 0.310524 0.0673658 0.00409613 0.000561859 0.00138341 0.986981 0.991729 -2.97848e-06 -85.6643 0.0930175 31186.5 302.646 0.983513 0.319147 0.73234 0.732336 9.99958 2.98262e-06 1.19304e-05 0.131433 0.982417 0.931682 -0.0132927 4.90753e-06 0.504096 -1.91384e-20 7.06569e-24 -1.91313e-20 0.00139557 0.997817 8.59603e-05 0.152613 2.85207 0.00139557 0.997821 0.724626 0.00105385 0.00188023 0.000859603 0.455562 0.00188023 0.439538 0.000129117 1.02 0.88791 0.534616 0.286372 1.71735e-07 3.06639e-09 2383.75 3114.76 -0.0553521 0.482149 0.277495 0.253208 -0.593388 -0.169524 0.496903 -0.267436 -0.229476 1.879 1 0 297.836 0 2.12282 1.877 0.000299797 0.853045 0.665215 0.368438 0.415855 2.12303 133.159 83.9315 18.7215 60.8716 0.00402486 0 -40 10
0.978 2.83278e-08 2.53905e-06 0.11159 0.111589 0.012037 1.28763e-05 0.00115411 0.139488 0.000658064 0.140141 0.88747 101.793 0.242683 0.758942 4.20724 0.0573173 0.0396909 0.960309 0.0197772 0.00432066 0.0190401 0.00414911 0.00522283 0.00595992 0.208913 0.238397 58.0002 -87.8962 126.26 15.9643 145.02 0.000141173 0.267167 192.854 0.310524 0.0673658 0.00409613 0.00056186 0.00138341 0.986981 0.991729 -2.9785e-06 -85.6643 0.0930176 31186.4 302.653 0.983513 0.319147 0.732337 0.732333 9.99958 2.98262e-06 1.19304e-05 0.131436 0.98242 0.931682 -0.0132927 4.90756e-06 0.504107 -1.91394e-20 7.06609e-24 -1.91323e-20 0.00139557 0.997817 8.59603e-05 0.152613 2.85207 0.00139557 0.997821 0.724722 0.00105387 0.00188024 0.000859603 0.455562 0.00188023 0.439546 0.00012912 1.02 0.887911 0.534616 0.286373 1.71736e-07 3.06641e-09 2383.73 3114.75 -0.0553523 0.482149 0.277495 0.253207 -0.593388 -0.169524 0.496901 -0.267434 -0.229477 1.88 1 0 297.836 0 2.12297 1.878 0.000299797 0.853041 0.665263 0.368318 0.415881 2.12318 133.167 83.9317 18.7215 60.8717 0.00402485 0 -40 10
0.979 2.83567e-08 2.53905e-06 0.111652 0.11165 0.012037 1.28894e-05 0.00115411 0.139565 0.000658066 0.140218 0.887541 101.792 0.242674 0.759049 4.20751 0.0573259 0.0396935 0.960306 0.0197769 0.0043209 0.0190398 0.00414932 0.00522313 0.00596022 0.208925 0.238409 58.0003 -87.8962 126.26 15.9642 145.02 0.000141173 0.267167 192.854 0.310524 0.0673657 0.00409613 0.00056186 0.00138342 0.986981 0.991729 -2.97851e-06 -85.6643 0.0930177 31186.4 302.66 0.983513 0.319147 0.732334 0.73233 9.99958 2.98263e-06 1.19304e-05 0.131438 0.982424 0.931683 -0.0132927 4.90759e-06 0.504117 -1.91403e-20 7.06649e-24 -1.91333e-20 0.00139557 0.997817 8.59604e-05 0.152613 2.85208 0.00139557 0.997821 0.724818 0.00105388 0.00188024 0.000859604 0.455562 0.00188024 0.439553 0.000129123 1.02 0.887912 0.534615 0.286375 1.71736e-07 3.06643e-09 2383.72 3114.73 -0.0553525 0.482149 0.277495 0.253206 -0.593388 -0.169524 0.4969 -0.267432 -0.229477 1.881 1 0 297.836 0 2.12312 1.879 0.000299796 0.853038 0.665311 0.368199 0.415906 2.12333 133.176 83.9318 18.7215 60.8717 0.00402484 0 -40 10
0.98 2.83856e-08 2.53905e-06 0.111713 0.111712 0.012037 1.29026e-05 0.00115411 0.139642 0.000658067 0.140295 0.887612 101.792 0.242666 0.759157 4.20779 0.0573345 0.0396961 0.960304 0.0197766 0.00432115 0.0190395 0.00414953 0.00522343 0.00596052 0.208937 0.238421 58.0003 -87.8962 126.26 15.9642 145.02 0.000141172 0.267167 192.854 0.310523 0.0673657 0.00409614 0.000561861 0.00138342 0.986981 0.991729 -2.97853e-06 -85.6643 0.0930178 31186.4 302.666 0.983513 0.319147 0.732331 0.732327 9.99958 2.98263e-06 1.19304e-05 0.131441 0.982427 0.931684 -0.0132927 4.90762e-06 0.504127 -1.91413e-20 7.06689e-24 -1.91342e-20 0.00139557 0.997817 8.59605e-05 0.152613 2.85208 0.00139557 0.997821 0.724914 0.0010539 0.00188024 0.000859605 0.455561 0.00188024 0.439561 0.000129126 1.02 0.887914 0.534615 0.286376 1.71736e-07 3.06645e-09 2383.7 3114.72 -0.0553528 0.482149 0.277495 0.253205 -0.593388 -0.169524 0.496898 -0.26743 -0.229478 1.882 1 0 297.836 0 2.12328 1.88 0.000299796 0.853035 0.665359 0.36808 0.415932 2.12349 133.184 83.932 18.7216 60.8718 0.00402484 0 -40 10
0.981 2.84146e-08 2.53905e-06 0.111775 0.111773 0.012037 1.29157e-05 0.00115411 0.139719 0.000658069 0.140372 0.887684 101.792 0.242657 0.759264 4.20806 0.057343 0.0396987 0.960301 0.0197763 0.00432139 0.0190392 0.00414973 0.00522373 0.00596082 0.208949 0.238433 58.0004 -87.8962 126.26 15.9642 145.02 0.000141172 0.267168 192.854 0.310523 0.0673656 0.00409614 0.000561862 0.00138342 0.986981 0.991729 -2.97854e-06 -85.6643 0.0930179 31186.4 302.673 0.983513 0.319147 0.732328 0.732324 9.99958 2.98264e-06 1.19304e-05 0.131443 0.98243 0.931685 -0.0132927 4.90765e-06 0.504138 -1.91423e-20 7.06729e-24 -1.91352e-20 0.00139557 0.997817 8.59606e-05 0.152613 2.85208 0.00139557 0.997821 0.725009 0.00105392 0.00188024 0.000859606 0.455561 0.00188024 0.439568 0.000129129 1.02 0.887915 0.534615 0.286378 1.71737e-07 3.06648e-09 2383.68 3114.71 -0.055353 0.48215 0.277494 0.253204 -0.593388 -0.169524 0.496896 -0.267428 -0.229478 1.883 1 0 297.836 0 2.12343 1.881 0.000299795 0.853031 0.665407 0.367961 0.415957 2.12364 133.192 83.9321 18.7216 60.8719 0.00402483 0 -40 10
0.982 2.84435e-08 2.53905e-06 0.111836 0.111835 0.012037 1.29289e-05 0.00115412 0.139796 0.000658071 0.140449 0.887755 101.792 0.242648 0.759371 4.20834 0.0573516 0.0397013 0.960299 0.019776 0.00432164 0.0190389 0.00414994 0.00522403 0.00596113 0.208961 0.238445 58.0005 -87.8962 126.26 15.9641 145.02 0.000141171 0.267168 192.854 0.310522 0.0673656 0.00409614 0.000561862 0.00138342 0.986981 0.991729 -2.97856e-06 -85.6643 0.093018 31186.4 302.68 0.983513 0.319147 0.732325 0.732321 9.99958 2.98264e-06 1.19305e-05 0.131446 0.982434 0.931686 -0.0132927 4.90768e-06 0.504148 -1.91432e-20 7.06769e-24 -1.91362e-20 0.00139557 0.997817 8.59607e-05 0.152613 2.85208 0.00139557 0.997821 0.725105 0.00105394 0.00188024 0.000859607 0.455561 0.00188024 0.439576 0.000129132 1.02 0.887916 0.534614 0.286379 1.71737e-07 3.0665e-09 2383.67 3114.69 -0.0553533 0.48215 0.277494 0.253203 -0.593389 -0.169524 0.496895 -0.267425 -0.229478 1.884 1 0 297.836 0 2.12358 1.882 0.000299794 0.853028 0.665455 0.367842 0.415983 2.12379 133.2 83.9323 18.7216 60.8719 0.00402482 0 -40 10
0.983 2.84724e-08 2.53905e-06 0.111898 0.111896 0.0120369 1.2942e-05 0.00115412 0.139872 0.000658073 0.140526 0.887827 101.791 0.24264 0.759479 4.20862 0.0573602 0.0397039 0.960296 0.0197757 0.00432189 0.0190386 0.00415015 0.00522434 0.00596143 0.208973 0.238457 58.0005 -87.8963 126.26 15.9641 145.02 0.000141171 0.267168 192.854 0.310522 0.0673655 0.00409615 0.000561863 0.00138342 0.986981 0.991729 -2.97857e-06 -85.6643 0.0930181 31186.3 302.686 0.983513 0.319147 0.732322 0.732318 9.99958 2.98265e-06 1.19305e-05 0.131448 0.982437 0.931687 -0.0132927 4.90771e-06 0.504159 -1.91442e-20 7.0681e-24 -1.91371e-20 0.00139557 0.997817 8.59607e-05 0.152614 2.85208 0.00139557 0.997821 0.7252 0.00105396 0.00188024 0.000859607 0.455561 0.00188024 0.439584 0.000129135 1.02 0.887917 0.534614 0.286381 1.71737e-07 3.06652e-09 2383.65 3114.68 -0.0553536 0.48215 0.277494 0.253203 -0.593389 -0.169524 0.496893 -0.267423 -0.229479 1.885 1 0 297.836 0 2.12374 1.883 0.000299794 0.853025 0.665503 0.367724 0.416008 2.12395 133.208 83.9324 18.7216 60.872 0.00402482 0 -40 10
0.984 2.85013e-08 2.53905e-06 0.111959 0.111958 0.0120369 1.29551e-05 0.00115412 0.139949 0.000658074 0.140603 0.887899 101.791 0.242631 0.759586 4.20889 0.0573688 0.0397065 0.960293 0.0197754 0.00432213 0.0190383 0.00415035 0.00522464 0.00596173 0.208986 0.238469 58.0006 -87.8963 126.26 15.964 145.02 0.00014117 0.267168 192.853 0.310521 0.0673655 0.00409615 0.000561864 0.00138343 0.986981 0.991729 -2.97859e-06 -85.6643 0.0930182 31186.3 302.693 0.983513 0.319147 0.732319 0.732315 9.99958 2.98265e-06 1.19305e-05 0.131451 0.982441 0.931687 -0.0132927 4.90774e-06 0.504169 -1.91452e-20 7.0685e-24 -1.91381e-20 0.00139558 0.997817 8.59608e-05 0.152614 2.85208 0.00139558 0.997821 0.725296 0.00105398 0.00188024 0.000859608 0.455561 0.00188024 0.439591 0.000129139 1.02 0.887918 0.534614 0.286382 1.71737e-07 3.06655e-09 2383.63 3114.67 -0.0553539 0.48215 0.277493 0.253202 -0.593389 -0.169525 0.496891 -0.267421 -0.229479 1.886 1 0 297.837 0 2.12389 1.884 0.000299793 0.853022 0.665551 0.367606 0.416034 2.1241 133.217 83.9325 18.7216 60.8721 0.00402481 0 -40 10
0.985 2.85302e-08 2.53906e-06 0.112021 0.112019 0.0120369 1.29683e-05 0.00115412 0.140026 0.000658076 0.140679 0.88797 101.791 0.242623 0.759694 4.20917 0.0573774 0.0397092 0.960291 0.0197751 0.00432238 0.019038 0.00415056 0.00522494 0.00596204 0.208998 0.238482 58.0007 -87.8963 126.26 15.964 145.02 0.000141169 0.267168 192.853 0.310521 0.0673654 0.00409615 0.000561864 0.00138343 0.986981 0.991729 -2.9786e-06 -85.6642 0.0930182 31186.3 302.7 0.983513 0.319147 0.732317 0.732312 9.99958 2.98266e-06 1.19305e-05 0.131453 0.982444 0.931688 -0.0132927 4.90777e-06 0.504179 -1.91461e-20 7.0689e-24 -1.91391e-20 0.00139558 0.997817 8.59609e-05 0.152614 2.85208 0.00139558 0.997821 0.725392 0.001054 0.00188025 0.000859609 0.45556 0.00188024 0.439599 0.000129142 1.02 0.887919 0.534614 0.286384 1.71738e-07 3.06657e-09 2383.62 3114.65 -0.0553542 0.48215 0.277493 0.253201 -0.593389 -0.169525 0.496889 -0.267419 -0.229479 1.887 1 0 297.837 0 2.12404 1.885 0.000299793 0.85302 0.665599 0.367488 0.416059 2.12425 133.225 83.9327 18.7216 60.8721 0.00402481 0 -40 10
0.986 2.85592e-08 2.53906e-06 0.112082 0.11208 0.0120369 1.29814e-05 0.00115412 0.140102 0.000658078 0.140756 0.888042 101.791 0.242614 0.759802 4.20945 0.057386 0.0397118 0.960288 0.0197748 0.00432263 0.0190377 0.00415077 0.00522525 0.00596234 0.20901 0.238494 58.0007 -87.8963 126.26 15.964 145.02 0.000141169 0.267169 192.853 0.310521 0.0673654 0.00409615 0.000561865 0.00138343 0.986981 0.991729 -2.97862e-06 -85.6642 0.0930183 31186.3 302.706 0.983513 0.319147 0.732314 0.732309 9.99958 2.98266e-06 1.19305e-05 0.131456 0.982447 0.931689 -0.0132927 4.9078e-06 0.50419 -1.91471e-20 7.0693e-24 -1.914e-20 0.00139558 0.997817 8.5961e-05 0.152614 2.85208 0.00139558 0.997821 0.725487 0.00105402 0.00188025 0.00085961 0.45556 0.00188025 0.439606 0.000129145 1.02 0.88792 0.534613 0.286385 1.71738e-07 3.06659e-09 2383.6 3114.64 -0.0553545 0.48215 0.277493 0.2532 -0.593389 -0.169525 0.496887 -0.267417 -0.229479 1.888 1 0 297.837 0 2.12419 1.886 0.000299792 0.853017 0.665647 0.36737 0.416084 2.1244 133.233 83.9328 18.7216 60.8722 0.0040248 0 -40 10
0.987 2.85881e-08 2.53906e-06 0.112143 0.112141 0.0120369 1.29946e-05 0.00115412 0.140179 0.000658079 0.140832 0.888114 101.79 0.242605 0.759909 4.20973 0.0573946 0.0397144 0.960286 0.0197744 0.00432288 0.0190373 0.00415098 0.00522555 0.00596265 0.209022 0.238506 58.0008 -87.8963 126.26 15.9639 145.02 0.000141168 0.267169 192.853 0.31052 0.0673653 0.00409616 0.000561866 0.00138343 0.986981 0.991729 -2.97863e-06 -85.6642 0.0930184 31186.2 302.713 0.983513 0.319147 0.732311 0.732307 9.99958 2.98266e-06 1.19306e-05 0.131458 0.982451 0.93169 -0.0132927 4.90782e-06 0.5042 -1.91481e-20 7.0697e-24 -1.9141e-20 0.00139558 0.997817 8.59611e-05 0.152614 2.85208 0.00139558 0.997821 0.725583 0.00105404 0.00188025 0.000859611 0.45556 0.00188025 0.439614 0.000129148 1.02 0.887921 0.534613 0.286387 1.71738e-07 3.06661e-09 2383.58 3114.63 -0.0553549 0.48215 0.277493 0.2532 -0.593389 -0.169525 0.496885 -0.267415 -0.22948 1.889 1 0 297.837 0 2.12435 1.887 0.000299792 0.853014 0.665695 0.367252 0.41611 2.12456 133.241 83.933 18.7216 60.8723 0.0040248 0 -40 10
0.988 2.8617e-08 2.53906e-06 0.112204 0.112203 0.0120369 1.30077e-05 0.00115412 0.140255 0.000658081 0.140909 0.888185 101.79 0.242597 0.760017 4.21001 0.0574032 0.039717 0.960283 0.0197741 0.00432312 0.019037 0.00415119 0.00522586 0.00596296 0.209034 0.238518 58.0009 -87.8963 126.261 15.9639 145.02 0.000141168 0.267169 192.853 0.31052 0.0673653 0.00409616 0.000561866 0.00138344 0.986981 0.991729 -2.97865e-06 -85.6642 0.0930185 31186.2 302.72 0.983513 0.319147 0.732309 0.732304 9.99958 2.98267e-06 1.19306e-05 0.131461 0.982454 0.931691 -0.0132927 4.90785e-06 0.504211 -1.91491e-20 7.0701e-24 -1.9142e-20 0.00139558 0.997817 8.59611e-05 0.152614 2.85208 0.00139558 0.997821 0.725678 0.00105405 0.00188025 0.000859611 0.45556 0.00188025 0.439622 0.000129151 1.02 0.887922 0.534613 0.286388 1.71738e-07 3.06664e-09 2383.57 3114.62 -0.0553553 0.48215 0.277492 0.253199 -0.593389 -0.169525 0.496883 -0.267413 -0.22948 1.89 1 0 297.837 0 2.1245 1.888 0.000299791 0.853012 0.665742 0.367135 0.416135 2.12471 133.249 83.9331 18.7216 60.8723 0.00402479 0 -40 10
0.989 2.86459e-08 2.53906e-06 0.112265 0.112264 0.0120369 1.30209e-05 0.00115412 0.140332 0.000658083 0.140985 0.888257 101.79 0.242588 0.760125 4.21029 0.0574118 0.0397197 0.96028 0.0197738 0.00432337 0.0190367 0.0041514 0.00522616 0.00596326 0.209047 0.23853 58.0009 -87.8963 126.261 15.9638 145.02 0.000141167 0.267169 192.853 0.310519 0.0673652 0.00409616 0.000561867 0.00138344 0.98698 0.991729 -2.97866e-06 -85.6642 0.0930186 31186.2 302.727 0.983513 0.319147 0.732306 0.732302 9.99958 2.98267e-06 1.19306e-05 0.131463 0.982457 0.931691 -0.0132927 4.90788e-06 0.504221 -1.915e-20 7.07051e-24 -1.9143e-20 0.00139558 0.997817 8.59612e-05 0.152614 2.85208 0.00139558 0.997821 0.725773 0.00105407 0.00188025 0.000859612 0.455559 0.00188025 0.439629 0.000129154 1.02 0.887923 0.534612 0.28639 1.71739e-07 3.06666e-09 2383.55 3114.61 -0.0553556 0.48215 0.277492 0.253198 -0.593389 -0.169525 0.496881 -0.267411 -0.22948 1.891 1 0 297.837 0 2.12465 1.889 0.000299791 0.853009 0.66579 0.367018 0.416161 2.12486 133.258 83.9332 18.7216 60.8724 0.00402479 0 -40 10
0.99 2.86748e-08 2.53906e-06 0.112326 0.112325 0.0120368 1.3034e-05 0.00115412 0.140408 0.000658084 0.141062 0.888329 101.789 0.24258 0.760233 4.21057 0.0574204 0.0397223 0.960278 0.0197735 0.00432362 0.0190364 0.00415161 0.00522647 0.00596357 0.209059 0.238543 58.001 -87.8963 126.261 15.9638 145.02 0.000141167 0.267169 192.852 0.310519 0.0673652 0.00409617 0.000561868 0.00138344 0.98698 0.991729 -2.97868e-06 -85.6642 0.0930187 31186.2 302.733 0.983513 0.319147 0.732303 0.732299 9.99958 2.98268e-06 1.19306e-05 0.131466 0.98246 0.931692 -0.0132927 4.90791e-06 0.504232 -1.9151e-20 7.07091e-24 -1.91439e-20 0.00139558 0.997817 8.59613e-05 0.152615 2.85209 0.00139558 0.997821 0.725869 0.00105409 0.00188025 0.000859613 0.455559 0.00188025 0.439637 0.000129157 1.02 0.887924 0.534612 0.286391 1.71739e-07 3.06668e-09 2383.53 3114.59 -0.055356 0.48215 0.277492 0.253198 -0.593389 -0.169525 0.496879 -0.267409 -0.22948 1.892 1 0 297.837 0 2.12481 1.89 0.00029979 0.853007 0.665838 0.366901 0.416186 2.12501 133.266 83.9333 18.7216 60.8725 0.00402478 0 -40 10
0.991 2.87037e-08 2.53906e-06 0.112387 0.112386 0.0120368 1.30472e-05 0.00115412 0.140484 0.000658086 0.141138 0.888401 101.789 0.242571 0.760341 4.21085 0.057429 0.039725 0.960275 0.0197732 0.00432387 0.0190361 0.00415182 0.00522677 0.00596388 0.209071 0.238555 58.001 -87.8963 126.261 15.9638 145.02 0.000141166 0.26717 192.852 0.310518 0.0673651 0.00409617 0.000561868 0.00138344 0.98698 0.991729 -2.97869e-06 -85.6642 0.0930188 31186.2 302.74 0.983513 0.319147 0.732301 0.732297 9.99958 2.98268e-06 1.19306e-05 0.131468 0.982464 0.931693 -0.0132927 4.90794e-06 0.504242 -1.9152e-20 7.07131e-24 -1.91449e-20 0.00139558 0.997817 8.59614e-05 0.152615 2.85209 0.00139558 0.997821 0.725964 0.00105411 0.00188025 0.000859614 0.455559 0.00188025 0.439644 0.00012916 1.02 0.887926 0.534612 0.286393 1.71739e-07 3.06671e-09 2383.52 3114.58 -0.0553565 0.48215 0.277491 0.253197 -0.59339 -0.169525 0.496877 -0.267407 -0.22948 1.893 1 0 297.837 0 2.12496 1.891 0.00029979 0.853005 0.665886 0.366785 0.416211 2.12517 133.274 83.9335 18.7216 60.8725 0.00402478 0 -40 10
0.992 2.87327e-08 2.53906e-06 0.112448 0.112447 0.0120368 1.30603e-05 0.00115412 0.140561 0.000658088 0.141214 0.888473 101.789 0.242562 0.760448 4.21113 0.0574376 0.0397276 0.960272 0.0197729 0.00432412 0.0190358 0.00415203 0.00522708 0.00596418 0.209083 0.238567 58.0011 -87.8963 126.261 15.9637 145.02 0.000141166 0.26717 192.852 0.310518 0.0673651 0.00409617 0.000561869 0.00138344 0.98698 0.991729 -2.97871e-06 -85.6642 0.0930188 31186.1 302.747 0.983513 0.319147 0.732298 0.732294 9.99958 2.98269e-06 1.19307e-05 0.131471 0.982467 0.931694 -0.0132927 4.90797e-06 0.504253 -1.9153e-20 7.07172e-24 -1.91459e-20 0.00139558 0.997817 8.59615e-05 0.152615 2.85209 0.00139558 0.997821 0.726059 0.00105413 0.00188026 0.000859615 0.455559 0.00188026 0.439652 0.000129163 1.02 0.887927 0.534611 0.286394 1.71739e-07 3.06673e-09 2383.5 3114.57 -0.0553569 0.48215 0.277491 0.253196 -0.59339 -0.169525 0.496875 -0.267404 -0.22948 1.894 1 0 297.837 0 2.12511 1.892 0.000299789 0.853003 0.665934 0.366669 0.416237 2.12532 133.282 83.9336 18.7216 60.8726 0.00402477 0 -40 10
0.993 2.87616e-08 2.53906e-06 0.112509 0.112508 0.0120368 1.30734e-05 0.00115412 0.140637 0.000658089 0.14129 0.888545 101.789 0.242554 0.760557 4.21141 0.0574463 0.0397303 0.96027 0.0197726 0.00432437 0.0190355 0.00415224 0.00522739 0.00596449 0.209096 0.23858 58.0012 -87.8963 126.261 15.9637 145.02 0.000141166 0.26717 192.852 0.310518 0.067365 0.00409618 0.00056187 0.00138345 0.98698 0.991729 -2.97872e-06 -85.6642 0.0930189 31186.1 302.754 0.983513 0.319147 0.732296 0.732292 9.99958 2.98269e-06 1.19307e-05 0.131473 0.98247 0.931694 -0.0132927 4.908e-06 0.504263 -1.91539e-20 7.07212e-24 -1.91469e-20 0.00139559 0.997817 8.59615e-05 0.152615 2.85209 0.00139559 0.997821 0.726155 0.00105415 0.00188026 0.000859615 0.455559 0.00188026 0.43966 0.000129166 1.02 0.887928 0.534611 0.286396 1.7174e-07 3.06675e-09 2383.48 3114.56 -0.0553573 0.48215 0.277491 0.253196 -0.59339 -0.169525 0.496872 -0.267402 -0.229479 1.895 1 0 297.837 0 2.12526 1.893 0.000299788 0.853001 0.665981 0.366553 0.416262 2.12547 133.29 83.9337 18.7217 60.8726 0.00402477 0 -40 10
0.994 2.87905e-08 2.53906e-06 0.11257 0.112569 0.0120368 1.30866e-05 0.00115412 0.140713 0.000658091 0.141366 0.888617 101.788 0.242545 0.760665 4.21169 0.0574549 0.0397329 0.960267 0.0197723 0.00432462 0.0190352 0.00415245 0.0052277 0.0059648 0.209108 0.238592 58.0012 -87.8963 126.261 15.9637 145.02 0.000141165 0.26717 192.852 0.310517 0.067365 0.00409618 0.00056187 0.00138345 0.98698 0.991729 -2.97874e-06 -85.6642 0.093019 31186.1 302.76 0.983513 0.319147 0.732294 0.732289 9.99958 2.9827e-06 1.19307e-05 0.131476 0.982474 0.931695 -0.0132927 4.90803e-06 0.504274 -1.91549e-20 7.07252e-24 -1.91478e-20 0.00139559 0.997817 8.59616e-05 0.152615 2.85209 0.00139559 0.997821 0.72625 0.00105417 0.00188026 0.000859616 0.455558 0.00188026 0.439667 0.000129169 1.02 0.887929 0.534611 0.286398 1.7174e-07 3.06677e-09 2383.47 3114.55 -0.0553578 0.482151 0.277491 0.253195 -0.59339 -0.169525 0.49687 -0.2674 -0.229479 1.896 1 0 297.837 0 2.12542 1.894 0.000299788 0.852999 0.666029 0.366437 0.416287 2.12563 133.298 83.9338 18.7217 60.8727 0.00402476 0 -40 10
0.995 2.88194e-08 2.53906e-06 0.112631 0.112629 0.0120368 1.30997e-05 0.00115412 0.140789 0.000658093 0.141442 0.888688 101.788 0.242536 0.760773 4.21197 0.0574635 0.0397356 0.960264 0.019772 0.00432487 0.0190349 0.00415266 0.005228 0.00596511 0.20912 0.238604 58.0013 -87.8963 126.261 15.9636 145.02 0.000141165 0.26717 192.852 0.310517 0.0673649 0.00409618 0.000561871 0.00138345 0.98698 0.991729 -2.97875e-06 -85.6641 0.0930191 31186.1 302.767 0.983513 0.319147 0.732291 0.732287 9.99958 2.9827e-06 1.19307e-05 0.131479 0.982477 0.931696 -0.0132927 4.90806e-06 0.504285 -1.91559e-20 7.07293e-24 -1.91488e-20 0.00139559 0.997817 8.59617e-05 0.152615 2.85209 0.00139559 0.997821 0.726345 0.00105419 0.00188026 0.000859617 0.455558 0.00188026 0.439675 0.000129173 1.02 0.88793 0.534611 0.286399 1.7174e-07 3.0668e-09 2383.45 3114.54 -0.0553583 0.482151 0.27749 0.253194 -0.59339 -0.169525 0.496868 -0.267398 -0.229479 1.897 1 0 297.836 0 2.12557 1.895 0.000299787 0.852997 0.666077 0.366321 0.416313 2.12578 133.307 83.9339 18.7217 60.8727 0.00402476 0 -40 10
0.996 2.88483e-08 2.53906e-06 0.112692 0.11269 0.0120368 1.31129e-05 0.00115412 0.140865 0.000658094 0.141518 0.888761 101.788 0.242528 0.760881 4.21225 0.0574722 0.0397382 0.960262 0.0197717 0.00432512 0.0190346 0.00415287 0.00522831 0.00596542 0.209132 0.238617 58.0014 -87.8963 126.261 15.9636 145.02 0.000141164 0.26717 192.851 0.310516 0.0673649 0.00409618 0.000561872 0.00138345 0.98698 0.991729 -2.97877e-06 -85.6641 0.0930192 31186 302.774 0.983513 0.319147 0.732289 0.732285 9.99958 2.98271e-06 1.19307e-05 0.131481 0.98248 0.931697 -0.0132927 4.90809e-06 0.504295 -1.91569e-20 7.07333e-24 -1.91498e-20 0.00139559 0.997817 8.59618e-05 0.152615 2.85209 0.00139559 0.997821 0.72644 0.0010542 0.00188026 0.000859618 0.455558 0.00188026 0.439682 0.000129176 1.02 0.887931 0.53461 0.286401 1.71741e-07 3.06682e-09 2383.43 3114.53 -0.0553588 0.482151 0.27749 0.253194 -0.59339 -0.169525 0.496865 -0.267396 -0.229479 1.898 1 0 297.836 0 2.12572 1.896 0.000299787 0.852995 0.666125 0.366206 0.416338 2.12593 133.315 83.934 18.7217 60.8728 0.00402475 0 -40 10
0.997 2.88772e-08 2.53906e-06 0.112753 0.112751 0.0120368 1.3126e-05 0.00115412 0.140941 0.000658096 0.141594 0.888833 101.787 0.242519 0.760989 4.21254 0.0574808 0.0397409 0.960259 0.0197714 0.00432537 0.0190343 0.00415308 0.00522862 0.00596573 0.209145 0.238629 58.0014 -87.8963 126.261 15.9635 145.02 0.000141164 0.267171 192.851 0.310516 0.0673648 0.00409619 0.000561872 0.00138345 0.98698 0.991728 -2.97878e-06 -85.6641 0.0930193 31186 302.781 0.983513 0.319147 0.732287 0.732283 9.99958 2.98271e-06 1.19307e-05 0.131484 0.982483 0.931697 -0.0132927 4.90812e-06 0.504306 -1.91578e-20 7.07374e-24 -1.91508e-20 0.00139559 0.997817 8.59619e-05 0.152616 2.85209 0.00139559 0.997821 0.726535 0.00105422 0.00188026 0.000859619 0.455558 0.00188026 0.43969 0.000129179 1.02 0.887932 0.53461 0.286402 1.71741e-07 3.06684e-09 2383.42 3114.52 -0.0553593 0.482151 0.27749 0.253193 -0.59339 -0.169525 0.496863 -0.267394 -0.229478 1.899 1 0 297.836 0 2.12587 1.897 0.000299786 0.852994 0.666173 0.366091 0.416363 2.12608 133.323 83.9341 18.7217 60.8728 0.00402475 0 -40 10
0.998 2.89062e-08 2.53906e-06 0.112813 0.112812 0.0120367 1.31392e-05 0.00115412 0.141017 0.000658098 0.14167 0.888905 101.787 0.242511 0.761097 4.21282 0.0574895 0.0397436 0.960256 0.0197711 0.00432562 0.019034 0.00415329 0.00522893 0.00596604 0.209157 0.238641 58.0015 -87.8963 126.261 15.9635 145.02 0.000141163 0.267171 192.851 0.310515 0.0673648 0.00409619 0.000561873 0.00138346 0.98698 0.991728 -2.9788e-06 -85.6641 0.0930194 31186 302.787 0.983513 0.319147 0.732285 0.732281 9.99958 2.98272e-06 1.19308e-05 0.131486 0.982487 0.931698 -0.0132927 4.90815e-06 0.504316 -1.91588e-20 7.07414e-24 -1.91518e-20 0.00139559 0.997817 8.59619e-05 0.152616 2.85209 0.00139559 0.997821 0.72663 0.00105424 0.00188027 0.000859619 0.455557 0.00188026 0.439697 0.000129182 1.02 0.887933 0.53461 0.286404 1.71741e-07 3.06686e-09 2383.4 3114.51 -0.0553598 0.482151 0.277489 0.253193 -0.59339 -0.169525 0.49686 -0.267392 -0.229478 1.9 1 0 297.836 0 2.12603 1.898 0.000299786 0.852992 0.66622 0.365976 0.416389 2.12623 133.331 83.9343 18.7217 60.8729 0.00402474 0 -40 10
0.999 2.89351e-08 2.53906e-06 0.112874 0.112872 0.0120367 1.31523e-05 0.00115412 0.141092 0.000658099 0.141746 0.888977 101.787 0.242502 0.761206 4.2131 0.0574981 0.0397463 0.960254 0.0197708 0.00432587 0.0190337 0.0041535 0.00522924 0.00596635 0.209169 0.238654 58.0016 -87.8963 126.261 15.9635 145.02 0.000141163 0.267171 192.851 0.310515 0.0673647 0.00409619 0.000561874 0.00138346 0.98698 0.991728 -2.97881e-06 -85.6641 0.0930195 31186 302.794 0.983513 0.319147 0.732283 0.732278 9.99958 2.98272e-06 1.19308e-05 0.131489 0.98249 0.931699 -0.0132927 4.90818e-06 0.504327 -1.91598e-20 7.07455e-24 -1.91527e-20 0.00139559 0.997817 8.5962e-05 0.152616 2.85209 0.00139559 0.997821 0.726726 0.00105426 0.00188027 0.00085962 0.455557 0.00188027 0.439705 0.000129185 1.02 0.887934 0.534609 0.286405 1.71741e-07 3.06689e-09 2383.38 3114.5 -0.0553604 0.482151 0.277489 0.253192 -0.59339 -0.169525 0.496858 -0.26739 -0.229477 1.901 1 0 297.836 0 2.12618 1.899 0.000299785 0.852991 0.666268 0.365861 0.416414 2.12639 133.339 83.9344 18.7217 60.8729 0.00402474 0 -40 10
1 2.8964e-08 2.53907e-06 0.112935 0.112933 0.0120367 1.31655e-05 0.00115412 0.141168 0.000658101 0.141822 0.889049 101.787 0.242493 0.761314 4.21339 0.0575068 0.0397489 0.960251 0.0197705 0.00432612 0.0190333 0.00415371 0.00522955 0.00596666 0.209182 0.238666 58.0016 -87.8963 126.261 15.9634 145.021 0.000141163 0.267171 192.851 0.310515 0.0673646 0.0040962 0.000561874 0.00138346 0.98698 0.991728 -2.97883e-06 -85.6641 0.0930195 31186 302.801 0.983513 0.319147 0.732281 0.732276 9.99958 2.98273e-06 1.19308e-05 0.131491 0.982493 0.9317 -0.0132927 4.90821e-06 0.504338 -1.91608e-20 7.07495e-24 -1.91537e-20 0.00139559 0.997817 8.59621e-05 0.152616 2.85209 0.00139559 0.99782 0.726821 0.00105428 0.00188027 0.000859621 0.455557 0.00188027 0.439712 0.000129188 1.02 0.887935 0.534609 0.286407 1.71742e-07 3.06691e-09 2383.37 3114.49 -0.0553609 0.482151 0.277489 0.253192 -0.59339 -0.169526 0.496855 -0.267388 -0.229477 1.902 1 0 297.836 0 2.12633 1.9 0.000299785 0.852989 0.666316 0.365747 0.416439 2.12654 133.347 83.9345 18.7217 60.873 0.00402473 0 -40 10
1.001 2.89929e-08 2.53907e-06 0.112995 0.112993 0.0120367 1.31786e-05 0.00115412 0.141244 0.000658103 0.141897 0.889121 101.786 0.242485 0.761423 4.21367 0.0575155 0.0397516 0.960248 0.0197701 0.00432638 0.019033 0.00415393 0.00522986 0.00596697 0.209194 0.238679 58.0017 -87.8963 126.261 15.9634 145.021 0.000141162 0.267171 192.851 0.310514 0.0673646 0.0040962 0.000561875 0.00138346 0.98698 0.991728 -2.97884e-06 -85.6641 0.0930196 31185.9 302.808 0.983513 0.319147 0.732279 0.732274 9.99958 2.98273e-06 1.19308e-05 0.131494 0.982496 0.9317 -0.0132927 4.90824e-06 0.504348 -1.91618e-20 7.07536e-24 -1.91547e-20 0.00139559 0.997817 8.59622e-05 0.152616 2.8521 0.00139559 0.99782 0.726916 0.0010543 0.00188027 0.000859622 0.455557 0.00188027 0.43972 0.000129191 1.02 0.887937 0.534609 0.286408 1.71742e-07 3.06693e-09 2383.35 3114.48 -0.0553615 0.482151 0.277489 0.253191 -0.59339 -0.169526 0.496852 -0.267385 -0.229476 1.903 1 0 297.836 0 2.12648 1.901 0.000299784 0.852988 0.666363 0.365632 0.416465 2.12669 133.356 83.9346 18.7217 60.873 0.00402473 0 -40 10
1.002 2.90218e-08 2.53907e-06 0.113056 0.113054 0.0120367 1.31917e-05 0.00115412 0.141319 0.000658104 0.141973 0.889193 101.786 0.242476 0.761531 4.21396 0.0575241 0.0397543 0.960246 0.0197698 0.00432663 0.0190327 0.00415414 0.00523017 0.00596728 0.209207 0.238691 58.0017 -87.8963 126.261 15.9634 145.021 0.000141162 0.267172 192.851 0.310514 0.0673645 0.0040962 0.000561876 0.00138347 0.98698 0.991728 -2.97886e-06 -85.6641 0.0930197 31185.9 302.815 0.983513 0.319147 0.732277 0.732272 9.99958 2.98274e-06 1.19308e-05 0.131497 0.982499 0.931701 -0.0132927 4.90827e-06 0.504359 -1.91627e-20 7.07576e-24 -1.91557e-20 0.0013956 0.997817 8.59623e-05 0.152616 2.8521 0.0013956 0.99782 0.727011 0.00105432 0.00188027 0.000859623 0.455557 0.00188027 0.439728 0.000129194 1.02 0.887938 0.534608 0.28641 1.71742e-07 3.06696e-09 2383.33 3114.47 -0.0553621 0.482151 0.277488 0.25319 -0.59339 -0.169526 0.49685 -0.267383 -0.229476 1.904 1 0 297.835 0 2.12664 1.902 0.000299784 0.852987 0.666411 0.365518 0.41649 2.12684 133.364 83.9347 18.7217 60.8731 0.00402473 0 -40 10
1.003 2.90507e-08 2.53907e-06 0.113116 0.113114 0.0120367 1.32049e-05 0.00115412 0.141395 0.000658106 0.142049 0.889266 101.786 0.242467 0.76164 4.21424 0.0575328 0.039757 0.960243 0.0197695 0.00432688 0.0190324 0.00415435 0.00523048 0.00596759 0.209219 0.238704 58.0018 -87.8963 126.261 15.9633 145.021 0.000141161 0.267172 192.85 0.310513 0.0673645 0.00409621 0.000561876 0.00138347 0.98698 0.991728 -2.97887e-06 -85.6641 0.0930198 31185.9 302.822 0.983513 0.319147 0.732275 0.732271 9.99958 2.98274e-06 1.19309e-05 0.131499 0.982503 0.931702 -0.0132927 4.9083e-06 0.50437 -1.91637e-20 7.07617e-24 -1.91567e-20 0.0013956 0.997817 8.59623e-05 0.152617 2.8521 0.0013956 0.99782 0.727105 0.00105434 0.00188027 0.000859623 0.455556 0.00188027 0.439735 0.000129197 1.02 0.887939 0.534608 0.286411 1.71742e-07 3.06698e-09 2383.32 3114.46 -0.0553627 0.482151 0.277488 0.25319 -0.593391 -0.169526 0.496847 -0.267381 -0.229475 1.905 1 0 297.835 0 2.12679 1.903 0.000299783 0.852986 0.666459 0.365405 0.416515 2.127 133.372 83.9347 18.7217 60.8731 0.00402472 0 -40 10
1.004 2.90797e-08 2.53907e-06 0.113176 0.113175 0.0120367 1.3218e-05 0.00115412 0.141471 0.000658107 0.142124 0.889338 101.785 0.242459 0.761748 4.21453 0.0575415 0.0397597 0.96024 0.0197692 0.00432713 0.0190321 0.00415457 0.00523079 0.00596791 0.209232 0.238716 58.0019 -87.8963 126.261 15.9633 145.021 0.000141161 0.267172 192.85 0.310513 0.0673644 0.00409621 0.000561877 0.00138347 0.98698 0.991728 -2.97889e-06 -85.6641 0.0930199 31185.9 302.829 0.983513 0.319147 0.732273 0.732269 9.99958 2.98275e-06 1.19309e-05 0.131502 0.982506 0.931702 -0.0132927 4.90833e-06 0.50438 -1.91647e-20 7.07658e-24 -1.91576e-20 0.0013956 0.997817 8.59624e-05 0.152617 2.8521 0.0013956 0.99782 0.7272 0.00105436 0.00188027 0.000859624 0.455556 0.00188027 0.439743 0.0001292 1.02 0.88794 0.534608 0.286413 1.71743e-07 3.067e-09 2383.3 3114.46 -0.0553633 0.482151 0.277488 0.253189 -0.593391 -0.169526 0.496844 -0.267379 -0.229474 1.906 1 0 297.835 0 2.12694 1.904 0.000299782 0.852985 0.666506 0.365291 0.41654 2.12715 133.38 83.9348 18.7217 60.8732 0.00402472 0 -40 10
1.005 2.91086e-08 2.53907e-06 0.113237 0.113235 0.0120366 1.32312e-05 0.00115412 0.141546 0.000658109 0.142199 0.88941 101.785 0.24245 0.761857 4.21482 0.0575502 0.0397624 0.960238 0.0197689 0.00432739 0.0190318 0.00415478 0.0052311 0.00596822 0.209244 0.238729 58.0019 -87.8963 126.261 15.9632 145.021 0.000141161 0.267172 192.85 0.310512 0.0673644 0.00409621 0.000561878 0.00138347 0.98698 0.991728 -2.9789e-06 -85.6641 0.09302 31185.8 302.835 0.983513 0.319147 0.732271 0.732267 9.99958 2.98275e-06 1.19309e-05 0.131504 0.982509 0.931703 -0.0132927 4.90836e-06 0.504391 -1.91657e-20 7.07698e-24 -1.91586e-20 0.0013956 0.997817 8.59625e-05 0.152617 2.8521 0.0013956 0.99782 0.727295 0.00105437 0.00188028 0.000859625 0.455556 0.00188027 0.43975 0.000129203 1.02 0.887941 0.534607 0.286414 1.71743e-07 3.06702e-09 2383.28 3114.45 -0.055364 0.482151 0.277487 0.253189 -0.593391 -0.169526 0.496841 -0.267377 -0.229474 1.907 1 0 297.835 0 2.12709 1.905 0.000299782 0.852984 0.666554 0.365178 0.416566 2.1273 133.388 83.9349 18.7217 60.8732 0.00402471 0 -40 10
1.006 2.91375e-08 2.53907e-06 0.113297 0.113295 0.0120366 1.32443e-05 0.00115412 0.141621 0.000658111 0.142275 0.889483 101.785 0.242441 0.761966 4.2151 0.0575588 0.0397651 0.960235 0.0197686 0.00432764 0.0190315 0.00415499 0.00523141 0.00596853 0.209257 0.238741 58.002 -87.8963 126.261 15.9632 145.021 0.00014116 0.267172 192.85 0.310512 0.0673643 0.00409621 0.000561878 0.00138347 0.98698 0.991728 -2.97892e-06 -85.664 0.0930201 31185.8 302.842 0.983513 0.319147 0.732269 0.732265 9.99958 2.98276e-06 1.19309e-05 0.131507 0.982512 0.931704 -0.0132927 4.90839e-06 0.504402 -1.91667e-20 7.07739e-24 -1.91596e-20 0.0013956 0.997817 8.59626e-05 0.152617 2.8521 0.0013956 0.99782 0.72739 0.00105439 0.00188028 0.000859626 0.455556 0.00188028 0.439758 0.000129206 1.02 0.887942 0.534607 0.286416 1.71743e-07 3.06705e-09 2383.27 3114.44 -0.0553646 0.482151 0.277487 0.253189 -0.593391 -0.169526 0.496839 -0.267375 -0.229473 1.908 1 0 297.835 0 2.12724 1.906 0.000299781 0.852983 0.666602 0.365065 0.416591 2.12745 133.396 83.935 18.7217 60.8733 0.00402471 0 -40 10
1.007 2.91664e-08 2.53907e-06 0.113357 0.113356 0.0120366 1.32575e-05 0.00115412 0.141697 0.000658112 0.14235 0.889555 101.785 0.242432 0.762075 4.21539 0.0575675 0.0397678 0.960232 0.0197683 0.00432789 0.0190312 0.00415521 0.00523173 0.00596884 0.209269 0.238754 58.0021 -87.8963 126.261 15.9632 145.021 0.00014116 0.267173 192.85 0.310512 0.0673643 0.00409622 0.000561879 0.00138348 0.98698 0.991728 -2.97893e-06 -85.664 0.0930201 31185.8 302.849 0.983513 0.319147 0.732268 0.732263 9.99958 2.98276e-06 1.19309e-05 0.13151 0.982515 0.931704 -0.0132927 4.90842e-06 0.504412 -1.91677e-20 7.0778e-24 -1.91606e-20 0.0013956 0.997817 8.59627e-05 0.152617 2.8521 0.0013956 0.99782 0.727485 0.00105441 0.00188028 0.000859627 0.455555 0.00188028 0.439765 0.000129209 1.02 0.887943 0.534607 0.286417 1.71743e-07 3.06707e-09 2383.25 3114.43 -0.0553653 0.482151 0.277487 0.253188 -0.593391 -0.169526 0.496836 -0.267373 -0.229472 1.909 1 0 297.834 0 2.1274 1.907 0.000299781 0.852983 0.666649 0.364952 0.416616 2.1276 133.404 83.9351 18.7217 60.8733 0.00402471 0 -40 10
1.008 2.91953e-08 2.53907e-06 0.113418 0.113416 0.0120366 1.32706e-05 0.00115412 0.141772 0.000658114 0.142425 0.889628 101.784 0.242424 0.762184 4.21568 0.0575762 0.0397705 0.960229 0.019768 0.00432815 0.0190308 0.00415542 0.00523204 0.00596916 0.209282 0.238766 58.0021 -87.8963 126.261 15.9631 145.021 0.00014116 0.267173 192.85 0.310511 0.0673642 0.00409622 0.00056188 0.00138348 0.98698 0.991728 -2.97895e-06 -85.664 0.0930202 31185.8 302.856 0.983513 0.319147 0.732266 0.732262 9.99958 2.98277e-06 1.1931e-05 0.131512 0.982518 0.931705 -0.0132927 4.90845e-06 0.504423 -1.91687e-20 7.07821e-24 -1.91616e-20 0.0013956 0.997817 8.59627e-05 0.152617 2.8521 0.0013956 0.99782 0.72758 0.00105443 0.00188028 0.000859627 0.455555 0.00188028 0.439773 0.000129213 1.02 0.887944 0.534607 0.286419 1.71744e-07 3.06709e-09 2383.23 3114.42 -0.055366 0.482152 0.277487 0.253188 -0.593391 -0.169526 0.496833 -0.267371 -0.229471 1.91 1 0 297.834 0 2.12755 1.908 0.00029978 0.852982 0.666697 0.364839 0.416641 2.12776 133.413 83.9352 18.7217 60.8733 0.0040247 0 -40 10
1.009 2.92242e-08 2.53907e-06 0.113478 0.113476 0.0120366 1.32837e-05 0.00115412 0.141847 0.000658116 0.142501 0.8897 101.784 0.242415 0.762293 4.21596 0.0575849 0.0397733 0.960227 0.0197676 0.0043284 0.0190305 0.00415564 0.00523235 0.00596947 0.209294 0.238779 58.0022 -87.8963 126.261 15.9631 145.021 0.000141159 0.267173 192.849 0.310511 0.0673642 0.00409622 0.00056188 0.00138348 0.98698 0.991728 -2.97896e-06 -85.664 0.0930203 31185.8 302.863 0.983513 0.319147 0.732264 0.73226 9.99958 2.98277e-06 1.1931e-05 0.131515 0.982521 0.931706 -0.0132927 4.90848e-06 0.504434 -1.91696e-20 7.07862e-24 -1.91626e-20 0.0013956 0.997817 8.59628e-05 0.152617 2.8521 0.0013956 0.99782 0.727674 0.00105445 0.00188028 0.000859628 0.455555 0.00188028 0.43978 0.000129216 1.02 0.887945 0.534606 0.28642 1.71744e-07 3.06712e-09 2383.22 3114.42 -0.0553667 0.482152 0.277486 0.253187 -0.593391 -0.169526 0.49683 -0.267369 -0.22947 1.911 1 0 297.834 0 2.1277 1.909 0.00029978 0.852982 0.666745 0.364727 0.416667 2.12791 133.421 83.9353 18.7217 60.8734 0.0040247 0 -40 10
1.01 2.92531e-08 2.53907e-06 0.113538 0.113536 0.0120366 1.32969e-05 0.00115412 0.141922 0.000658117 0.142576 0.889773 101.784 0.242406 0.762402 4.21625 0.0575936 0.039776 0.960224 0.0197673 0.00432866 0.0190302 0.00415585 0.00523267 0.00596979 0.209307 0.238792 58.0023 -87.8964 126.261 15.9631 145.021 0.000141159 0.267173 192.849 0.31051 0.0673641 0.00409623 0.000561881 0.00138348 0.98698 0.991728 -2.97897e-06 -85.664 0.0930204 31185.7 302.87 0.983513 0.319147 0.732263 0.732259 9.99958 2.98278e-06 1.1931e-05 0.131517 0.982524 0.931706 -0.0132927 4.9085e-06 0.504445 -1.91706e-20 7.07902e-24 -1.91636e-20 0.00139561 0.997817 8.59629e-05 0.152618 2.8521 0.00139561 0.99782 0.727769 0.00105447 0.00188028 0.000859629 0.455555 0.00188028 0.439788 0.000129219 1.02 0.887946 0.534606 0.286422 1.71744e-07 3.06714e-09 2383.2 3114.41 -0.0553674 0.482152 0.277486 0.253187 -0.593391 -0.169526 0.496827 -0.267366 -0.229469 1.912 1 0 297.833 0 2.12785 1.91 0.000299779 0.852981 0.666792 0.364615 0.416692 2.12806 133.429 83.9353 18.7218 60.8734 0.0040247 0 -40 10
1.011 2.92821e-08 2.53907e-06 0.113598 0.113596 0.0120366 1.331e-05 0.00115412 0.141997 0.000658119 0.142651 0.889845 101.783 0.242398 0.762511 4.21654 0.0576024 0.0397787 0.960221 0.019767 0.00432891 0.0190299 0.00415607 0.00523298 0.0059701 0.209319 0.238804 58.0023 -87.8964 126.261 15.963 145.021 0.000141159 0.267173 192.849 0.31051 0.0673641 0.00409623 0.000561882 0.00138348 0.98698 0.991728 -2.97899e-06 -85.664 0.0930205 31185.7 302.877 0.983513 0.319147 0.732261 0.732257 9.99958 2.98278e-06 1.1931e-05 0.13152 0.982528 0.931707 -0.0132927 4.90853e-06 0.504456 -1.91716e-20 7.07943e-24 -1.91645e-20 0.00139561 0.997817 8.5963e-05 0.152618 2.8521 0.00139561 0.99782 0.727864 0.00105449 0.00188028 0.00085963 0.455555 0.00188028 0.439795 0.000129222 1.02 0.887947 0.534606 0.286423 1.71745e-07 3.06716e-09 2383.18 3114.4 -0.0553681 0.482152 0.277486 0.253186 -0.593391 -0.169526 0.496823 -0.267364 -0.229468 1.913 1 0 297.833 0 2.128 1.911 0.000299779 0.852981 0.66684 0.364503 0.416717 2.12821 133.437 83.9354 18.7218 60.8735 0.00402469 0 -40 10
1.012 2.9311e-08 2.53907e-06 0.113658 0.113656 0.0120366 1.33232e-05 0.00115412 0.142072 0.00065812 0.142726 0.889918 101.783 0.242389 0.76262 4.21683 0.0576111 0.0397814 0.960219 0.0197667 0.00432917 0.0190296 0.00415628 0.00523329 0.00597042 0.209332 0.238817 58.0024 -87.8964 126.261 15.963 145.021 0.000141159 0.267174 192.849 0.31051 0.067364 0.00409623 0.000561882 0.00138349 0.98698 0.991728 -2.979e-06 -85.664 0.0930206 31185.7 302.884 0.983513 0.319147 0.73226 0.732256 9.99958 2.98279e-06 1.1931e-05 0.131523 0.982531 0.931708 -0.0132927 4.90856e-06 0.504466 -1.91726e-20 7.07984e-24 -1.91655e-20 0.00139561 0.997817 8.59631e-05 0.152618 2.85211 0.00139561 0.99782 0.727958 0.00105451 0.00188029 0.000859631 0.455554 0.00188028 0.439803 0.000129225 1.02 0.887949 0.534605 0.286425 1.71745e-07 3.06718e-09 2383.17 3114.39 -0.0553688 0.482152 0.277485 0.253186 -0.593391 -0.169526 0.49682 -0.267362 -0.229467 1.914 1 0 297.833 0 2.12816 1.912 0.000299778 0.852981 0.666887 0.364391 0.416742 2.12836 133.445 83.9355 18.7218 60.8735 0.00402469 0 -40 10
1.013 2.93399e-08 2.53907e-06 0.113718 0.113716 0.0120365 1.33363e-05 0.00115412 0.142147 0.000658122 0.142801 0.88999 101.783 0.24238 0.762729 4.21712 0.0576198 0.0397842 0.960216 0.0197664 0.00432943 0.0190293 0.0041565 0.00523361 0.00597073 0.209344 0.238829 58.0024 -87.8964 126.261 15.9629 145.021 0.000141158 0.267174 192.849 0.310509 0.067364 0.00409624 0.000561883 0.00138349 0.98698 0.991728 -2.97902e-06 -85.664 0.0930207 31185.7 302.891 0.983513 0.319147 0.732259 0.732254 9.99958 2.98279e-06 1.19311e-05 0.131525 0.982534 0.931708 -0.0132927 4.90859e-06 0.504477 -1.91736e-20 7.08025e-24 -1.91665e-20 0.00139561 0.997817 8.59631e-05 0.152618 2.85211 0.00139561 0.99782 0.728053 0.00105452 0.00188029 0.000859631 0.455554 0.00188029 0.43981 0.000129228 1.02 0.88795 0.534605 0.286426 1.71745e-07 3.06721e-09 2383.15 3114.39 -0.0553696 0.482152 0.277485 0.253186 -0.593391 -0.169526 0.496817 -0.26736 -0.229466 1.915 1 0 297.832 0 2.12831 1.913 0.000299777 0.852981 0.666935 0.364279 0.416768 2.12852 133.453 83.9356 18.7218 60.8735 0.00402469 0 -40 10
1.014 2.93688e-08 2.53907e-06 0.113778 0.113776 0.0120365 1.33495e-05 0.00115412 0.142222 0.000658124 0.142876 0.890063 101.783 0.242371 0.762838 4.21741 0.0576285 0.0397869 0.960213 0.0197661 0.00432968 0.0190289 0.00415671 0.00523392 0.00597105 0.209357 0.238842 58.0025 -87.8964 126.261 15.9629 145.021 0.000141158 0.267174 192.849 0.310509 0.0673639 0.00409624 0.000561884 0.00138349 0.98698 0.991728 -2.97903e-06 -85.664 0.0930208 31185.6 302.898 0.983513 0.319147 0.732257 0.732253 9.99958 2.9828e-06 1.19311e-05 0.131528 0.982537 0.931709 -0.0132927 4.90862e-06 0.504488 -1.91746e-20 7.08066e-24 -1.91675e-20 0.00139561 0.997817 8.59632e-05 0.152618 2.85211 0.00139561 0.99782 0.728148 0.00105454 0.00188029 0.000859632 0.455554 0.00188029 0.439818 0.000129231 1.02 0.887951 0.534605 0.286428 1.71745e-07 3.06723e-09 2383.13 3114.38 -0.0553704 0.482152 0.277485 0.253185 -0.593391 -0.169526 0.496814 -0.267358 -0.229465 1.916 1 0 297.832 0 2.12846 1.914 0.000299777 0.852981 0.666982 0.364168 0.416793 2.12867 133.461 83.9356 18.7218 60.8736 0.00402469 0 -40 10
1.015 2.93977e-08 2.53908e-06 0.113838 0.113836 0.0120365 1.33626e-05 0.00115413 0.142297 0.000658125 0.142951 0.890136 101.782 0.242363 0.762947 4.2177 0.0576372 0.0397896 0.96021 0.0197658 0.00432994 0.0190286 0.00415693 0.00523424 0.00597137 0.20937 0.238855 58.0026 -87.8964 126.261 15.9629 145.021 0.000141158 0.267174 192.848 0.310508 0.0673639 0.00409624 0.000561884 0.00138349 0.98698 0.991728 -2.97905e-06 -85.664 0.0930208 31185.6 302.905 0.983513 0.319147 0.732256 0.732251 9.99958 2.9828e-06 1.19311e-05 0.13153 0.98254 0.93171 -0.0132927 4.90865e-06 0.504499 -1.91756e-20 7.08107e-24 -1.91685e-20 0.00139561 0.997817 8.59633e-05 0.152618 2.85211 0.00139561 0.99782 0.728242 0.00105456 0.00188029 0.000859633 0.455554 0.00188029 0.439825 0.000129234 1.02 0.887952 0.534604 0.286429 1.71746e-07 3.06725e-09 2383.12 3114.37 -0.0553712 0.482152 0.277485 0.253185 -0.593391 -0.169527 0.496811 -0.267356 -0.229464 1.917 1 0 297.832 0 2.12861 1.915 0.000299776 0.852981 0.66703 0.364057 0.416818 2.12882 133.47 83.9357 18.7218 60.8736 0.00402468 0 -40 10
1.016 2.94266e-08 2.53908e-06 0.113897 0.113896 0.0120365 1.33757e-05 0.00115413 0.142372 0.000658127 0.143025 0.890209 101.782 0.242354 0.763056 4.21799 0.057646 0.0397924 0.960208 0.0197654 0.00433019 0.0190283 0.00415715 0.00523455 0.00597169 0.209382 0.238867 58.0026 -87.8964 126.261 15.9628 145.021 0.000141157 0.267174 192.848 0.310508 0.0673638 0.00409625 0.000561885 0.0013835 0.98698 0.991728 -2.97906e-06 -85.664 0.0930209 31185.6 302.912 0.983512 0.319147 0.732254 0.73225 9.99958 2.98281e-06 1.19311e-05 0.131533 0.982543 0.93171 -0.0132927 4.90868e-06 0.50451 -1.91766e-20 7.08148e-24 -1.91695e-20 0.00139561 0.997817 8.59634e-05 0.152619 2.85211 0.00139561 0.99782 0.728337 0.00105458 0.00188029 0.000859634 0.455553 0.00188029 0.439833 0.000129237 1.02 0.887953 0.534604 0.286431 1.71746e-07 3.06727e-09 2383.1 3114.37 -0.055372 0.482152 0.277484 0.253184 -0.593391 -0.169527 0.496807 -0.267354 -0.229463 1.918 1 0 297.831 0 2.12876 1.916 0.000299776 0.852981 0.667077 0.363946 0.416843 2.12897 133.478 83.9358 18.7218 60.8736 0.00402468 0 -40 10
1.017 2.94556e-08 2.53908e-06 0.113957 0.113956 0.0120365 1.33889e-05 0.00115413 0.142446 0.000658128 0.1431 0.890281 101.782 0.242345 0.763166 4.21828 0.0576547 0.0397951 0.960205 0.0197651 0.00433045 0.019028 0.00415736 0.00523487 0.005972 0.209395 0.23888 58.0027 -87.8964 126.262 15.9628 145.021 0.000141157 0.267174 192.848 0.310507 0.0673638 0.00409625 0.000561886 0.0013835 0.98698 0.991728 -2.97908e-06 -85.6639 0.093021 31185.6 302.919 0.983512 0.319147 0.732253 0.732249 9.99958 2.98281e-06 1.19311e-05 0.131536 0.982546 0.931711 -0.0132927 4.90871e-06 0.504521 -1.91776e-20 7.08189e-24 -1.91705e-20 0.00139561 0.997817 8.59635e-05 0.152619 2.85211 0.00139561 0.99782 0.728431 0.0010546 0.00188029 0.000859635 0.455553 0.00188029 0.43984 0.00012924 1.02 0.887954 0.534604 0.286432 1.71746e-07 3.0673e-09 2383.08 3114.36 -0.0553728 0.482152 0.277484 0.253184 -0.593391 -0.169527 0.496804 -0.267352 -0.229462 1.919 1 0 297.831 0 2.12891 1.917 0.000299775 0.852981 0.667125 0.363835 0.416868 2.12912 133.486 83.9358 18.7218 60.8737 0.00402468 0 -40 10
1.018 2.94845e-08 2.53908e-06 0.114017 0.114015 0.0120365 1.3402e-05 0.00115413 0.142521 0.00065813 0.143175 0.890354 101.781 0.242337 0.763275 4.21858 0.0576635 0.0397979 0.960202 0.0197648 0.00433071 0.0190277 0.00415758 0.00523519 0.00597232 0.209408 0.238893 58.0028 -87.8964 126.262 15.9627 145.021 0.000141157 0.267175 192.848 0.310507 0.0673637 0.00409625 0.000561886 0.0013835 0.98698 0.991728 -2.97909e-06 -85.6639 0.0930211 31185.6 302.925 0.983512 0.319147 0.732252 0.732248 9.99958 2.98282e-06 1.19312e-05 0.131538 0.982549 0.931712 -0.0132927 4.90874e-06 0.504532 -1.91786e-20 7.0823e-24 -1.91715e-20 0.00139561 0.997817 8.59635e-05 0.152619 2.85211 0.00139561 0.99782 0.728526 0.00105462 0.0018803 0.000859635 0.455553 0.00188029 0.439848 0.000129243 1.02 0.887955 0.534603 0.286434 1.71746e-07 3.06732e-09 2383.07 3114.36 -0.0553736 0.482152 0.277484 0.253184 -0.593391 -0.169527 0.496801 -0.26735 -0.22946 1.92 1 0 297.83 0 2.12907 1.918 0.000299775 0.852981 0.667172 0.363725 0.416893 2.12927 133.494 83.9359 18.7218 60.8737 0.00402468 0 -40 10
1.019 2.95134e-08 2.53908e-06 0.114077 0.114075 0.0120365 1.34152e-05 0.00115413 0.142596 0.000658132 0.143249 0.890427 101.781 0.242328 0.763385 4.21887 0.0576722 0.0398007 0.960199 0.0197645 0.00433097 0.0190274 0.0041578 0.0052355 0.00597264 0.20942 0.238906 58.0028 -87.8964 126.262 15.9627 145.021 0.000141157 0.267175 192.848 0.310507 0.0673637 0.00409625 0.000561887 0.0013835 0.98698 0.991728 -2.97911e-06 -85.6639 0.0930212 31185.5 302.932 0.983512 0.319147 0.732251 0.732247 9.99958 2.98282e-06 1.19312e-05 0.131541 0.982552 0.931712 -0.0132927 4.90877e-06 0.504542 -1.91796e-20 7.08271e-24 -1.91725e-20 0.00139562 0.997817 8.59636e-05 0.152619 2.85211 0.00139562 0.99782 0.72862 0.00105464 0.0018803 0.000859636 0.455553 0.0018803 0.439855 0.000129246 1.02 0.887956 0.534603 0.286435 1.71747e-07 3.06734e-09 2383.05 3114.35 -0.0553745 0.482152 0.277483 0.253183 -0.593391 -0.169527 0.496797 -0.267347 -0.229459 1.921 1 0 297.83 0 2.12922 1.919 0.000299774 0.852982 0.66722 0.363615 0.416919 2.12943 133.502 83.9359 18.7218 60.8737 0.00402467 0 -40 10
1.02 2.95423e-08 2.53908e-06 0.114136 0.114135 0.0120364 1.34283e-05 0.00115413 0.14267 0.000658133 0.143324 0.8905 101.781 0.242319 0.763494 4.21916 0.057681 0.0398034 0.960197 0.0197642 0.00433123 0.019027 0.00415801 0.00523582 0.00597296 0.209433 0.238918 58.0029 -87.8964 126.262 15.9627 145.021 0.000141157 0.267175 192.848 0.310506 0.0673636 0.00409626 0.000561888 0.0013835 0.98698 0.991728 -2.97912e-06 -85.6639 0.0930213 31185.5 302.939 0.983512 0.319147 0.73225 0.732245 9.99958 2.98283e-06 1.19312e-05 0.131544 0.982555 0.931713 -0.0132927 4.9088e-06 0.504553 -1.91806e-20 7.08312e-24 -1.91735e-20 0.00139562 0.997817 8.59637e-05 0.152619 2.85211 0.00139562 0.99782 0.728714 0.00105466 0.0018803 0.000859637 0.455552 0.0018803 0.439863 0.000129249 1.02 0.887957 0.534603 0.286437 1.71747e-07 3.06737e-09 2383.03 3114.35 -0.0553753 0.482152 0.277483 0.253183 -0.593391 -0.169527 0.496794 -0.267345 -0.229458 1.922 1 0 297.829 0 2.12937 1.92 0.000299773 0.852982 0.667267 0.363505 0.416944 2.12958 133.51 83.936 18.7218 60.8737 0.00402467 0 -40 10
1.021 2.95712e-08 2.53908e-06 0.114196 0.114194 0.0120364 1.34415e-05 0.00115413 0.142745 0.000658135 0.143398 0.890573 101.781 0.24231 0.763604 4.21945 0.0576897 0.0398062 0.960194 0.0197639 0.00433148 0.0190267 0.00415823 0.00523614 0.00597328 0.209446 0.238931 58.003 -87.8964 126.262 15.9626 145.021 0.000141156 0.267175 192.847 0.310506 0.0673635 0.00409626 0.000561888 0.00138351 0.98698 0.991728 -2.97914e-06 -85.6639 0.0930214 31185.5 302.946 0.983512 0.319147 0.732249 0.732244 9.99958 2.98283e-06 1.19312e-05 0.131546 0.982558 0.931713 -0.0132927 4.90883e-06 0.504564 -1.91816e-20 7.08353e-24 -1.91745e-20 0.00139562 0.997817 8.59638e-05 0.152619 2.85211 0.00139562 0.99782 0.728809 0.00105467 0.0018803 0.000859638 0.455552 0.0018803 0.43987 0.000129252 1.02 0.887958 0.534603 0.286438 1.71747e-07 3.06739e-09 2383.02 3114.34 -0.0553762 0.482153 0.277483 0.253183 -0.593391 -0.169527 0.49679 -0.267343 -0.229456 1.923 1 0 297.829 0 2.12952 1.921 0.000299773 0.852983 0.667315 0.363395 0.416969 2.12973 133.518 83.936 18.7218 60.8738 0.00402467 0 -40 10
1.022 2.96001e-08 2.53908e-06 0.114255 0.114254 0.0120364 1.34546e-05 0.00115413 0.142819 0.000658136 0.143473 0.890646 101.78 0.242302 0.763713 4.21975 0.0576985 0.0398089 0.960191 0.0197635 0.00433174 0.0190264 0.00415845 0.00523646 0.0059736 0.209458 0.238944 58.003 -87.8964 126.262 15.9626 145.021 0.000141156 0.267175 192.847 0.310505 0.0673635 0.00409626 0.000561889 0.00138351 0.98698 0.991728 -2.97915e-06 -85.6639 0.0930215 31185.5 302.954 0.983512 0.319147 0.732248 0.732243 9.99958 2.98284e-06 1.19312e-05 0.131549 0.982561 0.931714 -0.0132927 4.90886e-06 0.504575 -1.91826e-20 7.08394e-24 -1.91755e-20 0.00139562 0.997817 8.59639e-05 0.152619 2.85211 0.00139562 0.99782 0.728903 0.00105469 0.0018803 0.000859639 0.455552 0.0018803 0.439878 0.000129255 1.02 0.887959 0.534602 0.28644 1.71747e-07 3.06741e-09 2383 3114.34 -0.0553771 0.482153 0.277483 0.253183 -0.593391 -0.169527 0.496786 -0.267341 -0.229455 1.924 1 0 297.828 0 2.12967 1.922 0.000299772 0.852984 0.667362 0.363285 0.416994 2.12988 133.526 83.9361 18.7218 60.8738 0.00402467 0 -40 10
1.023 2.9629e-08 2.53908e-06 0.114315 0.114313 0.0120364 1.34677e-05 0.00115413 0.142893 0.000658138 0.143547 0.890719 101.78 0.242293 0.763823 4.22004 0.0577072 0.0398117 0.960188 0.0197632 0.004332 0.0190261 0.00415867 0.00523678 0.00597392 0.209471 0.238957 58.0031 -87.8964 126.262 15.9626 145.021 0.000141156 0.267176 192.847 0.310505 0.0673634 0.00409627 0.00056189 0.00138351 0.98698 0.991728 -2.97917e-06 -85.6639 0.0930215 31185.4 302.961 0.983512 0.319147 0.732247 0.732242 9.99958 2.98284e-06 1.19313e-05 0.131551 0.982564 0.931715 -0.0132927 4.90889e-06 0.504586 -1.91835e-20 7.08436e-24 -1.91765e-20 0.00139562 0.997817 8.59639e-05 0.15262 2.85212 0.00139562 0.99782 0.728997 0.00105471 0.0018803 0.000859639 0.455552 0.0018803 0.439885 0.000129258 1.02 0.887961 0.534602 0.286442 1.71748e-07 3.06743e-09 2382.98 3114.33 -0.055378 0.482153 0.277482 0.253182 -0.593391 -0.169527 0.496783 -0.267339 -0.229453 1.925 1 0 297.828 0 2.12982 1.923 0.000299772 0.852985 0.66741 0.363176 0.417019 2.13003 133.535 83.9361 18.7218 60.8738 0.00402466 0 -40 10
1.024 2.96579e-08 2.53908e-06 0.114374 0.114373 0.0120364 1.34809e-05 0.00115413 0.142968 0.000658139 0.143621 0.890792 101.78 0.242284 0.763933 4.22034 0.057716 0.0398145 0.960185 0.0197629 0.00433226 0.0190258 0.00415889 0.0052371 0.00597424 0.209484 0.23897 58.0031 -87.8964 126.262 15.9625 145.021 0.000141156 0.267176 192.847 0.310504 0.0673634 0.00409627 0.00056189 0.00138351 0.98698 0.991728 -2.97918e-06 -85.6639 0.0930216 31185.4 302.968 0.983512 0.319147 0.732246 0.732241 9.99958 2.98285e-06 1.19313e-05 0.131554 0.982567 0.931715 -0.0132927 4.90892e-06 0.504597 -1.91845e-20 7.08477e-24 -1.91775e-20 0.00139562 0.997817 8.5964e-05 0.15262 2.85212 0.00139562 0.99782 0.729091 0.00105473 0.0018803 0.00085964 0.455552 0.0018803 0.439893 0.000129261 1.02 0.887962 0.534602 0.286443 1.71748e-07 3.06746e-09 2382.97 3114.33 -0.0553789 0.482153 0.277482 0.253182 -0.593391 -0.169527 0.496779 -0.267337 -0.229452 1.926 1 0 297.827 0 2.12998 1.924 0.000299771 0.852985 0.667457 0.363067 0.417044 2.13018 133.543 83.9362 18.7218 60.8738 0.00402466 0 -40 10
1.025 2.96869e-08 2.53908e-06 0.114434 0.114432 0.0120364 1.3494e-05 0.00115413 0.143042 0.000658141 0.143696 0.890865 101.779 0.242275 0.764043 4.22063 0.0577248 0.0398173 0.960183 0.0197626 0.00433252 0.0190254 0.00415911 0.00523742 0.00597456 0.209497 0.238982 58.0032 -87.8964 126.262 15.9625 145.021 0.000141156 0.267176 192.847 0.310504 0.0673633 0.00409627 0.000561891 0.00138351 0.98698 0.991728 -2.9792e-06 -85.6639 0.0930217 31185.4 302.975 0.983512 0.319147 0.732245 0.732241 9.99958 2.98285e-06 1.19313e-05 0.131557 0.98257 0.931716 -0.0132927 4.90895e-06 0.504608 -1.91855e-20 7.08518e-24 -1.91785e-20 0.00139562 0.997817 8.59641e-05 0.15262 2.85212 0.00139562 0.99782 0.729186 0.00105475 0.00188031 0.000859641 0.455551 0.0018803 0.4399 0.000129265 1.02 0.887963 0.534601 0.286445 1.71748e-07 3.06748e-09 2382.95 3114.32 -0.0553798 0.482153 0.277482 0.253182 -0.593391 -0.169527 0.496775 -0.267335 -0.22945 1.927 1 0 297.827 0 2.13013 1.925 0.000299771 0.852986 0.667505 0.362958 0.417069 2.13033 133.551 83.9362 18.7218 60.8739 0.00402466 0 -40 10
1.026 2.97158e-08 2.53908e-06 0.114493 0.114491 0.0120364 1.35072e-05 0.00115413 0.143116 0.000658143 0.14377 0.890938 101.779 0.242266 0.764152 4.22093 0.0577336 0.0398201 0.96018 0.0197623 0.00433278 0.0190251 0.00415933 0.00523774 0.00597488 0.209509 0.238995 58.0033 -87.8964 126.262 15.9624 145.021 0.000141155 0.267176 192.847 0.310504 0.0673633 0.00409628 0.000561892 0.00138352 0.986979 0.991728 -2.97921e-06 -85.6639 0.0930218 31185.4 302.982 0.983512 0.319147 0.732244 0.73224 9.99958 2.98286e-06 1.19313e-05 0.131559 0.982573 0.931716 -0.0132927 4.90898e-06 0.504619 -1.91865e-20 7.08559e-24 -1.91795e-20 0.00139562 0.997817 8.59642e-05 0.15262 2.85212 0.00139562 0.99782 0.72928 0.00105477 0.00188031 0.000859642 0.455551 0.00188031 0.439907 0.000129268 1.02 0.887964 0.534601 0.286446 1.71749e-07 3.0675e-09 2382.93 3114.32 -0.0553808 0.482153 0.277481 0.253182 -0.593392 -0.169527 0.496772 -0.267333 -0.229448 1.928 1 0 297.826 0 2.13028 1.926 0.00029977 0.852987 0.667552 0.362849 0.417095 2.13049 133.559 83.9363 18.7218 60.8739 0.00402466 0 -40 10
1.027 2.97447e-08 2.53908e-06 0.114552 0.114551 0.0120364 1.35203e-05 0.00115413 0.14319 0.000658144 0.143844 0.891011 101.779 0.242258 0.764262 4.22122 0.0577423 0.0398229 0.960177 0.0197619 0.00433304 0.0190248 0.00415955 0.00523806 0.0059752 0.209522 0.239008 58.0033 -87.8964 126.262 15.9624 145.021 0.000141155 0.267176 192.846 0.310503 0.0673632 0.00409628 0.000561892 0.00138352 0.986979 0.991728 -2.97923e-06 -85.6639 0.0930219 31185.4 302.989 0.983512 0.319147 0.732243 0.732239 9.99958 2.98286e-06 1.19313e-05 0.131562 0.982576 0.931717 -0.0132926 4.90901e-06 0.50463 -1.91875e-20 7.08601e-24 -1.91805e-20 0.00139562 0.997817 8.59643e-05 0.15262 2.85212 0.00139562 0.99782 0.729374 0.00105479 0.00188031 0.000859643 0.455551 0.00188031 0.439915 0.000129271 1.02 0.887965 0.534601 0.286448 1.71749e-07 3.06753e-09 2382.91 3114.31 -0.0553818 0.482153 0.277481 0.253181 -0.593392 -0.169527 0.496768 -0.267331 -0.229447 1.929 1 0 297.826 0 2.13043 1.927 0.000299769 0.852989 0.667599 0.362741 0.41712 2.13064 133.567 83.9363 18.7218 60.8739 0.00402466 0 -40 10
1.028 2.97736e-08 2.53908e-06 0.114611 0.11461 0.0120363 1.35335e-05 0.00115413 0.143264 0.000658146 0.143918 0.891084 101.778 0.242249 0.764372 4.22152 0.0577511 0.0398257 0.960174 0.0197616 0.0043333 0.0190245 0.00415977 0.00523838 0.00597552 0.209535 0.239021 58.0034 -87.8964 126.262 15.9624 145.021 0.000141155 0.267177 192.846 0.310503 0.0673632 0.00409628 0.000561893 0.00138352 0.986979 0.991728 -2.97924e-06 -85.6638 0.093022 31185.3 302.996 0.983512 0.319147 0.732243 0.732238 9.99958 2.98287e-06 1.19314e-05 0.131565 0.982579 0.931717 -0.0132926 4.90904e-06 0.504641 -1.91885e-20 7.08642e-24 -1.91815e-20 0.00139563 0.997817 8.59643e-05 0.15262 2.85212 0.00139563 0.99782 0.729468 0.00105481 0.00188031 0.000859643 0.455551 0.00188031 0.439922 0.000129274 1.02 0.887966 0.5346 0.286449 1.71749e-07 3.06755e-09 2382.9 3114.31 -0.0553827 0.482153 0.277481 0.253181 -0.593392 -0.169527 0.496764 -0.267328 -0.229445 1.93 1 0 297.825 0 2.13058 1.928 0.000299769 0.85299 0.667647 0.362633 0.417145 2.13079 133.575 83.9363 18.7218 60.8739 0.00402466 0 -40 10
1.029 2.98025e-08 2.53909e-06 0.114671 0.114669 0.0120363 1.35466e-05 0.00115413 0.143338 0.000658147 0.143992 0.891157 101.778 0.24224 0.764482 4.22182 0.0577599 0.0398285 0.960172 0.0197613 0.00433356 0.0190242 0.00415999 0.0052387 0.00597585 0.209548 0.239034 58.0035 -87.8964 126.262 15.9623 145.021 0.000141155 0.267177 192.846 0.310502 0.0673631 0.00409628 0.000561894 0.00138352 0.986979 0.991728 -2.97926e-06 -85.6638 0.0930221 31185.3 303.003 0.983512 0.319147 0.732242 0.732237 9.99958 2.98287e-06 1.19314e-05 0.131567 0.982582 0.931718 -0.0132926 4.90907e-06 0.504652 -1.91896e-20 7.08683e-24 -1.91825e-20 0.00139563 0.997817 8.59644e-05 0.152621 2.85212 0.00139563 0.99782 0.729562 0.00105482 0.00188031 0.000859644 0.45555 0.00188031 0.43993 0.000129277 1.02 0.887967 0.5346 0.286451 1.71749e-07 3.06757e-09 2382.88 3114.31 -0.0553837 0.482153 0.277481 0.253181 -0.593392 -0.169527 0.49676 -0.267326 -0.229443 1.931 1 0 297.825 0 2.13073 1.929 0.000299768 0.852991 0.667694 0.362524 0.41717 2.13094 133.583 83.9364 18.7218 60.8739 0.00402465 0 -40 10
1.03 2.98314e-08 2.53909e-06 0.11473 0.114728 0.0120363 1.35597e-05 0.00115413 0.143412 0.000658149 0.144066 0.891231 101.778 0.242231 0.764592 4.22211 0.0577687 0.0398313 0.960169 0.019761 0.00433382 0.0190238 0.00416021 0.00523902 0.00597617 0.209561 0.239047 58.0035 -87.8964 126.262 15.9623 145.021 0.000141155 0.267177 192.846 0.310502 0.0673631 0.00409629 0.000561894 0.00138353 0.986979 0.991728 -2.97927e-06 -85.6638 0.0930221 31185.3 303.01 0.983512 0.319147 0.732241 0.732237 9.99958 2.98288e-06 1.19314e-05 0.13157 0.982584 0.931719 -0.0132926 4.9091e-06 0.504663 -1.91906e-20 7.08725e-24 -1.91835e-20 0.00139563 0.997817 8.59645e-05 0.152621 2.85212 0.00139563 0.99782 0.729656 0.00105484 0.00188031 0.000859645 0.45555 0.00188031 0.439937 0.00012928 1.02 0.887968 0.5346 0.286452 1.7175e-07 3.06759e-09 2382.86 3114.3 -0.0553847 0.482153 0.27748 0.253181 -0.593392 -0.169527 0.496756 -0.267324 -0.229441 1.932 1 0 297.824 0 2.13088 1.93 0.000299768 0.852993 0.667742 0.362417 0.417195 2.13109 133.591 83.9364 18.7218 60.8739 0.00402465 0 -40 10
1.031 2.98603e-08 2.53909e-06 0.114789 0.114787 0.0120363 1.35729e-05 0.00115413 0.143486 0.00065815 0.14414 0.891304 101.778 0.242222 0.764702 4.22241 0.0577775 0.0398341 0.960166 0.0197607 0.00433409 0.0190235 0.00416043 0.00523934 0.00597649 0.209574 0.23906 58.0036 -87.8964 126.262 15.9623 145.021 0.000141155 0.267177 192.846 0.310501 0.067363 0.00409629 0.000561895 0.00138353 0.986979 0.991728 -2.97929e-06 -85.6638 0.0930222 31185.3 303.017 0.983512 0.319147 0.732241 0.732236 9.99958 2.98288e-06 1.19314e-05 0.131573 0.982587 0.931719 -0.0132926 4.90913e-06 0.504674 -1.91916e-20 7.08766e-24 -1.91845e-20 0.00139563 0.997817 8.59646e-05 0.152621 2.85212 0.00139563 0.99782 0.72975 0.00105486 0.00188031 0.000859646 0.45555 0.00188031 0.439945 0.000129283 1.02 0.887969 0.534599 0.286454 1.7175e-07 3.06762e-09 2382.85 3114.3 -0.0553857 0.482153 0.27748 0.253181 -0.593392 -0.169528 0.496752 -0.267322 -0.229439 1.933 1 0 297.823 0 2.13103 1.931 0.000299767 0.852994 0.667789 0.362309 0.41722 2.13124 133.599 83.9364 18.7218 60.874 0.00402465 0 -40 10
1.032 2.98893e-08 2.53909e-06 0.114848 0.114846 0.0120363 1.3586e-05 0.00115413 0.14356 0.000658152 0.144214 0.891377 101.777 0.242214 0.764813 4.22271 0.0577863 0.0398369 0.960163 0.0197603 0.00433435 0.0190232 0.00416065 0.00523966 0.00597682 0.209586 0.239073 58.0037 -87.8964 126.262 15.9622 145.021 0.000141155 0.267177 192.846 0.310501 0.067363 0.00409629 0.000561896 0.00138353 0.986979 0.991728 -2.9793e-06 -85.6638 0.0930223 31185.2 303.024 0.983512 0.319147 0.73224 0.732236 9.99958 2.98289e-06 1.19314e-05 0.131575 0.98259 0.93172 -0.0132926 4.90916e-06 0.504685 -1.91926e-20 7.08808e-24 -1.91855e-20 0.00139563 0.997817 8.59647e-05 0.152621 2.85212 0.00139563 0.99782 0.729844 0.00105488 0.00188032 0.000859647 0.45555 0.00188031 0.439952 0.000129286 1.02 0.88797 0.534599 0.286455 1.7175e-07 3.06764e-09 2382.83 3114.3 -0.0553868 0.482153 0.27748 0.253181 -0.593392 -0.169528 0.496748 -0.26732 -0.229437 1.934 1 0 297.823 0 2.13119 1.932 0.000299767 0.852996 0.667836 0.362202 0.417245 2.13139 133.608 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.033 2.99182e-08 2.53909e-06 0.114907 0.114905 0.0120363 1.35992e-05 0.00115413 0.143634 0.000658153 0.144287 0.89145 101.777 0.242205 0.764923 4.22301 0.0577951 0.0398397 0.96016 0.01976 0.00433461 0.0190229 0.00416087 0.00523998 0.00597714 0.209599 0.239086 58.0037 -87.8964 126.262 15.9622 145.021 0.000141155 0.267178 192.845 0.310501 0.0673629 0.0040963 0.000561896 0.00138353 0.986979 0.991728 -2.97932e-06 -85.6638 0.0930224 31185.2 303.031 0.983512 0.319147 0.732239 0.732235 9.99958 2.98289e-06 1.19315e-05 0.131578 0.982593 0.93172 -0.0132926 4.90918e-06 0.504697 -1.91936e-20 7.08849e-24 -1.91865e-20 0.00139563 0.997817 8.59647e-05 0.152621 2.85212 0.00139563 0.99782 0.729938 0.0010549 0.00188032 0.000859647 0.45555 0.00188032 0.439959 0.000129289 1.02 0.887972 0.534599 0.286457 1.7175e-07 3.06766e-09 2382.81 3114.29 -0.0553878 0.482153 0.277479 0.25318 -0.593392 -0.169528 0.496744 -0.267318 -0.229435 1.935 1 0 297.822 0 2.13134 1.933 0.000299766 0.852997 0.667884 0.362094 0.41727 2.13154 133.616 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.034 2.99471e-08 2.53909e-06 0.114966 0.114964 0.0120363 1.36123e-05 0.00115413 0.143707 0.000658155 0.144361 0.891524 101.777 0.242196 0.765033 4.22331 0.0578039 0.0398425 0.960157 0.0197597 0.00433487 0.0190225 0.00416109 0.00524031 0.00597746 0.209612 0.239099 58.0038 -87.8964 126.262 15.9621 145.021 0.000141155 0.267178 192.845 0.3105 0.0673629 0.0040963 0.000561897 0.00138353 0.986979 0.991728 -2.97933e-06 -85.6638 0.0930225 31185.2 303.038 0.983512 0.319147 0.732239 0.732235 9.99958 2.9829e-06 1.19315e-05 0.131581 0.982596 0.931721 -0.0132926 4.90921e-06 0.504708 -1.91946e-20 7.08891e-24 -1.91875e-20 0.00139563 0.997817 8.59648e-05 0.152621 2.85213 0.00139563 0.99782 0.730032 0.00105492 0.00188032 0.000859648 0.455549 0.00188032 0.439967 0.000129292 1.02 0.887973 0.534599 0.286458 1.71751e-07 3.06769e-09 2382.8 3114.29 -0.0553889 0.482154 0.277479 0.25318 -0.593392 -0.169528 0.49674 -0.267316 -0.229434 1.936 1 0 297.822 0 2.13149 1.934 0.000299765 0.852999 0.667931 0.361987 0.417295 2.13169 133.624 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.035 2.9976e-08 2.53909e-06 0.115025 0.115023 0.0120362 1.36255e-05 0.00115413 0.143781 0.000658157 0.144435 0.891597 101.776 0.242187 0.765143 4.22361 0.0578127 0.0398453 0.960155 0.0197594 0.00433513 0.0190222 0.00416131 0.00524063 0.00597779 0.209625 0.239112 58.0038 -87.8964 126.262 15.9621 145.021 0.000141154 0.267178 192.845 0.3105 0.0673628 0.0040963 0.000561898 0.00138354 0.986979 0.991728 -2.97935e-06 -85.6638 0.0930226 31185.2 303.046 0.983512 0.319147 0.732239 0.732234 9.99958 2.9829e-06 1.19315e-05 0.131584 0.982599 0.931721 -0.0132926 4.90924e-06 0.504719 -1.91956e-20 7.08932e-24 -1.91885e-20 0.00139563 0.997817 8.59649e-05 0.152621 2.85213 0.00139563 0.99782 0.730126 0.00105494 0.00188032 0.000859649 0.455549 0.00188032 0.439974 0.000129295 1.02 0.887974 0.534598 0.28646 1.71751e-07 3.06771e-09 2382.78 3114.29 -0.05539 0.482154 0.277479 0.25318 -0.593392 -0.169528 0.496736 -0.267314 -0.229431 1.937 1 0 297.821 0 2.13164 1.935 0.000299765 0.853001 0.667978 0.36188 0.41732 2.13185 133.632 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.036 3.00049e-08 2.53909e-06 0.115084 0.115082 0.0120362 1.36386e-05 0.00115413 0.143855 0.000658158 0.144508 0.891671 101.776 0.242178 0.765254 4.22391 0.0578216 0.0398482 0.960152 0.019759 0.0043354 0.0190219 0.00416153 0.00524095 0.00597811 0.209638 0.239125 58.0039 -87.8965 126.262 15.9621 145.021 0.000141154 0.267178 192.845 0.310499 0.0673628 0.00409631 0.000561898 0.00138354 0.986979 0.991728 -2.97936e-06 -85.6638 0.0930227 31185.2 303.053 0.983512 0.319147 0.732238 0.732234 9.99958 2.98291e-06 1.19315e-05 0.131586 0.982602 0.931722 -0.0132926 4.90927e-06 0.50473 -1.91966e-20 7.08974e-24 -1.91895e-20 0.00139563 0.997817 8.5965e-05 0.152622 2.85213 0.00139563 0.99782 0.73022 0.00105496 0.00188032 0.00085965 0.455549 0.00188032 0.439982 0.000129298 1.02 0.887975 0.534598 0.286461 1.71751e-07 3.06773e-09 2382.76 3114.28 -0.0553911 0.482154 0.277479 0.25318 -0.593392 -0.169528 0.496732 -0.267312 -0.229429 1.938 1 0 297.82 0 2.13179 1.936 0.000299764 0.853003 0.668025 0.361774 0.417345 2.132 133.64 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.037 3.00338e-08 2.53909e-06 0.115143 0.115141 0.0120362 1.36517e-05 0.00115413 0.143928 0.00065816 0.144582 0.891744 101.776 0.24217 0.765364 4.22421 0.0578304 0.039851 0.960149 0.0197587 0.00433566 0.0190216 0.00416176 0.00524128 0.00597844 0.209651 0.239138 58.004 -87.8965 126.262 15.962 145.021 0.000141154 0.267178 192.845 0.310499 0.0673627 0.00409631 0.000561899 0.00138354 0.986979 0.991728 -2.97938e-06 -85.6638 0.0930228 31185.1 303.06 0.983512 0.319146 0.732238 0.732233 9.99958 2.98291e-06 1.19315e-05 0.131589 0.982605 0.931722 -0.0132926 4.9093e-06 0.504741 -1.91976e-20 7.09015e-24 -1.91905e-20 0.00139564 0.997817 8.59651e-05 0.152622 2.85213 0.00139564 0.99782 0.730313 0.00105497 0.00188032 0.000859651 0.455549 0.00188032 0.439989 0.000129301 1.02 0.887976 0.534598 0.286463 1.71752e-07 3.06775e-09 2382.75 3114.28 -0.0553922 0.482154 0.277478 0.25318 -0.593392 -0.169528 0.496727 -0.26731 -0.229427 1.939 1 0 297.819 0 2.13194 1.937 0.000299764 0.853005 0.668073 0.361667 0.41737 2.13215 133.648 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.038 3.00627e-08 2.53909e-06 0.115201 0.1152 0.0120362 1.36649e-05 0.00115413 0.144002 0.000658161 0.144655 0.891818 101.775 0.242161 0.765475 4.22451 0.0578392 0.0398538 0.960146 0.0197584 0.00433593 0.0190212 0.00416198 0.0052416 0.00597877 0.209664 0.239151 58.004 -87.8965 126.262 15.962 145.021 0.000141154 0.267178 192.845 0.310498 0.0673627 0.00409631 0.0005619 0.00138354 0.986979 0.991728 -2.97939e-06 -85.6637 0.0930228 31185.1 303.067 0.983512 0.319146 0.732237 0.732233 9.99958 2.98292e-06 1.19316e-05 0.131592 0.982607 0.931723 -0.0132926 4.90933e-06 0.504752 -1.91986e-20 7.09057e-24 -1.91915e-20 0.00139564 0.997817 8.59651e-05 0.152622 2.85213 0.00139564 0.99782 0.730407 0.00105499 0.00188032 0.000859651 0.455548 0.00188032 0.439997 0.000129304 1.02 0.887977 0.534597 0.286464 1.71752e-07 3.06778e-09 2382.73 3114.28 -0.0553933 0.482154 0.277478 0.25318 -0.593392 -0.169528 0.496723 -0.267307 -0.229425 1.94 1 0 297.819 0 2.13209 1.938 0.000299763 0.853007 0.66812 0.361561 0.417395 2.1323 133.656 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.039 3.00916e-08 2.53909e-06 0.11526 0.115259 0.0120362 1.3678e-05 0.00115413 0.144075 0.000658163 0.144729 0.891891 101.775 0.242152 0.765585 4.22481 0.0578481 0.0398567 0.960143 0.0197581 0.00433619 0.0190209 0.0041622 0.00524193 0.00597909 0.209677 0.239164 58.0041 -87.8965 126.262 15.9619 145.021 0.000141154 0.267179 192.844 0.310498 0.0673626 0.00409631 0.0005619 0.00138355 0.986979 0.991728 -2.97941e-06 -85.6637 0.0930229 31185.1 303.074 0.983512 0.319146 0.732237 0.732233 9.99958 2.98292e-06 1.19316e-05 0.131594 0.98261 0.931723 -0.0132926 4.90936e-06 0.504763 -1.91996e-20 7.09099e-24 -1.91925e-20 0.00139564 0.997817 8.59652e-05 0.152622 2.85213 0.00139564 0.99782 0.730501 0.00105501 0.00188033 0.000859652 0.455548 0.00188032 0.440004 0.000129307 1.02 0.887978 0.534597 0.286466 1.71752e-07 3.0678e-09 2382.71 3114.28 -0.0553944 0.482154 0.277478 0.25318 -0.593392 -0.169528 0.496719 -0.267305 -0.229423 1.941 1 0 297.818 0 2.13224 1.939 0.000299763 0.853009 0.668167 0.361455 0.417421 2.13245 133.664 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.04 3.01206e-08 2.53909e-06 0.115319 0.115317 0.0120362 1.36912e-05 0.00115413 0.144148 0.000658164 0.144802 0.891965 101.775 0.242143 0.765696 4.22511 0.0578569 0.0398595 0.96014 0.0197577 0.00433645 0.0190206 0.00416243 0.00524225 0.00597942 0.20969 0.239177 58.0042 -87.8965 126.262 15.9619 145.021 0.000141154 0.267179 192.844 0.310498 0.0673625 0.00409632 0.000561901 0.00138355 0.986979 0.991728 -2.97942e-06 -85.6637 0.093023 31185.1 303.081 0.983512 0.319146 0.732237 0.732233 9.99958 2.98293e-06 1.19316e-05 0.131597 0.982613 0.931724 -0.0132926 4.90939e-06 0.504775 -1.92006e-20 7.0914e-24 -1.91935e-20 0.00139564 0.997817 8.59653e-05 0.152622 2.85213 0.00139564 0.99782 0.730595 0.00105503 0.00188033 0.000859653 0.455548 0.00188033 0.440011 0.00012931 1.02 0.887979 0.534597 0.286467 1.71752e-07 3.06782e-09 2382.7 3114.28 -0.0553956 0.482154 0.277477 0.25318 -0.593392 -0.169528 0.496714 -0.267303 -0.229421 1.942 1 0 297.817 0 2.13239 1.94 0.000299762 0.853012 0.668215 0.361349 0.417446 2.1326 133.672 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.041 3.01495e-08 2.53909e-06 0.115377 0.115376 0.0120362 1.37043e-05 0.00115413 0.144222 0.000658166 0.144875 0.892038 101.775 0.242134 0.765806 4.22541 0.0578657 0.0398624 0.960138 0.0197574 0.00433672 0.0190203 0.00416265 0.00524258 0.00597975 0.209703 0.23919 58.0042 -87.8965 126.262 15.9619 145.021 0.000141154 0.267179 192.844 0.310497 0.0673625 0.00409632 0.000561902 0.00138355 0.986979 0.991728 -2.97944e-06 -85.6637 0.0930231 31185 303.088 0.983512 0.319146 0.732237 0.732232 9.99958 2.98293e-06 1.19316e-05 0.1316 0.982616 0.931724 -0.0132926 4.90942e-06 0.504786 -1.92016e-20 7.09182e-24 -1.91945e-20 0.00139564 0.997817 8.59654e-05 0.152622 2.85213 0.00139564 0.99782 0.730688 0.00105505 0.00188033 0.000859654 0.455548 0.00188033 0.440019 0.000129313 1.02 0.88798 0.534596 0.286469 1.71753e-07 3.06784e-09 2382.68 3114.28 -0.0553967 0.482154 0.277477 0.25318 -0.593391 -0.169528 0.49671 -0.267301 -0.229418 1.943 1 0 297.817 0 2.13254 1.941 0.000299761 0.853014 0.668262 0.361244 0.417471 2.13275 133.68 83.9366 18.7218 60.874 0.00402464 0 -40 10
1.042 3.01784e-08 2.53909e-06 0.115436 0.115434 0.0120361 1.37174e-05 0.00115413 0.144295 0.000658167 0.144948 0.892112 101.774 0.242125 0.765917 4.22571 0.0578746 0.0398652 0.960135 0.0197571 0.00433698 0.0190199 0.00416287 0.00524291 0.00598007 0.209716 0.239203 58.0043 -87.8965 126.262 15.9618 145.021 0.000141154 0.267179 192.844 0.310497 0.0673624 0.00409632 0.000561902 0.00138355 0.986979 0.991728 -2.97945e-06 -85.6637 0.0930232 31185 303.096 0.983512 0.319146 0.732237 0.732232 9.99958 2.98294e-06 1.19316e-05 0.131602 0.982619 0.931725 -0.0132926 4.90945e-06 0.504797 -1.92026e-20 7.09224e-24 -1.91956e-20 0.00139564 0.997817 8.59655e-05 0.152623 2.85213 0.00139564 0.99782 0.730782 0.00105507 0.00188033 0.000859655 0.455548 0.00188033 0.440026 0.000129316 1.02 0.887981 0.534596 0.28647 1.71753e-07 3.06787e-09 2382.66 3114.27 -0.0553979 0.482154 0.277477 0.25318 -0.593391 -0.169528 0.496706 -0.267299 -0.229416 1.944 1 0 297.816 0 2.1327 1.942 0.000299761 0.853016 0.668309 0.361138 0.417496 2.1329 133.688 83.9366 18.7218 60.874 0.00402464 0 -40 10
1.043 3.02073e-08 2.5391e-06 0.115494 0.115493 0.0120361 1.37306e-05 0.00115413 0.144368 0.000658169 0.145022 0.892186 101.774 0.242117 0.766028 4.22602 0.0578834 0.0398681 0.960132 0.0197568 0.00433725 0.0190196 0.0041631 0.00524323 0.0059804 0.209729 0.239216 58.0044 -87.8965 126.262 15.9618 145.021 0.000141154 0.267179 192.844 0.310496 0.0673624 0.00409633 0.000561903 0.00138355 0.986979 0.991728 -2.97947e-06 -85.6637 0.0930233 31185 303.103 0.983512 0.319146 0.732237 0.732232 9.99958 2.98294e-06 1.19317e-05 0.131605 0.982621 0.931725 -0.0132926 4.90948e-06 0.504808 -1.92037e-20 7.09265e-24 -1.91966e-20 0.00139564 0.997817 8.59655e-05 0.152623 2.85213 0.00139564 0.99782 0.730876 0.00105509 0.00188033 0.000859655 0.455547 0.00188033 0.440034 0.000129319 1.02 0.887983 0.534596 0.286472 1.71753e-07 3.06789e-09 2382.65 3114.27 -0.0553991 0.482154 0.277477 0.25318 -0.593391 -0.169528 0.496701 -0.267297 -0.229414 1.945 1 0 297.815 0 2.13285 1.943 0.00029976 0.853019 0.668356 0.361033 0.417521 2.13305 133.697 83.9366 18.7218 60.8741 0.00402464 0 -40 10
1.044 3.02362e-08 2.5391e-06 0.115553 0.115551 0.0120361 1.37437e-05 0.00115413 0.144441 0.00065817 0.145095 0.892259 101.774 0.242108 0.766139 4.22632 0.0578923 0.0398709 0.960129 0.0197564 0.00433751 0.0190193 0.00416332 0.00524356 0.00598073 0.209742 0.239229 58.0044 -87.8965 126.262 15.9618 145.021 0.000141154 0.26718 192.844 0.310496 0.0673623 0.00409633 0.000561904 0.00138356 0.986979 0.991728 -2.97948e-06 -85.6637 0.0930234 31185 303.11 0.983512 0.319146 0.732237 0.732232 9.99958 2.98295e-06 1.19317e-05 0.131608 0.982624 0.931726 -0.0132926 4.90951e-06 0.50482 -1.92047e-20 7.09307e-24 -1.91976e-20 0.00139564 0.997817 8.59656e-05 0.152623 2.85213 0.00139564 0.99782 0.730969 0.00105511 0.00188033 0.000859656 0.455547 0.00188033 0.440041 0.000129322 1.02 0.887984 0.534595 0.286473 1.71753e-07 3.06791e-09 2382.63 3114.27 -0.0554003 0.482154 0.277476 0.25318 -0.593391 -0.169528 0.496697 -0.267295 -0.229411 1.946 1 0 297.814 0 2.133 1.944 0.00029976 0.853022 0.668403 0.360928 0.417546 2.1332 133.705 83.9366 18.7218 60.8741 0.00402464 0 -40 10
1.045 3.02651e-08 2.5391e-06 0.115611 0.11561 0.0120361 1.37569e-05 0.00115414 0.144514 0.000658172 0.145168 0.892333 101.773 0.242099 0.76625 4.22662 0.0579012 0.0398738 0.960126 0.0197561 0.00433778 0.0190189 0.00416354 0.00524389 0.00598106 0.209755 0.239242 58.0045 -87.8965 126.262 15.9617 145.021 0.000141154 0.26718 192.843 0.310495 0.0673623 0.00409633 0.000561904 0.00138356 0.986979 0.991728 -2.9795e-06 -85.6637 0.0930235 31184.9 303.117 0.983512 0.319146 0.732236 0.732232 9.99958 2.98295e-06 1.19317e-05 0.131611 0.982627 0.931726 -0.0132926 4.90954e-06 0.504831 -1.92057e-20 7.09349e-24 -1.91986e-20 0.00139565 0.997817 8.59657e-05 0.152623 2.85214 0.00139564 0.99782 0.731063 0.00105512 0.00188034 0.000859657 0.455547 0.00188033 0.440048 0.000129325 1.02 0.887985 0.534595 0.286475 1.71754e-07 3.06794e-09 2382.61 3114.27 -0.0554015 0.482154 0.277476 0.25318 -0.593391 -0.169528 0.496692 -0.267293 -0.229409 1.947 1 0 297.813 0 2.13315 1.945 0.000299759 0.853024 0.668451 0.360823 0.417571 2.13335 133.713 83.9366 18.7218 60.8741 0.00402464 0 -40 10
1.046 3.0294e-08 2.5391e-06 0.11567 0.115668 0.0120361 1.377e-05 0.00115414 0.144587 0.000658173 0.145241 0.892407 101.773 0.24209 0.76636 4.22693 0.05791 0.0398767 0.960123 0.0197558 0.00433805 0.0190186 0.00416377 0.00524421 0.00598139 0.209769 0.239256 58.0045 -87.8965 126.262 15.9617 145.021 0.000141154 0.26718 192.843 0.310495 0.0673622 0.00409634 0.000561905 0.00138356 0.986979 0.991728 -2.97951e-06 -85.6637 0.0930235 31184.9 303.124 0.983512 0.319146 0.732237 0.732232 9.99958 2.98296e-06 1.19317e-05 0.131613 0.98263 0.931727 -0.0132926 4.90957e-06 0.504842 -1.92067e-20 7.09391e-24 -1.91996e-20 0.00139565 0.997817 8.59658e-05 0.152623 2.85214 0.00139565 0.99782 0.731156 0.00105514 0.00188034 0.000859658 0.455547 0.00188034 0.440056 0.000129328 1.02 0.887986 0.534595 0.286476 1.71754e-07 3.06796e-09 2382.6 3114.27 -0.0554027 0.482154 0.277476 0.25318 -0.593391 -0.169528 0.496688 -0.267291 -0.229406 1.948 1 0 297.813 0 2.1333 1.946 0.000299758 0.853027 0.668498 0.360719 0.417596 2.1335 133.721 83.9366 18.7218 60.8741 0.00402464 0 -40 10
1.047 3.03229e-08 2.5391e-06 0.115728 0.115727 0.0120361 1.37832e-05 0.00115414 0.14466 0.000658175 0.145314 0.892481 101.773 0.242081 0.766471 4.22723 0.0579189 0.0398795 0.96012 0.0197555 0.00433831 0.0190183 0.00416399 0.00524454 0.00598172 0.209782 0.239269 58.0046 -87.8965 126.262 15.9616 145.021 0.000141154 0.26718 192.843 0.310495 0.0673622 0.00409634 0.000561906 0.00138356 0.986979 0.991728 -2.97953e-06 -85.6637 0.0930236 31184.9 303.132 0.983512 0.319146 0.732237 0.732232 9.99958 2.98296e-06 1.19317e-05 0.131616 0.982633 0.931727 -0.0132926 4.9096e-06 0.504853 -1.92077e-20 7.09433e-24 -1.92006e-20 0.00139565 0.997817 8.59659e-05 0.152623 2.85214 0.00139565 0.99782 0.73125 0.00105516 0.00188034 0.000859659 0.455546 0.00188034 0.440063 0.000129331 1.02 0.887987 0.534595 0.286478 1.71754e-07 3.06798e-09 2382.58 3114.27 -0.0554039 0.482154 0.277475 0.25318 -0.593391 -0.169529 0.496683 -0.267288 -0.229404 1.949 1 0 297.812 0 2.13345 1.947 0.000299758 0.85303 0.668545 0.360615 0.41762 2.13365 133.729 83.9366 18.7218 60.8741 0.00402464 0 -40 10
1.048 3.03519e-08 2.5391e-06 0.115786 0.115785 0.0120361 1.37963e-05 0.00115414 0.144733 0.000658176 0.145387 0.892555 101.772 0.242072 0.766582 4.22754 0.0579278 0.0398824 0.960118 0.0197551 0.00433858 0.019018 0.00416422 0.00524487 0.00598205 0.209795 0.239282 58.0047 -87.8965 126.262 15.9616 145.021 0.000141154 0.26718 192.843 0.310494 0.0673621 0.00409634 0.000561906 0.00138356 0.986979 0.991728 -2.97954e-06 -85.6637 0.0930237 31184.9 303.139 0.983512 0.319146 0.732237 0.732232 9.99958 2.98297e-06 1.19318e-05 0.131619 0.982635 0.931728 -0.0132926 4.90963e-06 0.504865 -1.92087e-20 7.09475e-24 -1.92016e-20 0.00139565 0.997817 8.59659e-05 0.152623 2.85214 0.00139565 0.99782 0.731343 0.00105518 0.00188034 0.000859659 0.455546 0.00188034 0.44007 0.000129334 1.02 0.887988 0.534594 0.286479 1.71754e-07 3.068e-09 2382.56 3114.27 -0.0554052 0.482155 0.277475 0.25318 -0.593391 -0.169529 0.496678 -0.267286 -0.229401 1.95 1 0 297.811 0 2.1336 1.948 0.000299757 0.853033 0.668592 0.36051 0.417645 2.1338 133.737 83.9366 18.7218 60.874 0.00402464 0 -40 10
1.049 3.03808e-08 2.5391e-06 0.115845 0.115843 0.0120361 1.38094e-05 0.00115414 0.144806 0.000658178 0.145459 0.892628 101.772 0.242063 0.766693 4.22784 0.0579366 0.0398853 0.960115 0.0197548 0.00433885 0.0190176 0.00416445 0.0052452 0.00598238 0.209808 0.239295 58.0047 -87.8965 126.262 15.9616 145.022 0.000141154 0.267181 192.843 0.310494 0.0673621 0.00409634 0.000561907 0.00138357 0.986979 0.991728 -2.97956e-06 -85.6636 0.0930238 31184.9 303.146 0.983512 0.319146 0.732237 0.732232 9.99958 2.98297e-06 1.19318e-05 0.131621 0.982638 0.931728 -0.0132926 4.90966e-06 0.504876 -1.92098e-20 7.09517e-24 -1.92027e-20 0.00139565 0.997817 8.5966e-05 0.152624 2.85214 0.00139565 0.99782 0.731437 0.0010552 0.00188034 0.00085966 0.455546 0.00188034 0.440078 0.000129337 1.02 0.887989 0.534594 0.286481 1.71755e-07 3.06803e-09 2382.55 3114.27 -0.0554065 0.482155 0.277475 0.25318 -0.593391 -0.169529 0.496673 -0.267284 -0.229399 1.951 1 0 297.81 0 2.13375 1.949 0.000299757 0.853036 0.668639 0.360406 0.41767 2.13396 133.745 83.9366 18.7218 60.874 0.00402464 0 -40 10
1.05 3.04097e-08 2.5391e-06 0.115903 0.115901 0.012036 1.38226e-05 0.00115414 0.144879 0.000658179 0.145532 0.892702 101.772 0.242054 0.766805 4.22815 0.0579455 0.0398882 0.960112 0.0197545 0.00433912 0.0190173 0.00416467 0.00524553 0.00598271 0.209821 0.239308 58.0048 -87.8965 126.262 15.9615 145.022 0.000141154 0.267181 192.843 0.310493 0.067362 0.00409635 0.000561908 0.00138357 0.986979 0.991728 -2.97957e-06 -85.6636 0.0930239 31184.8 303.153 0.983512 0.319146 0.732237 0.732233 9.99958 2.98298e-06 1.19318e-05 0.131624 0.982641 0.931728 -0.0132926 4.90969e-06 0.504887 -1.92108e-20 7.09559e-24 -1.92037e-20 0.00139565 0.997817 8.59661e-05 0.152624 2.85214 0.00139565 0.997819 0.73153 0.00105522 0.00188034 0.000859661 0.455546 0.00188034 0.440085 0.00012934 1.02 0.88799 0.534594 0.286482 1.71755e-07 3.06805e-09 2382.53 3114.27 -0.0554077 0.482155 0.277475 0.25318 -0.593391 -0.169529 0.496669 -0.267282 -0.229396 1.952 1 0 297.809 0 2.1339 1.95 0.000299756 0.853039 0.668686 0.360303 0.417695 2.13411 133.753 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.051 3.04386e-08 2.5391e-06 0.115961 0.11596 0.012036 1.38357e-05 0.00115414 0.144951 0.000658181 0.145605 0.892776 101.772 0.242046 0.766916 4.22845 0.0579544 0.0398911 0.960109 0.0197541 0.00433938 0.019017 0.0041649 0.00524586 0.00598304 0.209834 0.239322 58.0049 -87.8965 126.262 15.9615 145.022 0.000141154 0.267181 192.842 0.310493 0.067362 0.00409635 0.000561908 0.00138357 0.986979 0.991728 -2.97959e-06 -85.6636 0.093024 31184.8 303.161 0.983512 0.319146 0.732237 0.732233 9.99958 2.98298e-06 1.19318e-05 0.131627 0.982644 0.931729 -0.0132926 4.90972e-06 0.504899 -1.92118e-20 7.09601e-24 -1.92047e-20 0.00139565 0.997817 8.59662e-05 0.152624 2.85214 0.00139565 0.997819 0.731623 0.00105524 0.00188034 0.000859662 0.455546 0.00188034 0.440093 0.000129344 1.02 0.887991 0.534593 0.286484 1.71755e-07 3.06807e-09 2382.51 3114.27 -0.055409 0.482155 0.277474 0.25318 -0.593391 -0.169529 0.496664 -0.26728 -0.229393 1.953 1 0 297.808 0 2.13405 1.951 0.000299755 0.853042 0.668734 0.360199 0.41772 2.13426 133.761 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.052 3.04675e-08 2.5391e-06 0.116019 0.116018 0.012036 1.38489e-05 0.00115414 0.145024 0.000658182 0.145678 0.89285 101.771 0.242037 0.767027 4.22876 0.0579633 0.039894 0.960106 0.0197538 0.00433965 0.0190166 0.00416512 0.00524619 0.00598337 0.209847 0.239335 58.0049 -87.8965 126.262 15.9615 145.022 0.000141154 0.267181 192.842 0.310492 0.0673619 0.00409635 0.000561909 0.00138357 0.986979 0.991728 -2.9796e-06 -85.6636 0.0930241 31184.8 303.168 0.983512 0.319146 0.732238 0.732233 9.99958 2.98299e-06 1.19318e-05 0.13163 0.982646 0.931729 -0.0132926 4.90975e-06 0.50491 -1.92128e-20 7.09643e-24 -1.92057e-20 0.00139565 0.997817 8.59663e-05 0.152624 2.85214 0.00139565 0.997819 0.731717 0.00105525 0.00188035 0.000859663 0.455545 0.00188034 0.4401 0.000129347 1.02 0.887992 0.534593 0.286486 1.71756e-07 3.0681e-09 2382.5 3114.27 -0.0554103 0.482155 0.277474 0.25318 -0.593391 -0.169529 0.496659 -0.267278 -0.229391 1.954 1 0 297.807 0 2.1342 1.952 0.000299755 0.853046 0.668781 0.360096 0.417745 2.13441 133.769 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.053 3.04964e-08 2.5391e-06 0.116077 0.116076 0.012036 1.3862e-05 0.00115414 0.145097 0.000658184 0.14575 0.892924 101.771 0.242028 0.767138 4.22907 0.0579722 0.0398969 0.960103 0.0197535 0.00433992 0.0190163 0.00416535 0.00524652 0.00598371 0.209861 0.239348 58.005 -87.8965 126.262 15.9614 145.022 0.000141154 0.267181 192.842 0.310492 0.0673619 0.00409636 0.00056191 0.00138358 0.986979 0.991728 -2.97962e-06 -85.6636 0.0930241 31184.8 303.175 0.983512 0.319146 0.732238 0.732234 9.99958 2.98299e-06 1.19319e-05 0.131632 0.982649 0.93173 -0.0132926 4.90978e-06 0.504921 -1.92138e-20 7.09685e-24 -1.92067e-20 0.00139565 0.997817 8.59663e-05 0.152624 2.85214 0.00139565 0.997819 0.73181 0.00105527 0.00188035 0.000859663 0.455545 0.00188035 0.440107 0.00012935 1.02 0.887993 0.534593 0.286487 1.71756e-07 3.06812e-09 2382.48 3114.27 -0.0554117 0.482155 0.277474 0.25318 -0.593391 -0.169529 0.496654 -0.267276 -0.229388 1.955 1 0 297.806 0 2.13435 1.953 0.000299754 0.853049 0.668828 0.359992 0.41777 2.13456 133.777 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.054 3.05253e-08 2.5391e-06 0.116135 0.116134 0.012036 1.38751e-05 0.00115414 0.145169 0.000658185 0.145823 0.892998 101.771 0.242019 0.767249 4.22937 0.0579811 0.0398998 0.9601 0.0197532 0.00434019 0.019016 0.00416558 0.00524685 0.00598404 0.209874 0.239362 58.0051 -87.8965 126.262 15.9614 145.022 0.000141154 0.267182 192.842 0.310492 0.0673618 0.00409636 0.00056191 0.00138358 0.986979 0.991728 -2.97963e-06 -85.6636 0.0930242 31184.7 303.183 0.983512 0.319146 0.732238 0.732234 9.99958 2.983e-06 1.19319e-05 0.131635 0.982652 0.93173 -0.0132926 4.90981e-06 0.504933 -1.92149e-20 7.09727e-24 -1.92078e-20 0.00139566 0.997817 8.59664e-05 0.152624 2.85214 0.00139566 0.997819 0.731903 0.00105529 0.00188035 0.000859664 0.455545 0.00188035 0.440115 0.000129353 1.02 0.887995 0.534592 0.286489 1.71756e-07 3.06814e-09 2382.46 3114.27 -0.055413 0.482155 0.277473 0.25318 -0.593391 -0.169529 0.496649 -0.267274 -0.229385 1.956 1 0 297.806 0 2.1345 1.954 0.000299754 0.853053 0.668875 0.359889 0.417795 2.13471 133.785 83.9366 18.7218 60.874 0.00402465 0 -40 10
1.055 3.05542e-08 2.5391e-06 0.116193 0.116192 0.012036 1.38883e-05 0.00115414 0.145242 0.000658187 0.145895 0.893072 101.77 0.24201 0.767361 4.22968 0.05799 0.0399027 0.960097 0.0197528 0.00434046 0.0190156 0.0041658 0.00524718 0.00598437 0.209887 0.239375 58.0051 -87.8965 126.262 15.9613 145.022 0.000141154 0.267182 192.842 0.310491 0.0673618 0.00409636 0.000561911 0.00138358 0.986979 0.991728 -2.97965e-06 -85.6636 0.0930243 31184.7 303.19 0.983512 0.319146 0.732239 0.732234 9.99958 2.983e-06 1.19319e-05 0.131638 0.982654 0.931731 -0.0132926 4.90984e-06 0.504944 -1.92159e-20 7.09769e-24 -1.92088e-20 0.00139566 0.997817 8.59665e-05 0.152625 2.85214 0.00139566 0.997819 0.731996 0.00105531 0.00188035 0.000859665 0.455545 0.00188035 0.440122 0.000129356 1.02 0.887996 0.534592 0.28649 1.71756e-07 3.06816e-09 2382.45 3114.27 -0.0554143 0.482155 0.277473 0.25318 -0.593391 -0.169529 0.496644 -0.267272 -0.229382 1.957 1 0 297.805 0 2.13465 1.955 0.000299753 0.853056 0.668922 0.359787 0.41782 2.13486 133.793 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.056 3.05831e-08 2.53911e-06 0.116251 0.11625 0.012036 1.39014e-05 0.00115414 0.145314 0.000658188 0.145968 0.893147 101.77 0.242001 0.767472 4.22999 0.0579989 0.0399056 0.960094 0.0197525 0.00434073 0.0190153 0.00416603 0.00524751 0.0059847 0.2099 0.239388 58.0052 -87.8965 126.262 15.9613 145.022 0.000141155 0.267182 192.842 0.310491 0.0673617 0.00409637 0.000561912 0.00138358 0.986979 0.991728 -2.97966e-06 -85.6636 0.0930244 31184.7 303.197 0.983512 0.319146 0.732239 0.732235 9.99958 2.98301e-06 1.19319e-05 0.131641 0.982657 0.931731 -0.0132926 4.90987e-06 0.504956 -1.92169e-20 7.09811e-24 -1.92098e-20 0.00139566 0.997817 8.59666e-05 0.152625 2.85215 0.00139566 0.997819 0.73209 0.00105533 0.00188035 0.000859666 0.455544 0.00188035 0.440129 0.000129359 1.02 0.887997 0.534592 0.286492 1.71757e-07 3.06819e-09 2382.43 3114.27 -0.0554157 0.482155 0.277473 0.25318 -0.593391 -0.169529 0.496639 -0.267269 -0.229379 1.958 1 0 297.804 0 2.1348 1.956 0.000299752 0.85306 0.668969 0.359684 0.417845 2.13501 133.801 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.057 3.06121e-08 2.53911e-06 0.116309 0.116308 0.0120359 1.39146e-05 0.00115414 0.145386 0.00065819 0.14604 0.893221 101.77 0.241992 0.767584 4.2303 0.0580078 0.0399085 0.960092 0.0197522 0.004341 0.019015 0.00416626 0.00524784 0.00598504 0.209914 0.239402 58.0052 -87.8965 126.262 15.9613 145.022 0.000141155 0.267182 192.842 0.31049 0.0673617 0.00409637 0.000561912 0.00138358 0.986979 0.991728 -2.97968e-06 -85.6636 0.0930245 31184.7 303.205 0.983512 0.319146 0.73224 0.732235 9.99958 2.98301e-06 1.19319e-05 0.131643 0.98266 0.931731 -0.0132926 4.9099e-06 0.504967 -1.92179e-20 7.09853e-24 -1.92108e-20 0.00139566 0.997817 8.59667e-05 0.152625 2.85215 0.00139566 0.997819 0.732183 0.00105535 0.00188035 0.000859667 0.455544 0.00188035 0.440137 0.000129362 1.02 0.887998 0.534591 0.286493 1.71757e-07 3.06821e-09 2382.41 3114.28 -0.0554171 0.482155 0.277473 0.25318 -0.593391 -0.169529 0.496634 -0.267267 -0.229376 1.959 1 0 297.803 0 2.13495 1.957 0.000299752 0.853063 0.669016 0.359582 0.41787 2.13516 133.809 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.058 3.0641e-08 2.53911e-06 0.116367 0.116365 0.0120359 1.39277e-05 0.00115414 0.145459 0.000658191 0.146112 0.893295 101.769 0.241983 0.767695 4.23061 0.0580167 0.0399114 0.960089 0.0197518 0.00434127 0.0190146 0.00416649 0.00524817 0.00598537 0.209927 0.239415 58.0053 -87.8965 126.262 15.9612 145.022 0.000141155 0.267182 192.841 0.31049 0.0673616 0.00409637 0.000561913 0.00138359 0.986979 0.991728 -2.97969e-06 -85.6636 0.0930246 31184.7 303.212 0.983512 0.319146 0.73224 0.732236 9.99958 2.98301e-06 1.1932e-05 0.131646 0.982662 0.931732 -0.0132926 4.90992e-06 0.504979 -1.92189e-20 7.09895e-24 -1.92118e-20 0.00139566 0.997817 8.59668e-05 0.152625 2.85215 0.00139566 0.997819 0.732276 0.00105537 0.00188035 0.000859668 0.455544 0.00188035 0.440144 0.000129365 1.02 0.887999 0.534591 0.286495 1.71757e-07 3.06823e-09 2382.4 3114.28 -0.0554185 0.482155 0.277472 0.253181 -0.593391 -0.169529 0.496629 -0.267265 -0.229373 1.96 1 0 297.802 0 2.1351 1.958 0.000299751 0.853067 0.669063 0.359479 0.417895 2.13531 133.817 83.9365 18.7218 60.874 0.00402465 0 -40 10
1.059 3.06699e-08 2.53911e-06 0.116425 0.116423 0.0120359 1.39409e-05 0.00115414 0.145531 0.000658193 0.146184 0.893369 101.769 0.241974 0.767807 4.23092 0.0580257 0.0399143 0.960086 0.0197515 0.00434154 0.0190143 0.00416672 0.00524851 0.00598571 0.20994 0.239428 58.0054 -87.8965 126.262 15.9612 145.022 0.000141155 0.267182 192.841 0.310489 0.0673616 0.00409638 0.000561914 0.00138359 0.986979 0.991727 -2.97971e-06 -85.6636 0.0930247 31184.6 303.219 0.983512 0.319146 0.732241 0.732236 9.99958 2.98302e-06 1.1932e-05 0.131649 0.982665 0.931732 -0.0132926 4.90995e-06 0.50499 -1.922e-20 7.09937e-24 -1.92129e-20 0.00139566 0.997817 8.59668e-05 0.152625 2.85215 0.00139566 0.997819 0.732369 0.00105539 0.00188036 0.000859668 0.455544 0.00188035 0.440151 0.000129368 1.02 0.888 0.534591 0.286496 1.71757e-07 3.06826e-09 2382.38 3114.28 -0.0554199 0.482155 0.277472 0.253181 -0.593391 -0.169529 0.496624 -0.267263 -0.22937 1.961 1 0 297.801 0 2.13525 1.959 0.000299751 0.853071 0.66911 0.359377 0.41792 2.13546 133.826 83.9364 18.7218 60.874 0.00402465 0 -40 10
1.06 3.06988e-08 2.53911e-06 0.116482 0.116481 0.0120359 1.3954e-05 0.00115414 0.145603 0.000658194 0.146257 0.893443 101.769 0.241965 0.767918 4.23123 0.0580346 0.0399173 0.960083 0.0197512 0.00434181 0.019014 0.00416694 0.00524884 0.00598604 0.209954 0.239442 58.0054 -87.8965 126.262 15.9612 145.022 0.000141155 0.267183 192.841 0.310489 0.0673615 0.00409638 0.000561914 0.00138359 0.986979 0.991727 -2.97972e-06 -85.6635 0.0930248 31184.6 303.227 0.983512 0.319146 0.732241 0.732237 9.99958 2.98302e-06 1.1932e-05 0.131652 0.982668 0.931733 -0.0132926 4.90998e-06 0.505001 -1.9221e-20 7.0998e-24 -1.92139e-20 0.00139566 0.997817 8.59669e-05 0.152625 2.85215 0.00139566 0.997819 0.732462 0.0010554 0.00188036 0.000859669 0.455543 0.00188036 0.440159 0.000129371 1.02 0.888001 0.534591 0.286498 1.71758e-07 3.06828e-09 2382.36 3114.28 -0.0554213 0.482155 0.277472 0.253181 -0.593391 -0.169529 0.496619 -0.267261 -0.229367 1.962 1 0 297.8 0 2.1354 1.96 0.00029975 0.853075 0.669157 0.359276 0.417945 2.13561 133.834 83.9364 18.7218 60.8739 0.00402465 0 -40 10
1.061 3.07277e-08 2.53911e-06 0.11654 0.116539 0.0120359 1.39671e-05 0.00115414 0.145675 0.000658196 0.146329 0.893518 101.768 0.241956 0.76803 4.23154 0.0580435 0.0399202 0.96008 0.0197508 0.00434208 0.0190136 0.00416717 0.00524917 0.00598638 0.209967 0.239455 58.0055 -87.8965 126.262 15.9611 145.022 0.000141155 0.267183 192.841 0.310489 0.0673614 0.00409638 0.000561915 0.00138359 0.986979 0.991727 -2.97974e-06 -85.6635 0.0930248 31184.6 303.234 0.983512 0.319146 0.732242 0.732238 9.99958 2.98303e-06 1.1932e-05 0.131654 0.98267 0.931733 -0.0132926 4.91001e-06 0.505013 -1.9222e-20 7.10022e-24 -1.92149e-20 0.00139566 0.997817 8.5967e-05 0.152625 2.85215 0.00139566 0.997819 0.732555 0.00105542 0.00188036 0.00085967 0.455543 0.00188036 0.440166 0.000129374 1.02 0.888002 0.53459 0.286499 1.71758e-07 3.0683e-09 2382.35 3114.28 -0.0554227 0.482156 0.277471 0.253181 -0.593391 -0.169529 0.496614 -0.267259 -0.229364 1.963 1 0 297.799 0 2.13555 1.961 0.000299749 0.853079 0.669204 0.359174 0.417969 2.13576 133.842 83.9364 18.7218 60.8739 0.00402466 0 -40 10
1.062 3.07566e-08 2.53911e-06 0.116598 0.116596 0.0120359 1.39803e-05 0.00115414 0.145747 0.000658197 0.146401 0.893592 101.768 0.241948 0.768142 4.23185 0.0580525 0.0399231 0.960077 0.0197505 0.00434235 0.0190133 0.0041674 0.00524951 0.00598671 0.20998 0.239469 58.0056 -87.8965 126.262 15.9611 145.022 0.000141155 0.267183 192.841 0.310488 0.0673614 0.00409638 0.000561916 0.00138359 0.986979 0.991727 -2.97975e-06 -85.6635 0.0930249 31184.6 303.241 0.983512 0.319146 0.732243 0.732238 9.99958 2.98303e-06 1.1932e-05 0.131657 0.982673 0.931733 -0.0132926 4.91004e-06 0.505024 -1.9223e-20 7.10064e-24 -1.92159e-20 0.00139566 0.997817 8.59671e-05 0.152626 2.85215 0.00139566 0.997819 0.732648 0.00105544 0.00188036 0.000859671 0.455543 0.00188036 0.440173 0.000129377 1.02 0.888003 0.53459 0.286501 1.71758e-07 3.06832e-09 2382.33 3114.29 -0.0554241 0.482156 0.277471 0.253181 -0.593391 -0.16953 0.496609 -0.267257 -0.229361 1.964 1 0 297.798 0 2.1357 1.962 0.000299749 0.853083 0.669251 0.359073 0.417994 2.13591 133.85 83.9363 18.7218 60.8739 0.00402466 0 -40 10
1.063 3.07855e-08 2.53911e-06 0.116655 0.116654 0.0120359 1.39934e-05 0.00115414 0.145819 0.000658199 0.146473 0.893666 101.768 0.241939 0.768254 4.23216 0.0580614 0.0399261 0.960074 0.0197502 0.00434262 0.019013 0.00416763 0.00524984 0.00598705 0.209994 0.239482 58.0056 -87.8966 126.262 15.961 145.022 0.000141155 0.267183 192.841 0.310488 0.0673613 0.00409639 0.000561916 0.0013836 0.986978 0.991727 -2.97977e-06 -85.6635 0.093025 31184.5 303.249 0.983512 0.319146 0.732243 0.732239 9.99958 2.98304e-06 1.19321e-05 0.13166 0.982676 0.931734 -0.0132926 4.91007e-06 0.505036 -1.92241e-20 7.10107e-24 -1.9217e-20 0.00139567 0.997817 8.59672e-05 0.152626 2.85215 0.00139567 0.997819 0.732741 0.00105546 0.00188036 0.000859672 0.455543 0.00188036 0.440181 0.00012938 1.02 0.888004 0.53459 0.286502 1.71759e-07 3.06835e-09 2382.31 3114.29 -0.0554256 0.482156 0.277471 0.253181 -0.593391 -0.16953 0.496603 -0.267255 -0.229358 1.965 1 0 297.797 0 2.13585 1.963 0.000299748 0.853087 0.669298 0.358971 0.418019 2.13606 133.858 83.9363 18.7218 60.8739 0.00402466 0 -40 10
1.064 3.08144e-08 2.53911e-06 0.116713 0.116711 0.0120359 1.40066e-05 0.00115414 0.145891 0.0006582 0.146545 0.893741 101.768 0.24193 0.768365 4.23247 0.0580703 0.039929 0.960071 0.0197498 0.00434289 0.0190126 0.00416786 0.00525018 0.00598739 0.210007 0.239495 58.0057 -87.8966 126.262 15.961 145.022 0.000141155 0.267183 192.84 0.310487 0.0673613 0.00409639 0.000561917 0.0013836 0.986978 0.991727 -2.97978e-06 -85.6635 0.0930251 31184.5 303.256 0.983512 0.319146 0.732244 0.73224 9.99958 2.98304e-06 1.19321e-05 0.131663 0.982678 0.931734 -0.0132926 4.9101e-06 0.505047 -1.92251e-20 7.10149e-24 -1.9218e-20 0.00139567 0.997817 8.59672e-05 0.152626 2.85215 0.00139567 0.997819 0.732834 0.00105548 0.00188036 0.000859672 0.455543 0.00188036 0.440188 0.000129383 1.02 0.888006 0.534589 0.286504 1.71759e-07 3.06837e-09 2382.3 3114.29 -0.0554271 0.482156 0.277471 0.253182 -0.593391 -0.16953 0.496598 -0.267253 -0.229355 1.966 1 0 297.796 0 2.136 1.964 0.000299748 0.853092 0.669345 0.35887 0.418044 2.13621 133.866 83.9363 18.7218 60.8739 0.00402466 0 -40 10
1.065 3.08433e-08 2.53911e-06 0.11677 0.116769 0.0120358 1.40197e-05 0.00115414 0.145963 0.000658201 0.146617 0.893815 101.767 0.241921 0.768477 4.23279 0.0580793 0.039932 0.960068 0.0197495 0.00434317 0.0190123 0.00416809 0.00525051 0.00598772 0.21002 0.239509 58.0058 -87.8966 126.262 15.961 145.022 0.000141156 0.267184 192.84 0.310487 0.0673612 0.00409639 0.000561918 0.0013836 0.986978 0.991727 -2.9798e-06 -85.6635 0.0930252 31184.5 303.263 0.983511 0.319146 0.732245 0.732241 9.99958 2.98305e-06 1.19321e-05 0.131666 0.982681 0.931735 -0.0132926 4.91013e-06 0.505059 -1.92261e-20 7.10191e-24 -1.9219e-20 0.00139567 0.997817 8.59673e-05 0.152626 2.85215 0.00139567 0.997819 0.732927 0.0010555 0.00188036 0.000859673 0.455542 0.00188036 0.440195 0.000129386 1.02 0.888007 0.534589 0.286505 1.71759e-07 3.06839e-09 2382.28 3114.29 -0.0554285 0.482156 0.27747 0.253182 -0.59339 -0.16953 0.496593 -0.26725 -0.229352 1.967 1 0 297.795 0 2.13615 1.965 0.000299747 0.853096 0.669392 0.358769 0.418069 2.13636 133.874 83.9362 18.7218 60.8739 0.00402466 0 -40 10
1.066 3.08722e-08 2.53911e-06 0.116828 0.116826 0.0120358 1.40328e-05 0.00115414 0.146035 0.000658203 0.146688 0.89389 101.767 0.241912 0.768589 4.2331 0.0580882 0.0399349 0.960065 0.0197492 0.00434344 0.0190119 0.00416832 0.00525085 0.00598806 0.210034 0.239522 58.0058 -87.8966 126.262 15.9609 145.022 0.000141156 0.267184 192.84 0.310486 0.0673612 0.0040964 0.000561918 0.0013836 0.986978 0.991727 -2.97981e-06 -85.6635 0.0930253 31184.5 303.271 0.983511 0.319146 0.732246 0.732241 9.99958 2.98305e-06 1.19321e-05 0.131668 0.982683 0.931735 -0.0132926 4.91016e-06 0.505071 -1.92272e-20 7.10234e-24 -1.92201e-20 0.00139567 0.997817 8.59674e-05 0.152626 2.85215 0.00139567 0.997819 0.73302 0.00105552 0.00188037 0.000859674 0.455542 0.00188036 0.440202 0.000129389 1.02 0.888008 0.534589 0.286507 1.71759e-07 3.06842e-09 2382.26 3114.3 -0.05543 0.482156 0.27747 0.253182 -0.59339 -0.16953 0.496587 -0.267248 -0.229348 1.968 1 0 297.793 0 2.1363 1.966 0.000299746 0.8531 0.669439 0.358669 0.418094 2.13651 133.882 83.9362 18.7218 60.8738 0.00402466 0 -40 10
1.067 3.09012e-08 2.53911e-06 0.116885 0.116884 0.0120358 1.4046e-05 0.00115414 0.146107 0.000658204 0.14676 0.893964 101.767 0.241903 0.768701 4.23341 0.0580972 0.0399379 0.960062 0.0197488 0.00434371 0.0190116 0.00416855 0.00525118 0.0059884 0.210047 0.239536 58.0059 -87.8966 126.262 15.9609 145.022 0.000141156 0.267184 192.84 0.310486 0.0673611 0.0040964 0.000561919 0.00138361 0.986978 0.991727 -2.97983e-06 -85.6635 0.0930254 31184.5 303.278 0.983511 0.319146 0.732247 0.732242 9.99958 2.98306e-06 1.19321e-05 0.131671 0.982686 0.931735 -0.0132926 4.91019e-06 0.505082 -1.92282e-20 7.10276e-24 -1.92211e-20 0.00139567 0.997817 8.59675e-05 0.152626 2.85216 0.00139567 0.997819 0.733112 0.00105553 0.00188037 0.000859675 0.455542 0.00188037 0.44021 0.000129392 1.02 0.888009 0.534588 0.286508 1.7176e-07 3.06844e-09 2382.25 3114.3 -0.0554315 0.482156 0.27747 0.253182 -0.59339 -0.16953 0.496582 -0.267246 -0.229345 1.969 1 0 297.792 0 2.13645 1.967 0.000299746 0.853105 0.669486 0.358568 0.418119 2.13666 133.89 83.9361 18.7218 60.8738 0.00402466 0 -40 10
1.068 3.09301e-08 2.53911e-06 0.116943 0.116941 0.0120358 1.40591e-05 0.00115414 0.146178 0.000658206 0.146832 0.894039 101.766 0.241894 0.768813 4.23373 0.0581061 0.0399408 0.960059 0.0197485 0.00434399 0.0190113 0.00416878 0.00525152 0.00598874 0.210061 0.239549 58.0059 -87.8966 126.262 15.9608 145.022 0.000141156 0.267184 192.84 0.310486 0.0673611 0.0040964 0.00056192 0.00138361 0.986978 0.991727 -2.97984e-06 -85.6635 0.0930255 31184.4 303.286 0.983511 0.319146 0.732248 0.732243 9.99958 2.98306e-06 1.19321e-05 0.131674 0.982689 0.931736 -0.0132926 4.91022e-06 0.505094 -1.92292e-20 7.10319e-24 -1.92221e-20 0.00139567 0.997817 8.59676e-05 0.152627 2.85216 0.00139567 0.997819 0.733205 0.00105555 0.00188037 0.000859676 0.455542 0.00188037 0.440217 0.000129395 1.02 0.88801 0.534588 0.28651 1.7176e-07 3.06846e-09 2382.23 3114.3 -0.055433 0.482156 0.277469 0.253183 -0.59339 -0.16953 0.496576 -0.267244 -0.229342 1.97 1 0 297.791 0 2.1366 1.968 0.000299745 0.85311 0.669533 0.358468 0.418143 2.13681 133.898 83.9361 18.7218 60.8738 0.00402467 0 -40 10
1.069 3.0959e-08 2.53911e-06 0.117 0.116999 0.0120358 1.40723e-05 0.00115414 0.14625 0.000658207 0.146904 0.894113 101.766 0.241885 0.768925 4.23404 0.0581151 0.0399438 0.960056 0.0197481 0.00434426 0.0190109 0.00416901 0.00525185 0.00598907 0.210074 0.239563 58.006 -87.8966 126.262 15.9608 145.022 0.000141156 0.267184 192.84 0.310485 0.067361 0.00409641 0.00056192 0.00138361 0.986978 0.991727 -2.97986e-06 -85.6635 0.0930255 31184.4 303.293 0.983511 0.319146 0.732249 0.732244 9.99958 2.98307e-06 1.19322e-05 0.131677 0.982691 0.931736 -0.0132926 4.91025e-06 0.505105 -1.92303e-20 7.10361e-24 -1.92232e-20 0.00139567 0.997817 8.59676e-05 0.152627 2.85216 0.00139567 0.997819 0.733298 0.00105557 0.00188037 0.000859676 0.455541 0.00188037 0.440224 0.000129398 1.02 0.888011 0.534588 0.286511 1.7176e-07 3.06848e-09 2382.21 3114.31 -0.0554346 0.482156 0.277469 0.253183 -0.59339 -0.16953 0.496571 -0.267242 -0.229338 1.971 1 0 297.79 0 2.13675 1.969 0.000299745 0.853114 0.66958 0.358368 0.418168 2.13696 133.906 83.9361 18.7218 60.8738 0.00402467 0 -40 10
1.07 3.09879e-08 2.53912e-06 0.117057 0.117056 0.0120358 1.40854e-05 0.00115414 0.146322 0.000658209 0.146975 0.894188 101.766 0.241876 0.769037 4.23436 0.0581241 0.0399467 0.960053 0.0197478 0.00434453 0.0190106 0.00416925 0.00525219 0.00598941 0.210088 0.239577 58.0061 -87.8966 126.262 15.9608 145.022 0.000141157 0.267185 192.839 0.310485 0.067361 0.00409641 0.000561921 0.00138361 0.986978 0.991727 -2.97987e-06 -85.6634 0.0930256 31184.4 303.3 0.983511 0.319146 0.73225 0.732245 9.99958 2.98307e-06 1.19322e-05 0.13168 0.982694 0.931736 -0.0132926 4.91028e-06 0.505117 -1.92313e-20 7.10404e-24 -1.92242e-20 0.00139567 0.997817 8.59677e-05 0.152627 2.85216 0.00139567 0.997819 0.733391 0.00105559 0.00188037 0.000859677 0.455541 0.00188037 0.440232 0.000129401 1.02 0.888012 0.534587 0.286513 1.7176e-07 3.06851e-09 2382.2 3114.31 -0.0554361 0.482156 0.277469 0.253183 -0.59339 -0.16953 0.496565 -0.26724 -0.229335 1.972 1 0 297.789 0 2.1369 1.97 0.000299744 0.853119 0.669627 0.358268 0.418193 2.13711 133.914 83.936 18.7218 60.8737 0.00402467 0 -40 10
1.071 3.10168e-08 2.53912e-06 0.117115 0.117113 0.0120358 1.40985e-05 0.00115414 0.146393 0.00065821 0.147047 0.894262 101.765 0.241867 0.76915 4.23467 0.058133 0.0399497 0.96005 0.0197475 0.00434481 0.0190102 0.00416948 0.00525253 0.00598975 0.210101 0.23959 58.0061 -87.8966 126.262 15.9607 145.022 0.000141157 0.267185 192.839 0.310484 0.0673609 0.00409641 0.000561922 0.00138361 0.986978 0.991727 -2.97989e-06 -85.6634 0.0930257 31184.4 303.308 0.983511 0.319146 0.732251 0.732246 9.99958 2.98308e-06 1.19322e-05 0.131682 0.982696 0.931737 -0.0132926 4.91031e-06 0.505129 -1.92323e-20 7.10446e-24 -1.92252e-20 0.00139567 0.997817 8.59678e-05 0.152627 2.85216 0.00139567 0.997819 0.733483 0.00105561 0.00188037 0.000859678 0.455541 0.00188037 0.440239 0.000129404 1.02 0.888013 0.534587 0.286514 1.71761e-07 3.06853e-09 2382.18 3114.31 -0.0554377 0.482156 0.277469 0.253183 -0.59339 -0.16953 0.49656 -0.267238 -0.229331 1.973 1 0 297.788 0 2.13705 1.971 0.000299743 0.853124 0.669674 0.358168 0.418218 2.13726 133.922 83.936 18.7218 60.8737 0.00402467 0 -40 10
1.072 3.10457e-08 2.53912e-06 0.117172 0.11717 0.0120357 1.41117e-05 0.00115414 0.146465 0.000658212 0.147118 0.894337 101.765 0.241858 0.769262 4.23499 0.058142 0.0399527 0.960047 0.0197471 0.00434508 0.0190099 0.00416971 0.00525287 0.00599009 0.210115 0.239604 58.0062 -87.8966 126.262 15.9607 145.022 0.000141157 0.267185 192.839 0.310484 0.0673609 0.00409641 0.000561922 0.00138362 0.986978 0.991727 -2.9799e-06 -85.6634 0.0930258 31184.3 303.315 0.983511 0.319146 0.732252 0.732247 9.99958 2.98308e-06 1.19322e-05 0.131685 0.982699 0.931737 -0.0132926 4.91034e-06 0.50514 -1.92334e-20 7.10489e-24 -1.92263e-20 0.00139568 0.997817 8.59679e-05 0.152627 2.85216 0.00139568 0.997819 0.733576 0.00105563 0.00188038 0.000859679 0.455541 0.00188037 0.440246 0.000129407 1.02 0.888014 0.534587 0.286516 1.71761e-07 3.06855e-09 2382.16 3114.32 -0.0554392 0.482156 0.277468 0.253184 -0.59339 -0.16953 0.496554 -0.267236 -0.229328 1.974 1 0 297.787 0 2.1372 1.972 0.000299743 0.853129 0.669721 0.358069 0.418243 2.13741 133.93 83.9359 18.7218 60.8737 0.00402467 0 -40 10
1.073 3.10746e-08 2.53912e-06 0.117229 0.117227 0.0120357 1.41248e-05 0.00115414 0.146536 0.000658213 0.14719 0.894412 101.765 0.241849 0.769374 4.2353 0.058151 0.0399557 0.960044 0.0197468 0.00434536 0.0190096 0.00416994 0.0052532 0.00599043 0.210128 0.239617 58.0063 -87.8966 126.262 15.9607 145.022 0.000141157 0.267185 192.839 0.310483 0.0673608 0.00409642 0.000561923 0.00138362 0.986978 0.991727 -2.97992e-06 -85.6634 0.0930259 31184.3 303.323 0.983511 0.319146 0.732253 0.732248 9.99958 2.98309e-06 1.19322e-05 0.131688 0.982701 0.931737 -0.0132926 4.91037e-06 0.505152 -1.92344e-20 7.10531e-24 -1.92273e-20 0.00139568 0.997817 8.5968e-05 0.152627 2.85216 0.00139568 0.997819 0.733669 0.00105565 0.00188038 0.00085968 0.455541 0.00188038 0.440254 0.00012941 1.02 0.888015 0.534587 0.286517 1.71761e-07 3.06858e-09 2382.15 3114.32 -0.0554408 0.482156 0.277468 0.253184 -0.59339 -0.16953 0.496548 -0.267234 -0.229324 1.975 1 0 297.786 0 2.13735 1.973 0.000299742 0.853134 0.669768 0.357969 0.418268 2.13756 133.938 83.9358 18.7218 60.8737 0.00402468 0 -40 10
1.074 3.11035e-08 2.53912e-06 0.117286 0.117284 0.0120357 1.4138e-05 0.00115414 0.146607 0.000658214 0.147261 0.894486 101.764 0.24184 0.769486 4.23562 0.05816 0.0399587 0.960041 0.0197465 0.00434563 0.0190092 0.00417017 0.00525354 0.00599077 0.210142 0.239631 58.0063 -87.8966 126.262 15.9606 145.022 0.000141157 0.267185 192.839 0.310483 0.0673608 0.00409642 0.000561924 0.00138362 0.986978 0.991727 -2.97993e-06 -85.6634 0.093026 31184.3 303.33 0.983511 0.319146 0.732254 0.73225 9.99958 2.98309e-06 1.19323e-05 0.131691 0.982704 0.931738 -0.0132926 4.9104e-06 0.505163 -1.92354e-20 7.10574e-24 -1.92283e-20 0.00139568 0.997817 8.5968e-05 0.152627 2.85216 0.00139568 0.997819 0.733761 0.00105566 0.00188038 0.00085968 0.45554 0.00188038 0.440261 0.000129413 1.02 0.888016 0.534586 0.286519 1.71761e-07 3.0686e-09 2382.13 3114.33 -0.0554424 0.482157 0.277468 0.253184 -0.59339 -0.16953 0.496543 -0.267231 -0.229321 1.976 1 0 297.784 0 2.1375 1.974 0.000299742 0.853139 0.669815 0.35787 0.418292 2.13771 133.946 83.9358 18.7218 60.8736 0.00402468 0 -40 10
1.075 3.11324e-08 2.53912e-06 0.117343 0.117342 0.0120357 1.41511e-05 0.00115415 0.146679 0.000658216 0.147332 0.894561 101.764 0.241831 0.769599 4.23593 0.058169 0.0399617 0.960038 0.0197461 0.00434591 0.0190089 0.00417041 0.00525388 0.00599111 0.210155 0.239645 58.0064 -87.8966 126.261 15.9606 145.022 0.000141158 0.267186 192.839 0.310483 0.0673607 0.00409642 0.000561924 0.00138362 0.986978 0.991727 -2.97995e-06 -85.6634 0.0930261 31184.3 303.338 0.983511 0.319146 0.732255 0.732251 9.99958 2.9831e-06 1.19323e-05 0.131694 0.982706 0.931738 -0.0132926 4.91043e-06 0.505175 -1.92365e-20 7.10617e-24 -1.92294e-20 0.00139568 0.997817 8.59681e-05 0.152628 2.85216 0.00139568 0.997819 0.733854 0.00105568 0.00188038 0.000859681 0.45554 0.00188038 0.440268 0.000129416 1.02 0.888018 0.534586 0.28652 1.71762e-07 3.06862e-09 2382.11 3114.33 -0.055444 0.482157 0.277467 0.253185 -0.59339 -0.16953 0.496537 -0.267229 -0.229317 1.977 1 0 297.783 0 2.13765 1.975 0.000299741 0.853144 0.669862 0.357771 0.418317 2.13786 133.954 83.9357 18.7218 60.8736 0.00402468 0 -40 10
1.076 3.11613e-08 2.53912e-06 0.1174 0.117399 0.0120357 1.41642e-05 0.00115415 0.14675 0.000658217 0.147404 0.894636 101.764 0.241822 0.769711 4.23625 0.058178 0.0399646 0.960035 0.0197458 0.00434618 0.0190085 0.00417064 0.00525422 0.00599146 0.210169 0.239658 58.0064 -87.8966 126.261 15.9605 145.022 0.000141158 0.267186 192.838 0.310482 0.0673607 0.00409643 0.000561925 0.00138363 0.986978 0.991727 -2.97996e-06 -85.6634 0.0930261 31184.3 303.345 0.983511 0.319146 0.732256 0.732252 9.99958 2.9831e-06 1.19323e-05 0.131696 0.982709 0.931738 -0.0132926 4.91046e-06 0.505187 -1.92375e-20 7.1066e-24 -1.92304e-20 0.00139568 0.997817 8.59682e-05 0.152628 2.85216 0.00139568 0.997819 0.733946 0.0010557 0.00188038 0.000859682 0.45554 0.00188038 0.440275 0.000129419 1.02 0.888019 0.534586 0.286522 1.71762e-07 3.06864e-09 2382.1 3114.33 -0.0554456 0.482157 0.277467 0.253185 -0.59339 -0.16953 0.496531 -0.267227 -0.229313 1.978 1 0 297.782 0 2.1378 1.976 0.00029974 0.853149 0.669908 0.357672 0.418342 2.13801 133.962 83.9357 18.7218 60.8736 0.00402468 0 -40 10
1.077 3.11902e-08 2.53912e-06 0.117457 0.117456 0.0120357 1.41774e-05 0.00115415 0.146821 0.000658219 0.147475 0.894711 101.763 0.241813 0.769824 4.23657 0.058187 0.0399676 0.960032 0.0197454 0.00434646 0.0190082 0.00417087 0.00525456 0.0059918 0.210182 0.239672 58.0065 -87.8966 126.261 15.9605 145.022 0.000141158 0.267186 192.838 0.310482 0.0673606 0.00409643 0.000561926 0.00138363 0.986978 0.991727 -2.97998e-06 -85.6634 0.0930262 31184.2 303.353 0.983511 0.319146 0.732258 0.732253 9.99958 2.98311e-06 1.19323e-05 0.131699 0.982711 0.931739 -0.0132926 4.91049e-06 0.505199 -1.92385e-20 7.10702e-24 -1.92314e-20 0.00139568 0.997817 8.59683e-05 0.152628 2.85217 0.00139568 0.997819 0.734039 0.00105572 0.00188038 0.000859683 0.45554 0.00188038 0.440283 0.000129422 1.02 0.88802 0.534585 0.286523 1.71762e-07 3.06867e-09 2382.08 3114.34 -0.0554472 0.482157 0.277467 0.253185 -0.593389 -0.16953 0.496525 -0.267225 -0.22931 1.979 1 0 297.781 0 2.13795 1.977 0.00029974 0.853154 0.669955 0.357574 0.418367 2.13816 133.97 83.9356 18.7218 60.8735 0.00402469 0 -40 10
1.078 3.12192e-08 2.53912e-06 0.117514 0.117512 0.0120357 1.41905e-05 0.00115415 0.146892 0.00065822 0.147546 0.894786 101.763 0.241804 0.769936 4.23689 0.058196 0.0399706 0.960029 0.0197451 0.00434674 0.0190079 0.00417111 0.0052549 0.00599214 0.210196 0.239686 58.0066 -87.8966 126.261 15.9605 145.022 0.000141158 0.267186 192.838 0.310481 0.0673606 0.00409643 0.000561926 0.00138363 0.986978 0.991727 -2.97999e-06 -85.6634 0.0930263 31184.2 303.36 0.983511 0.319146 0.732259 0.732255 9.99958 2.98311e-06 1.19323e-05 0.131702 0.982714 0.931739 -0.0132926 4.91052e-06 0.50521 -1.92396e-20 7.10745e-24 -1.92325e-20 0.00139568 0.997817 8.59684e-05 0.152628 2.85217 0.00139568 0.997819 0.734131 0.00105574 0.00188038 0.000859684 0.455539 0.00188038 0.44029 0.000129425 1.02 0.888021 0.534585 0.286525 1.71763e-07 3.06869e-09 2382.06 3114.34 -0.0554489 0.482157 0.277467 0.253186 -0.593389 -0.169531 0.49652 -0.267223 -0.229306 1.98 1 0 297.78 0 2.1381 1.978 0.000299739 0.85316 0.670002 0.357475 0.418392 2.1383 133.978 83.9355 18.7218 60.8735 0.00402469 0 -40 10
1.079 3.12481e-08 2.53912e-06 0.117571 0.117569 0.0120356 1.42037e-05 0.00115415 0.146963 0.000658222 0.147617 0.89486 101.763 0.241795 0.770049 4.23721 0.058205 0.0399736 0.960026 0.0197448 0.00434701 0.0190075 0.00417134 0.00525524 0.00599248 0.21021 0.239699 58.0066 -87.8966 126.261 15.9604 145.022 0.000141159 0.267186 192.838 0.310481 0.0673605 0.00409644 0.000561927 0.00138363 0.986978 0.991727 -2.98001e-06 -85.6634 0.0930264 31184.2 303.368 0.983511 0.319146 0.73226 0.732256 9.99958 2.98312e-06 1.19324e-05 0.131705 0.982716 0.931739 -0.0132926 4.91055e-06 0.505222 -1.92406e-20 7.10788e-24 -1.92335e-20 0.00139568 0.997817 8.59684e-05 0.152628 2.85217 0.00139568 0.997819 0.734224 0.00105576 0.00188039 0.000859684 0.455539 0.00188038 0.440297 0.000129428 1.02 0.888022 0.534585 0.286527 1.71763e-07 3.06871e-09 2382.05 3114.35 -0.0554505 0.482157 0.277466 0.253186 -0.593389 -0.169531 0.496514 -0.267221 -0.229302 1.981 1 0 297.778 0 2.13825 1.979 0.000299739 0.853165 0.670049 0.357377 0.418416 2.13845 133.986 83.9355 18.7218 60.8735 0.00402469 0 -40 10
1.08 3.1277e-08 2.53912e-06 0.117628 0.117626 0.0120356 1.42168e-05 0.00115415 0.147034 0.000658223 0.147688 0.894935 101.762 0.241786 0.770161 4.23753 0.058214 0.0399767 0.960023 0.0197444 0.00434729 0.0190072 0.00417157 0.00525558 0.00599282 0.210223 0.239713 58.0067 -87.8966 126.261 15.9604 145.022 0.000141159 0.267186 192.838 0.31048 0.0673605 0.00409644 0.000561928 0.00138363 0.986978 0.991727 -2.98002e-06 -85.6634 0.0930265 31184.2 303.375 0.983511 0.319146 0.732262 0.732257 9.99958 2.98312e-06 1.19324e-05 0.131708 0.982719 0.93174 -0.0132926 4.91058e-06 0.505234 -1.92417e-20 7.10831e-24 -1.92346e-20 0.00139569 0.997817 8.59685e-05 0.152628 2.85217 0.00139568 0.997819 0.734316 0.00105578 0.00188039 0.000859685 0.455539 0.00188039 0.440304 0.000129431 1.02 0.888023 0.534584 0.286528 1.71763e-07 3.06874e-09 2382.03 3114.35 -0.0554522 0.482157 0.277466 0.253186 -0.593389 -0.169531 0.496508 -0.267219 -0.229298 1.982 1 0 297.777 0 2.1384 1.98 0.000299738 0.853171 0.670096 0.357279 0.418441 2.1386 133.994 83.9354 18.7218 60.8735 0.0040247 0 -40 10
1.081 3.13059e-08 2.53912e-06 0.117684 0.117683 0.0120356 1.42299e-05 0.00115415 0.147105 0.000658224 0.147759 0.89501 101.762 0.241777 0.770274 4.23784 0.058223 0.0399797 0.96002 0.0197441 0.00434757 0.0190068 0.00417181 0.00525592 0.00599317 0.210237 0.239727 58.0068 -87.8966 126.261 15.9604 145.022 0.000141159 0.267187 192.838 0.31048 0.0673604 0.00409644 0.000561928 0.00138364 0.986978 0.991727 -2.98004e-06 -85.6633 0.0930266 31184.1 303.383 0.983511 0.319146 0.732263 0.732259 9.99958 2.98313e-06 1.19324e-05 0.131711 0.982721 0.93174 -0.0132926 4.91061e-06 0.505245 -1.92427e-20 7.10873e-24 -1.92356e-20 0.00139569 0.997817 8.59686e-05 0.152629 2.85217 0.00139569 0.997819 0.734409 0.00105579 0.00188039 0.000859686 0.455539 0.00188039 0.440312 0.000129434 1.02 0.888024 0.534584 0.28653 1.71763e-07 3.06876e-09 2382.01 3114.36 -0.0554539 0.482157 0.277466 0.253187 -0.593389 -0.169531 0.496502 -0.267217 -0.229295 1.983 1 0 297.776 0 2.13855 1.981 0.000299737 0.853176 0.670143 0.357181 0.418466 2.13875 134.002 83.9353 18.7217 60.8734 0.0040247 0 -40 10
1.082 3.13348e-08 2.53912e-06 0.117741 0.11774 0.0120356 1.42431e-05 0.00115415 0.147176 0.000658226 0.14783 0.895085 101.762 0.241768 0.770387 4.23816 0.058232 0.0399827 0.960017 0.0197437 0.00434784 0.0190065 0.00417204 0.00525626 0.00599351 0.210251 0.23974 58.0068 -87.8966 126.261 15.9603 145.022 0.000141159 0.267187 192.837 0.31048 0.0673603 0.00409644 0.000561929 0.00138364 0.986978 0.991727 -2.98005e-06 -85.6633 0.0930267 31184.1 303.39 0.983511 0.319146 0.732265 0.73226 9.99958 2.98313e-06 1.19324e-05 0.131713 0.982724 0.93174 -0.0132926 4.91064e-06 0.505257 -1.92438e-20 7.10916e-24 -1.92366e-20 0.00139569 0.997817 8.59687e-05 0.152629 2.85217 0.00139569 0.997819 0.734501 0.00105581 0.00188039 0.000859687 0.455539 0.00188039 0.440319 0.000129437 1.02 0.888025 0.534584 0.286531 1.71764e-07 3.06878e-09 2382 3114.36 -0.0554555 0.482157 0.277465 0.253187 -0.593389 -0.169531 0.496496 -0.267215 -0.229291 1.984 1 0 297.775 0 2.1387 1.982 0.000299737 0.853182 0.670189 0.357084 0.418491 2.1389 134.01 83.9353 18.7217 60.8734 0.0040247 0 -40 10
1.083 3.13637e-08 2.53913e-06 0.117798 0.117796 0.0120356 1.42562e-05 0.00115415 0.147247 0.000658227 0.147901 0.89516 101.762 0.241759 0.7705 4.23848 0.058241 0.0399857 0.960014 0.0197434 0.00434812 0.0190061 0.00417228 0.00525661 0.00599386 0.210264 0.239754 58.0069 -87.8966 126.261 15.9603 145.022 0.00014116 0.267187 192.837 0.310479 0.0673603 0.00409645 0.00056193 0.00138364 0.986978 0.991727 -2.98007e-06 -85.6633 0.0930268 31184.1 303.398 0.983511 0.319146 0.732266 0.732262 9.99958 2.98314e-06 1.19324e-05 0.131716 0.982726 0.93174 -0.0132926 4.91066e-06 0.505269 -1.92448e-20 7.10959e-24 -1.92377e-20 0.00139569 0.997817 8.59688e-05 0.152629 2.85217 0.00139569 0.997819 0.734593 0.00105583 0.00188039 0.000859688 0.455538 0.00188039 0.440326 0.00012944 1.02 0.888026 0.534584 0.286533 1.71764e-07 3.0688e-09 2381.98 3114.37 -0.0554572 0.482157 0.277465 0.253188 -0.593389 -0.169531 0.49649 -0.267212 -0.229287 1.985 1 0 297.773 0 2.13885 1.983 0.000299736 0.853188 0.670236 0.356986 0.418515 2.13905 134.018 83.9352 18.7217 60.8733 0.0040247 0 -40 10
1.084 3.13926e-08 2.53913e-06 0.117854 0.117853 0.0120356 1.42694e-05 0.00115415 0.147318 0.000658229 0.147972 0.895235 101.761 0.24175 0.770612 4.23881 0.05825 0.0399887 0.960011 0.0197431 0.0043484 0.0190058 0.00417251 0.00525695 0.0059942 0.210278 0.239768 58.007 -87.8966 126.261 15.9602 145.022 0.00014116 0.267187 192.837 0.310479 0.0673602 0.00409645 0.00056193 0.00138364 0.986978 0.991727 -2.98008e-06 -85.6633 0.0930268 31184.1 303.405 0.983511 0.319146 0.732268 0.732263 9.99958 2.98314e-06 1.19325e-05 0.131719 0.982729 0.931741 -0.0132926 4.91069e-06 0.505281 -1.92458e-20 7.11002e-24 -1.92387e-20 0.00139569 0.997817 8.59688e-05 0.152629 2.85217 0.00139569 0.997819 0.734685 0.00105585 0.00188039 0.000859688 0.455538 0.00188039 0.440333 0.000129443 1.02 0.888027 0.534583 0.286534 1.71764e-07 3.06883e-09 2381.96 3114.38 -0.055459 0.482157 0.277465 0.253188 -0.593389 -0.169531 0.496484 -0.26721 -0.229283 1.986 1 0 297.772 0 2.139 1.984 0.000299735 0.853194 0.670283 0.356889 0.41854 2.1392 134.026 83.9351 18.7217 60.8733 0.00402471 0 -40 10
1.085 3.14215e-08 2.53913e-06 0.117911 0.11791 0.0120356 1.42825e-05 0.00115415 0.147389 0.00065823 0.148042 0.89531 101.761 0.241741 0.770725 4.23913 0.0582591 0.0399918 0.960008 0.0197427 0.00434868 0.0190055 0.00417275 0.00525729 0.00599455 0.210292 0.239782 58.007 -87.8966 126.261 15.9602 145.022 0.00014116 0.267187 192.837 0.310478 0.0673602 0.00409645 0.000561931 0.00138364 0.986978 0.991727 -2.9801e-06 -85.6633 0.0930269 31184.1 303.413 0.983511 0.319146 0.732269 0.732265 9.99958 2.98315e-06 1.19325e-05 0.131722 0.982731 0.931741 -0.0132926 4.91072e-06 0.505293 -1.92469e-20 7.11045e-24 -1.92398e-20 0.00139569 0.997817 8.59689e-05 0.152629 2.85217 0.00139569 0.997819 0.734778 0.00105587 0.00188039 0.000859689 0.455538 0.00188039 0.440341 0.000129446 1.02 0.888029 0.534583 0.286536 1.71764e-07 3.06885e-09 2381.95 3114.38 -0.0554607 0.482157 0.277465 0.253188 -0.593389 -0.169531 0.496478 -0.267208 -0.229279 1.987 1 0 297.771 0 2.13915 1.985 0.000299735 0.8532 0.67033 0.356792 0.418565 2.13935 134.034 83.935 18.7217 60.8733 0.00402471 0 -40 10
1.086 3.14504e-08 2.53913e-06 0.117968 0.117966 0.0120356 1.42956e-05 0.00115415 0.147459 0.000658231 0.148113 0.895386 101.761 0.241732 0.770838 4.23945 0.0582681 0.0399948 0.960005 0.0197424 0.00434896 0.0190051 0.00417298 0.00525763 0.00599489 0.210305 0.239796 58.0071 -87.8966 126.261 15.9602 145.022 0.000141161 0.267188 192.837 0.310478 0.0673601 0.00409646 0.000561932 0.00138365 0.986978 0.991727 -2.98011e-06 -85.6633 0.093027 31184 303.42 0.983511 0.319146 0.732271 0.732266 9.99958 2.98315e-06 1.19325e-05 0.131725 0.982734 0.931741 -0.0132926 4.91075e-06 0.505304 -1.92479e-20 7.11088e-24 -1.92408e-20 0.00139569 0.997817 8.5969e-05 0.152629 2.85217 0.00139569 0.997819 0.73487 0.00105589 0.0018804 0.00085969 0.455538 0.00188039 0.440348 0.000129449 1.02 0.88803 0.534583 0.286537 1.71765e-07 3.06887e-09 2381.93 3114.39 -0.0554624 0.482157 0.277464 0.253189 -0.593389 -0.169531 0.496472 -0.267206 -0.229275 1.988 1 0 297.769 0 2.1393 1.986 0.000299734 0.853205 0.670377 0.356695 0.41859 2.1395 134.042 83.935 18.7217 60.8732 0.00402471 0 -40 10
1.087 3.14793e-08 2.53913e-06 0.118024 0.118023 0.0120355 1.43088e-05 0.00115415 0.14753 0.000658233 0.148184 0.895461 101.76 0.241723 0.770951 4.23977 0.0582771 0.0399978 0.960002 0.019742 0.00434924 0.0190048 0.00417322 0.00525798 0.00599524 0.210319 0.239809 58.0071 -87.8966 126.261 15.9601 145.022 0.000141161 0.267188 192.837 0.310477 0.0673601 0.00409646 0.000561932 0.00138365 0.986978 0.991727 -2.98013e-06 -85.6633 0.0930271 31184 303.428 0.983511 0.319146 0.732272 0.732268 9.99958 2.98316e-06 1.19325e-05 0.131728 0.982736 0.931742 -0.0132926 4.91078e-06 0.505316 -1.9249e-20 7.11131e-24 -1.92419e-20 0.00139569 0.997817 8.59691e-05 0.152629 2.85217 0.00139569 0.997819 0.734962 0.00105591 0.0018804 0.000859691 0.455537 0.0018804 0.440355 0.000129452 1.02 0.888031 0.534582 0.286539 1.71765e-07 3.06889e-09 2381.91 3114.39 -0.0554642 0.482157 0.277464 0.253189 -0.593388 -0.169531 0.496465 -0.267204 -0.229271 1.989 1 0 297.768 0 2.13945 1.987 0.000299734 0.853212 0.670423 0.356598 0.418614 2.13965 134.05 83.9349 18.7217 60.8732 0.00402472 0 -40 10
1.088 3.15082e-08 2.53913e-06 0.11808 0.118079 0.0120355 1.43219e-05 0.00115415 0.147601 0.000658234 0.148254 0.895536 101.76 0.241714 0.771064 4.24009 0.0582862 0.0400009 0.959999 0.0197417 0.00434952 0.0190044 0.00417346 0.00525832 0.00599558 0.210333 0.239823 58.0072 -87.8966 126.261 15.9601 145.022 0.000141161 0.267188 192.836 0.310477 0.06736 0.00409646 0.000561933 0.00138365 0.986978 0.991727 -2.98014e-06 -85.6633 0.0930272 31184 303.436 0.983511 0.319146 0.732274 0.73227 9.99958 2.98316e-06 1.19325e-05 0.13173 0.982739 0.931742 -0.0132926 4.91081e-06 0.505328 -1.925e-20 7.11174e-24 -1.92429e-20 0.00139569 0.997817 8.59692e-05 0.15263 2.85218 0.00139569 0.997819 0.735054 0.00105592 0.0018804 0.000859692 0.455537 0.0018804 0.440362 0.000129455 1.02 0.888032 0.534582 0.28654 1.71765e-07 3.06892e-09 2381.9 3114.4 -0.0554659 0.482158 0.277464 0.25319 -0.593388 -0.169531 0.496459 -0.267202 -0.229267 1.99 1 0 297.767 0 2.1396 1.988 0.000299733 0.853218 0.67047 0.356501 0.418639 2.1398 134.058 83.9348 18.7217 60.8732 0.00402472 0 -40 10
1.089 3.15371e-08 2.53913e-06 0.118137 0.118135 0.0120355 1.43351e-05 0.00115415 0.147671 0.000658236 0.148325 0.895611 101.76 0.241705 0.771177 4.24042 0.0582952 0.0400039 0.959996 0.0197413 0.0043498 0.0190041 0.00417369 0.00525866 0.00599593 0.210347 0.239837 58.0073 -87.8967 126.261 15.9601 145.022 0.000141162 0.267188 192.836 0.310477 0.06736 0.00409647 0.000561934 0.00138365 0.986978 0.991727 -2.98016e-06 -85.6633 0.0930273 31184 303.443 0.983511 0.319146 0.732276 0.732271 9.99958 2.98317e-06 1.19326e-05 0.131733 0.982741 0.931742 -0.0132926 4.91084e-06 0.50534 -1.92511e-20 7.11217e-24 -1.9244e-20 0.0013957 0.997817 8.59692e-05 0.15263 2.85218 0.0013957 0.997819 0.735146 0.00105594 0.0018804 0.000859692 0.455537 0.0018804 0.44037 0.000129458 1.02 0.888033 0.534582 0.286542 1.71765e-07 3.06894e-09 2381.88 3114.41 -0.0554677 0.482158 0.277463 0.25319 -0.593388 -0.169531 0.496453 -0.2672 -0.229263 1.991 1 0 297.765 0 2.13974 1.989 0.000299732 0.853224 0.670517 0.356405 0.418664 2.13995 134.066 83.9347 18.7217 60.8731 0.00402472 0 -40 10
1.09 3.15661e-08 2.53913e-06 0.118193 0.118192 0.0120355 1.43482e-05 0.00115415 0.147742 0.000658237 0.148395 0.895686 101.759 0.241696 0.77129 4.24074 0.0583043 0.040007 0.959993 0.019741 0.00435008 0.0190037 0.00417393 0.00525901 0.00599628 0.21036 0.239851 58.0073 -87.8967 126.261 15.96 145.022 0.000141162 0.267188 192.836 0.310476 0.0673599 0.00409647 0.000561934 0.00138366 0.986978 0.991727 -2.98017e-06 -85.6633 0.0930274 31183.9 303.451 0.983511 0.319146 0.732278 0.732273 9.99958 2.98317e-06 1.19326e-05 0.131736 0.982743 0.931742 -0.0132926 4.91087e-06 0.505352 -1.92521e-20 7.1126e-24 -1.9245e-20 0.0013957 0.997817 8.59693e-05 0.15263 2.85218 0.0013957 0.997819 0.735238 0.00105596 0.0018804 0.000859693 0.455537 0.0018804 0.440377 0.000129461 1.02 0.888034 0.534581 0.286543 1.71766e-07 3.06896e-09 2381.86 3114.41 -0.0554695 0.482158 0.277463 0.253191 -0.593388 -0.169531 0.496447 -0.267198 -0.229258 1.992 1 0 297.764 0 2.13989 1.99 0.000299732 0.85323 0.670564 0.356308 0.418688 2.1401 134.074 83.9346 18.7217 60.8731 0.00402473 0 -40 10
1.091 3.1595e-08 2.53913e-06 0.11825 0.118248 0.0120355 1.43613e-05 0.00115415 0.147812 0.000658238 0.148466 0.895762 101.759 0.241687 0.771403 4.24106 0.0583133 0.04001 0.95999 0.0197406 0.00435036 0.0190034 0.00417417 0.00525935 0.00599662 0.210374 0.239865 58.0074 -87.8967 126.261 15.96 145.022 0.000141162 0.267189 192.836 0.310476 0.0673599 0.00409647 0.000561935 0.00138366 0.986978 0.991727 -2.98019e-06 -85.6633 0.0930275 31183.9 303.458 0.983511 0.319146 0.732279 0.732275 9.99958 2.98318e-06 1.19326e-05 0.131739 0.982746 0.931743 -0.0132926 4.9109e-06 0.505364 -1.92532e-20 7.11304e-24 -1.92461e-20 0.0013957 0.997817 8.59694e-05 0.15263 2.85218 0.0013957 0.997819 0.735331 0.00105598 0.0018804 0.000859694 0.455536 0.0018804 0.440384 0.000129464 1.02 0.888035 0.534581 0.286545 1.71766e-07 3.06899e-09 2381.85 3114.42 -0.0554713 0.482158 0.277463 0.253191 -0.593388 -0.169531 0.49644 -0.267196 -0.229254 1.993 1 0 297.763 0 2.14004 1.991 0.000299731 0.853236 0.67061 0.356212 0.418713 2.14025 134.082 83.9345 18.7217 60.873 0.00402473 0 -40 10
1.092 3.16239e-08 2.53913e-06 0.118306 0.118304 0.0120355 1.43745e-05 0.00115415 0.147882 0.00065824 0.148536 0.895837 101.759 0.241678 0.771517 4.24139 0.0583224 0.0400131 0.959987 0.0197403 0.00435064 0.019003 0.0041744 0.0052597 0.00599697 0.210388 0.239879 58.0075 -87.8967 126.261 15.9599 145.022 0.000141163 0.267189 192.836 0.310475 0.0673598 0.00409648 0.000561936 0.00138366 0.986978 0.991727 -2.9802e-06 -85.6632 0.0930275 31183.9 303.466 0.983511 0.319146 0.732281 0.732277 9.99958 2.98318e-06 1.19326e-05 0.131742 0.982748 0.931743 -0.0132926 4.91093e-06 0.505376 -1.92542e-20 7.11347e-24 -1.92471e-20 0.0013957 0.997817 8.59695e-05 0.15263 2.85218 0.0013957 0.997819 0.735423 0.001056 0.0018804 0.000859695 0.455536 0.0018804 0.440391 0.000129467 1.02 0.888036 0.534581 0.286546 1.71766e-07 3.06901e-09 2381.83 3114.43 -0.0554731 0.482158 0.277463 0.253192 -0.593388 -0.169531 0.496434 -0.267193 -0.22925 1.994 1 0 297.761 0 2.14019 1.992 0.00029973 0.853243 0.670657 0.356116 0.418738 2.14039 134.09 83.9344 18.7217 60.873 0.00402474 0 -40 10
1.093 3.16528e-08 2.53913e-06 0.118362 0.118361 0.0120355 1.43876e-05 0.00115415 0.147953 0.000658241 0.148606 0.895912 101.758 0.241669 0.77163 4.24171 0.0583314 0.0400161 0.959984 0.01974 0.00435092 0.0190027 0.00417464 0.00526004 0.00599732 0.210402 0.239893 58.0075 -87.8967 126.261 15.9599 145.022 0.000141163 0.267189 192.836 0.310475 0.0673598 0.00409648 0.000561936 0.00138366 0.986978 0.991727 -2.98022e-06 -85.6632 0.0930276 31183.9 303.474 0.983511 0.319146 0.732283 0.732279 9.99958 2.98319e-06 1.19326e-05 0.131745 0.982751 0.931743 -0.0132926 4.91096e-06 0.505388 -1.92553e-20 7.1139e-24 -1.92482e-20 0.0013957 0.997817 8.59696e-05 0.15263 2.85218 0.0013957 0.997819 0.735514 0.00105602 0.00188041 0.000859696 0.455536 0.00188041 0.440398 0.00012947 1.02 0.888037 0.53458 0.286548 1.71767e-07 3.06903e-09 2381.81 3114.44 -0.0554749 0.482158 0.277462 0.253192 -0.593388 -0.169531 0.496428 -0.267191 -0.229246 1.995 1 0 297.76 0 2.14034 1.993 0.00029973 0.853249 0.670704 0.356021 0.418762 2.14054 134.098 83.9343 18.7217 60.8729 0.00402474 0 -40 10
1.094 3.16817e-08 2.53913e-06 0.118418 0.118417 0.0120354 1.44008e-05 0.00115415 0.148023 0.000658243 0.148676 0.895988 101.758 0.241659 0.771743 4.24204 0.0583405 0.0400192 0.959981 0.0197396 0.0043512 0.0190023 0.00417488 0.00526039 0.00599767 0.210416 0.239907 58.0076 -87.8967 126.261 15.9599 145.022 0.000141163 0.267189 192.835 0.310474 0.0673597 0.00409648 0.000561937 0.00138366 0.986978 0.991727 -2.98023e-06 -85.6632 0.0930277 31183.8 303.481 0.983511 0.319146 0.732285 0.732281 9.99958 2.98319e-06 1.19327e-05 0.131748 0.982753 0.931743 -0.0132926 4.91099e-06 0.5054 -1.92563e-20 7.11433e-24 -1.92492e-20 0.0013957 0.997817 8.59696e-05 0.152631 2.85218 0.0013957 0.997819 0.735606 0.00105603 0.00188041 0.000859696 0.455536 0.00188041 0.440406 0.000129473 1.02 0.888038 0.53458 0.286549 1.71767e-07 3.06905e-09 2381.8 3114.44 -0.0554767 0.482158 0.277462 0.253193 -0.593388 -0.169532 0.496421 -0.267189 -0.229241 1.996 1 0 297.758 0 2.14049 1.994 0.000299729 0.853256 0.67075 0.355925 0.418787 2.14069 134.106 83.9342 18.7217 60.8729 0.00402474 0 -40 10
1.095 3.17106e-08 2.53914e-06 0.118474 0.118473 0.0120354 1.44139e-05 0.00115415 0.148093 0.000658244 0.148747 0.896063 101.758 0.24165 0.771857 4.24236 0.0583496 0.0400223 0.959978 0.0197393 0.00435148 0.019002 0.00417512 0.00526074 0.00599802 0.210429 0.239921 58.0077 -87.8967 126.261 15.9598 145.022 0.000141164 0.267189 192.835 0.310474 0.0673597 0.00409648 0.000561938 0.00138367 0.986978 0.991727 -2.98025e-06 -85.6632 0.0930278 31183.8 303.489 0.983511 0.319146 0.732287 0.732283 9.99958 2.9832e-06 1.19327e-05 0.131751 0.982755 0.931744 -0.0132926 4.91102e-06 0.505412 -1.92574e-20 7.11477e-24 -1.92503e-20 0.0013957 0.997817 8.59697e-05 0.152631 2.85218 0.0013957 0.997819 0.735698 0.00105605 0.00188041 0.000859697 0.455536 0.00188041 0.440413 0.000129476 1.02 0.88804 0.53458 0.286551 1.71767e-07 3.06908e-09 2381.78 3114.45 -0.0554786 0.482158 0.277462 0.253193 -0.593388 -0.169532 0.496415 -0.267187 -0.229237 1.997 1 0 297.757 0 2.14064 1.995 0.000299729 0.853263 0.670797 0.35583 0.418812 2.14084 134.114 83.9342 18.7217 60.8729 0.00402475 0 -40 10
1.096 3.17395e-08 2.53914e-06 0.118531 0.118529 0.0120354 1.4427e-05 0.00115415 0.148163 0.000658245 0.148817 0.896138 101.757 0.241641 0.77197 4.24269 0.0583587 0.0400254 0.959975 0.0197389 0.00435176 0.0190016 0.00417536 0.00526108 0.00599837 0.210443 0.239935 58.0077 -87.8967 126.261 15.9598 145.022 0.000141164 0.26719 192.835 0.310474 0.0673596 0.00409649 0.000561938 0.00138367 0.986978 0.991727 -2.98026e-06 -85.6632 0.0930279 31183.8 303.496 0.983511 0.319146 0.732289 0.732285 9.99958 2.9832e-06 1.19327e-05 0.131753 0.982758 0.931744 -0.0132925 4.91105e-06 0.505423 -1.92584e-20 7.1152e-24 -1.92513e-20 0.0013957 0.997817 8.59698e-05 0.152631 2.85218 0.0013957 0.997819 0.73579 0.00105607 0.00188041 0.000859698 0.455535 0.00188041 0.44042 0.000129479 1.02 0.888041 0.53458 0.286552 1.71767e-07 3.0691e-09 2381.76 3114.46 -0.0554804 0.482158 0.277461 0.253194 -0.593387 -0.169532 0.496408 -0.267185 -0.229233 1.998 1 0 297.755 0 2.14079 1.996 0.000299728 0.853269 0.670844 0.355735 0.418836 2.14099 134.122 83.9341 18.7217 60.8728 0.00402475 0 -40 10
1.097 3.17684e-08 2.53914e-06 0.118587 0.118585 0.0120354 1.44402e-05 0.00115415 0.148233 0.000658247 0.148887 0.896214 101.757 0.241632 0.772083 4.24301 0.0583677 0.0400284 0.959972 0.0197386 0.00435204 0.0190013 0.00417559 0.00526143 0.00599872 0.210457 0.239949 58.0078 -87.8967 126.261 15.9597 145.022 0.000141165 0.26719 192.835 0.310473 0.0673596 0.00409649 0.000561939 0.00138367 0.986978 0.991727 -2.98028e-06 -85.6632 0.093028 31183.8 303.504 0.983511 0.319146 0.732291 0.732287 9.99958 2.98321e-06 1.19327e-05 0.131756 0.98276 0.931744 -0.0132925 4.91108e-06 0.505435 -1.92595e-20 7.11563e-24 -1.92524e-20 0.0013957 0.997817 8.59699e-05 0.152631 2.85218 0.0013957 0.997819 0.735882 0.00105609 0.00188041 0.000859699 0.455535 0.00188041 0.440427 0.000129482 1.02 0.888042 0.534579 0.286554 1.71768e-07 3.06912e-09 2381.75 3114.47 -0.0554823 0.482158 0.277461 0.253194 -0.593387 -0.169532 0.496402 -0.267183 -0.229228 1.999 1 0 297.754 0 2.14094 1.997 0.000299727 0.853276 0.67089 0.35564 0.418861 2.14114 134.13 83.934 18.7217 60.8728 0.00402475 0 -40 10
1.098 3.17973e-08 2.53914e-06 0.118643 0.118641 0.0120354 1.44533e-05 0.00115415 0.148303 0.000658248 0.148957 0.896289 101.757 0.241623 0.772197 4.24334 0.0583768 0.0400315 0.959968 0.0197382 0.00435233 0.0190009 0.00417583 0.00526178 0.00599907 0.210471 0.239963 58.0078 -87.8967 126.261 15.9597 145.023 0.000141165 0.26719 192.835 0.310473 0.0673595 0.00409649 0.00056194 0.00138367 0.986978 0.991727 -2.98029e-06 -85.6632 0.0930281 31183.8 303.512 0.983511 0.319146 0.732293 0.732289 9.99958 2.98321e-06 1.19327e-05 0.131759 0.982762 0.931744 -0.0132925 4.91111e-06 0.505447 -1.92605e-20 7.11606e-24 -1.92534e-20 0.00139571 0.997817 8.597e-05 0.152631 2.85218 0.00139571 0.997819 0.735974 0.00105611 0.00188041 0.0008597 0.455535 0.00188041 0.440434 0.000129485 1.02 0.888043 0.534579 0.286555 1.71768e-07 3.06915e-09 2381.73 3114.47 -0.0554842 0.482158 0.277461 0.253195 -0.593387 -0.169532 0.496395 -0.267181 -0.229224 2 1 0 297.753 0 2.14109 1.998 0.000299727 0.853283 0.670937 0.355545 0.418886 2.14129 134.138 83.9339 18.7217 60.8727 0.00402476 0 -40 10
1.099 3.18262e-08 2.53914e-06 0.118699 0.118697 0.0120354 1.44665e-05 0.00115415 0.148373 0.00065825 0.149027 0.896365 101.756 0.241614 0.77231 4.24367 0.0583859 0.0400346 0.959965 0.0197379 0.00435261 0.0190006 0.00417607 0.00526213 0.00599942 0.210485 0.239977 58.0079 -87.8967 126.261 15.9597 145.023 0.000141165 0.26719 192.835 0.310472 0.0673595 0.0040965 0.00056194 0.00138367 0.986978 0.991727 -2.98031e-06 -85.6632 0.0930282 31183.7 303.519 0.983511 0.319146 0.732295 0.732291 9.99958 2.98322e-06 1.19328e-05 0.131762 0.982765 0.931745 -0.0132925 4.91114e-06 0.505459 -1.92616e-20 7.1165e-24 -1.92545e-20 0.00139571 0.997817 8.597e-05 0.152631 2.85219 0.00139571 0.997819 0.736066 0.00105613 0.00188042 0.0008597 0.455535 0.00188041 0.440442 0.000129488 1.02 0.888044 0.534579 0.286557 1.71768e-07 3.06917e-09 2381.71 3114.48 -0.0554861 0.482158 0.277461 0.253195 -0.593387 -0.169532 0.496389 -0.267179 -0.229219 2.001 1 0 297.751 0 2.14123 1.999 0.000299726 0.85329 0.670984 0.35545 0.41891 2.14144 134.146 83.9337 18.7217 60.8727 0.00402476 0 -40 10
1.1 3.18551e-08 2.53914e-06 0.118754 0.118753 0.0120354 1.44796e-05 0.00115415 0.148443 0.000658251 0.149097 0.89644 101.756 0.241605 0.772424 4.244 0.058395 0.0400377 0.959962 0.0197375 0.00435289 0.0190002 0.00417631 0.00526247 0.00599977 0.210499 0.239991 58.008 -87.8967 126.261 15.9596 145.023 0.000141166 0.26719 192.834 0.310472 0.0673594 0.0040965 0.000561941 0.00138368 0.986977 0.991727 -2.98032e-06 -85.6632 0.0930282 31183.7 303.527 0.983511 0.319146 0.732297 0.732293 9.99958 2.98322e-06 1.19328e-05 0.131765 0.982767 0.931745 -0.0132925 4.91117e-06 0.505471 -1.92627e-20 7.11693e-24 -1.92555e-20 0.00139571 0.997817 8.59701e-05 0.152631 2.85219 0.00139571 0.997819 0.736157 0.00105615 0.00188042 0.000859701 0.455534 0.00188042 0.440449 0.000129491 1.02 0.888045 0.534578 0.286558 1.71768e-07 3.06919e-09 2381.7 3114.49 -0.055488 0.482158 0.27746 0.253196 -0.593387 -0.169532 0.496382 -0.267177 -0.229215 2.002 1 0 297.75 0 2.14138 2 0.000299725 0.853297 0.67103 0.355356 0.418935 2.14159 134.154 83.9336 18.7217 60.8726 0.00402477 0 -40 10
1.101 3.1884e-08 2.53914e-06 0.11881 0.118809 0.0120354 1.44927e-05 0.00115415 0.148513 0.000658252 0.149167 0.896516 101.756 0.241596 0.772538 4.24432 0.0584041 0.0400408 0.959959 0.0197372 0.00435318 0.0189999 0.00417655 0.00526282 0.00600012 0.210513 0.240005 58.008 -87.8967 126.261 15.9596 145.023 0.000141166 0.26719 192.834 0.310472 0.0673593 0.0040965 0.000561942 0.00138368 0.986977 0.991727 -2.98034e-06 -85.6632 0.0930283 31183.7 303.535 0.983511 0.319146 0.732299 0.732295 9.99958 2.98323e-06 1.19328e-05 0.131768 0.982769 0.931745 -0.0132925 4.9112e-06 0.505483 -1.92637e-20 7.11737e-24 -1.92566e-20 0.00139571 0.997817 8.59702e-05 0.152632 2.85219 0.00139571 0.997819 0.736249 0.00105616 0.00188042 0.000859702 0.455534 0.00188042 0.440456 0.000129493 1.02 0.888046 0.534578 0.28656 1.71769e-07 3.06921e-09 2381.68 3114.5 -0.0554899 0.482159 0.27746 0.253197 -0.593387 -0.169532 0.496376 -0.267174 -0.22921 2.003 1 0 297.748 0 2.14153 2.001 0.000299725 0.853304 0.671077 0.355261 0.41896 2.14174 134.162 83.9335 18.7216 60.8726 0.00402477 0 -40 10
1.102 3.19129e-08 2.53914e-06 0.118866 0.118865 0.0120353 1.45059e-05 0.00115415 0.148583 0.000658254 0.149236 0.896592 101.755 0.241587 0.772651 4.24465 0.0584132 0.0400439 0.959956 0.0197368 0.00435346 0.0189995 0.00417679 0.00526317 0.00600047 0.210527 0.240019 58.0081 -87.8967 126.261 15.9596 145.023 0.000141167 0.267191 192.834 0.310471 0.0673593 0.00409651 0.000561942 0.00138368 0.986977 0.991727 -2.98035e-06 -85.6631 0.0930284 31183.7 303.543 0.983511 0.319146 0.732302 0.732297 9.99958 2.98323e-06 1.19328e-05 0.131771 0.982772 0.931745 -0.0132925 4.91123e-06 0.505496 -1.92648e-20 7.1178e-24 -1.92577e-20 0.00139571 0.997817 8.59703e-05 0.152632 2.85219 0.00139571 0.997819 0.736341 0.00105618 0.00188042 0.000859703 0.455534 0.00188042 0.440463 0.000129496 1.02 0.888047 0.534578 0.286561 1.71769e-07 3.06924e-09 2381.66 3114.51 -0.0554918 0.482159 0.27746 0.253197 -0.593387 -0.169532 0.496369 -0.267172 -0.229206 2.004 1 0 297.747 0 2.14168 2.002 0.000299724 0.853311 0.671124 0.355167 0.418984 2.14188 134.17 83.9334 18.7216 60.8725 0.00402478 0 -40 10
1.103 3.19418e-08 2.53914e-06 0.118922 0.118921 0.0120353 1.4519e-05 0.00115416 0.148652 0.000658255 0.149306 0.896667 101.755 0.241578 0.772765 4.24498 0.0584223 0.040047 0.959953 0.0197365 0.00435374 0.0189992 0.00417703 0.00526352 0.00600082 0.210541 0.240033 58.0082 -87.8967 126.261 15.9595 145.023 0.000141167 0.267191 192.834 0.310471 0.0673592 0.00409651 0.000561943 0.00138368 0.986977 0.991727 -2.98037e-06 -85.6631 0.0930285 31183.6 303.55 0.983511 0.319146 0.732304 0.732299 9.99958 2.98324e-06 1.19328e-05 0.131774 0.982774 0.931745 -0.0132925 4.91126e-06 0.505508 -1.92658e-20 7.11824e-24 -1.92587e-20 0.00139571 0.997817 8.59704e-05 0.152632 2.85219 0.00139571 0.997819 0.736433 0.0010562 0.00188042 0.000859704 0.455534 0.00188042 0.44047 0.000129499 1.02 0.888048 0.534577 0.286563 1.71769e-07 3.06926e-09 2381.65 3114.52 -0.0554937 0.482159 0.277459 0.253198 -0.593386 -0.169532 0.496362 -0.26717 -0.229201 2.005 1 0 297.745 0 2.14183 2.003 0.000299723 0.853318 0.67117 0.355073 0.419009 2.14203 134.178 83.9333 18.7216 60.8724 0.00402478 0 -40 10
1.104 3.19707e-08 2.53914e-06 0.118978 0.118976 0.0120353 1.45322e-05 0.00115416 0.148722 0.000658256 0.149376 0.896743 101.755 0.241569 0.772879 4.24531 0.0584314 0.0400501 0.95995 0.0197361 0.00435403 0.0189988 0.00417727 0.00526387 0.00600117 0.210555 0.240047 58.0082 -87.8967 126.261 15.9595 145.023 0.000141167 0.267191 192.834 0.31047 0.0673592 0.00409651 0.000561944 0.00138369 0.986977 0.991727 -2.98038e-06 -85.6631 0.0930286 31183.6 303.558 0.983511 0.319146 0.732306 0.732302 9.99958 2.98324e-06 1.19329e-05 0.131777 0.982776 0.931746 -0.0132925 4.91129e-06 0.50552 -1.92669e-20 7.11867e-24 -1.92598e-20 0.00139571 0.997817 8.59704e-05 0.152632 2.85219 0.00139571 0.997819 0.736524 0.00105622 0.00188042 0.000859704 0.455534 0.00188042 0.440477 0.000129502 1.02 0.888049 0.534577 0.286565 1.7177e-07 3.06928e-09 2381.63 3114.53 -0.0554957 0.482159 0.277459 0.253198 -0.593386 -0.169532 0.496355 -0.267168 -0.229197 2.006 1 0 297.744 0 2.14198 2.004 0.000299723 0.853326 0.671217 0.354979 0.419034 2.14218 134.186 83.9332 18.7216 60.8724 0.00402479 0 -40 10
1.105 3.19997e-08 2.53914e-06 0.119033 0.119032 0.0120353 1.45453e-05 0.00115416 0.148792 0.000658258 0.149445 0.896819 101.754 0.24156 0.772993 4.24564 0.0584405 0.0400532 0.959947 0.0197358 0.00435431 0.0189985 0.00417751 0.00526422 0.00600153 0.210569 0.240061 58.0083 -87.8967 126.261 15.9594 145.023 0.000141168 0.267191 192.834 0.31047 0.0673591 0.00409651 0.000561944 0.00138369 0.986977 0.991727 -2.9804e-06 -85.6631 0.0930287 31183.6 303.566 0.983511 0.319146 0.732308 0.732304 9.99958 2.98325e-06 1.19329e-05 0.13178 0.982779 0.931746 -0.0132925 4.91132e-06 0.505532 -1.92679e-20 7.11911e-24 -1.92608e-20 0.00139571 0.997817 8.59705e-05 0.152632 2.85219 0.00139571 0.997819 0.736616 0.00105624 0.00188042 0.000859705 0.455533 0.00188042 0.440485 0.000129505 1.02 0.88805 0.534577 0.286566 1.7177e-07 3.06931e-09 2381.61 3114.53 -0.0554976 0.482159 0.277459 0.253199 -0.593386 -0.169532 0.496349 -0.267166 -0.229192 2.007 1 0 297.742 0 2.14213 2.005 0.000299722 0.853333 0.671263 0.354886 0.419058 2.14233 134.194 83.9331 18.7216 60.8723 0.00402479 0 -40 10
1.106 3.20286e-08 2.53914e-06 0.119089 0.119088 0.0120353 1.45584e-05 0.00115416 0.148861 0.000658259 0.149515 0.896894 101.754 0.24155 0.773107 4.24597 0.0584496 0.0400563 0.959944 0.0197354 0.0043546 0.0189981 0.00417775 0.00526457 0.00600188 0.210583 0.240075 58.0084 -87.8967 126.26 15.9594 145.023 0.000141168 0.267191 192.833 0.310469 0.0673591 0.00409652 0.000561945 0.00138369 0.986977 0.991727 -2.98041e-06 -85.6631 0.0930288 31183.6 303.573 0.983511 0.319146 0.732311 0.732306 9.99958 2.98325e-06 1.19329e-05 0.131782 0.982781 0.931746 -0.0132925 4.91135e-06 0.505544 -1.9269e-20 7.11954e-24 -1.92619e-20 0.00139571 0.997817 8.59706e-05 0.152632 2.85219 0.00139571 0.997819 0.736707 0.00105626 0.00188043 0.000859706 0.455533 0.00188042 0.440492 0.000129508 1.02 0.888052 0.534576 0.286568 1.7177e-07 3.06933e-09 2381.6 3114.54 -0.0554996 0.482159 0.277459 0.2532 -0.593386 -0.169532 0.496342 -0.267164 -0.229187 2.008 1 0 297.74 0 2.14228 2.006 0.000299722 0.853341 0.67131 0.354792 0.419083 2.14248 134.202 83.933 18.7216 60.8723 0.0040248 0 -40 10
1.107 3.20575e-08 2.53914e-06 0.119145 0.119143 0.0120353 1.45716e-05 0.00115416 0.148931 0.00065826 0.149584 0.89697 101.754 0.241541 0.773221 4.2463 0.0584587 0.0400595 0.959941 0.0197351 0.00435488 0.0189978 0.00417799 0.00526492 0.00600223 0.210597 0.240089 58.0084 -87.8967 126.26 15.9594 145.023 0.000141169 0.267192 192.833 0.310469 0.067359 0.00409652 0.000561946 0.00138369 0.986977 0.991727 -2.98042e-06 -85.6631 0.0930288 31183.6 303.581 0.983511 0.319146 0.732313 0.732309 9.99958 2.98326e-06 1.19329e-05 0.131785 0.982783 0.931746 -0.0132925 4.91138e-06 0.505556 -1.92701e-20 7.11998e-24 -1.9263e-20 0.00139572 0.997817 8.59707e-05 0.152632 2.85219 0.00139572 0.997819 0.736799 0.00105627 0.00188043 0.000859707 0.455533 0.00188043 0.440499 0.000129511 1.02 0.888053 0.534576 0.286569 1.7177e-07 3.06935e-09 2381.58 3114.55 -0.0555016 0.482159 0.277458 0.2532 -0.593386 -0.169532 0.496335 -0.267162 -0.229182 2.009 1 0 297.739 0 2.14243 2.007 0.000299721 0.853348 0.671357 0.354699 0.419107 2.14263 134.21 83.9329 18.7216 60.8722 0.0040248 0 -40 10
1.108 3.20864e-08 2.53915e-06 0.1192 0.119199 0.0120353 1.45847e-05 0.00115416 0.149 0.000658262 0.149654 0.897046 101.753 0.241532 0.773335 4.24663 0.0584678 0.0400626 0.959937 0.0197347 0.00435517 0.0189974 0.00417824 0.00526528 0.00600259 0.210611 0.240104 58.0085 -87.8967 126.26 15.9593 145.023 0.000141169 0.267192 192.833 0.310469 0.067359 0.00409652 0.000561946 0.00138369 0.986977 0.991727 -2.98044e-06 -85.6631 0.0930289 31183.5 303.589 0.983511 0.319146 0.732315 0.732311 9.99958 2.98326e-06 1.19329e-05 0.131788 0.982785 0.931746 -0.0132925 4.91141e-06 0.505568 -1.92711e-20 7.12042e-24 -1.9264e-20 0.00139572 0.997817 8.59708e-05 0.152633 2.85219 0.00139572 0.997819 0.73689 0.00105629 0.00188043 0.000859708 0.455533 0.00188043 0.440506 0.000129514 1.02 0.888054 0.534576 0.286571 1.71771e-07 3.06937e-09 2381.56 3114.56 -0.0555036 0.482159 0.277458 0.253201 -0.593386 -0.169532 0.496328 -0.26716 -0.229178 2.01 1 0 297.737 0 2.14257 2.008 0.00029972 0.853356 0.671403 0.354606 0.419132 2.14278 134.218 83.9327 18.7216 60.8722 0.0040248 0 -40 10
1.109 3.21153e-08 2.53915e-06 0.119256 0.119254 0.0120352 1.45979e-05 0.00115416 0.14907 0.000658263 0.149723 0.897122 101.753 0.241523 0.773449 4.24697 0.058477 0.0400657 0.959934 0.0197344 0.00435546 0.0189971 0.00417848 0.00526563 0.00600294 0.210625 0.240118 58.0085 -87.8967 126.26 15.9593 145.023 0.00014117 0.267192 192.833 0.310468 0.0673589 0.00409653 0.000561947 0.0013837 0.986977 0.991727 -2.98045e-06 -85.6631 0.093029 31183.5 303.597 0.983511 0.319146 0.732318 0.732314 9.99958 2.98327e-06 1.1933e-05 0.131791 0.982788 0.931747 -0.0132925 4.91144e-06 0.50558 -1.92722e-20 7.12085e-24 -1.92651e-20 0.00139572 0.997817 8.59709e-05 0.152633 2.85219 0.00139572 0.997819 0.736982 0.00105631 0.00188043 0.000859709 0.455532 0.00188043 0.440513 0.000129517 1.02 0.888055 0.534576 0.286572 1.71771e-07 3.0694e-09 2381.55 3114.57 -0.0555056 0.482159 0.277458 0.253202 -0.593386 -0.169533 0.496321 -0.267158 -0.229173 2.011 1 0 297.736 0 2.14272 2.009 0.00029972 0.853363 0.67145 0.354513 0.419157 2.14292 134.226 83.9326 18.7216 60.8721 0.00402481 0 -40 10
1.11 3.21442e-08 2.53915e-06 0.119311 0.11931 0.0120352 1.4611e-05 0.00115416 0.149139 0.000658264 0.149793 0.897198 101.753 0.241514 0.773563 4.2473 0.0584861 0.0400689 0.959931 0.019734 0.00435574 0.0189967 0.00417872 0.00526598 0.0060033 0.210639 0.240132 58.0086 -87.8967 126.26 15.9593 145.023 0.00014117 0.267192 192.833 0.310468 0.0673589 0.00409653 0.000561948 0.0013837 0.986977 0.991727 -2.98047e-06 -85.6631 0.0930291 31183.5 303.604 0.983511 0.319146 0.73232 0.732316 9.99958 2.98327e-06 1.1933e-05 0.131794 0.98279 0.931747 -0.0132925 4.91146e-06 0.505592 -1.92733e-20 7.12129e-24 -1.92661e-20 0.00139572 0.997817 8.59709e-05 0.152633 2.8522 0.00139572 0.997819 0.737073 0.00105633 0.00188043 0.000859709 0.455532 0.00188043 0.44052 0.00012952 1.02 0.888056 0.534575 0.286574 1.71771e-07 3.06942e-09 2381.53 3114.58 -0.0555076 0.482159 0.277457 0.253202 -0.593385 -0.169533 0.496314 -0.267155 -0.229168 2.012 1 0 297.734 0 2.14287 2.01 0.000299719 0.853371 0.671496 0.35442 0.419181 2.14307 134.234 83.9325 18.7216 60.8721 0.00402481 0 -40 10
1.111 3.21731e-08 2.53915e-06 0.119367 0.119365 0.0120352 1.46241e-05 0.00115416 0.149208 0.000658266 0.149862 0.897274 101.752 0.241505 0.773677 4.24763 0.0584952 0.040072 0.959928 0.0197337 0.00435603 0.0189963 0.00417896 0.00526633 0.00600365 0.210653 0.240146 58.0087 -87.8967 126.26 15.9592 145.023 0.000141171 0.267192 192.833 0.310467 0.0673588 0.00409653 0.000561948 0.0013837 0.986977 0.991727 -2.98048e-06 -85.6631 0.0930292 31183.5 303.612 0.983511 0.319146 0.732323 0.732319 9.99958 2.98328e-06 1.1933e-05 0.131797 0.982792 0.931747 -0.0132925 4.91149e-06 0.505605 -1.92743e-20 7.12173e-24 -1.92672e-20 0.00139572 0.997817 8.5971e-05 0.152633 2.8522 0.00139572 0.997819 0.737165 0.00105635 0.00188043 0.00085971 0.455532 0.00188043 0.440528 0.000129523 1.02 0.888057 0.534575 0.286575 1.71771e-07 3.06944e-09 2381.51 3114.59 -0.0555096 0.482159 0.277457 0.253203 -0.593385 -0.169533 0.496307 -0.267153 -0.229163 2.013 1 0 297.733 0 2.14302 2.011 0.000299718 0.853379 0.671543 0.354327 0.419206 2.14322 134.242 83.9324 18.7216 60.872 0.00402482 0 -40 10
1.112 3.2202e-08 2.53915e-06 0.119422 0.119421 0.0120352 1.46373e-05 0.00115416 0.149277 0.000658267 0.149931 0.89735 101.752 0.241496 0.773791 4.24796 0.0585044 0.0400751 0.959925 0.0197333 0.00435632 0.018996 0.00417921 0.00526668 0.00600401 0.210667 0.24016 58.0087 -87.8967 126.26 15.9592 145.023 0.000141171 0.267193 192.832 0.310467 0.0673588 0.00409654 0.000561949 0.0013837 0.986977 0.991727 -2.9805e-06 -85.6631 0.0930293 31183.4 303.62 0.983511 0.319146 0.732325 0.732321 9.99958 2.98328e-06 1.1933e-05 0.1318 0.982794 0.931747 -0.0132925 4.91152e-06 0.505617 -1.92754e-20 7.12217e-24 -1.92683e-20 0.00139572 0.997817 8.59711e-05 0.152633 2.8522 0.00139572 0.997819 0.737256 0.00105637 0.00188043 0.000859711 0.455532 0.00188043 0.440535 0.000129526 1.02 0.888058 0.534575 0.286577 1.71772e-07 3.06947e-09 2381.5 3114.6 -0.0555116 0.482159 0.277457 0.253204 -0.593385 -0.169533 0.4963 -0.267151 -0.229158 2.014 1 0 297.731 0 2.14317 2.012 0.000299718 0.853387 0.671589 0.354235 0.41923 2.14337 134.25 83.9322 18.7216 60.8719 0.00402483 0 -40 10
1.113 3.22309e-08 2.53915e-06 0.119477 0.119476 0.0120352 1.46504e-05 0.00115416 0.149347 0.000658268 0.15 0.897426 101.752 0.241486 0.773905 4.2483 0.0585135 0.0400783 0.959922 0.019733 0.0043566 0.0189956 0.00417945 0.00526704 0.00600436 0.210682 0.240175 58.0088 -87.8967 126.26 15.9591 145.023 0.000141172 0.267193 192.832 0.310466 0.0673587 0.00409654 0.00056195 0.00138371 0.986977 0.991727 -2.98051e-06 -85.663 0.0930294 31183.4 303.628 0.983511 0.319146 0.732328 0.732324 9.99958 2.98329e-06 1.1933e-05 0.131803 0.982797 0.931747 -0.0132925 4.91155e-06 0.505629 -1.92765e-20 7.1226e-24 -1.92693e-20 0.00139572 0.997817 8.59712e-05 0.152633 2.8522 0.00139572 0.997819 0.737347 0.00105639 0.00188044 0.000859712 0.455532 0.00188043 0.440542 0.000129529 1.02 0.888059 0.534574 0.286578 1.71772e-07 3.06949e-09 2381.48 3114.61 -0.0555137 0.482159 0.277457 0.253204 -0.593385 -0.169533 0.496293 -0.267149 -0.229153 2.015 1 0 297.729 0 2.14332 2.013 0.000299717 0.853395 0.671636 0.354143 0.419255 2.14352 134.258 83.9321 18.7216 60.8719 0.00402483 0 -40 10
1.114 3.22598e-08 2.53915e-06 0.119533 0.119531 0.0120352 1.46635e-05 0.00115416 0.149416 0.00065827 0.150069 0.897502 101.751 0.241477 0.774019 4.24863 0.0585226 0.0400814 0.959919 0.0197326 0.00435689 0.0189953 0.00417969 0.00526739 0.00600472 0.210696 0.240189 58.0089 -87.8967 126.26 15.9591 145.023 0.000141172 0.267193 192.832 0.310466 0.0673587 0.00409654 0.00056195 0.00138371 0.986977 0.991727 -2.98053e-06 -85.663 0.0930295 31183.4 303.636 0.983511 0.319146 0.732331 0.732326 9.99958 2.98329e-06 1.19331e-05 0.131806 0.982799 0.931747 -0.0132925 4.91158e-06 0.505641 -1.92775e-20 7.12304e-24 -1.92704e-20 0.00139572 0.997817 8.59713e-05 0.152634 2.8522 0.00139572 0.997819 0.737439 0.0010564 0.00188044 0.000859713 0.455531 0.00188044 0.440549 0.000129532 1.02 0.88806 0.534574 0.28658 1.71772e-07 3.06951e-09 2381.46 3114.62 -0.0555157 0.482159 0.277456 0.253205 -0.593385 -0.169533 0.496286 -0.267147 -0.229148 2.016 1 0 297.728 0 2.14346 2.014 0.000299716 0.853403 0.671682 0.354051 0.41928 2.14367 134.266 83.932 18.7216 60.8718 0.00402484 0 -40 10
1.115 3.22887e-08 2.53915e-06 0.119588 0.119586 0.0120352 1.46767e-05 0.00115416 0.149485 0.000658271 0.150138 0.897578 101.751 0.241468 0.774134 4.24897 0.0585318 0.0400846 0.959915 0.0197323 0.00435718 0.0189949 0.00417994 0.00526775 0.00600508 0.21071 0.240203 58.0089 -87.8967 126.26 15.9591 145.023 0.000141173 0.267193 192.832 0.310466 0.0673586 0.00409654 0.000561951 0.00138371 0.986977 0.991727 -2.98054e-06 -85.663 0.0930295 31183.4 303.643 0.98351 0.319146 0.732333 0.732329 9.99958 2.9833e-06 1.19331e-05 0.131809 0.982801 0.931747 -0.0132925 4.91161e-06 0.505653 -1.92786e-20 7.12348e-24 -1.92715e-20 0.00139573 0.997817 8.59713e-05 0.152634 2.8522 0.00139572 0.997819 0.73753 0.00105642 0.00188044 0.000859713 0.455531 0.00188044 0.440556 0.000129535 1.02 0.888061 0.534574 0.286581 1.71772e-07 3.06953e-09 2381.45 3114.63 -0.0555178 0.48216 0.277456 0.253206 -0.593385 -0.169533 0.496279 -0.267145 -0.229143 2.017 1 0 297.726 0 2.14361 2.015 0.000299716 0.853411 0.671729 0.353959 0.419304 2.14382 134.274 83.9319 18.7215 60.8717 0.00402484 0 -40 10
1.116 3.23176e-08 2.53915e-06 0.119643 0.119642 0.0120352 1.46898e-05 0.00115416 0.149554 0.000658272 0.150207 0.897654 101.751 0.241459 0.774248 4.2493 0.0585409 0.0400877 0.959912 0.0197319 0.00435747 0.0189946 0.00418018 0.0052681 0.00600543 0.210724 0.240217 58.009 -87.8968 126.26 15.959 145.023 0.000141173 0.267193 192.832 0.310465 0.0673586 0.00409655 0.000561952 0.00138371 0.986977 0.991727 -2.98056e-06 -85.663 0.0930296 31183.4 303.651 0.98351 0.319146 0.732336 0.732332 9.99958 2.9833e-06 1.19331e-05 0.131812 0.982803 0.931748 -0.0132925 4.91164e-06 0.505666 -1.92797e-20 7.12392e-24 -1.92725e-20 0.00139573 0.997817 8.59714e-05 0.152634 2.8522 0.00139573 0.997819 0.737621 0.00105644 0.00188044 0.000859714 0.455531 0.00188044 0.440563 0.000129538 1.02 0.888063 0.534573 0.286583 1.71773e-07 3.06956e-09 2381.43 3114.64 -0.0555199 0.48216 0.277456 0.253206 -0.593384 -0.169533 0.496272 -0.267143 -0.229138 2.018 1 0 297.724 0 2.14376 2.016 0.000299715 0.853419 0.671775 0.353867 0.419329 2.14396 134.282 83.9317 18.7215 60.8717 0.00402485 0 -40 10
1.117 3.23465e-08 2.53915e-06 0.119698 0.119697 0.0120351 1.4703e-05 0.00115416 0.149623 0.000658274 0.150276 0.89773 101.75 0.24145 0.774362 4.24964 0.0585501 0.0400909 0.959909 0.0197315 0.00435775 0.0189942 0.00418042 0.00526845 0.00600579 0.210738 0.240232 58.0091 -87.8968 126.26 15.959 145.023 0.000141174 0.267194 192.832 0.310465 0.0673585 0.00409655 0.000561952 0.00138371 0.986977 0.991727 -2.98057e-06 -85.663 0.0930297 31183.3 303.659 0.98351 0.319146 0.732339 0.732334 9.99958 2.98331e-06 1.19331e-05 0.131815 0.982806 0.931748 -0.0132925 4.91167e-06 0.505678 -1.92807e-20 7.12436e-24 -1.92736e-20 0.00139573 0.997817 8.59715e-05 0.152634 2.8522 0.00139573 0.997819 0.737712 0.00105646 0.00188044 0.000859715 0.455531 0.00188044 0.44057 0.000129541 1.02 0.888064 0.534573 0.286584 1.71773e-07 3.06958e-09 2381.41 3114.66 -0.055522 0.48216 0.277455 0.253207 -0.593384 -0.169533 0.496264 -0.267141 -0.229133 2.019 1 0 297.723 0 2.14391 2.017 0.000299714 0.853427 0.671822 0.353775 0.419353 2.14411 134.289 83.9316 18.7215 60.8716 0.00402485 0 -40 10
1.118 3.23754e-08 2.53915e-06 0.119753 0.119752 0.0120351 1.47161e-05 0.00115416 0.149692 0.000658275 0.150345 0.897806 101.75 0.241441 0.774477 4.24997 0.0585593 0.0400941 0.959906 0.0197312 0.00435804 0.0189939 0.00418067 0.00526881 0.00600615 0.210752 0.240246 58.0091 -87.8968 126.26 15.959 145.023 0.000141174 0.267194 192.831 0.310464 0.0673585 0.00409655 0.000561953 0.00138372 0.986977 0.991727 -2.98059e-06 -85.663 0.0930298 31183.3 303.667 0.98351 0.319146 0.732341 0.732337 9.99958 2.98331e-06 1.19331e-05 0.131818 0.982808 0.931748 -0.0132925 4.9117e-06 0.50569 -1.92818e-20 7.1248e-24 -1.92747e-20 0.00139573 0.997817 8.59716e-05 0.152634 2.8522 0.00139573 0.997818 0.737804 0.00105648 0.00188044 0.000859716 0.45553 0.00188044 0.440578 0.000129544 1.02 0.888065 0.534573 0.286586 1.71773e-07 3.0696e-09 2381.4 3114.67 -0.0555241 0.48216 0.277455 0.253208 -0.593384 -0.169533 0.496257 -0.267139 -0.229128 2.02 1 0 297.721 0 2.14406 2.018 0.000299714 0.853435 0.671868 0.353684 0.419378 2.14426 134.297 83.9315 18.7215 60.8716 0.00402486 0 -40 10
1.119 3.24043e-08 2.53915e-06 0.119808 0.119807 0.0120351 1.47292e-05 0.00115416 0.14976 0.000658276 0.150414 0.897882 101.75 0.241432 0.774591 4.25031 0.0585684 0.0400972 0.959903 0.0197308 0.00435833 0.0189935 0.00418091 0.00526917 0.00600651 0.210767 0.24026 58.0092 -87.8968 126.26 15.9589 145.023 0.000141175 0.267194 192.831 0.310464 0.0673584 0.00409656 0.000561954 0.00138372 0.986977 0.991727 -2.9806e-06 -85.663 0.0930299 31183.3 303.675 0.98351 0.319146 0.732344 0.73234 9.99958 2.98332e-06 1.19332e-05 0.131821 0.98281 0.931748 -0.0132925 4.91173e-06 0.505702 -1.92829e-20 7.12524e-24 -1.92758e-20 0.00139573 0.997817 8.59717e-05 0.152634 2.8522 0.00139573 0.997818 0.737895 0.0010565 0.00188045 0.000859717 0.45553 0.00188044 0.440585 0.000129547 1.02 0.888066 0.534572 0.286587 1.71774e-07 3.06963e-09 2381.38 3114.68 -0.0555262 0.48216 0.277455 0.253209 -0.593384 -0.169533 0.49625 -0.267136 -0.229123 2.021 1 0 297.719 0 2.14421 2.019 0.000299713 0.853444 0.671915 0.353592 0.419402 2.14441 134.305 83.9313 18.7215 60.8715 0.00402486 0 -40 10
1.12 3.24332e-08 2.53916e-06 0.119863 0.119862 0.0120351 1.47424e-05 0.00115416 0.149829 0.000658278 0.150483 0.897958 101.749 0.241422 0.774706 4.25064 0.0585776 0.0401004 0.9599 0.0197305 0.00435862 0.0189931 0.00418116 0.00526952 0.00600687 0.210781 0.240275 58.0092 -87.8968 126.26 15.9589 145.023 0.000141175 0.267194 192.831 0.310463 0.0673583 0.00409656 0.000561954 0.00138372 0.986977 0.991727 -2.98062e-06 -85.663 0.09303 31183.3 303.682 0.98351 0.319146 0.732347 0.732343 9.99958 2.98332e-06 1.19332e-05 0.131824 0.982812 0.931748 -0.0132925 4.91176e-06 0.505715 -1.9284e-20 7.12568e-24 -1.92768e-20 0.00139573 0.997817 8.59717e-05 0.152634 2.8522 0.00139573 0.997818 0.737986 0.00105651 0.00188045 0.000859717 0.45553 0.00188045 0.440592 0.00012955 1.02 0.888067 0.534572 0.286589 1.71774e-07 3.06965e-09 2381.36 3114.69 -0.0555283 0.48216 0.277455 0.253209 -0.593384 -0.169533 0.496243 -0.267134 -0.229118 2.022 1 0 297.718 0 2.14436 2.02 0.000299712 0.853452 0.671961 0.353501 0.419427 2.14456 134.313 83.9312 18.7215 60.8714 0.00402487 0 -40 10
1.121 3.24621e-08 2.53916e-06 0.119918 0.119917 0.0120351 1.47555e-05 0.00115416 0.149898 0.000658279 0.150552 0.898034 101.749 0.241413 0.774821 4.25098 0.0585868 0.0401036 0.959896 0.0197301 0.00435891 0.0189928 0.0041814 0.00526988 0.00600723 0.210795 0.240289 58.0093 -87.8968 126.26 15.9588 145.023 0.000141176 0.267194 192.831 0.310463 0.0673583 0.00409656 0.000561955 0.00138372 0.986977 0.991726 -2.98063e-06 -85.663 0.0930301 31183.2 303.69 0.98351 0.319146 0.73235 0.732346 9.99958 2.98333e-06 1.19332e-05 0.131826 0.982814 0.931748 -0.0132925 4.91179e-06 0.505727 -1.9285e-20 7.12612e-24 -1.92779e-20 0.00139573 0.997817 8.59718e-05 0.152635 2.85221 0.00139573 0.997818 0.738077 0.00105653 0.00188045 0.000859718 0.45553 0.00188045 0.440599 0.000129553 1.02 0.888068 0.534572 0.28659 1.71774e-07 3.06967e-09 2381.35 3114.7 -0.0555304 0.48216 0.277454 0.25321 -0.593384 -0.169533 0.496235 -0.267132 -0.229113 2.023 1 0 297.716 0 2.1445 2.021 0.000299712 0.85346 0.672007 0.35341 0.419451 2.1447 134.321 83.931 18.7215 60.8714 0.00402487 0 -40 10
1.122 3.2491e-08 2.53916e-06 0.119973 0.119972 0.0120351 1.47687e-05 0.00115416 0.149967 0.00065828 0.15062 0.898111 101.749 0.241404 0.774935 4.25132 0.0585959 0.0401068 0.959893 0.0197298 0.0043592 0.0189924 0.00418165 0.00527023 0.00600759 0.210809 0.240303 58.0094 -87.8968 126.26 15.9588 145.023 0.000141176 0.267194 192.831 0.310463 0.0673582 0.00409657 0.000561956 0.00138372 0.986977 0.991726 -2.98065e-06 -85.663 0.0930302 31183.2 303.698 0.98351 0.319146 0.732353 0.732348 9.99958 2.98333e-06 1.19332e-05 0.131829 0.982817 0.931748 -0.0132925 4.91182e-06 0.505739 -1.92861e-20 7.12656e-24 -1.9279e-20 0.00139573 0.997817 8.59719e-05 0.152635 2.85221 0.00139573 0.997818 0.738168 0.00105655 0.00188045 0.000859719 0.455529 0.00188045 0.440606 0.000129556 1.02 0.888069 0.534572 0.286592 1.71774e-07 3.06969e-09 2381.33 3114.71 -0.0555326 0.48216 0.277454 0.253211 -0.593383 -0.169533 0.496228 -0.26713 -0.229107 2.024 1 0 297.714 0 2.14465 2.022 0.000299711 0.853469 0.672054 0.35332 0.419476 2.14485 134.329 83.9309 18.7215 60.8713 0.00402488 0 -40 10
1.123 3.25199e-08 2.53916e-06 0.120028 0.120027 0.0120351 1.47818e-05 0.00115416 0.150035 0.000658282 0.150689 0.898187 101.748 0.241395 0.77505 4.25166 0.0586051 0.04011 0.95989 0.0197294 0.00435949 0.0189921 0.00418189 0.00527059 0.00600795 0.210824 0.240318 58.0094 -87.8968 126.26 15.9588 145.023 0.000141177 0.267195 192.831 0.310462 0.0673582 0.00409657 0.000561956 0.00138373 0.986977 0.991726 -2.98066e-06 -85.663 0.0930302 31183.2 303.706 0.98351 0.319146 0.732356 0.732351 9.99958 2.98334e-06 1.19332e-05 0.131832 0.982819 0.931749 -0.0132925 4.91185e-06 0.505752 -1.92872e-20 7.127e-24 -1.928e-20 0.00139573 0.997817 8.5972e-05 0.152635 2.85221 0.00139573 0.997818 0.738259 0.00105657 0.00188045 0.00085972 0.455529 0.00188045 0.440613 0.000129559 1.02 0.88807 0.534571 0.286593 1.71775e-07 3.06972e-09 2381.31 3114.72 -0.0555347 0.48216 0.277454 0.253212 -0.593383 -0.169533 0.496221 -0.267128 -0.229102 2.025 1 0 297.712 0 2.1448 2.023 0.000299711 0.853478 0.6721 0.353229 0.4195 2.145 134.337 83.9308 18.7215 60.8712 0.00402489 0 -40 10
1.124 3.25488e-08 2.53916e-06 0.120083 0.120082 0.012035 1.47949e-05 0.00115416 0.150104 0.000658283 0.150758 0.898263 101.748 0.241386 0.775165 4.252 0.0586143 0.0401132 0.959887 0.0197291 0.00435978 0.0189917 0.00418214 0.00527095 0.00600831 0.210838 0.240332 58.0095 -87.8968 126.26 15.9587 145.023 0.000141178 0.267195 192.831 0.310462 0.0673581 0.00409657 0.000561957 0.00138373 0.986977 0.991726 -2.98068e-06 -85.6629 0.0930303 31183.2 303.714 0.98351 0.319146 0.732359 0.732354 9.99958 2.98334e-06 1.19333e-05 0.131835 0.982821 0.931749 -0.0132925 4.91188e-06 0.505764 -1.92883e-20 7.12744e-24 -1.92811e-20 0.00139574 0.997817 8.59721e-05 0.152635 2.85221 0.00139574 0.997818 0.73835 0.00105659 0.00188045 0.000859721 0.455529 0.00188045 0.44062 0.000129562 1.02 0.888071 0.534571 0.286595 1.71775e-07 3.06974e-09 2381.29 3114.73 -0.0555369 0.48216 0.277453 0.253213 -0.593383 -0.169533 0.496213 -0.267126 -0.229097 2.026 1 0 297.711 0 2.14495 2.024 0.00029971 0.853486 0.672147 0.353138 0.419525 2.14515 134.345 83.9306 18.7215 60.8711 0.00402489 0 -40 10
1.125 3.25778e-08 2.53916e-06 0.120138 0.120137 0.012035 1.48081e-05 0.00115416 0.150172 0.000658284 0.150826 0.89834 101.748 0.241377 0.775279 4.25233 0.0586235 0.0401164 0.959884 0.0197287 0.00436007 0.0189913 0.00418238 0.00527131 0.00600867 0.210852 0.240347 58.0096 -87.8968 126.26 15.9587 145.023 0.000141178 0.267195 192.83 0.310461 0.0673581 0.00409658 0.000561958 0.00138373 0.986977 0.991726 -2.98069e-06 -85.6629 0.0930304 31183.2 303.722 0.98351 0.319146 0.732362 0.732357 9.99958 2.98335e-06 1.19333e-05 0.131838 0.982823 0.931749 -0.0132925 4.91191e-06 0.505776 -1.92893e-20 7.12788e-24 -1.92822e-20 0.00139574 0.997817 8.59721e-05 0.152635 2.85221 0.00139574 0.997818 0.738441 0.00105661 0.00188045 0.000859721 0.455529 0.00188045 0.440627 0.000129565 1.02 0.888072 0.534571 0.286596 1.71775e-07 3.06976e-09 2381.28 3114.75 -0.0555391 0.48216 0.277453 0.253213 -0.593383 -0.169534 0.496206 -0.267124 -0.229091 2.027 1 0 297.709 0 2.1451 2.025 0.000299709 0.853495 0.672193 0.353048 0.419549 2.1453 134.353 83.9305 18.7215 60.8711 0.0040249 0 -40 10
1.126 3.26067e-08 2.53916e-06 0.120193 0.120191 0.012035 1.48212e-05 0.00115416 0.150241 0.000658286 0.150894 0.898416 101.747 0.241367 0.775394 4.25267 0.0586327 0.0401196 0.95988 0.0197283 0.00436036 0.018991 0.00418263 0.00527166 0.00600903 0.210867 0.240361 58.0096 -87.8968 126.259 15.9586 145.023 0.000141179 0.267195 192.83 0.310461 0.067358 0.00409658 0.000561958 0.00138373 0.986977 0.991726 -2.98071e-06 -85.6629 0.0930305 31183.1 303.73 0.98351 0.319146 0.732365 0.73236 9.99958 2.98335e-06 1.19333e-05 0.131841 0.982825 0.931749 -0.0132925 4.91194e-06 0.505789 -1.92904e-20 7.12832e-24 -1.92833e-20 0.00139574 0.997817 8.59722e-05 0.152635 2.85221 0.00139574 0.997818 0.738532 0.00105662 0.00188046 0.000859722 0.455529 0.00188045 0.440634 0.000129568 1.02 0.888074 0.53457 0.286598 1.71775e-07 3.06979e-09 2381.26 3114.76 -0.0555413 0.48216 0.277453 0.253214 -0.593383 -0.169534 0.496198 -0.267122 -0.229086 2.028 1 0 297.707 0 2.14524 2.026 0.000299709 0.853504 0.67224 0.352958 0.419574 2.14545 134.361 83.9303 18.7215 60.871 0.0040249 0 -40 10
1.127 3.26356e-08 2.53916e-06 0.120247 0.120246 0.012035 1.48343e-05 0.00115416 0.150309 0.000658287 0.150963 0.898492 101.747 0.241358 0.775509 4.25301 0.0586419 0.0401228 0.959877 0.019728 0.00436065 0.0189906 0.00418288 0.00527202 0.00600939 0.210881 0.240376 58.0097 -87.8968 126.259 15.9586 145.023 0.000141179 0.267195 192.83 0.31046 0.067358 0.00409658 0.000561959 0.00138374 0.986977 0.991726 -2.98072e-06 -85.6629 0.0930306 31183.1 303.738 0.98351 0.319146 0.732368 0.732363 9.99958 2.98336e-06 1.19333e-05 0.131844 0.982827 0.931749 -0.0132925 4.91197e-06 0.505801 -1.92915e-20 7.12877e-24 -1.92844e-20 0.00139574 0.997817 8.59723e-05 0.152636 2.85221 0.00139574 0.997818 0.738623 0.00105664 0.00188046 0.000859723 0.455528 0.00188046 0.440641 0.00012957 1.02 0.888075 0.53457 0.286599 1.71776e-07 3.06981e-09 2381.24 3114.77 -0.0555435 0.48216 0.277453 0.253215 -0.593383 -0.169534 0.496191 -0.26712 -0.229081 2.029 1 0 297.705 0 2.14539 2.027 0.000299708 0.853513 0.672286 0.352868 0.419598 2.14559 134.369 83.9302 18.7215 60.8709 0.00402491 0 -40 10
1.128 3.26645e-08 2.53916e-06 0.120302 0.120301 0.012035 1.48475e-05 0.00115416 0.150378 0.000658288 0.151031 0.898569 101.747 0.241349 0.775624 4.25335 0.0586511 0.040126 0.959874 0.0197276 0.00436095 0.0189902 0.00418312 0.00527238 0.00600975 0.210895 0.24039 58.0098 -87.8968 126.259 15.9586 145.023 0.00014118 0.267196 192.83 0.31046 0.0673579 0.00409658 0.00056196 0.00138374 0.986977 0.991726 -2.98074e-06 -85.6629 0.0930307 31183.1 303.746 0.98351 0.319146 0.732371 0.732366 9.99958 2.98336e-06 1.19333e-05 0.131847 0.982829 0.931749 -0.0132925 4.912e-06 0.505813 -1.92926e-20 7.12921e-24 -1.92854e-20 0.00139574 0.997817 8.59724e-05 0.152636 2.85221 0.00139574 0.997818 0.738714 0.00105666 0.00188046 0.000859724 0.455528 0.00188046 0.440649 0.000129573 1.02 0.888076 0.53457 0.286601 1.71776e-07 3.06983e-09 2381.23 3114.78 -0.0555457 0.482161 0.277452 0.253216 -0.593382 -0.169534 0.496183 -0.267117 -0.229075 2.03 1 0 297.704 0 2.14554 2.028 0.000299707 0.853522 0.672332 0.352778 0.419623 2.14574 134.377 83.93 18.7214 60.8709 0.00402492 0 -40 10
1.129 3.26934e-08 2.53916e-06 0.120357 0.120355 0.012035 1.48606e-05 0.00115416 0.150446 0.00065829 0.151099 0.898645 101.746 0.24134 0.775739 4.25369 0.0586603 0.0401292 0.959871 0.0197273 0.00436124 0.0189899 0.00418337 0.00527274 0.00601011 0.21091 0.240405 58.0098 -87.8968 126.259 15.9585 145.023 0.000141181 0.267196 192.83 0.31046 0.0673579 0.00409659 0.00056196 0.00138374 0.986977 0.991726 -2.98075e-06 -85.6629 0.0930308 31183.1 303.753 0.98351 0.319146 0.732374 0.73237 9.99958 2.98337e-06 1.19334e-05 0.13185 0.982832 0.931749 -0.0132925 4.91203e-06 0.505826 -1.92936e-20 7.12965e-24 -1.92865e-20 0.00139574 0.997817 8.59725e-05 0.152636 2.85221 0.00139574 0.997818 0.738804 0.00105668 0.00188046 0.000859725 0.455528 0.00188046 0.440656 0.000129576 1.02 0.888077 0.534569 0.286603 1.71776e-07 3.06985e-09 2381.21 3114.8 -0.0555479 0.482161 0.277452 0.253217 -0.593382 -0.169534 0.496176 -0.267115 -0.22907 2.031 1 0 297.702 0 2.14569 2.029 0.000299707 0.853531 0.672379 0.352688 0.419647 2.14589 134.385 83.9299 18.7214 60.8708 0.00402492 0 -40 10
1.13 3.27223e-08 2.53916e-06 0.120411 0.12041 0.012035 1.48738e-05 0.00115417 0.150514 0.000658291 0.151168 0.898722 101.746 0.241331 0.775854 4.25403 0.0586695 0.0401324 0.959868 0.0197269 0.00436153 0.0189895 0.00418362 0.0052731 0.00601048 0.210924 0.240419 58.0099 -87.8968 126.259 15.9585 145.023 0.000141181 0.267196 192.83 0.310459 0.0673578 0.00409659 0.000561961 0.00138374 0.986977 0.991726 -2.98077e-06 -85.6629 0.0930309 31183 303.761 0.98351 0.319146 0.732377 0.732373 9.99958 2.98337e-06 1.19334e-05 0.131853 0.982834 0.931749 -0.0132925 4.91206e-06 0.505838 -1.92947e-20 7.13009e-24 -1.92876e-20 0.00139574 0.997817 8.59725e-05 0.152636 2.85221 0.00139574 0.997818 0.738895 0.0010567 0.00188046 0.000859725 0.455528 0.00188046 0.440663 0.000129579 1.02 0.888078 0.534569 0.286604 1.71777e-07 3.06988e-09 2381.19 3114.81 -0.0555501 0.482161 0.277452 0.253218 -0.593382 -0.169534 0.496168 -0.267113 -0.229064 2.032 1 0 297.7 0 2.14584 2.03 0.000299706 0.85354 0.672425 0.352599 0.419672 2.14604 134.393 83.9297 18.7214 60.8707 0.00402493 0 -40 10
1.131 3.27512e-08 2.53916e-06 0.120466 0.120464 0.0120349 1.48869e-05 0.00115417 0.150582 0.000658292 0.151236 0.898798 101.746 0.241321 0.775969 4.25438 0.0586787 0.0401356 0.959864 0.0197265 0.00436182 0.0189892 0.00418387 0.00527346 0.00601084 0.210938 0.240434 58.0099 -87.8968 126.259 15.9585 145.023 0.000141182 0.267196 192.829 0.310459 0.0673578 0.00409659 0.000561962 0.00138374 0.986977 0.991726 -2.98078e-06 -85.6629 0.0930309 31183 303.769 0.98351 0.319146 0.73238 0.732376 9.99958 2.98338e-06 1.19334e-05 0.131856 0.982836 0.931749 -0.0132925 4.91209e-06 0.505851 -1.92958e-20 7.13054e-24 -1.92887e-20 0.00139574 0.997817 8.59726e-05 0.152636 2.85221 0.00139574 0.997818 0.738986 0.00105672 0.00188046 0.000859726 0.455527 0.00188046 0.44067 0.000129582 1.02 0.888079 0.534569 0.286606 1.71777e-07 3.0699e-09 2381.18 3114.82 -0.0555524 0.482161 0.277451 0.253218 -0.593382 -0.169534 0.49616 -0.267111 -0.229059 2.033 1 0 297.698 0 2.14598 2.031 0.000299705 0.853549 0.672471 0.35251 0.419696 2.14619 134.401 83.9295 18.7214 60.8706 0.00402494 0 -40 10
1.132 3.27801e-08 2.53917e-06 0.12052 0.120519 0.0120349 1.49e-05 0.00115417 0.15065 0.000658293 0.151304 0.898875 101.745 0.241312 0.776084 4.25472 0.0586879 0.0401388 0.959861 0.0197262 0.00436212 0.0189888 0.00418412 0.00527382 0.0060112 0.210953 0.240448 58.01 -87.8968 126.259 15.9584 145.023 0.000141182 0.267196 192.829 0.310458 0.0673577 0.0040966 0.000561962 0.00138375 0.986977 0.991726 -2.9808e-06 -85.6629 0.093031 31183 303.777 0.98351 0.319146 0.732383 0.732379 9.99958 2.98338e-06 1.19334e-05 0.131859 0.982838 0.931749 -0.0132925 4.91212e-06 0.505863 -1.92969e-20 7.13098e-24 -1.92898e-20 0.00139574 0.997817 8.59727e-05 0.152636 2.85222 0.00139574 0.997818 0.739077 0.00105673 0.00188046 0.000859727 0.455527 0.00188046 0.440677 0.000129585 1.02 0.88808 0.534568 0.286607 1.71777e-07 3.06992e-09 2381.16 3114.83 -0.0555546 0.482161 0.277451 0.253219 -0.593382 -0.169534 0.496153 -0.267109 -0.229053 2.034 1 0 297.696 0 2.14613 2.032 0.000299705 0.853558 0.672518 0.35242 0.419721 2.14633 134.409 83.9294 18.7214 60.8706 0.00402494 0 -40 10
1.133 3.2809e-08 2.53917e-06 0.120575 0.120573 0.0120349 1.49132e-05 0.00115417 0.150718 0.000658295 0.151372 0.898952 101.745 0.241303 0.776199 4.25506 0.0586971 0.0401421 0.959858 0.0197258 0.00436241 0.0189884 0.00418436 0.00527418 0.00601157 0.210967 0.240463 58.0101 -87.8968 126.259 15.9584 145.023 0.000141183 0.267197 192.829 0.310458 0.0673577 0.0040966 0.000561963 0.00138375 0.986977 0.991726 -2.98081e-06 -85.6629 0.0930311 31183 303.785 0.98351 0.319146 0.732387 0.732382 9.99958 2.98339e-06 1.19334e-05 0.131862 0.98284 0.93175 -0.0132925 4.91215e-06 0.505876 -1.9298e-20 7.13143e-24 -1.92908e-20 0.00139575 0.997817 8.59728e-05 0.152636 2.85222 0.00139575 0.997818 0.739167 0.00105675 0.00188047 0.000859728 0.455527 0.00188046 0.440684 0.000129588 1.02 0.888081 0.534568 0.286609 1.71777e-07 3.06995e-09 2381.14 3114.85 -0.0555569 0.482161 0.277451 0.25322 -0.593381 -0.169534 0.496145 -0.267107 -0.229048 2.035 1 0 297.694 0 2.14628 2.033 0.000299704 0.853567 0.672564 0.352331 0.419745 2.14648 134.417 83.9292 18.7214 60.8705 0.00402495 0 -40 10
1.134 3.28379e-08 2.53917e-06 0.120629 0.120628 0.0120349 1.49263e-05 0.00115417 0.150786 0.000658296 0.15144 0.899028 101.745 0.241294 0.776314 4.2554 0.0587064 0.0401453 0.959855 0.0197255 0.0043627 0.0189881 0.00418461 0.00527454 0.00601193 0.210982 0.240477 58.0101 -87.8968 126.259 15.9583 145.023 0.000141184 0.267197 192.829 0.310457 0.0673576 0.0040966 0.000561964 0.00138375 0.986977 0.991726 -2.98083e-06 -85.6628 0.0930312 31182.9 303.793 0.98351 0.319146 0.73239 0.732386 9.99958 2.98339e-06 1.19335e-05 0.131865 0.982842 0.93175 -0.0132925 4.91218e-06 0.505888 -1.92991e-20 7.13187e-24 -1.92919e-20 0.00139575 0.997817 8.59729e-05 0.152637 2.85222 0.00139575 0.997818 0.739258 0.00105677 0.00188047 0.000859729 0.455527 0.00188047 0.440691 0.000129591 1.02 0.888082 0.534568 0.28661 1.71778e-07 3.06997e-09 2381.13 3114.86 -0.0555591 0.482161 0.277451 0.253221 -0.593381 -0.169534 0.496137 -0.267105 -0.229042 2.036 1 0 297.693 0 2.14643 2.034 0.000299703 0.853577 0.67261 0.352242 0.41977 2.14663 134.424 83.9291 18.7214 60.8704 0.00402496 0 -40 10
1.135 3.28668e-08 2.53917e-06 0.120683 0.120682 0.0120349 1.49394e-05 0.00115417 0.150854 0.000658297 0.151508 0.899105 101.744 0.241284 0.77643 4.25575 0.0587156 0.0401486 0.959851 0.0197251 0.004363 0.0189877 0.00418486 0.00527491 0.0060123 0.210996 0.240492 58.0102 -87.8968 126.259 15.9583 145.023 0.000141184 0.267197 192.829 0.310457 0.0673576 0.00409661 0.000561964 0.00138375 0.986977 0.991726 -2.98084e-06 -85.6628 0.0930313 31182.9 303.801 0.98351 0.319146 0.732393 0.732389 9.99958 2.9834e-06 1.19335e-05 0.131868 0.982844 0.93175 -0.0132925 4.91221e-06 0.505901 -1.93001e-20 7.13231e-24 -1.9293e-20 0.00139575 0.997817 8.59729e-05 0.152637 2.85222 0.00139575 0.997818 0.739349 0.00105679 0.00188047 0.000859729 0.455527 0.00188047 0.440698 0.000129594 1.02 0.888083 0.534568 0.286612 1.71778e-07 3.06999e-09 2381.11 3114.87 -0.0555614 0.482161 0.27745 0.253222 -0.593381 -0.169534 0.49613 -0.267103 -0.229036 2.037 1 0 297.691 0 2.14658 2.035 0.000299703 0.853586 0.672657 0.352154 0.419794 2.14678 134.432 83.9289 18.7214 60.8703 0.00402496 0 -40 10
1.136 3.28957e-08 2.53917e-06 0.120738 0.120737 0.0120349 1.49526e-05 0.00115417 0.150922 0.000658299 0.151576 0.899181 101.744 0.241275 0.776545 4.25609 0.0587248 0.0401518 0.959848 0.0197247 0.00436329 0.0189873 0.00418511 0.00527527 0.00601266 0.211011 0.240506 58.0103 -87.8968 126.259 15.9583 145.023 0.000141185 0.267197 192.829 0.310457 0.0673575 0.00409661 0.000561965 0.00138375 0.986977 0.991726 -2.98086e-06 -85.6628 0.0930314 31182.9 303.809 0.98351 0.319146 0.732397 0.732392 9.99958 2.9834e-06 1.19335e-05 0.131871 0.982846 0.93175 -0.0132925 4.91224e-06 0.505913 -1.93012e-20 7.13276e-24 -1.92941e-20 0.00139575 0.997817 8.5973e-05 0.152637 2.85222 0.00139575 0.997818 0.739439 0.00105681 0.00188047 0.00085973 0.455526 0.00188047 0.440705 0.000129597 1.02 0.888085 0.534567 0.286613 1.71778e-07 3.07001e-09 2381.09 3114.89 -0.0555637 0.482161 0.27745 0.253223 -0.593381 -0.169534 0.496122 -0.267101 -0.229031 2.038 1 0 297.689 0 2.14672 2.036 0.000299702 0.853596 0.672703 0.352065 0.419818 2.14692 134.44 83.9287 18.7214 60.8702 0.00402497 0 -40 10
1.137 3.29246e-08 2.53917e-06 0.120792 0.120791 0.0120349 1.49657e-05 0.00115417 0.15099 0.0006583 0.151644 0.899258 101.744 0.241266 0.77666 4.25643 0.058734 0.040155 0.959845 0.0197244 0.00436359 0.018987 0.00418536 0.00527563 0.00601303 0.211025 0.240521 58.0103 -87.8968 126.259 15.9582 145.023 0.000141186 0.267197 192.828 0.310456 0.0673575 0.00409661 0.000561966 0.00138376 0.986976 0.991726 -2.98087e-06 -85.6628 0.0930315 31182.9 303.817 0.98351 0.319146 0.7324 0.732396 9.99958 2.98341e-06 1.19335e-05 0.131874 0.982848 0.93175 -0.0132925 4.91227e-06 0.505926 -1.93023e-20 7.1332e-24 -1.92952e-20 0.00139575 0.997817 8.59731e-05 0.152637 2.85222 0.00139575 0.997818 0.73953 0.00105683 0.00188047 0.000859731 0.455526 0.00188047 0.440712 0.0001296 1.02 0.888086 0.534567 0.286615 1.71778e-07 3.07004e-09 2381.08 3114.9 -0.055566 0.482161 0.27745 0.253224 -0.593381 -0.169534 0.496114 -0.267098 -0.229025 2.039 1 0 297.687 0 2.14687 2.037 0.000299701 0.853605 0.672749 0.351977 0.419843 2.14707 134.448 83.9286 18.7214 60.8702 0.00402498 0 -40 10
1.138 3.29535e-08 2.53917e-06 0.120846 0.120845 0.0120349 1.49789e-05 0.00115417 0.151058 0.000658301 0.151712 0.899335 101.743 0.241257 0.776776 4.25678 0.0587433 0.0401583 0.959842 0.019724 0.00436388 0.0189866 0.00418561 0.00527599 0.00601339 0.21104 0.240536 58.0104 -87.8968 126.259 15.9582 145.023 0.000141186 0.267198 192.828 0.310456 0.0673574 0.00409661 0.000561966 0.00138376 0.986976 0.991726 -2.98089e-06 -85.6628 0.0930316 31182.9 303.825 0.98351 0.319146 0.732403 0.732399 9.99958 2.98341e-06 1.19335e-05 0.131877 0.98285 0.93175 -0.0132925 4.91229e-06 0.505938 -1.93034e-20 7.13365e-24 -1.92963e-20 0.00139575 0.997817 8.59732e-05 0.152637 2.85222 0.00139575 0.997818 0.73962 0.00105684 0.00188047 0.000859732 0.455526 0.00188047 0.440719 0.000129603 1.02 0.888087 0.534567 0.286616 1.71779e-07 3.07006e-09 2381.06 3114.92 -0.0555683 0.482161 0.277449 0.253225 -0.59338 -0.169534 0.496106 -0.267096 -0.229019 2.04 1 0 297.685 0 2.14702 2.038 0.000299701 0.853615 0.672796 0.351888 0.419867 2.14722 134.456 83.9284 18.7213 60.8701 0.00402498 0 -40 10
1.139 3.29824e-08 2.53917e-06 0.120901 0.120899 0.0120348 1.4992e-05 0.00115417 0.151126 0.000658303 0.151779 0.899412 101.743 0.241247 0.776891 4.25712 0.0587525 0.0401615 0.959838 0.0197236 0.00436418 0.0189862 0.00418586 0.00527636 0.00601376 0.211054 0.24055 58.0105 -87.8968 126.259 15.9582 145.023 0.000141187 0.267198 192.828 0.310455 0.0673573 0.00409662 0.000561967 0.00138376 0.986976 0.991726 -2.9809e-06 -85.6628 0.0930316 31182.8 303.833 0.98351 0.319146 0.732407 0.732402 9.99958 2.98342e-06 1.19336e-05 0.13188 0.982853 0.93175 -0.0132925 4.91232e-06 0.505951 -1.93045e-20 7.1341e-24 -1.92973e-20 0.00139575 0.997817 8.59733e-05 0.152637 2.85222 0.00139575 0.997818 0.739711 0.00105686 0.00188047 0.000859733 0.455526 0.00188047 0.440726 0.000129606 1.02 0.888088 0.534566 0.286618 1.71779e-07 3.07008e-09 2381.04 3114.93 -0.0555706 0.482161 0.277449 0.253226 -0.59338 -0.169534 0.496098 -0.267094 -0.229013 2.041 1 0 297.683 0 2.14717 2.039 0.0002997 0.853624 0.672842 0.3518 0.419892 2.14737 134.464 83.9282 18.7213 60.87 0.00402499 0 -40 10
1.14 3.30113e-08 2.53917e-06 0.120955 0.120953 0.0120348 1.50051e-05 0.00115417 0.151193 0.000658304 0.151847 0.899488 101.743 0.241238 0.777006 4.25747 0.0587618 0.0401648 0.959835 0.0197233 0.00436447 0.0189859 0.00418611 0.00527672 0.00601412 0.211069 0.240565 58.0105 -87.8968 126.259 15.9581 145.023 0.000141188 0.267198 192.828 0.310455 0.0673573 0.00409662 0.000561968 0.00138376 0.986976 0.991726 -2.98092e-06 -85.6628 0.0930317 31182.8 303.841 0.98351 0.319146 0.73241 0.732406 9.99958 2.98342e-06 1.19336e-05 0.131883 0.982855 0.93175 -0.0132925 4.91235e-06 0.505963 -1.93056e-20 7.13454e-24 -1.92984e-20 0.00139575 0.997817 8.59733e-05 0.152638 2.85222 0.00139575 0.997818 0.739801 0.00105688 0.00188048 0.000859733 0.455525 0.00188048 0.440733 0.000129609 1.02 0.888089 0.534566 0.286619 1.71779e-07 3.07011e-09 2381.03 3114.94 -0.055573 0.482161 0.277449 0.253226 -0.59338 -0.169535 0.49609 -0.267092 -0.229008 2.042 1 0 297.681 0 2.14731 2.04 0.000299699 0.853634 0.672888 0.351712 0.419916 2.14752 134.472 83.928 18.7213 60.8699 0.004025 0 -40 10
1.141 3.30402e-08 2.53917e-06 0.121009 0.121008 0.0120348 1.50183e-05 0.00115417 0.151261 0.000658305 0.151915 0.899565 101.742 0.241229 0.777122 4.25782 0.058771 0.0401681 0.959832 0.0197229 0.00436477 0.0189855 0.00418636 0.00527708 0.00601449 0.211083 0.24058 58.0106 -87.8968 126.259 15.9581 145.023 0.000141188 0.267198 192.828 0.310454 0.0673572 0.00409662 0.000561968 0.00138377 0.986976 0.991726 -2.98093e-06 -85.6628 0.0930318 31182.8 303.849 0.98351 0.319146 0.732414 0.732409 9.99958 2.98343e-06 1.19336e-05 0.131886 0.982857 0.93175 -0.0132925 4.91238e-06 0.505976 -1.93067e-20 7.13499e-24 -1.92995e-20 0.00139575 0.997817 8.59734e-05 0.152638 2.85222 0.00139575 0.997818 0.739892 0.0010569 0.00188048 0.000859734 0.455525 0.00188048 0.44074 0.000129612 1.02 0.88809 0.534566 0.286621 1.71779e-07 3.07013e-09 2381.01 3114.96 -0.0555753 0.482162 0.277449 0.253227 -0.59338 -0.169535 0.496082 -0.26709 -0.229002 2.043 1 0 297.679 0 2.14746 2.041 0.000299699 0.853644 0.672934 0.351625 0.419941 2.14766 134.48 83.9279 18.7213 60.8698 0.004025 0 -40 10
1.142 3.30691e-08 2.53917e-06 0.121063 0.121062 0.0120348 1.50314e-05 0.00115417 0.151329 0.000658306 0.151982 0.899642 101.742 0.24122 0.777237 4.25816 0.0587803 0.0401713 0.959829 0.0197226 0.00436506 0.0189851 0.00418661 0.00527745 0.00601486 0.211098 0.240594 58.0106 -87.8968 126.259 15.958 145.023 0.000141189 0.267198 192.828 0.310454 0.0673572 0.00409663 0.000561969 0.00138377 0.986976 0.991726 -2.98095e-06 -85.6628 0.0930319 31182.8 303.857 0.98351 0.319146 0.732417 0.732413 9.99958 2.98343e-06 1.19336e-05 0.131889 0.982859 0.93175 -0.0132925 4.91241e-06 0.505988 -1.93077e-20 7.13543e-24 -1.93006e-20 0.00139576 0.997817 8.59735e-05 0.152638 2.85222 0.00139576 0.997818 0.739982 0.00105692 0.00188048 0.000859735 0.455525 0.00188048 0.440747 0.000129615 1.02 0.888091 0.534565 0.286622 1.7178e-07 3.07015e-09 2380.99 3114.97 -0.0555777 0.482162 0.277448 0.253228 -0.59338 -0.169535 0.496074 -0.267088 -0.228996 2.044 1 0 297.677 0 2.14761 2.042 0.000299698 0.853654 0.672981 0.351537 0.419965 2.14781 134.488 83.9277 18.7213 60.8697 0.00402501 0 -40 10
1.143 3.3098e-08 2.53917e-06 0.121117 0.121116 0.0120348 1.50446e-05 0.00115417 0.151396 0.000658308 0.15205 0.899719 101.741 0.24121 0.777353 4.25851 0.0587895 0.0401746 0.959825 0.0197222 0.00436536 0.0189848 0.00418686 0.00527781 0.00601523 0.211112 0.240609 58.0107 -87.8969 126.258 15.958 145.023 0.00014119 0.267198 192.827 0.310454 0.0673571 0.00409663 0.00056197 0.00138377 0.986976 0.991726 -2.98096e-06 -85.6628 0.093032 31182.7 303.865 0.98351 0.319146 0.732421 0.732416 9.99958 2.98344e-06 1.19336e-05 0.131892 0.982861 0.93175 -0.0132925 4.91244e-06 0.506001 -1.93088e-20 7.13588e-24 -1.93017e-20 0.00139576 0.997817 8.59736e-05 0.152638 2.85223 0.00139576 0.997818 0.740073 0.00105694 0.00188048 0.000859736 0.455525 0.00188048 0.440754 0.000129618 1.02 0.888092 0.534565 0.286624 1.7178e-07 3.07017e-09 2380.98 3114.99 -0.05558 0.482162 0.277448 0.253229 -0.593379 -0.169535 0.496066 -0.267086 -0.22899 2.045 1 0 297.676 0 2.14776 2.043 0.000299697 0.853664 0.673027 0.35145 0.419989 2.14796 134.496 83.9275 18.7213 60.8697 0.00402502 0 -40 10
1.144 3.31269e-08 2.53918e-06 0.121171 0.12117 0.0120348 1.50577e-05 0.00115417 0.151464 0.000658309 0.152117 0.899796 101.741 0.241201 0.777469 4.25886 0.0587988 0.0401779 0.959822 0.0197218 0.00436566 0.0189844 0.00418711 0.00527818 0.0060156 0.211127 0.240624 58.0108 -87.8969 126.258 15.958 145.023 0.00014119 0.267199 192.827 0.310453 0.0673571 0.00409663 0.00056197 0.00138377 0.986976 0.991726 -2.98098e-06 -85.6628 0.0930321 31182.7 303.873 0.98351 0.319146 0.732424 0.73242 9.99958 2.98344e-06 1.19337e-05 0.131895 0.982863 0.93175 -0.0132925 4.91247e-06 0.506014 -1.93099e-20 7.13633e-24 -1.93028e-20 0.00139576 0.997817 8.59737e-05 0.152638 2.85223 0.00139576 0.997818 0.740163 0.00105695 0.00188048 0.000859737 0.455525 0.00188048 0.440761 0.00012962 1.02 0.888093 0.534565 0.286625 1.7178e-07 3.0702e-09 2380.96 3115 -0.0555824 0.482162 0.277448 0.25323 -0.593379 -0.169535 0.496058 -0.267084 -0.228984 2.046 1 0 297.674 0 2.14791 2.044 0.000299697 0.853674 0.673073 0.351362 0.420014 2.14811 134.504 83.9273 18.7213 60.8696 0.00402503 0 -40 10
1.145 3.31558e-08 2.53918e-06 0.121225 0.121223 0.0120348 1.50708e-05 0.00115417 0.151531 0.00065831 0.152185 0.899873 101.741 0.241192 0.777584 4.2592 0.058808 0.0401812 0.959819 0.0197215 0.00436595 0.018984 0.00418736 0.00527854 0.00601596 0.211142 0.240639 58.0108 -87.8969 126.258 15.9579 145.023 0.000141191 0.267199 192.827 0.310453 0.067357 0.00409664 0.000561971 0.00138377 0.986976 0.991726 -2.98099e-06 -85.6627 0.0930322 31182.7 303.881 0.98351 0.319146 0.732428 0.732424 9.99958 2.98345e-06 1.19337e-05 0.131898 0.982865 0.93175 -0.0132925 4.9125e-06 0.506026 -1.9311e-20 7.13678e-24 -1.93039e-20 0.00139576 0.997817 8.59737e-05 0.152638 2.85223 0.00139576 0.997818 0.740253 0.00105697 0.00188048 0.000859737 0.455524 0.00188048 0.440768 0.000129623 1.02 0.888094 0.534564 0.286627 1.71781e-07 3.07022e-09 2380.94 3115.02 -0.0555848 0.482162 0.277447 0.253231 -0.593379 -0.169535 0.49605 -0.267082 -0.228978 2.047 1 0 297.672 0 2.14805 2.045 0.000299696 0.853684 0.673119 0.351275 0.420038 2.14825 134.512 83.9272 18.7213 60.8695 0.00402503 0 -40 10
1.146 3.31847e-08 2.53918e-06 0.121279 0.121277 0.0120347 1.5084e-05 0.00115417 0.151598 0.000658311 0.152252 0.89995 101.74 0.241183 0.7777 4.25955 0.0588173 0.0401844 0.959816 0.0197211 0.00436625 0.0189837 0.00418762 0.00527891 0.00601633 0.211156 0.240653 58.0109 -87.8969 126.258 15.9579 145.023 0.000141192 0.267199 192.827 0.310452 0.067357 0.00409664 0.000561972 0.00138378 0.986976 0.991726 -2.98101e-06 -85.6627 0.0930323 31182.7 303.889 0.98351 0.319146 0.732432 0.732427 9.99958 2.98345e-06 1.19337e-05 0.131901 0.982867 0.93175 -0.0132925 4.91253e-06 0.506039 -1.93121e-20 7.13722e-24 -1.9305e-20 0.00139576 0.997817 8.59738e-05 0.152638 2.85223 0.00139576 0.997818 0.740344 0.00105699 0.00188049 0.000859738 0.455524 0.00188048 0.440776 0.000129626 1.02 0.888095 0.534564 0.286628 1.71781e-07 3.07024e-09 2380.93 3115.03 -0.0555872 0.482162 0.277447 0.253232 -0.593379 -0.169535 0.496042 -0.267079 -0.228972 2.048 1 0 297.67 0 2.1482 2.046 0.000299695 0.853694 0.673165 0.351188 0.420062 2.1484 134.519 83.927 18.7213 60.8694 0.00402504 0 -40 10
1.147 3.32136e-08 2.53918e-06 0.121332 0.121331 0.0120347 1.50971e-05 0.00115417 0.151666 0.000658313 0.152319 0.900027 101.74 0.241173 0.777816 4.2599 0.0588266 0.0401877 0.959812 0.0197207 0.00436655 0.0189833 0.00418787 0.00527927 0.0060167 0.211171 0.240668 58.011 -87.8969 126.258 15.9579 145.024 0.000141192 0.267199 192.827 0.310452 0.0673569 0.00409664 0.000561972 0.00138378 0.986976 0.991726 -2.98102e-06 -85.6627 0.0930323 31182.7 303.898 0.98351 0.319146 0.732435 0.732431 9.99958 2.98345e-06 1.19337e-05 0.131905 0.982869 0.93175 -0.0132925 4.91256e-06 0.506051 -1.93132e-20 7.13767e-24 -1.93061e-20 0.00139576 0.997817 8.59739e-05 0.152639 2.85223 0.00139576 0.997818 0.740434 0.00105701 0.00188049 0.000859739 0.455524 0.00188049 0.440783 0.000129629 1.02 0.888097 0.534564 0.28663 1.71781e-07 3.07027e-09 2380.91 3115.05 -0.0555896 0.482162 0.277447 0.253233 -0.593379 -0.169535 0.496034 -0.267077 -0.228966 2.049 1 0 297.668 0 2.14835 2.047 0.000299695 0.853704 0.673212 0.351101 0.420087 2.14855 134.527 83.9268 18.7213 60.8693 0.00402505 0 -40 10
1.148 3.32425e-08 2.53918e-06 0.121386 0.121385 0.0120347 1.51102e-05 0.00115417 0.151733 0.000658314 0.152387 0.900104 101.74 0.241164 0.777932 4.26025 0.0588359 0.040191 0.959809 0.0197204 0.00436685 0.0189829 0.00418812 0.00527964 0.00601707 0.211186 0.240683 58.011 -87.8969 126.258 15.9578 145.024 0.000141193 0.267199 192.827 0.310451 0.0673569 0.00409665 0.000561973 0.00138378 0.986976 0.991726 -2.98104e-06 -85.6627 0.0930324 31182.6 303.906 0.98351 0.319146 0.732439 0.732435 9.99958 2.98346e-06 1.19337e-05 0.131908 0.982871 0.93175 -0.0132925 4.91259e-06 0.506064 -1.93143e-20 7.13812e-24 -1.93072e-20 0.00139576 0.997817 8.5974e-05 0.152639 2.85223 0.00139576 0.997818 0.740524 0.00105703 0.00188049 0.00085974 0.455524 0.00188049 0.44079 0.000129632 1.02 0.888098 0.534564 0.286631 1.71781e-07 3.07029e-09 2380.89 3115.06 -0.055592 0.482162 0.277447 0.253234 -0.593378 -0.169535 0.496026 -0.267075 -0.22896 2.05 1 0 297.666 0 2.1485 2.048 0.000299694 0.853714 0.673258 0.351014 0.420111 2.1487 134.535 83.9266 18.7212 60.8692 0.00402506 0 -40 10
1.149 3.32714e-08 2.53918e-06 0.12144 0.121439 0.0120347 1.51234e-05 0.00115417 0.1518 0.000658315 0.152454 0.900181 101.739 0.241155 0.778048 4.2606 0.0588451 0.0401943 0.959806 0.01972 0.00436714 0.0189826 0.00418837 0.00528001 0.00601744 0.2112 0.240698 58.0111 -87.8969 126.258 15.9578 145.024 0.000141194 0.2672 192.826 0.310451 0.0673568 0.00409665 0.000561974 0.00138378 0.986976 0.991726 -2.98105e-06 -85.6627 0.0930325 31182.6 303.914 0.98351 0.319146 0.732443 0.732439 9.99958 2.98346e-06 1.19338e-05 0.131911 0.982873 0.93175 -0.0132925 4.91262e-06 0.506077 -1.93154e-20 7.13857e-24 -1.93083e-20 0.00139576 0.997817 8.59741e-05 0.152639 2.85223 0.00139576 0.997818 0.740614 0.00105705 0.00188049 0.000859741 0.455523 0.00188049 0.440797 0.000129635 1.02 0.888099 0.534563 0.286633 1.71782e-07 3.07031e-09 2380.88 3115.08 -0.0555944 0.482162 0.277446 0.253235 -0.593378 -0.169535 0.496018 -0.267073 -0.228954 2.051 1 0 297.664 0 2.14864 2.049 0.000299693 0.853725 0.673304 0.350928 0.420136 2.14884 134.543 83.9264 18.7212 60.8691 0.00402506 0 -40 10
1.15 3.33003e-08 2.53918e-06 0.121494 0.121493 0.0120347 1.51365e-05 0.00115417 0.151867 0.000658316 0.152521 0.900258 101.739 0.241146 0.778163 4.26095 0.0588544 0.0401976 0.959802 0.0197196 0.00436744 0.0189822 0.00418863 0.00528037 0.00601781 0.211215 0.240712 58.0111 -87.8969 126.258 15.9577 145.024 0.000141195 0.2672 192.826 0.310451 0.0673568 0.00409665 0.000561974 0.00138379 0.986976 0.991726 -2.98107e-06 -85.6627 0.0930326 31182.6 303.922 0.98351 0.319146 0.732447 0.732442 9.99958 2.98347e-06 1.19338e-05 0.131914 0.982875 0.93175 -0.0132925 4.91265e-06 0.506089 -1.93165e-20 7.13902e-24 -1.93094e-20 0.00139577 0.997817 8.59741e-05 0.152639 2.85223 0.00139577 0.997818 0.740704 0.00105706 0.00188049 0.000859741 0.455523 0.00188049 0.440804 0.000129638 1.02 0.8881 0.534563 0.286634 1.71782e-07 3.07034e-09 2380.86 3115.09 -0.0555968 0.482162 0.277446 0.253236 -0.593378 -0.169535 0.49601 -0.267071 -0.228948 2.052 1 0 297.662 0 2.14879 2.05 0.000299693 0.853735 0.67335 0.350841 0.42016 2.14899 134.551 83.9262 18.7212 60.869 0.00402507 0 -40 10
1.151 3.33292e-08 2.53918e-06 0.121547 0.121546 0.0120347 1.51496e-05 0.00115417 0.151934 0.000658318 0.152588 0.900335 101.739 0.241136 0.778279 4.2613 0.0588637 0.0402009 0.959799 0.0197193 0.00436774 0.0189818 0.00418888 0.00528074 0.00601818 0.21123 0.240727 58.0112 -87.8969 126.258 15.9577 145.024 0.000141195 0.2672 192.826 0.31045 0.0673567 0.00409665 0.000561975 0.00138379 0.986976 0.991726 -2.98108e-06 -85.6627 0.0930327 31182.6 303.93 0.98351 0.319146 0.73245 0.732446 9.99958 2.98347e-06 1.19338e-05 0.131917 0.982877 0.93175 -0.0132925 4.91268e-06 0.506102 -1.93176e-20 7.13947e-24 -1.93105e-20 0.00139577 0.997817 8.59742e-05 0.152639 2.85223 0.00139577 0.997818 0.740795 0.00105708 0.00188049 0.000859742 0.455523 0.00188049 0.440811 0.000129641 1.02 0.888101 0.534563 0.286636 1.71782e-07 3.07036e-09 2380.84 3115.11 -0.0555993 0.482162 0.277446 0.253237 -0.593378 -0.169535 0.496001 -0.267069 -0.228942 2.053 1 0 297.66 0 2.14894 2.051 0.000299692 0.853746 0.673396 0.350755 0.420184 2.14914 134.559 83.9261 18.7212 60.869 0.00402508 0 -40 10
1.152 3.33581e-08 2.53918e-06 0.121601 0.1216 0.0120347 1.51628e-05 0.00115417 0.152001 0.000658319 0.152655 0.900413 101.738 0.241127 0.778395 4.26165 0.058873 0.0402042 0.959796 0.0197189 0.00436804 0.0189814 0.00418913 0.00528111 0.00601855 0.211244 0.240742 58.0113 -87.8969 126.258 15.9577 145.024 0.000141196 0.2672 192.826 0.31045 0.0673567 0.00409666 0.000561976 0.00138379 0.986976 0.991726 -2.9811e-06 -85.6627 0.0930328 31182.5 303.938 0.98351 0.319146 0.732454 0.73245 9.99958 2.98348e-06 1.19338e-05 0.13192 0.982879 0.93175 -0.0132925 4.91271e-06 0.506115 -1.93187e-20 7.13992e-24 -1.93116e-20 0.00139577 0.997817 8.59743e-05 0.152639 2.85223 0.00139577 0.997818 0.740885 0.0010571 0.00188049 0.000859743 0.455523 0.00188049 0.440818 0.000129644 1.02 0.888102 0.534562 0.286637 1.71782e-07 3.07038e-09 2380.83 3115.12 -0.0556017 0.482162 0.277446 0.253238 -0.593377 -0.169535 0.495993 -0.267067 -0.228936 2.054 1 0 297.658 0 2.14908 2.052 0.000299691 0.853756 0.673443 0.350669 0.420209 2.14928 134.567 83.9259 18.7212 60.8689 0.00402509 0 -40 10
1.153 3.3387e-08 2.53918e-06 0.121655 0.121653 0.0120347 1.51759e-05 0.00115417 0.152068 0.00065832 0.152722 0.90049 101.738 0.241118 0.778511 4.262 0.0588823 0.0402076 0.959792 0.0197185 0.00436834 0.0189811 0.00418939 0.00528148 0.00601893 0.211259 0.240757 58.0113 -87.8969 126.258 15.9576 145.024 0.000141197 0.2672 192.826 0.310449 0.0673566 0.00409666 0.000561976 0.00138379 0.986976 0.991726 -2.98111e-06 -85.6627 0.0930329 31182.5 303.946 0.98351 0.319146 0.732458 0.732454 9.99958 2.98348e-06 1.19338e-05 0.131923 0.982881 0.93175 -0.0132925 4.91274e-06 0.506128 -1.93198e-20 7.14037e-24 -1.93127e-20 0.00139577 0.997817 8.59744e-05 0.15264 2.85223 0.00139577 0.997818 0.740975 0.00105712 0.0018805 0.000859744 0.455522 0.00188049 0.440825 0.000129647 1.02 0.888103 0.534562 0.286639 1.71783e-07 3.0704e-09 2380.81 3115.14 -0.0556042 0.482162 0.277445 0.253239 -0.593377 -0.169535 0.495985 -0.267065 -0.228929 2.055 1 0 297.656 0 2.14923 2.053 0.000299691 0.853767 0.673489 0.350583 0.420233 2.14943 134.575 83.9257 18.7212 60.8688 0.0040251 0 -40 10
1.154 3.34159e-08 2.53918e-06 0.121708 0.121707 0.0120346 1.51891e-05 0.00115417 0.152135 0.000658321 0.152789 0.900567 101.738 0.241108 0.778628 4.26235 0.0588916 0.0402109 0.959789 0.0197182 0.00436864 0.0189807 0.00418964 0.00528185 0.0060193 0.211274 0.240772 58.0114 -87.8969 126.258 15.9576 145.024 0.000141198 0.267201 192.826 0.310449 0.0673566 0.00409666 0.000561977 0.00138379 0.986976 0.991726 -2.98113e-06 -85.6627 0.0930329 31182.5 303.954 0.98351 0.319146 0.732462 0.732458 9.99958 2.98349e-06 1.19339e-05 0.131926 0.982883 0.93175 -0.0132925 4.91277e-06 0.50614 -1.93209e-20 7.14082e-24 -1.93138e-20 0.00139577 0.997817 8.59745e-05 0.15264 2.85224 0.00139577 0.997818 0.741065 0.00105714 0.0018805 0.000859745 0.455522 0.0018805 0.440832 0.00012965 1.02 0.888104 0.534562 0.286641 1.71783e-07 3.07043e-09 2380.79 3115.15 -0.0556067 0.482163 0.277445 0.25324 -0.593377 -0.169535 0.495976 -0.267063 -0.228923 2.056 1 0 297.654 0 2.14938 2.054 0.00029969 0.853777 0.673535 0.350497 0.420257 2.14958 134.583 83.9255 18.7212 60.8687 0.0040251 0 -40 10
1.155 3.34448e-08 2.53918e-06 0.121762 0.12176 0.0120346 1.52022e-05 0.00115417 0.152202 0.000658323 0.152856 0.900644 101.737 0.241099 0.778744 4.2627 0.0589009 0.0402142 0.959786 0.0197178 0.00436894 0.0189803 0.00418989 0.00528222 0.00601967 0.211289 0.240787 58.0115 -87.8969 126.258 15.9575 145.024 0.000141198 0.267201 192.825 0.310448 0.0673565 0.00409667 0.000561978 0.0013838 0.986976 0.991726 -2.98114e-06 -85.6627 0.093033 31182.5 303.962 0.98351 0.319146 0.732466 0.732462 9.99958 2.98349e-06 1.19339e-05 0.131929 0.982885 0.93175 -0.0132925 4.9128e-06 0.506153 -1.9322e-20 7.14127e-24 -1.93149e-20 0.00139577 0.997817 8.59746e-05 0.15264 2.85224 0.00139577 0.997818 0.741155 0.00105716 0.0018805 0.000859746 0.455522 0.0018805 0.440839 0.000129653 1.02 0.888105 0.534561 0.286642 1.71783e-07 3.07045e-09 2380.78 3115.17 -0.0556092 0.482163 0.277445 0.253241 -0.593377 -0.169535 0.495968 -0.26706 -0.228917 2.057 1 0 297.651 0 2.14953 2.055 0.000299689 0.853788 0.673581 0.350412 0.420282 2.14973 134.591 83.9253 18.7212 60.8686 0.00402511 0 -40 10
1.156 3.34737e-08 2.53919e-06 0.121815 0.121814 0.0120346 1.52153e-05 0.00115418 0.152269 0.000658324 0.152923 0.900721 101.737 0.24109 0.77886 4.26306 0.0589102 0.0402175 0.959782 0.0197174 0.00436924 0.01898 0.00419015 0.00528259 0.00602004 0.211303 0.240802 58.0115 -87.8969 126.258 15.9575 145.024 0.000141199 0.267201 192.825 0.310448 0.0673565 0.00409667 0.000561978 0.0013838 0.986976 0.991726 -2.98116e-06 -85.6626 0.0930331 31182.5 303.971 0.98351 0.319146 0.73247 0.732466 9.99958 2.9835e-06 1.19339e-05 0.131932 0.982887 0.93175 -0.0132925 4.91283e-06 0.506166 -1.93231e-20 7.14172e-24 -1.9316e-20 0.00139577 0.997817 8.59746e-05 0.15264 2.85224 0.00139577 0.997818 0.741245 0.00105717 0.0018805 0.000859746 0.455522 0.0018805 0.440846 0.000129656 1.02 0.888106 0.534561 0.286644 1.71784e-07 3.07047e-09 2380.76 3115.19 -0.0556116 0.482163 0.277444 0.253243 -0.593377 -0.169536 0.49596 -0.267058 -0.228911 2.058 1 0 297.649 0 2.14967 2.056 0.000299688 0.853799 0.673627 0.350326 0.420306 2.14987 134.598 83.9251 18.7212 60.8685 0.00402512 0 -40 10
1.157 3.35026e-08 2.53919e-06 0.121869 0.121867 0.0120346 1.52285e-05 0.00115418 0.152336 0.000658325 0.152989 0.900799 101.737 0.241081 0.778976 4.26341 0.0589195 0.0402208 0.959779 0.019717 0.00436954 0.0189796 0.0041904 0.00528295 0.00602042 0.211318 0.240817 58.0116 -87.8969 126.257 15.9575 145.024 0.0001412 0.267201 192.825 0.310448 0.0673564 0.00409667 0.000561979 0.0013838 0.986976 0.991726 -2.98117e-06 -85.6626 0.0930332 31182.4 303.979 0.98351 0.319146 0.732474 0.73247 9.99958 2.9835e-06 1.19339e-05 0.131935 0.982889 0.93175 -0.0132925 4.91286e-06 0.506179 -1.93242e-20 7.14217e-24 -1.93171e-20 0.00139577 0.997816 8.59747e-05 0.15264 2.85224 0.00139577 0.997818 0.741335 0.00105719 0.0018805 0.000859747 0.455522 0.0018805 0.440853 0.000129659 1.02 0.888108 0.534561 0.286645 1.71784e-07 3.0705e-09 2380.74 3115.2 -0.0556141 0.482163 0.277444 0.253244 -0.593376 -0.169536 0.495951 -0.267056 -0.228904 2.059 1 0 297.647 0 2.14982 2.057 0.000299688 0.853809 0.673673 0.350241 0.42033 2.15002 134.606 83.9249 18.7211 60.8684 0.00402513 0 -40 10
1.158 3.35315e-08 2.53919e-06 0.121922 0.121921 0.0120346 1.52416e-05 0.00115418 0.152402 0.000658326 0.153056 0.900876 101.736 0.241071 0.779092 4.26376 0.0589288 0.0402242 0.959776 0.0197167 0.00436984 0.0189792 0.00419066 0.00528333 0.00602079 0.211333 0.240832 58.0117 -87.8969 126.257 15.9574 145.024 0.000141201 0.267201 192.825 0.310447 0.0673563 0.00409668 0.00056198 0.0013838 0.986976 0.991726 -2.98119e-06 -85.6626 0.0930333 31182.4 303.987 0.98351 0.319146 0.732478 0.732474 9.99958 2.98351e-06 1.19339e-05 0.131938 0.982891 0.93175 -0.0132925 4.91289e-06 0.506191 -1.93253e-20 7.14262e-24 -1.93182e-20 0.00139577 0.997816 8.59748e-05 0.15264 2.85224 0.00139577 0.997818 0.741425 0.00105721 0.0018805 0.000859748 0.455521 0.0018805 0.44086 0.000129661 1.02 0.888109 0.53456 0.286647 1.71784e-07 3.07052e-09 2380.73 3115.22 -0.0556167 0.482163 0.277444 0.253245 -0.593376 -0.169536 0.495943 -0.267054 -0.228898 2.06 1 0 297.645 0 2.14997 2.058 0.000299687 0.85382 0.673719 0.350155 0.420355 2.15017 134.614 83.9247 18.7211 60.8683 0.00402514 0 -40 10
1.159 3.35604e-08 2.53919e-06 0.121975 0.121974 0.0120346 1.52547e-05 0.00115418 0.152469 0.000658328 0.153123 0.900954 101.736 0.241062 0.779209 4.26412 0.0589381 0.0402275 0.959772 0.0197163 0.00437014 0.0189788 0.00419091 0.0052837 0.00602116 0.211348 0.240847 58.0117 -87.8969 126.257 15.9574 145.024 0.000141201 0.267202 192.825 0.310447 0.0673563 0.00409668 0.00056198 0.0013838 0.986976 0.991726 -2.9812e-06 -85.6626 0.0930334 31182.4 303.995 0.98351 0.319146 0.732482 0.732478 9.99958 2.98351e-06 1.1934e-05 0.131941 0.982892 0.93175 -0.0132925 4.91292e-06 0.506204 -1.93264e-20 7.14307e-24 -1.93193e-20 0.00139578 0.997816 8.59749e-05 0.15264 2.85224 0.00139578 0.997818 0.741514 0.00105723 0.0018805 0.000859749 0.455521 0.0018805 0.440867 0.000129664 1.02 0.88811 0.53456 0.286648 1.71784e-07 3.07054e-09 2380.71 3115.23 -0.0556192 0.482163 0.277444 0.253246 -0.593376 -0.169536 0.495934 -0.267052 -0.228892 2.061 1 0 297.643 0 2.15012 2.059 0.000299686 0.853831 0.673765 0.35007 0.420379 2.15032 134.622 83.9245 18.7211 60.8682 0.00402514 0 -40 10
1.16 3.35893e-08 2.53919e-06 0.122029 0.122027 0.0120346 1.52679e-05 0.00115418 0.152536 0.000658329 0.153189 0.901031 101.736 0.241053 0.779325 4.26447 0.0589474 0.0402309 0.959769 0.0197159 0.00437044 0.0189785 0.00419117 0.00528407 0.00602154 0.211363 0.240862 58.0118 -87.8969 126.257 15.9574 145.024 0.000141202 0.267202 192.825 0.310446 0.0673562 0.00409668 0.000561981 0.00138381 0.986976 0.991726 -2.98122e-06 -85.6626 0.0930335 31182.4 304.003 0.98351 0.319146 0.732486 0.732482 9.99958 2.98352e-06 1.1934e-05 0.131944 0.982894 0.93175 -0.0132925 4.91295e-06 0.506217 -1.93275e-20 7.14353e-24 -1.93204e-20 0.00139578 0.997816 8.5975e-05 0.152641 2.85224 0.00139578 0.997818 0.741604 0.00105725 0.00188051 0.00085975 0.455521 0.0018805 0.440874 0.000129667 1.02 0.888111 0.53456 0.28665 1.71785e-07 3.07056e-09 2380.69 3115.25 -0.0556217 0.482163 0.277443 0.253247 -0.593376 -0.169536 0.495926 -0.26705 -0.228885 2.062 1 0 297.641 0 2.15026 2.06 0.000299686 0.853842 0.673812 0.349985 0.420403 2.15046 134.63 83.9243 18.7211 60.8681 0.00402515 0 -40 10
1.161 3.36182e-08 2.53919e-06 0.122082 0.122081 0.0120345 1.5281e-05 0.00115418 0.152602 0.00065833 0.153256 0.901108 101.735 0.241043 0.779441 4.26483 0.0589568 0.0402342 0.959766 0.0197156 0.00437075 0.0189781 0.00419142 0.00528444 0.00602191 0.211378 0.240877 58.0118 -87.8969 126.257 15.9573 145.024 0.000141203 0.267202 192.824 0.310446 0.0673562 0.00409668 0.000561982 0.00138381 0.986976 0.991726 -2.98123e-06 -85.6626 0.0930336 31182.3 304.011 0.98351 0.319146 0.73249 0.732486 9.99958 2.98352e-06 1.1934e-05 0.131947 0.982896 0.93175 -0.0132925 4.91298e-06 0.50623 -1.93286e-20 7.14398e-24 -1.93215e-20 0.00139578 0.997816 8.5975e-05 0.152641 2.85224 0.00139578 0.997818 0.741694 0.00105727 0.00188051 0.00085975 0.455521 0.00188051 0.44088 0.00012967 1.02 0.888112 0.53456 0.286651 1.71785e-07 3.07059e-09 2380.68 3115.27 -0.0556242 0.482163 0.277443 0.253248 -0.593375 -0.169536 0.495917 -0.267048 -0.228879 2.063 1 0 297.639 0 2.15041 2.061 0.000299685 0.853853 0.673858 0.349901 0.420428 2.15061 134.638 83.9241 18.7211 60.868 0.00402516 0 -40 10
1.162 3.36471e-08 2.53919e-06 0.122135 0.122134 0.0120345 1.52942e-05 0.00115418 0.152669 0.000658331 0.153322 0.901186 101.735 0.241034 0.779558 4.26518 0.0589661 0.0402376 0.959762 0.0197152 0.00437105 0.0189777 0.00419168 0.00528481 0.00602229 0.211392 0.240892 58.0119 -87.8969 126.257 15.9573 145.024 0.000141204 0.267202 192.824 0.310445 0.0673561 0.00409669 0.000561982 0.00138381 0.986976 0.991726 -2.98125e-06 -85.6626 0.0930336 31182.3 304.02 0.98351 0.319146 0.732494 0.73249 9.99958 2.98353e-06 1.1934e-05 0.13195 0.982898 0.93175 -0.0132925 4.91301e-06 0.506243 -1.93297e-20 7.14443e-24 -1.93226e-20 0.00139578 0.997816 8.59751e-05 0.152641 2.85224 0.00139578 0.997818 0.741784 0.00105728 0.00188051 0.000859751 0.45552 0.00188051 0.440887 0.000129673 1.02 0.888113 0.534559 0.286653 1.71785e-07 3.07061e-09 2380.66 3115.29 -0.0556268 0.482163 0.277443 0.253249 -0.593375 -0.169536 0.495909 -0.267046 -0.228872 2.064 1 0 297.637 0 2.15056 2.062 0.000299684 0.853864 0.673904 0.349816 0.420452 2.15076 134.646 83.9239 18.7211 60.8679 0.00402517 0 -40 10
1.163 3.3676e-08 2.53919e-06 0.122188 0.122187 0.0120345 1.53073e-05 0.00115418 0.152735 0.000658333 0.153389 0.901263 101.734 0.241025 0.779674 4.26554 0.0589754 0.0402409 0.959759 0.0197148 0.00437135 0.0189773 0.00419194 0.00528518 0.00602266 0.211407 0.240907 58.012 -87.8969 126.257 15.9572 145.024 0.000141205 0.267202 192.824 0.310445 0.0673561 0.00409669 0.000561983 0.00138381 0.986976 0.991726 -2.98126e-06 -85.6626 0.0930337 31182.3 304.028 0.98351 0.319146 0.732499 0.732494 9.99958 2.98353e-06 1.1934e-05 0.131954 0.9829 0.93175 -0.0132925 4.91304e-06 0.506256 -1.93308e-20 7.14488e-24 -1.93237e-20 0.00139578 0.997816 8.59752e-05 0.152641 2.85224 0.00139578 0.997818 0.741874 0.0010573 0.00188051 0.000859752 0.45552 0.00188051 0.440894 0.000129676 1.02 0.888114 0.534559 0.286654 1.71785e-07 3.07063e-09 2380.64 3115.3 -0.0556293 0.482163 0.277442 0.25325 -0.593375 -0.169536 0.4959 -0.267044 -0.228866 2.065 1 0 297.635 0 2.1507 2.063 0.000299684 0.853876 0.67395 0.349732 0.420476 2.1509 134.654 83.9237 18.7211 60.8678 0.00402518 0 -40 10
1.164 3.37049e-08 2.53919e-06 0.122241 0.12224 0.0120345 1.53204e-05 0.00115418 0.152802 0.000658334 0.153455 0.901341 101.734 0.241015 0.779791 4.26589 0.0589847 0.0402443 0.959756 0.0197144 0.00437165 0.018977 0.00419219 0.00528555 0.00602304 0.211422 0.240922 58.012 -87.8969 126.257 15.9572 145.024 0.000141205 0.267202 192.824 0.310445 0.067356 0.00409669 0.000561984 0.00138382 0.986976 0.991726 -2.98128e-06 -85.6626 0.0930338 31182.3 304.036 0.983509 0.319146 0.732503 0.732498 9.99958 2.98354e-06 1.1934e-05 0.131957 0.982902 0.93175 -0.0132925 4.91307e-06 0.506269 -1.93319e-20 7.14534e-24 -1.93248e-20 0.00139578 0.997816 8.59753e-05 0.152641 2.85225 0.00139578 0.997818 0.741963 0.00105732 0.00188051 0.000859753 0.45552 0.00188051 0.440901 0.000129679 1.02 0.888115 0.534559 0.286656 1.71786e-07 3.07066e-09 2380.63 3115.32 -0.0556319 0.482163 0.277442 0.253251 -0.593375 -0.169536 0.495892 -0.267041 -0.228859 2.066 1 0 297.633 0 2.15085 2.064 0.000299683 0.853887 0.673996 0.349647 0.4205 2.15105 134.662 83.9235 18.7211 60.8677 0.00402519 0 -40 10
1.165 3.37338e-08 2.53919e-06 0.122294 0.122293 0.0120345 1.53336e-05 0.00115418 0.152868 0.000658335 0.153522 0.901418 101.734 0.241006 0.779907 4.26625 0.0589941 0.0402476 0.959752 0.0197141 0.00437196 0.0189766 0.00419245 0.00528593 0.00602342 0.211437 0.240937 58.0121 -87.8969 126.257 15.9572 145.024 0.000141206 0.267203 192.824 0.310444 0.067356 0.0040967 0.000561984 0.00138382 0.986976 0.991726 -2.98129e-06 -85.6626 0.0930339 31182.3 304.044 0.983509 0.319146 0.732507 0.732503 9.99958 2.98354e-06 1.19341e-05 0.13196 0.982904 0.93175 -0.0132925 4.9131e-06 0.506281 -1.9333e-20 7.14579e-24 -1.93259e-20 0.00139578 0.997816 8.59754e-05 0.152641 2.85225 0.00139578 0.997818 0.742053 0.00105734 0.00188051 0.000859754 0.45552 0.00188051 0.440908 0.000129682 1.02 0.888116 0.534558 0.286657 1.71786e-07 3.07068e-09 2380.61 3115.34 -0.0556345 0.482163 0.277442 0.253253 -0.593374 -0.169536 0.495883 -0.267039 -0.228853 2.067 1 0 297.63 0 2.151 2.065 0.000299682 0.853898 0.674042 0.349563 0.420525 2.1512 134.669 83.9233 18.7211 60.8676 0.00402519 0 -40 10
1.166 3.37627e-08 2.53919e-06 0.122347 0.122346 0.0120345 1.53467e-05 0.00115418 0.152934 0.000658336 0.153588 0.901496 101.733 0.240997 0.780024 4.26661 0.0590034 0.040251 0.959749 0.0197137 0.00437226 0.0189762 0.00419271 0.0052863 0.00602379 0.211452 0.240952 58.0122 -87.8969 126.257 15.9571 145.024 0.000141207 0.267203 192.824 0.310444 0.0673559 0.0040967 0.000561985 0.00138382 0.986976 0.991726 -2.98131e-06 -85.6625 0.093034 31182.2 304.052 0.983509 0.319146 0.732511 0.732507 9.99958 2.98355e-06 1.19341e-05 0.131963 0.982906 0.93175 -0.0132924 4.91313e-06 0.506294 -1.93342e-20 7.14625e-24 -1.9327e-20 0.00139578 0.997816 8.59754e-05 0.152642 2.85225 0.00139578 0.997818 0.742143 0.00105736 0.00188052 0.000859754 0.45552 0.00188051 0.440915 0.000129685 1.02 0.888117 0.534558 0.286659 1.71786e-07 3.0707e-09 2380.59 3115.35 -0.0556371 0.482163 0.277442 0.253254 -0.593374 -0.169536 0.495874 -0.267037 -0.228846 2.068 1 0 297.628 0 2.15115 2.066 0.000299682 0.853909 0.674088 0.349479 0.420549 2.15134 134.677 83.9231 18.721 60.8675 0.0040252 0 -40 10
1.167 3.37916e-08 2.53919e-06 0.1224 0.122399 0.0120345 1.53598e-05 0.00115418 0.153 0.000658337 0.153654 0.901574 101.733 0.240987 0.780141 4.26696 0.0590128 0.0402544 0.959746 0.0197133 0.00437256 0.0189758 0.00419296 0.00528667 0.00602417 0.211467 0.240967 58.0122 -87.8969 126.257 15.9571 145.024 0.000141208 0.267203 192.823 0.310443 0.0673559 0.0040967 0.000561986 0.00138382 0.986976 0.991726 -2.98132e-06 -85.6625 0.0930341 31182.2 304.061 0.983509 0.319146 0.732516 0.732511 9.99958 2.98355e-06 1.19341e-05 0.131966 0.982908 0.93175 -0.0132924 4.91315e-06 0.506307 -1.93353e-20 7.1467e-24 -1.93281e-20 0.00139578 0.997816 8.59755e-05 0.152642 2.85225 0.00139578 0.997818 0.742232 0.00105737 0.00188052 0.000859755 0.455519 0.00188052 0.440922 0.000129688 1.02 0.888119 0.534558 0.28666 1.71787e-07 3.07072e-09 2380.58 3115.37 -0.0556397 0.482163 0.277441 0.253255 -0.593374 -0.169536 0.495865 -0.267035 -0.22884 2.069 1 0 297.626 0 2.15129 2.067 0.000299681 0.853921 0.674134 0.349395 0.420573 2.15149 134.685 83.9228 18.721 60.8674 0.00402521 0 -40 10
1.168 3.38205e-08 2.5392e-06 0.122453 0.122452 0.0120344 1.5373e-05 0.00115418 0.153067 0.000658339 0.15372 0.901651 101.733 0.240978 0.780257 4.26732 0.0590221 0.0402578 0.959742 0.019713 0.00437287 0.0189755 0.00419322 0.00528705 0.00602455 0.211482 0.240982 58.0123 -87.8969 126.257 15.9571 145.024 0.000141209 0.267203 192.823 0.310443 0.0673558 0.00409671 0.000561986 0.00138382 0.986976 0.991726 -2.98134e-06 -85.6625 0.0930342 31182.2 304.069 0.983509 0.319146 0.73252 0.732515 9.99958 2.98356e-06 1.19341e-05 0.131969 0.98291 0.93175 -0.0132924 4.91318e-06 0.50632 -1.93364e-20 7.14715e-24 -1.93292e-20 0.00139579 0.997816 8.59756e-05 0.152642 2.85225 0.00139579 0.997818 0.742322 0.00105739 0.00188052 0.000859756 0.455519 0.00188052 0.440929 0.000129691 1.02 0.88812 0.534557 0.286662 1.71787e-07 3.07075e-09 2380.56 3115.39 -0.0556423 0.482164 0.277441 0.253256 -0.593374 -0.169536 0.495857 -0.267033 -0.228833 2.07 1 0 297.624 0 2.15144 2.068 0.00029968 0.853932 0.67418 0.349311 0.420598 2.15164 134.693 83.9226 18.721 60.8673 0.00402522 0 -40 10
1.169 3.38494e-08 2.5392e-06 0.122506 0.122505 0.0120344 1.53861e-05 0.00115418 0.153133 0.00065834 0.153787 0.901729 101.732 0.240969 0.780374 4.26768 0.0590315 0.0402611 0.959739 0.0197126 0.00437317 0.0189751 0.00419348 0.00528742 0.00602493 0.211497 0.240997 58.0124 -87.897 126.257 15.957 145.024 0.000141209 0.267203 192.823 0.310442 0.0673558 0.00409671 0.000561987 0.00138383 0.986976 0.991726 -2.98135e-06 -85.6625 0.0930343 31182.2 304.077 0.983509 0.319146 0.732524 0.73252 9.99958 2.98356e-06 1.19341e-05 0.131972 0.982911 0.93175 -0.0132924 4.91321e-06 0.506333 -1.93375e-20 7.14761e-24 -1.93303e-20 0.00139579 0.997816 8.59757e-05 0.152642 2.85225 0.00139579 0.997818 0.742411 0.00105741 0.00188052 0.000859757 0.455519 0.00188052 0.440936 0.000129693 1.02 0.888121 0.534557 0.286663 1.71787e-07 3.07077e-09 2380.54 3115.41 -0.0556449 0.482164 0.277441 0.253257 -0.593373 -0.169536 0.495848 -0.267031 -0.228827 2.071 1 0 297.622 0 2.15159 2.069 0.00029968 0.853944 0.674226 0.349228 0.420622 2.15178 134.701 83.9224 18.721 60.8672 0.00402523 0 -40 10
1.17 3.38783e-08 2.5392e-06 0.122559 0.122558 0.0120344 1.53992e-05 0.00115418 0.153199 0.000658341 0.153853 0.901807 101.732 0.240959 0.780491 4.26804 0.0590408 0.0402645 0.959735 0.0197122 0.00437348 0.0189747 0.00419374 0.0052878 0.0060253 0.211512 0.241012 58.0124 -87.897 126.256 15.957 145.024 0.00014121 0.267204 192.823 0.310442 0.0673557 0.00409671 0.000561988 0.00138383 0.986976 0.991726 -2.98137e-06 -85.6625 0.0930343 31182.1 304.085 0.983509 0.319146 0.732529 0.732524 9.99958 2.98357e-06 1.19342e-05 0.131975 0.982913 0.93175 -0.0132924 4.91324e-06 0.506346 -1.93386e-20 7.14806e-24 -1.93314e-20 0.00139579 0.997816 8.59758e-05 0.152642 2.85225 0.00139579 0.997818 0.742501 0.00105743 0.00188052 0.000859758 0.455519 0.00188052 0.440943 0.000129696 1.02 0.888122 0.534557 0.286665 1.71787e-07 3.07079e-09 2380.53 3115.42 -0.0556475 0.482164 0.27744 0.253258 -0.593373 -0.169536 0.495839 -0.267029 -0.22882 2.072 1 0 297.62 0 2.15173 2.07 0.000299679 0.853955 0.674272 0.349144 0.420646 2.15193 134.709 83.9222 18.721 60.8671 0.00402524 0 -40 10
1.171 3.39072e-08 2.5392e-06 0.122612 0.122611 0.0120344 1.54124e-05 0.00115418 0.153265 0.000658342 0.153919 0.901884 101.732 0.24095 0.780608 4.2684 0.0590502 0.0402679 0.959732 0.0197118 0.00437378 0.0189743 0.004194 0.00528817 0.00602568 0.211527 0.241027 58.0125 -87.897 126.256 15.9569 145.024 0.000141211 0.267204 192.823 0.310442 0.0673557 0.00409671 0.000561988 0.00138383 0.986976 0.991726 -2.98138e-06 -85.6625 0.0930344 31182.1 304.094 0.983509 0.319146 0.732533 0.732529 9.99958 2.98357e-06 1.19342e-05 0.131978 0.982915 0.93175 -0.0132924 4.91327e-06 0.506359 -1.93397e-20 7.14852e-24 -1.93326e-20 0.00139579 0.997816 8.59758e-05 0.152642 2.85225 0.00139579 0.997818 0.742591 0.00105745 0.00188052 0.000859758 0.455518 0.00188052 0.44095 0.000129699 1.02 0.888123 0.534556 0.286666 1.71788e-07 3.07082e-09 2380.51 3115.44 -0.0556501 0.482164 0.27744 0.25326 -0.593373 -0.169536 0.49583 -0.267027 -0.228813 2.073 1 0 297.617 0 2.15188 2.071 0.000299678 0.853967 0.674318 0.349061 0.42067 2.15208 134.717 83.922 18.721 60.867 0.00402525 0 -40 10
1.172 3.39361e-08 2.5392e-06 0.122665 0.122663 0.0120344 1.54255e-05 0.00115418 0.153331 0.000658344 0.153985 0.901962 101.731 0.24094 0.780724 4.26876 0.0590595 0.0402713 0.959729 0.0197115 0.00437408 0.0189739 0.00419425 0.00528855 0.00602606 0.211542 0.241043 58.0125 -87.897 126.256 15.9569 145.024 0.000141212 0.267204 192.823 0.310441 0.0673556 0.00409672 0.000561989 0.00138383 0.986976 0.991726 -2.9814e-06 -85.6625 0.0930345 31182.1 304.102 0.983509 0.319146 0.732537 0.732533 9.99958 2.98358e-06 1.19342e-05 0.131982 0.982917 0.93175 -0.0132924 4.9133e-06 0.506372 -1.93408e-20 7.14898e-24 -1.93337e-20 0.00139579 0.997816 8.59759e-05 0.152642 2.85225 0.00139579 0.997818 0.74268 0.00105747 0.00188052 0.000859759 0.455518 0.00188052 0.440957 0.000129702 1.02 0.888124 0.534556 0.286668 1.71788e-07 3.07084e-09 2380.49 3115.46 -0.0556528 0.482164 0.27744 0.253261 -0.593373 -0.169537 0.495822 -0.267025 -0.228806 2.074 1 0 297.615 0 2.15203 2.072 0.000299677 0.853979 0.674364 0.348978 0.420695 2.15223 134.725 83.9218 18.721 60.8669 0.00402526 0 -40 10
1.173 3.3965e-08 2.5392e-06 0.122717 0.122716 0.0120344 1.54387e-05 0.00115418 0.153397 0.000658345 0.15405 0.90204 101.731 0.240931 0.780841 4.26912 0.0590689 0.0402747 0.959725 0.0197111 0.00437439 0.0189736 0.00419451 0.00528892 0.00602644 0.211557 0.241058 58.0126 -87.897 126.256 15.9569 145.024 0.000141213 0.267204 192.822 0.310441 0.0673556 0.00409672 0.00056199 0.00138383 0.986975 0.991726 -2.98141e-06 -85.6625 0.0930346 31182.1 304.11 0.983509 0.319146 0.732542 0.732537 9.99958 2.98358e-06 1.19342e-05 0.131985 0.982919 0.93175 -0.0132924 4.91333e-06 0.506385 -1.93419e-20 7.14943e-24 -1.93348e-20 0.00139579 0.997816 8.5976e-05 0.152643 2.85225 0.00139579 0.997818 0.742769 0.00105748 0.00188053 0.00085976 0.455518 0.00188052 0.440964 0.000129705 1.02 0.888125 0.534556 0.286669 1.71788e-07 3.07086e-09 2380.48 3115.48 -0.0556554 0.482164 0.27744 0.253262 -0.593372 -0.169537 0.495813 -0.267022 -0.2288 2.075 1 0 297.613 0 2.15217 2.073 0.000299677 0.85399 0.67441 0.348895 0.420719 2.15237 134.732 83.9215 18.721 60.8668 0.00402527 0 -40 10
1.174 3.39939e-08 2.5392e-06 0.12277 0.122769 0.0120344 1.54518e-05 0.00115418 0.153463 0.000658346 0.154116 0.902118 101.731 0.240922 0.780958 4.26948 0.0590783 0.0402781 0.959722 0.0197107 0.0043747 0.0189732 0.00419477 0.0052893 0.00602682 0.211572 0.241073 58.0127 -87.897 126.256 15.9568 145.024 0.000141214 0.267204 192.822 0.31044 0.0673555 0.00409672 0.00056199 0.00138384 0.986975 0.991726 -2.98143e-06 -85.6625 0.0930347 31182 304.119 0.983509 0.319146 0.732546 0.732542 9.99958 2.98359e-06 1.19342e-05 0.131988 0.982921 0.93175 -0.0132924 4.91336e-06 0.506398 -1.93431e-20 7.14989e-24 -1.93359e-20 0.00139579 0.997816 8.59761e-05 0.152643 2.85225 0.00139579 0.997818 0.742859 0.0010575 0.00188053 0.000859761 0.455518 0.00188053 0.440971 0.000129708 1.02 0.888126 0.534556 0.286671 1.71788e-07 3.07088e-09 2380.46 3115.5 -0.0556581 0.482164 0.277439 0.253263 -0.593372 -0.169537 0.495804 -0.26702 -0.228793 2.076 1 0 297.611 0 2.15232 2.074 0.000299676 0.854002 0.674456 0.348812 0.420743 2.15252 134.74 83.9213 18.7209 60.8667 0.00402527 0 -40 10
1.175 3.40228e-08 2.5392e-06 0.122823 0.122822 0.0120344 1.54649e-05 0.00115418 0.153528 0.000658347 0.154182 0.902196 101.73 0.240912 0.781075 4.26984 0.0590877 0.0402815 0.959718 0.0197103 0.004375 0.0189728 0.00419503 0.00528968 0.0060272 0.211587 0.241088 58.0127 -87.897 126.256 15.9568 145.024 0.000141215 0.267205 192.822 0.31044 0.0673555 0.00409673 0.000561991 0.00138384 0.986975 0.991726 -2.98144e-06 -85.6625 0.0930348 31182 304.127 0.983509 0.319146 0.732551 0.732546 9.99958 2.98359e-06 1.19343e-05 0.131991 0.982923 0.93175 -0.0132924 4.91339e-06 0.506411 -1.93442e-20 7.15034e-24 -1.9337e-20 0.00139579 0.997816 8.59762e-05 0.152643 2.85226 0.00139579 0.997818 0.742948 0.00105752 0.00188053 0.000859762 0.455518 0.00188053 0.440978 0.000129711 1.02 0.888127 0.534555 0.286672 1.71789e-07 3.07091e-09 2380.44 3115.52 -0.0556608 0.482164 0.277439 0.253264 -0.593372 -0.169537 0.495795 -0.267018 -0.228786 2.077 1 0 297.608 0 2.15247 2.075 0.000299675 0.854014 0.674502 0.348729 0.420767 2.15267 134.748 83.9211 18.7209 60.8666 0.00402528 0 -40 10
1.176 3.40517e-08 2.5392e-06 0.122875 0.122874 0.0120343 1.54781e-05 0.00115418 0.153594 0.000658348 0.154248 0.902273 101.73 0.240903 0.781192 4.2702 0.059097 0.0402849 0.959715 0.0197099 0.00437531 0.0189724 0.00419529 0.00529005 0.00602758 0.211602 0.241103 58.0128 -87.897 126.256 15.9568 145.024 0.000141216 0.267205 192.822 0.310439 0.0673554 0.00409673 0.000561992 0.00138384 0.986975 0.991726 -2.98146e-06 -85.6625 0.0930349 31182 304.135 0.983509 0.319146 0.732555 0.732551 9.99958 2.9836e-06 1.19343e-05 0.131994 0.982924 0.93175 -0.0132924 4.91342e-06 0.506424 -1.93453e-20 7.1508e-24 -1.93381e-20 0.00139579 0.997816 8.59762e-05 0.152643 2.85226 0.00139579 0.997818 0.743038 0.00105754 0.00188053 0.000859762 0.455517 0.00188053 0.440985 0.000129714 1.02 0.888128 0.534555 0.286674 1.71789e-07 3.07093e-09 2380.43 3115.53 -0.0556634 0.482164 0.277439 0.253266 -0.593372 -0.169537 0.495786 -0.267016 -0.228779 2.078 1 0 297.606 0 2.15261 2.076 0.000299675 0.854026 0.674548 0.348646 0.420791 2.15281 134.756 83.9209 18.7209 60.8665 0.00402529 0 -40 10
1.177 3.40806e-08 2.5392e-06 0.122928 0.122927 0.0120343 1.54912e-05 0.00115418 0.15366 0.00065835 0.154314 0.902351 101.729 0.240894 0.781309 4.27056 0.0591064 0.0402883 0.959712 0.0197096 0.00437561 0.018972 0.00419555 0.00529043 0.00602796 0.211617 0.241119 58.0129 -87.897 126.256 15.9567 145.024 0.000141216 0.267205 192.822 0.310439 0.0673553 0.00409673 0.000561993 0.00138384 0.986975 0.991726 -2.98147e-06 -85.6624 0.093035 31182 304.143 0.983509 0.319146 0.73256 0.732556 9.99958 2.9836e-06 1.19343e-05 0.131997 0.982926 0.931749 -0.0132924 4.91345e-06 0.506437 -1.93464e-20 7.15126e-24 -1.93393e-20 0.0013958 0.997816 8.59763e-05 0.152643 2.85226 0.0013958 0.997818 0.743127 0.00105756 0.00188053 0.000859763 0.455517 0.00188053 0.440992 0.000129717 1.02 0.88813 0.534555 0.286676 1.71789e-07 3.07095e-09 2380.41 3115.55 -0.0556661 0.482164 0.277438 0.253267 -0.593371 -0.169537 0.495777 -0.267014 -0.228772 2.079 1 0 297.604 0 2.15276 2.077 0.000299674 0.854038 0.674594 0.348564 0.420816 2.15296 134.764 83.9206 18.7209 60.8663 0.0040253 0 -40 10
1.178 3.41095e-08 2.5392e-06 0.12298 0.122979 0.0120343 1.55043e-05 0.00115418 0.153726 0.000658351 0.154379 0.902429 101.729 0.240884 0.781427 4.27093 0.0591158 0.0402918 0.959708 0.0197092 0.00437592 0.0189717 0.00419581 0.00529081 0.00602835 0.211632 0.241134 58.0129 -87.897 126.256 15.9567 145.024 0.000141217 0.267205 192.822 0.310439 0.0673553 0.00409674 0.000561993 0.00138385 0.986975 0.991726 -2.98149e-06 -85.6624 0.093035 31182 304.152 0.983509 0.319146 0.732565 0.73256 9.99958 2.98361e-06 1.19343e-05 0.132 0.982928 0.931749 -0.0132924 4.91348e-06 0.50645 -1.93475e-20 7.15172e-24 -1.93404e-20 0.0013958 0.997816 8.59764e-05 0.152643 2.85226 0.0013958 0.997818 0.743216 0.00105758 0.00188053 0.000859764 0.455517 0.00188053 0.440999 0.00012972 1.02 0.888131 0.534554 0.286677 1.71789e-07 3.07098e-09 2380.39 3115.57 -0.0556688 0.482164 0.277438 0.253268 -0.593371 -0.169537 0.495768 -0.267012 -0.228765 2.08 1 0 297.602 0 2.15291 2.078 0.000299673 0.85405 0.67464 0.348481 0.42084 2.15311 134.772 83.9204 18.7209 60.8662 0.00402531 0 -40 10
1.179 3.41384e-08 2.53921e-06 0.123033 0.123032 0.0120343 1.55175e-05 0.00115418 0.153791 0.000658352 0.154445 0.902507 101.729 0.240875 0.781544 4.27129 0.0591252 0.0402952 0.959705 0.0197088 0.00437623 0.0189713 0.00419607 0.00529118 0.00602873 0.211647 0.241149 58.013 -87.897 126.256 15.9566 145.024 0.000141218 0.267205 192.821 0.310438 0.0673552 0.00409674 0.000561994 0.00138385 0.986975 0.991726 -2.9815e-06 -85.6624 0.0930351 31181.9 304.16 0.983509 0.319146 0.732569 0.732565 9.99958 2.98361e-06 1.19343e-05 0.132003 0.98293 0.931749 -0.0132924 4.91351e-06 0.506463 -1.93486e-20 7.15217e-24 -1.93415e-20 0.0013958 0.997816 8.59765e-05 0.152644 2.85226 0.0013958 0.997818 0.743305 0.00105759 0.00188053 0.000859765 0.455517 0.00188053 0.441005 0.000129723 1.02 0.888132 0.534554 0.286679 1.7179e-07 3.071e-09 2380.38 3115.59 -0.0556715 0.482164 0.277438 0.253269 -0.593371 -0.169537 0.495759 -0.26701 -0.228759 2.081 1 0 297.599 0 2.15305 2.079 0.000299673 0.854062 0.674686 0.348399 0.420864 2.15325 134.78 83.9202 18.7209 60.8661 0.00402532 0 -40 10
1.18 3.41673e-08 2.53921e-06 0.123085 0.123084 0.0120343 1.55306e-05 0.00115418 0.153857 0.000658353 0.15451 0.902585 101.728 0.240865 0.781661 4.27165 0.0591346 0.0402986 0.959701 0.0197084 0.00437654 0.0189709 0.00419633 0.00529156 0.00602911 0.211663 0.241164 58.0131 -87.897 126.256 15.9566 145.024 0.000141219 0.267206 192.821 0.310438 0.0673552 0.00409674 0.000561995 0.00138385 0.986975 0.991726 -2.98152e-06 -85.6624 0.0930352 31181.9 304.168 0.983509 0.319146 0.732574 0.73257 9.99958 2.98362e-06 1.19344e-05 0.132007 0.982932 0.931749 -0.0132924 4.91354e-06 0.506476 -1.93498e-20 7.15263e-24 -1.93426e-20 0.0013958 0.997816 8.59766e-05 0.152644 2.85226 0.0013958 0.997818 0.743395 0.00105761 0.00188054 0.000859766 0.455516 0.00188053 0.441012 0.000129725 1.02 0.888133 0.534554 0.28668 1.7179e-07 3.07102e-09 2380.36 3115.61 -0.0556742 0.482164 0.277438 0.253271 -0.593371 -0.169537 0.49575 -0.267008 -0.228752 2.082 1 0 297.597 0 2.1532 2.08 0.000299672 0.854074 0.674732 0.348317 0.420888 2.1534 134.787 83.92 18.7209 60.866 0.00402533 0 -40 10
1.181 3.41962e-08 2.53921e-06 0.123138 0.123137 0.0120343 1.55437e-05 0.00115419 0.153922 0.000658354 0.154576 0.902663 101.728 0.240856 0.781778 4.27202 0.059144 0.040302 0.959698 0.0197081 0.00437684 0.0189705 0.00419659 0.00529194 0.00602949 0.211678 0.24118 58.0131 -87.897 126.256 15.9566 145.024 0.00014122 0.267206 192.821 0.310437 0.0673551 0.00409675 0.000561995 0.00138385 0.986975 0.991726 -2.98153e-06 -85.6624 0.0930353 31181.9 304.177 0.983509 0.319146 0.732579 0.732574 9.99958 2.98362e-06 1.19344e-05 0.13201 0.982934 0.931749 -0.0132924 4.91357e-06 0.506489 -1.93509e-20 7.15309e-24 -1.93437e-20 0.0013958 0.997816 8.59766e-05 0.152644 2.85226 0.0013958 0.997818 0.743484 0.00105763 0.00188054 0.000859766 0.455516 0.00188054 0.441019 0.000129728 1.02 0.888134 0.534553 0.286682 1.7179e-07 3.07104e-09 2380.34 3115.63 -0.055677 0.482165 0.277437 0.253272 -0.59337 -0.169537 0.495741 -0.267006 -0.228745 2.083 1 0 297.595 0 2.15335 2.081 0.000299671 0.854087 0.674778 0.348235 0.420913 2.15355 134.795 83.9197 18.7208 60.8659 0.00402534 0 -40 10
1.182 3.42251e-08 2.53921e-06 0.12319 0.123189 0.0120343 1.55569e-05 0.00115419 0.153988 0.000658356 0.154641 0.902741 101.728 0.240847 0.781895 4.27238 0.0591534 0.0403055 0.959695 0.0197077 0.00437715 0.0189701 0.00419686 0.00529232 0.00602987 0.211693 0.241195 58.0132 -87.897 126.255 15.9565 145.024 0.000141221 0.267206 192.821 0.310437 0.0673551 0.00409675 0.000561996 0.00138385 0.986975 0.991726 -2.98155e-06 -85.6624 0.0930354 31181.9 304.185 0.983509 0.319146 0.732583 0.732579 9.99958 2.98363e-06 1.19344e-05 0.132013 0.982935 0.931749 -0.0132924 4.9136e-06 0.506503 -1.9352e-20 7.15355e-24 -1.93449e-20 0.0013958 0.997816 8.59767e-05 0.152644 2.85226 0.0013958 0.997818 0.743573 0.00105765 0.00188054 0.000859767 0.455516 0.00188054 0.441026 0.000129731 1.02 0.888135 0.534553 0.286683 1.71791e-07 3.07107e-09 2380.33 3115.65 -0.0556797 0.482165 0.277437 0.253273 -0.59337 -0.169537 0.495732 -0.267003 -0.228738 2.084 1 0 297.592 0 2.15349 2.082 0.00029967 0.854099 0.674823 0.348153 0.420937 2.15369 134.803 83.9195 18.7208 60.8658 0.00402535 0 -40 10
1.183 3.4254e-08 2.53921e-06 0.123242 0.123241 0.0120342 1.557e-05 0.00115419 0.154053 0.000658357 0.154707 0.902819 101.727 0.240837 0.782013 4.27274 0.0591628 0.0403089 0.959691 0.0197073 0.00437746 0.0189697 0.00419712 0.0052927 0.00603026 0.211708 0.24121 58.0132 -87.897 126.255 15.9565 145.024 0.000141222 0.267206 192.821 0.310436 0.067355 0.00409675 0.000561997 0.00138386 0.986975 0.991725 -2.98156e-06 -85.6624 0.0930355 31181.8 304.194 0.983509 0.319146 0.732588 0.732584 9.99958 2.98363e-06 1.19344e-05 0.132016 0.982937 0.931749 -0.0132924 4.91363e-06 0.506516 -1.93531e-20 7.15401e-24 -1.9346e-20 0.0013958 0.997816 8.59768e-05 0.152644 2.85226 0.0013958 0.997818 0.743662 0.00105767 0.00188054 0.000859768 0.455516 0.00188054 0.441033 0.000129734 1.02 0.888136 0.534553 0.286685 1.71791e-07 3.07109e-09 2380.31 3115.67 -0.0556824 0.482165 0.277437 0.253274 -0.59337 -0.169537 0.495723 -0.267001 -0.228731 2.085 1 0 297.59 0 2.15364 2.083 0.00029967 0.854111 0.674869 0.348072 0.420961 2.15384 134.811 83.9193 18.7208 60.8657 0.00402536 0 -40 10
1.184 3.42829e-08 2.53921e-06 0.123295 0.123293 0.0120342 1.55831e-05 0.00115419 0.154118 0.000658358 0.154772 0.902898 101.727 0.240828 0.78213 4.27311 0.0591722 0.0403124 0.959688 0.0197069 0.00437777 0.0189694 0.00419738 0.00529308 0.00603064 0.211723 0.241226 58.0133 -87.897 126.255 15.9564 145.024 0.000141223 0.267206 192.821 0.310436 0.067355 0.00409675 0.000561997 0.00138386 0.986975 0.991725 -2.98158e-06 -85.6624 0.0930356 31181.8 304.202 0.983509 0.319146 0.732593 0.732588 9.99958 2.98364e-06 1.19344e-05 0.132019 0.982939 0.931749 -0.0132924 4.91366e-06 0.506529 -1.93543e-20 7.15447e-24 -1.93471e-20 0.0013958 0.997816 8.59769e-05 0.152644 2.85226 0.0013958 0.997818 0.743751 0.00105768 0.00188054 0.000859769 0.455515 0.00188054 0.44104 0.000129737 1.02 0.888137 0.534552 0.286686 1.71791e-07 3.07111e-09 2380.29 3115.69 -0.0556852 0.482165 0.277436 0.253276 -0.59337 -0.169537 0.495713 -0.266999 -0.228724 2.086 1 0 297.588 0 2.15379 2.084 0.000299669 0.854124 0.674915 0.34799 0.420985 2.15398 134.819 83.919 18.7208 60.8656 0.00402537 0 -40 10
1.185 3.43118e-08 2.53921e-06 0.123347 0.123346 0.0120342 1.55963e-05 0.00115419 0.154184 0.000658359 0.154837 0.902976 101.727 0.240818 0.782248 4.27347 0.0591816 0.0403158 0.959684 0.0197065 0.00437808 0.018969 0.00419764 0.00529346 0.00603103 0.211738 0.241241 58.0134 -87.897 126.255 15.9564 145.024 0.000141224 0.267207 192.82 0.310436 0.0673549 0.00409676 0.000561998 0.00138386 0.986975 0.991725 -2.98159e-06 -85.6624 0.0930357 31181.8 304.21 0.983509 0.319146 0.732598 0.732593 9.99958 2.98364e-06 1.19345e-05 0.132022 0.982941 0.931749 -0.0132924 4.91369e-06 0.506542 -1.93554e-20 7.15493e-24 -1.93482e-20 0.00139581 0.997816 8.5977e-05 0.152644 2.85226 0.00139581 0.997818 0.74384 0.0010577 0.00188054 0.00085977 0.455515 0.00188054 0.441047 0.00012974 1.02 0.888138 0.534552 0.286688 1.71791e-07 3.07114e-09 2380.28 3115.71 -0.0556879 0.482165 0.277436 0.253277 -0.593369 -0.169537 0.495704 -0.266997 -0.228716 2.087 1 0 297.585 0 2.15393 2.085 0.000299668 0.854136 0.674961 0.347909 0.421009 2.15413 134.827 83.9188 18.7208 60.8655 0.00402538 0 -40 10
1.186 3.43407e-08 2.53921e-06 0.123399 0.123398 0.0120342 1.56094e-05 0.00115419 0.154249 0.00065836 0.154903 0.903054 101.726 0.240809 0.782365 4.27384 0.059191 0.0403193 0.959681 0.0197062 0.00437839 0.0189686 0.0041979 0.00529384 0.00603141 0.211754 0.241256 58.0134 -87.897 126.255 15.9564 145.024 0.000141225 0.267207 192.82 0.310435 0.0673549 0.00409676 0.000561999 0.00138386 0.986975 0.991725 -2.98161e-06 -85.6624 0.0930357 31181.8 304.219 0.983509 0.319146 0.732602 0.732598 9.99958 2.98365e-06 1.19345e-05 0.132025 0.982942 0.931749 -0.0132924 4.91372e-06 0.506555 -1.93565e-20 7.15539e-24 -1.93494e-20 0.00139581 0.997816 8.5977e-05 0.152645 2.85227 0.00139581 0.997818 0.743929 0.00105772 0.00188054 0.00085977 0.455515 0.00188054 0.441054 0.000129743 1.02 0.888139 0.534552 0.286689 1.71792e-07 3.07116e-09 2380.26 3115.73 -0.0556907 0.482165 0.277436 0.253278 -0.593369 -0.169537 0.495695 -0.266995 -0.228709 2.088 1 0 297.583 0 2.15408 2.086 0.000299668 0.854149 0.675007 0.347828 0.421033 2.15428 134.835 83.9185 18.7208 60.8653 0.00402539 0 -40 10
1.187 3.43696e-08 2.53921e-06 0.123451 0.12345 0.0120342 1.56226e-05 0.00115419 0.154314 0.000658362 0.154968 0.903132 101.726 0.2408 0.782482 4.27421 0.0592004 0.0403227 0.959677 0.0197058 0.0043787 0.0189682 0.00419817 0.00529422 0.0060318 0.211769 0.241272 58.0135 -87.897 126.255 15.9563 145.024 0.000141225 0.267207 192.82 0.310435 0.0673548 0.00409676 0.000561999 0.00138387 0.986975 0.991725 -2.98162e-06 -85.6624 0.0930358 31181.8 304.227 0.983509 0.319146 0.732607 0.732603 9.99958 2.98365e-06 1.19345e-05 0.132029 0.982944 0.931748 -0.0132924 4.91375e-06 0.506568 -1.93576e-20 7.15585e-24 -1.93505e-20 0.00139581 0.997816 8.59771e-05 0.152645 2.85227 0.00139581 0.997818 0.744018 0.00105774 0.00188055 0.000859771 0.455515 0.00188055 0.441061 0.000129746 1.02 0.88814 0.534552 0.286691 1.71792e-07 3.07118e-09 2380.24 3115.75 -0.0556935 0.482165 0.277436 0.25328 -0.593369 -0.169538 0.495686 -0.266993 -0.228702 2.089 1 0 297.581 0 2.15423 2.087 0.000299667 0.854161 0.675053 0.347747 0.421058 2.15442 134.842 83.9183 18.7208 60.8652 0.0040254 0 -40 10
1.188 3.43985e-08 2.53921e-06 0.123503 0.123502 0.0120342 1.56357e-05 0.00115419 0.154379 0.000658363 0.155033 0.90321 101.725 0.24079 0.7826 4.27457 0.0592098 0.0403262 0.959674 0.0197054 0.00437901 0.0189678 0.00419843 0.0052946 0.00603218 0.211784 0.241287 58.0136 -87.897 126.255 15.9563 145.024 0.000141226 0.267207 192.82 0.310434 0.0673548 0.00409677 0.000562 0.00138387 0.986975 0.991725 -2.98164e-06 -85.6623 0.0930359 31181.7 304.235 0.983509 0.319146 0.732612 0.732608 9.99958 2.98366e-06 1.19345e-05 0.132032 0.982946 0.931748 -0.0132924 4.91378e-06 0.506582 -1.93588e-20 7.15631e-24 -1.93516e-20 0.00139581 0.997816 8.59772e-05 0.152645 2.85227 0.00139581 0.997818 0.744107 0.00105776 0.00188055 0.000859772 0.455515 0.00188055 0.441067 0.000129749 1.02 0.888142 0.534551 0.286692 1.71792e-07 3.0712e-09 2380.23 3115.77 -0.0556963 0.482165 0.277435 0.253281 -0.593368 -0.169538 0.495676 -0.266991 -0.228695 2.09 1 0 297.578 0 2.15437 2.088 0.000299666 0.854174 0.675099 0.347666 0.421082 2.15457 134.85 83.9181 18.7208 60.8651 0.00402541 0 -40 10
1.189 3.44274e-08 2.53921e-06 0.123555 0.123554 0.0120342 1.56488e-05 0.00115419 0.154444 0.000658364 0.155098 0.903289 101.725 0.240781 0.782718 4.27494 0.0592193 0.0403296 0.95967 0.019705 0.00437932 0.0189674 0.00419869 0.00529498 0.00603257 0.211799 0.241303 58.0136 -87.897 126.255 15.9563 145.024 0.000141227 0.267207 192.82 0.310434 0.0673547 0.00409677 0.000562001 0.00138387 0.986975 0.991725 -2.98165e-06 -85.6623 0.093036 31181.7 304.244 0.983509 0.319146 0.732617 0.732613 9.99958 2.98366e-06 1.19345e-05 0.132035 0.982948 0.931748 -0.0132924 4.91381e-06 0.506595 -1.93599e-20 7.15677e-24 -1.93527e-20 0.00139581 0.997816 8.59773e-05 0.152645 2.85227 0.00139581 0.997818 0.744196 0.00105778 0.00188055 0.000859773 0.455514 0.00188055 0.441074 0.000129751 1.02 0.888143 0.534551 0.286694 1.71792e-07 3.07123e-09 2380.21 3115.79 -0.0556991 0.482165 0.277435 0.253282 -0.593368 -0.169538 0.495667 -0.266989 -0.228688 2.091 1 0 297.576 0 2.15452 2.089 0.000299665 0.854187 0.675145 0.347585 0.421106 2.15472 134.858 83.9178 18.7207 60.865 0.00402542 0 -40 10
1.19 3.44563e-08 2.53922e-06 0.123607 0.123606 0.0120341 1.5662e-05 0.00115419 0.154509 0.000658365 0.155163 0.903367 101.725 0.240771 0.782835 4.27531 0.0592287 0.0403331 0.959667 0.0197046 0.00437963 0.018967 0.00419896 0.00529537 0.00603295 0.211815 0.241318 58.0137 -87.897 126.255 15.9562 145.024 0.000141228 0.267207 192.82 0.310433 0.0673547 0.00409677 0.000562001 0.00138387 0.986975 0.991725 -2.98167e-06 -85.6623 0.0930361 31181.7 304.252 0.983509 0.319146 0.732622 0.732618 9.99958 2.98367e-06 1.19346e-05 0.132038 0.98295 0.931748 -0.0132924 4.91384e-06 0.506608 -1.9361e-20 7.15723e-24 -1.93539e-20 0.00139581 0.997816 8.59774e-05 0.152645 2.85227 0.00139581 0.997818 0.744285 0.00105779 0.00188055 0.000859774 0.455514 0.00188055 0.441081 0.000129754 1.02 0.888144 0.534551 0.286695 1.71793e-07 3.07125e-09 2380.19 3115.81 -0.0557019 0.482165 0.277435 0.253284 -0.593368 -0.169538 0.495658 -0.266987 -0.228681 2.092 1 0 297.574 0 2.15466 2.09 0.000299665 0.854199 0.67519 0.347504 0.42113 2.15486 134.866 83.9176 18.7207 60.8649 0.00402543 0 -40 10
1.191 3.44852e-08 2.53922e-06 0.123659 0.123658 0.0120341 1.56751e-05 0.00115419 0.154574 0.000658366 0.155228 0.903445 101.724 0.240762 0.782953 4.27568 0.0592381 0.0403366 0.959663 0.0197043 0.00437994 0.0189667 0.00419922 0.00529575 0.00603334 0.21183 0.241334 58.0137 -87.897 126.255 15.9562 145.024 0.000141229 0.267208 192.819 0.310433 0.0673546 0.00409678 0.000562002 0.00138387 0.986975 0.991725 -2.98168e-06 -85.6623 0.0930362 31181.7 304.261 0.983509 0.319146 0.732627 0.732623 9.99958 2.98367e-06 1.19346e-05 0.132041 0.982951 0.931748 -0.0132924 4.91387e-06 0.506621 -1.93621e-20 7.15769e-24 -1.9355e-20 0.00139581 0.997816 8.59775e-05 0.152645 2.85227 0.00139581 0.997818 0.744374 0.00105781 0.00188055 0.000859775 0.455514 0.00188055 0.441088 0.000129757 1.02 0.888145 0.53455 0.286697 1.71793e-07 3.07127e-09 2380.18 3115.83 -0.0557047 0.482165 0.277434 0.253285 -0.593368 -0.169538 0.495648 -0.266984 -0.228673 2.093 1 0 297.571 0 2.15481 2.091 0.000299664 0.854212 0.675236 0.347424 0.421154 2.15501 134.874 83.9173 18.7207 60.8648 0.00402544 0 -40 10
1.192 3.45141e-08 2.53922e-06 0.123711 0.12371 0.0120341 1.56882e-05 0.00115419 0.154639 0.000658367 0.155293 0.903523 101.724 0.240752 0.783071 4.27605 0.0592475 0.0403401 0.95966 0.0197039 0.00438025 0.0189663 0.00419948 0.00529613 0.00603373 0.211845 0.241349 58.0138 -87.897 126.255 15.9561 145.024 0.00014123 0.267208 192.819 0.310433 0.0673546 0.00409678 0.000562003 0.00138388 0.986975 0.991725 -2.9817e-06 -85.6623 0.0930363 31181.6 304.269 0.983509 0.319146 0.732632 0.732628 9.99958 2.98368e-06 1.19346e-05 0.132044 0.982953 0.931748 -0.0132924 4.9139e-06 0.506634 -1.93633e-20 7.15815e-24 -1.93561e-20 0.00139581 0.997816 8.59775e-05 0.152646 2.85227 0.00139581 0.997818 0.744463 0.00105783 0.00188055 0.000859775 0.455514 0.00188055 0.441095 0.00012976 1.02 0.888146 0.53455 0.286698 1.71793e-07 3.0713e-09 2380.16 3115.85 -0.0557075 0.482165 0.277434 0.253286 -0.593367 -0.169538 0.495639 -0.266982 -0.228666 2.094 1 0 297.569 0 2.15496 2.092 0.000299663 0.854225 0.675282 0.347343 0.421178 2.15516 134.882 83.9171 18.7207 60.8646 0.00402545 0 -40 10
1.193 3.4543e-08 2.53922e-06 0.123763 0.123762 0.0120341 1.57014e-05 0.00115419 0.154704 0.000658369 0.155358 0.903602 101.724 0.240743 0.783188 4.27642 0.059257 0.0403435 0.959656 0.0197035 0.00438056 0.0189659 0.00419975 0.00529652 0.00603411 0.211861 0.241365 58.0139 -87.897 126.255 15.9561 145.024 0.000141231 0.267208 192.819 0.310432 0.0673545 0.00409678 0.000562003 0.00138388 0.986975 0.991725 -2.98171e-06 -85.6623 0.0930364 31181.6 304.278 0.983509 0.319146 0.732637 0.732633 9.99958 2.98368e-06 1.19346e-05 0.132048 0.982955 0.931748 -0.0132924 4.91393e-06 0.506648 -1.93644e-20 7.15862e-24 -1.93572e-20 0.00139581 0.997816 8.59776e-05 0.152646 2.85227 0.00139581 0.997818 0.744552 0.00105785 0.00188056 0.000859776 0.455513 0.00188055 0.441102 0.000129763 1.02 0.888147 0.53455 0.2867 1.71794e-07 3.07132e-09 2380.14 3115.87 -0.0557103 0.482165 0.277434 0.253288 -0.593367 -0.169538 0.49563 -0.26698 -0.228659 2.095 1 0 297.567 0 2.1551 2.093 0.000299663 0.854238 0.675328 0.347263 0.421202 2.1553 134.89 83.9168 18.7207 60.8645 0.00402546 0 -40 10
1.194 3.45719e-08 2.53922e-06 0.123815 0.123814 0.0120341 1.57145e-05 0.00115419 0.154769 0.00065837 0.155423 0.90368 101.723 0.240734 0.783306 4.27678 0.0592664 0.040347 0.959653 0.0197031 0.00438087 0.0189655 0.00420001 0.0052969 0.0060345 0.211876 0.24138 58.0139 -87.897 126.254 15.9561 145.024 0.000141232 0.267208 192.819 0.310432 0.0673545 0.00409678 0.000562004 0.00138388 0.986975 0.991725 -2.98173e-06 -85.6623 0.0930364 31181.6 304.286 0.983509 0.319146 0.732642 0.732638 9.99958 2.98369e-06 1.19346e-05 0.132051 0.982957 0.931748 -0.0132924 4.91396e-06 0.506661 -1.93655e-20 7.15908e-24 -1.93584e-20 0.00139582 0.997816 8.59777e-05 0.152646 2.85227 0.00139582 0.997818 0.74464 0.00105787 0.00188056 0.000859777 0.455513 0.00188056 0.441109 0.000129766 1.02 0.888148 0.534549 0.286701 1.71794e-07 3.07134e-09 2380.13 3115.89 -0.0557132 0.482166 0.277434 0.253289 -0.593367 -0.169538 0.49562 -0.266978 -0.228652 2.096 1 0 297.564 0 2.15525 2.094 0.000299662 0.854251 0.675374 0.347183 0.421227 2.15545 134.897 83.9166 18.7207 60.8644 0.00402547 0 -40 10
1.195 3.46008e-08 2.53922e-06 0.123867 0.123866 0.0120341 1.57276e-05 0.00115419 0.154834 0.000658371 0.155487 0.903759 101.723 0.240724 0.783424 4.27715 0.0592759 0.0403505 0.959649 0.0197027 0.00438118 0.0189651 0.00420028 0.00529728 0.00603489 0.211891 0.241396 58.014 -87.897 126.254 15.956 145.024 0.000141233 0.267208 192.819 0.310431 0.0673544 0.00409679 0.000562005 0.00138388 0.986975 0.991725 -2.98174e-06 -85.6623 0.0930365 31181.6 304.295 0.983509 0.319146 0.732647 0.732643 9.99958 2.98369e-06 1.19347e-05 0.132054 0.982958 0.931747 -0.0132924 4.91399e-06 0.506674 -1.93667e-20 7.15954e-24 -1.93595e-20 0.00139582 0.997816 8.59778e-05 0.152646 2.85227 0.00139582 0.997818 0.744729 0.00105788 0.00188056 0.000859778 0.455513 0.00188056 0.441116 0.000129769 1.02 0.888149 0.534549 0.286703 1.71794e-07 3.07136e-09 2380.11 3115.91 -0.055716 0.482166 0.277433 0.25329 -0.593367 -0.169538 0.495611 -0.266976 -0.228644 2.097 1 0 297.562 0 2.1554 2.095 0.000299661 0.854264 0.675419 0.347103 0.421251 2.15559 134.905 83.9163 18.7207 60.8643 0.00402548 0 -40 10
1.196 3.46297e-08 2.53922e-06 0.123919 0.123917 0.0120341 1.57408e-05 0.00115419 0.154898 0.000658372 0.155552 0.903837 101.722 0.240715 0.783542 4.27752 0.0592853 0.040354 0.959646 0.0197023 0.0043815 0.0189647 0.00420054 0.00529767 0.00603528 0.211907 0.241411 58.0141 -87.8971 126.254 15.956 145.025 0.000141234 0.267209 192.819 0.310431 0.0673543 0.00409679 0.000562005 0.00138388 0.986975 0.991725 -2.98176e-06 -85.6623 0.0930366 31181.6 304.303 0.983509 0.319146 0.732652 0.732648 9.99958 2.9837e-06 1.19347e-05 0.132057 0.98296 0.931747 -0.0132924 4.91401e-06 0.506688 -1.93678e-20 7.16e-24 -1.93606e-20 0.00139582 0.997816 8.59779e-05 0.152646 2.85227 0.00139582 0.997818 0.744818 0.0010579 0.00188056 0.000859779 0.455513 0.00188056 0.441122 0.000129772 1.02 0.88815 0.534549 0.286704 1.71794e-07 3.07139e-09 2380.09 3115.93 -0.0557189 0.482166 0.277433 0.253292 -0.593366 -0.169538 0.495601 -0.266974 -0.228637 2.098 1 0 297.559 0 2.15554 2.096 0.00029966 0.854277 0.675465 0.347023 0.421275 2.15574 134.913 83.9161 18.7206 60.8642 0.00402549 0 -40 10
1.197 3.46586e-08 2.53922e-06 0.12397 0.123969 0.0120341 1.57539e-05 0.00115419 0.154963 0.000658373 0.155617 0.903916 101.722 0.240705 0.78366 4.2779 0.0592948 0.0403575 0.959642 0.0197019 0.00438181 0.0189643 0.00420081 0.00529805 0.00603567 0.211922 0.241427 58.0141 -87.8971 126.254 15.956 145.025 0.000141235 0.267209 192.818 0.31043 0.0673543 0.00409679 0.000562006 0.00138389 0.986975 0.991725 -2.98177e-06 -85.6623 0.0930367 31181.5 304.312 0.983509 0.319146 0.732657 0.732653 9.99958 2.9837e-06 1.19347e-05 0.13206 0.982962 0.931747 -0.0132924 4.91404e-06 0.506701 -1.93689e-20 7.16047e-24 -1.93618e-20 0.00139582 0.997816 8.59779e-05 0.152646 2.85228 0.00139582 0.997818 0.744906 0.00105792 0.00188056 0.000859779 0.455513 0.00188056 0.441129 0.000129775 1.02 0.888151 0.534548 0.286706 1.71795e-07 3.07141e-09 2380.08 3115.95 -0.0557217 0.482166 0.277433 0.253293 -0.593366 -0.169538 0.495592 -0.266972 -0.228629 2.099 1 0 297.557 0 2.15569 2.097 0.00029966 0.85429 0.675511 0.346943 0.421299 2.15589 134.921 83.9158 18.7206 60.864 0.0040255 0 -40 10
1.198 3.46875e-08 2.53922e-06 0.124022 0.124021 0.012034 1.5767e-05 0.00115419 0.155028 0.000658374 0.155681 0.903994 101.722 0.240696 0.783778 4.27827 0.0593042 0.040361 0.959639 0.0197016 0.00438212 0.0189639 0.00420107 0.00529844 0.00603605 0.211937 0.241442 58.0142 -87.8971 126.254 15.9559 145.025 0.000141236 0.267209 192.818 0.31043 0.0673542 0.0040968 0.000562007 0.00138389 0.986975 0.991725 -2.98179e-06 -85.6622 0.0930368 31181.5 304.32 0.983509 0.319146 0.732662 0.732658 9.99958 2.98371e-06 1.19347e-05 0.132064 0.982963 0.931747 -0.0132924 4.91407e-06 0.506714 -1.93701e-20 7.16093e-24 -1.93629e-20 0.00139582 0.997816 8.5978e-05 0.152646 2.85228 0.00139582 0.997818 0.744995 0.00105794 0.00188056 0.00085978 0.455512 0.00188056 0.441136 0.000129777 1.02 0.888153 0.534548 0.286707 1.71795e-07 3.07143e-09 2380.06 3115.97 -0.0557246 0.482166 0.277432 0.253294 -0.593366 -0.169538 0.495582 -0.26697 -0.228622 2.1 1 0 297.554 0 2.15583 2.098 0.000299659 0.854303 0.675557 0.346863 0.421323 2.15603 134.929 83.9156 18.7206 60.8639 0.00402551 0 -40 10
1.199 3.47164e-08 2.53922e-06 0.124074 0.124073 0.012034 1.57802e-05 0.00115419 0.155092 0.000658376 0.155746 0.904073 101.721 0.240686 0.783896 4.27864 0.0593137 0.0403645 0.959635 0.0197012 0.00438244 0.0189636 0.00420134 0.00529882 0.00603644 0.211953 0.241458 58.0143 -87.8971 126.254 15.9559 145.025 0.000141237 0.267209 192.818 0.31043 0.0673542 0.0040968 0.000562007 0.00138389 0.986975 0.991725 -2.9818e-06 -85.6622 0.0930369 31181.5 304.328 0.983509 0.319146 0.732668 0.732663 9.99958 2.98371e-06 1.19347e-05 0.132067 0.982965 0.931747 -0.0132924 4.9141e-06 0.506728 -1.93712e-20 7.1614e-24 -1.93641e-20 0.00139582 0.997816 8.59781e-05 0.152647 2.85228 0.00139582 0.997818 0.745084 0.00105796 0.00188056 0.000859781 0.455512 0.00188056 0.441143 0.00012978 1.02 0.888154 0.534548 0.286709 1.71795e-07 3.07146e-09 2380.04 3116 -0.0557275 0.482166 0.277432 0.253296 -0.593365 -0.169538 0.495573 -0.266968 -0.228615 2.101 1 0 297.552 0 2.15598 2.099 0.000299658 0.854316 0.675603 0.346784 0.421347 2.15618 134.937 83.9153 18.7206 60.8638 0.00402552 0 -40 10
1.2 3.47453e-08 2.53922e-06 0.124125 0.124124 0.012034 1.57933e-05 0.00115419 0.155157 0.000658377 0.15581 0.904151 101.721 0.240677 0.784014 4.27901 0.0593231 0.040368 0.959632 0.0197008 0.00438275 0.0189632 0.0042016 0.00529921 0.00603683 0.211968 0.241473 58.0143 -87.8971 126.254 15.9558 145.025 0.000141238 0.267209 192.818 0.310429 0.0673541 0.0040968 0.000562008 0.00138389 0.986975 0.991725 -2.98182e-06 -85.6622 0.093037 31181.5 304.337 0.983509 0.319146 0.732673 0.732668 9.99958 2.98372e-06 1.19348e-05 0.13207 0.982967 0.931747 -0.0132924 4.91413e-06 0.506741 -1.93723e-20 7.16186e-24 -1.93652e-20 0.00139582 0.997816 8.59782e-05 0.152647 2.85228 0.00139582 0.997818 0.745172 0.00105797 0.00188057 0.000859782 0.455512 0.00188056 0.44115 0.000129783 1.02 0.888155 0.534548 0.286711 1.71795e-07 3.07148e-09 2380.03 3116.02 -0.0557304 0.482166 0.277432 0.253297 -0.593365 -0.169538 0.495563 -0.266965 -0.228607 2.102 1 0 297.55 0 2.15613 2.1 0.000299658 0.85433 0.675648 0.346704 0.421371 2.15632 134.944 83.9151 18.7206 60.8637 0.00402553 0 -40 10
1.201 3.47742e-08 2.53923e-06 0.124177 0.124176 0.012034 1.58064e-05 0.00115419 0.155221 0.000658378 0.155875 0.90423 101.721 0.240667 0.784132 4.27938 0.0593326 0.0403715 0.959628 0.0197004 0.00438306 0.0189628 0.00420187 0.00529959 0.00603722 0.211984 0.241489 58.0144 -87.8971 126.254 15.9558 145.025 0.000141239 0.26721 192.818 0.310429 0.0673541 0.00409681 0.000562009 0.0013839 0.986975 0.991725 -2.98183e-06 -85.6622 0.0930371 31181.4 304.346 0.983509 0.319146 0.732678 0.732674 9.99958 2.98372e-06 1.19348e-05 0.132073 0.982968 0.931747 -0.0132924 4.91416e-06 0.506754 -1.93735e-20 7.16232e-24 -1.93663e-20 0.00139582 0.997816 8.59783e-05 0.152647 2.85228 0.00139582 0.997818 0.745261 0.00105799 0.00188057 0.000859783 0.455512 0.00188057 0.441157 0.000129786 1.02 0.888156 0.534547 0.286712 1.71796e-07 3.0715e-09 2380.01 3116.04 -0.0557333 0.482166 0.277432 0.253299 -0.593365 -0.169538 0.495554 -0.266963 -0.2286 2.103 1 0 297.547 0 2.15627 2.101 0.000299657 0.854343 0.675694 0.346625 0.421395 2.15647 134.952 83.9148 18.7206 60.8635 0.00402554 0 -40 10
1.202 3.48031e-08 2.53923e-06 0.124228 0.124227 0.012034 1.58196e-05 0.00115419 0.155285 0.000658379 0.155939 0.904308 101.72 0.240658 0.78425 4.27976 0.0593421 0.0403751 0.959625 0.0197 0.00438338 0.0189624 0.00420214 0.00529998 0.00603761 0.211999 0.241505 58.0144 -87.8971 126.254 15.9558 145.025 0.00014124 0.26721 192.818 0.310428 0.067354 0.00409681 0.000562009 0.0013839 0.986975 0.991725 -2.98185e-06 -85.6622 0.0930371 31181.4 304.354 0.983509 0.319146 0.732683 0.732679 9.99958 2.98373e-06 1.19348e-05 0.132076 0.98297 0.931746 -0.0132924 4.91419e-06 0.506768 -1.93746e-20 7.16279e-24 -1.93675e-20 0.00139582 0.997816 8.59783e-05 0.152647 2.85228 0.00139582 0.997818 0.745349 0.00105801 0.00188057 0.000859783 0.455511 0.00188057 0.441163 0.000129789 1.02 0.888157 0.534547 0.286714 1.71796e-07 3.07152e-09 2379.99 3116.06 -0.0557362 0.482166 0.277431 0.2533 -0.593364 -0.169538 0.495544 -0.266961 -0.228592 2.104 1 0 297.545 0 2.15642 2.102 0.000299656 0.854356 0.67574 0.346546 0.421419 2.15662 134.96 83.9145 18.7205 60.8634 0.00402555 0 -40 10
1.203 3.4832e-08 2.53923e-06 0.12428 0.124279 0.012034 1.58327e-05 0.00115419 0.15535 0.00065838 0.156004 0.904387 101.72 0.240648 0.784368 4.28013 0.0593515 0.0403786 0.959621 0.0196996 0.00438369 0.018962 0.0042024 0.00530037 0.00603801 0.212015 0.24152 58.0145 -87.8971 126.254 15.9557 145.025 0.000141241 0.26721 192.818 0.310428 0.067354 0.00409681 0.00056201 0.0013839 0.986975 0.991725 -2.98186e-06 -85.6622 0.0930372 31181.4 304.363 0.983509 0.319146 0.732689 0.732684 9.99958 2.98373e-06 1.19348e-05 0.13208 0.982972 0.931746 -0.0132924 4.91422e-06 0.506781 -1.93758e-20 7.16326e-24 -1.93686e-20 0.00139583 0.997816 8.59784e-05 0.152647 2.85228 0.00139583 0.997818 0.745438 0.00105803 0.00188057 0.000859784 0.455511 0.00188057 0.44117 0.000129792 1.02 0.888158 0.534547 0.286715 1.71796e-07 3.07155e-09 2379.98 3116.08 -0.0557391 0.482166 0.277431 0.253301 -0.593364 -0.169539 0.495534 -0.266959 -0.228585 2.105 1 0 297.542 0 2.15657 2.103 0.000299655 0.85437 0.675786 0.346467 0.421444 2.15676 134.968 83.9143 18.7205 60.8633 0.00402556 0 -40 10
1.204 3.48609e-08 2.53923e-06 0.124331 0.12433 0.012034 1.58459e-05 0.00115419 0.155414 0.000658381 0.156068 0.904466 101.719 0.240639 0.784486 4.2805 0.059361 0.0403821 0.959618 0.0196992 0.00438401 0.0189616 0.00420267 0.00530075 0.0060384 0.21203 0.241536 58.0146 -87.8971 126.253 15.9557 145.025 0.000141242 0.26721 192.817 0.310427 0.0673539 0.00409682 0.000562011 0.0013839 0.986975 0.991725 -2.98188e-06 -85.6622 0.0930373 31181.4 304.371 0.983509 0.319146 0.732694 0.732689 9.99958 2.98374e-06 1.19348e-05 0.132083 0.982974 0.931746 -0.0132924 4.91425e-06 0.506794 -1.93769e-20 7.16372e-24 -1.93697e-20 0.00139583 0.997816 8.59785e-05 0.152647 2.85228 0.00139583 0.997818 0.745526 0.00105805 0.00188057 0.000859785 0.455511 0.00188057 0.441177 0.000129795 1.02 0.888159 0.534546 0.286717 1.71796e-07 3.07157e-09 2379.96 3116.1 -0.055742 0.482166 0.277431 0.253303 -0.593364 -0.169539 0.495525 -0.266957 -0.228577 2.106 1 0 297.54 0 2.15671 2.104 0.000299655 0.854383 0.675831 0.346388 0.421468 2.15691 134.976 83.914 18.7205 60.8632 0.00402557 0 -40 10
1.205 3.48898e-08 2.53923e-06 0.124383 0.124382 0.0120339 1.5859e-05 0.00115419 0.155478 0.000658382 0.156132 0.904544 101.719 0.24063 0.784605 4.28088 0.0593705 0.0403856 0.959614 0.0196989 0.00438432 0.0189612 0.00420294 0.00530114 0.00603879 0.212046 0.241552 58.0146 -87.8971 126.253 15.9557 145.025 0.000141243 0.26721 192.817 0.310427 0.0673539 0.00409682 0.000562011 0.0013839 0.986975 0.991725 -2.98189e-06 -85.6622 0.0930374 31181.4 304.38 0.983509 0.319146 0.732699 0.732695 9.99958 2.98374e-06 1.19349e-05 0.132086 0.982975 0.931746 -0.0132924 4.91428e-06 0.506808 -1.9378e-20 7.16419e-24 -1.93709e-20 0.00139583 0.997816 8.59786e-05 0.152648 2.85228 0.00139583 0.997818 0.745615 0.00105806 0.00188057 0.000859786 0.455511 0.00188057 0.441184 0.000129798 1.02 0.88816 0.534546 0.286718 1.71797e-07 3.07159e-09 2379.94 3116.13 -0.0557449 0.482166 0.27743 0.253304 -0.593364 -0.169539 0.495515 -0.266955 -0.228569 2.107 1 0 297.537 0 2.15686 2.105 0.000299654 0.854397 0.675877 0.34631 0.421492 2.15705 134.984 83.9138 18.7205 60.863 0.00402559 0 -40 10
1.206 3.49187e-08 2.53923e-06 0.124434 0.124433 0.0120339 1.58721e-05 0.0011542 0.155543 0.000658384 0.156196 0.904623 101.719 0.24062 0.784723 4.28125 0.05938 0.0403892 0.959611 0.0196985 0.00438464 0.0189608 0.00420321 0.00530153 0.00603918 0.212061 0.241567 58.0147 -87.8971 126.253 15.9556 145.025 0.000141244 0.267211 192.817 0.310427 0.0673538 0.00409682 0.000562012 0.00138391 0.986975 0.991725 -2.98191e-06 -85.6622 0.0930375 31181.3 304.388 0.983509 0.319146 0.732705 0.7327 9.99958 2.98375e-06 1.19349e-05 0.132089 0.982977 0.931746 -0.0132924 4.91431e-06 0.506821 -1.93792e-20 7.16465e-24 -1.9372e-20 0.00139583 0.997816 8.59787e-05 0.152648 2.85228 0.00139583 0.997818 0.745703 0.00105808 0.00188057 0.000859787 0.455511 0.00188057 0.441191 0.0001298 1.02 0.888161 0.534546 0.28672 1.71797e-07 3.07162e-09 2379.93 3116.15 -0.0557479 0.482166 0.27743 0.253306 -0.593363 -0.169539 0.495505 -0.266953 -0.228562 2.108 1 0 297.535 0 2.157 2.106 0.000299653 0.85441 0.675923 0.346231 0.421516 2.1572 134.991 83.9135 18.7205 60.8629 0.0040256 0 -40 10
1.207 3.49476e-08 2.53923e-06 0.124485 0.124484 0.0120339 1.58853e-05 0.0011542 0.155607 0.000658385 0.15626 0.904702 101.718 0.240611 0.784841 4.28163 0.0593895 0.0403927 0.959607 0.0196981 0.00438495 0.0189604 0.00420347 0.00530192 0.00603957 0.212077 0.241583 58.0148 -87.8971 126.253 15.9556 145.025 0.000141245 0.267211 192.817 0.310426 0.0673538 0.00409682 0.000562013 0.00138391 0.986975 0.991725 -2.98192e-06 -85.6622 0.0930376 31181.3 304.397 0.983509 0.319146 0.73271 0.732706 9.99958 2.98375e-06 1.19349e-05 0.132093 0.982979 0.931746 -0.0132924 4.91434e-06 0.506835 -1.93803e-20 7.16512e-24 -1.93732e-20 0.00139583 0.997816 8.59787e-05 0.152648 2.85228 0.00139583 0.997818 0.745792 0.0010581 0.00188058 0.000859787 0.45551 0.00188057 0.441198 0.000129803 1.02 0.888162 0.534545 0.286721 1.71797e-07 3.07164e-09 2379.91 3116.17 -0.0557508 0.482166 0.27743 0.253307 -0.593363 -0.169539 0.495495 -0.266951 -0.228554 2.109 1 0 297.532 0 2.15715 2.107 0.000299652 0.854424 0.675969 0.346153 0.42154 2.15735 134.999 83.9132 18.7205 60.8628 0.00402561 0 -40 10
1.208 3.49765e-08 2.53923e-06 0.124537 0.124535 0.0120339 1.58984e-05 0.0011542 0.155671 0.000658386 0.156325 0.904781 101.718 0.240601 0.78496 4.282 0.0593989 0.0403963 0.959604 0.0196977 0.00438527 0.01896 0.00420374 0.00530231 0.00603997 0.212092 0.241599 58.0148 -87.8971 126.253 15.9555 145.025 0.000141246 0.267211 192.817 0.310426 0.0673537 0.00409683 0.000562013 0.00138391 0.986975 0.991725 -2.98194e-06 -85.6622 0.0930377 31181.3 304.405 0.983509 0.319146 0.732715 0.732711 9.99958 2.98376e-06 1.19349e-05 0.132096 0.98298 0.931745 -0.0132924 4.91437e-06 0.506848 -1.93815e-20 7.16559e-24 -1.93743e-20 0.00139583 0.997816 8.59788e-05 0.152648 2.85229 0.00139583 0.997818 0.74588 0.00105812 0.00188058 0.000859788 0.45551 0.00188058 0.441204 0.000129806 1.02 0.888164 0.534545 0.286723 1.71798e-07 3.07166e-09 2379.89 3116.19 -0.0557538 0.482167 0.27743 0.253309 -0.593363 -0.169539 0.495486 -0.266949 -0.228546 2.11 1 0 297.53 0 2.15729 2.108 0.000299652 0.854438 0.676014 0.346074 0.421564 2.15749 135.007 83.913 18.7205 60.8626 0.00402562 0 -40 10
1.209 3.50054e-08 2.53923e-06 0.124588 0.124587 0.0120339 1.59115e-05 0.0011542 0.155735 0.000658387 0.156389 0.90486 101.718 0.240592 0.785078 4.28238 0.0594084 0.0403998 0.9596 0.0196973 0.00438558 0.0189596 0.00420401 0.00530269 0.00604036 0.212108 0.241614 58.0149 -87.8971 126.253 15.9555 145.025 0.000141247 0.267211 192.817 0.310425 0.0673537 0.00409683 0.000562014 0.00138391 0.986975 0.991725 -2.98195e-06 -85.6621 0.0930378 31181.3 304.414 0.983509 0.319146 0.732721 0.732716 9.99958 2.98376e-06 1.19349e-05 0.132099 0.982982 0.931745 -0.0132924 4.9144e-06 0.506862 -1.93826e-20 7.16605e-24 -1.93755e-20 0.00139583 0.997816 8.59789e-05 0.152648 2.85229 0.00139583 0.997818 0.745968 0.00105814 0.00188058 0.000859789 0.45551 0.00188058 0.441211 0.000129809 1.02 0.888165 0.534545 0.286724 1.71798e-07 3.07168e-09 2379.88 3116.21 -0.0557567 0.482167 0.277429 0.25331 -0.593362 -0.169539 0.495476 -0.266946 -0.228539 2.111 1 0 297.527 0 2.15744 2.109 0.000299651 0.854452 0.67606 0.345996 0.421588 2.15764 135.015 83.9127 18.7204 60.8625 0.00402563 0 -40 10
1.21 3.50343e-08 2.53923e-06 0.124639 0.124638 0.0120339 1.59247e-05 0.0011542 0.155799 0.000658388 0.156453 0.904938 101.717 0.240582 0.785196 4.28276 0.0594179 0.0404034 0.959597 0.0196969 0.0043859 0.0189592 0.00420428 0.00530308 0.00604075 0.212123 0.24163 58.015 -87.8971 126.253 15.9555 145.025 0.000141248 0.267211 192.816 0.310425 0.0673536 0.00409683 0.000562015 0.00138392 0.986974 0.991725 -2.98197e-06 -85.6621 0.0930378 31181.2 304.422 0.983509 0.319146 0.732726 0.732722 9.99958 2.98377e-06 1.1935e-05 0.132102 0.982984 0.931745 -0.0132924 4.91443e-06 0.506875 -1.93838e-20 7.16652e-24 -1.93766e-20 0.00139583 0.997816 8.5979e-05 0.152648 2.85229 0.00139583 0.997818 0.746057 0.00105816 0.00188058 0.00085979 0.45551 0.00188058 0.441218 0.000129812 1.02 0.888166 0.534544 0.286726 1.71798e-07 3.07171e-09 2379.86 3116.24 -0.0557597 0.482167 0.277429 0.253312 -0.593362 -0.169539 0.495466 -0.266944 -0.228531 2.112 1 0 297.525 0 2.15759 2.11 0.00029965 0.854465 0.676106 0.345918 0.421612 2.15778 135.023 83.9124 18.7204 60.8624 0.00402564 0 -40 10
1.211 3.50632e-08 2.53923e-06 0.12469 0.124689 0.0120339 1.59378e-05 0.0011542 0.155863 0.000658389 0.156516 0.905017 101.717 0.240573 0.785315 4.28313 0.0594274 0.0404069 0.959593 0.0196965 0.00438622 0.0189589 0.00420455 0.00530347 0.00604115 0.212139 0.241646 58.015 -87.8971 126.253 15.9554 145.025 0.000141249 0.267211 192.816 0.310424 0.0673536 0.00409684 0.000562015 0.00138392 0.986974 0.991725 -2.98198e-06 -85.6621 0.0930379 31181.2 304.431 0.983509 0.319146 0.732732 0.732727 9.99958 2.98377e-06 1.1935e-05 0.132105 0.982985 0.931745 -0.0132924 4.91446e-06 0.506889 -1.93849e-20 7.16699e-24 -1.93777e-20 0.00139583 0.997816 8.59791e-05 0.152648 2.85229 0.00139583 0.997818 0.746145 0.00105817 0.00188058 0.000859791 0.455509 0.00188058 0.441225 0.000129815 1.02 0.888167 0.534544 0.286727 1.71798e-07 3.07173e-09 2379.84 3116.26 -0.0557627 0.482167 0.277429 0.253313 -0.593362 -0.169539 0.495456 -0.266942 -0.228523 2.113 1 0 297.522 0 2.15773 2.111 0.00029965 0.854479 0.676151 0.34584 0.421636 2.15793 135.03 83.9121 18.7204 60.8623 0.00402565 0 -40 10
1.212 3.5092e-08 2.53924e-06 0.124741 0.12474 0.0120339 1.59509e-05 0.0011542 0.155927 0.00065839 0.15658 0.905096 101.716 0.240563 0.785433 4.28351 0.0594369 0.0404105 0.95959 0.0196961 0.00438653 0.0189585 0.00420482 0.00530386 0.00604154 0.212155 0.241662 58.0151 -87.8971 126.253 15.9554 145.025 0.000141251 0.267212 192.816 0.310424 0.0673535 0.00409684 0.000562016 0.00138392 0.986974 0.991725 -2.982e-06 -85.6621 0.093038 31181.2 304.44 0.983509 0.319146 0.732737 0.732733 9.99958 2.98378e-06 1.1935e-05 0.132109 0.982987 0.931745 -0.0132924 4.91449e-06 0.506902 -1.93861e-20 7.16746e-24 -1.93789e-20 0.00139584 0.997816 8.59791e-05 0.152649 2.85229 0.00139584 0.997818 0.746233 0.00105819 0.00188058 0.000859791 0.455509 0.00188058 0.441232 0.000129818 1.02 0.888168 0.534544 0.286729 1.71799e-07 3.07175e-09 2379.83 3116.28 -0.0557657 0.482167 0.277428 0.253315 -0.593361 -0.169539 0.495446 -0.26694 -0.228516 2.114 1 0 297.519 0 2.15788 2.112 0.000299649 0.854493 0.676197 0.345762 0.42166 2.15808 135.038 83.9119 18.7204 60.8621 0.00402566 0 -40 10
1.213 3.51209e-08 2.53924e-06 0.124792 0.124791 0.0120338 1.59641e-05 0.0011542 0.15599 0.000658392 0.156644 0.905175 101.716 0.240554 0.785552 4.28389 0.0594464 0.0404141 0.959586 0.0196957 0.00438685 0.0189581 0.00420509 0.00530425 0.00604194 0.21217 0.241677 58.0151 -87.8971 126.253 15.9554 145.025 0.000141252 0.267212 192.816 0.310424 0.0673535 0.00409684 0.000562017 0.00138392 0.986974 0.991725 -2.98201e-06 -85.6621 0.0930381 31181.2 304.448 0.983508 0.319146 0.732743 0.732738 9.99958 2.98378e-06 1.1935e-05 0.132112 0.982988 0.931744 -0.0132924 4.91452e-06 0.506916 -1.93872e-20 7.16792e-24 -1.938e-20 0.00139584 0.997816 8.59792e-05 0.152649 2.85229 0.00139584 0.997818 0.746321 0.00105821 0.00188059 0.000859792 0.455509 0.00188058 0.441238 0.000129821 1.02 0.888169 0.534544 0.28673 1.71799e-07 3.07178e-09 2379.81 3116.31 -0.0557687 0.482167 0.277428 0.253316 -0.593361 -0.169539 0.495436 -0.266938 -0.228508 2.115 1 0 297.517 0 2.15802 2.113 0.000299648 0.854507 0.676243 0.345685 0.421684 2.15822 135.046 83.9116 18.7204 60.862 0.00402567 0 -40 10
1.214 3.51498e-08 2.53924e-06 0.124843 0.124842 0.0120338 1.59772e-05 0.0011542 0.156054 0.000658393 0.156708 0.905254 101.716 0.240544 0.785671 4.28427 0.059456 0.0404176 0.959582 0.0196954 0.00438717 0.0189577 0.00420536 0.00530465 0.00604233 0.212186 0.241693 58.0152 -87.8971 126.252 15.9553 145.025 0.000141253 0.267212 192.816 0.310423 0.0673534 0.00409685 0.000562017 0.00138392 0.986974 0.991725 -2.98203e-06 -85.6621 0.0930382 31181.1 304.457 0.983508 0.319146 0.732748 0.732744 9.99958 2.98379e-06 1.1935e-05 0.132115 0.98299 0.931744 -0.0132924 4.91455e-06 0.506929 -1.93884e-20 7.16839e-24 -1.93812e-20 0.00139584 0.997816 8.59793e-05 0.152649 2.85229 0.00139584 0.997818 0.746409 0.00105823 0.00188059 0.000859793 0.455509 0.00188059 0.441245 0.000129823 1.02 0.88817 0.534543 0.286732 1.71799e-07 3.0718e-09 2379.79 3116.33 -0.0557717 0.482167 0.277428 0.253318 -0.593361 -0.169539 0.495426 -0.266936 -0.2285 2.116 1 0 297.514 0 2.15817 2.114 0.000299647 0.854521 0.676288 0.345607 0.421708 2.15837 135.054 83.9113 18.7204 60.8619 0.00402569 0 -40 10
1.215 3.51787e-08 2.53924e-06 0.124894 0.124893 0.0120338 1.59903e-05 0.0011542 0.156118 0.000658394 0.156772 0.905333 101.715 0.240535 0.785789 4.28465 0.0594655 0.0404212 0.959579 0.019695 0.00438749 0.0189573 0.00420563 0.00530504 0.00604273 0.212201 0.241709 58.0153 -87.8971 126.252 15.9553 145.025 0.000141254 0.267212 192.816 0.310423 0.0673533 0.00409685 0.000562018 0.00138393 0.986974 0.991725 -2.98204e-06 -85.6621 0.0930383 31181.1 304.466 0.983508 0.319146 0.732754 0.73275 9.99958 2.98379e-06 1.19351e-05 0.132118 0.982992 0.931744 -0.0132924 4.91458e-06 0.506943 -1.93895e-20 7.16886e-24 -1.93823e-20 0.00139584 0.997816 8.59794e-05 0.152649 2.85229 0.00139584 0.997818 0.746497 0.00105825 0.00188059 0.000859794 0.455508 0.00188059 0.441252 0.000129826 1.02 0.888171 0.534543 0.286733 1.71799e-07 3.07182e-09 2379.78 3116.35 -0.0557747 0.482167 0.277428 0.253319 -0.593361 -0.169539 0.495416 -0.266934 -0.228492 2.117 1 0 297.512 0 2.15832 2.115 0.000299647 0.854535 0.676334 0.34553 0.421732 2.15851 135.062 83.9111 18.7203 60.8617 0.0040257 0 -40 10
1.216 3.52076e-08 2.53924e-06 0.124945 0.124944 0.0120338 1.60035e-05 0.0011542 0.156182 0.000658395 0.156835 0.905412 101.715 0.240525 0.785908 4.28503 0.059475 0.0404248 0.959575 0.0196946 0.0043878 0.0189569 0.0042059 0.00530543 0.00604312 0.212217 0.241725 58.0153 -87.8971 126.252 15.9552 145.025 0.000141255 0.267212 192.815 0.310422 0.0673533 0.00409685 0.000562019 0.00138393 0.986974 0.991725 -2.98206e-06 -85.6621 0.0930384 31181.1 304.474 0.983508 0.319146 0.732759 0.732755 9.99958 2.9838e-06 1.19351e-05 0.132122 0.982993 0.931744 -0.0132924 4.91461e-06 0.506956 -1.93907e-20 7.16933e-24 -1.93835e-20 0.00139584 0.997816 8.59795e-05 0.152649 2.85229 0.00139584 0.997818 0.746586 0.00105826 0.00188059 0.000859795 0.455508 0.00188059 0.441259 0.000129829 1.02 0.888172 0.534543 0.286735 1.718e-07 3.07185e-09 2379.76 3116.37 -0.0557777 0.482167 0.277427 0.253321 -0.59336 -0.169539 0.495406 -0.266932 -0.228484 2.118 1 0 297.509 0 2.15846 2.116 0.000299646 0.854549 0.67638 0.345452 0.421756 2.15866 135.07 83.9108 18.7203 60.8616 0.00402571 0 -40 10
1.217 3.52365e-08 2.53924e-06 0.124996 0.124995 0.0120338 1.60166e-05 0.0011542 0.156245 0.000658396 0.156899 0.905491 101.715 0.240515 0.786027 4.28541 0.0594845 0.0404284 0.959572 0.0196942 0.00438812 0.0189565 0.00420617 0.00530582 0.00604352 0.212233 0.241741 58.0154 -87.8971 126.252 15.9552 145.025 0.000141256 0.267213 192.815 0.310422 0.0673532 0.00409685 0.000562019 0.00138393 0.986974 0.991725 -2.98207e-06 -85.6621 0.0930384 31181.1 304.483 0.983508 0.319146 0.732765 0.732761 9.99958 2.9838e-06 1.19351e-05 0.132125 0.982995 0.931744 -0.0132924 4.91464e-06 0.50697 -1.93918e-20 7.1698e-24 -1.93846e-20 0.00139584 0.997816 8.59795e-05 0.152649 2.85229 0.00139584 0.997818 0.746674 0.00105828 0.00188059 0.000859795 0.455508 0.00188059 0.441266 0.000129832 1.02 0.888173 0.534542 0.286736 1.718e-07 3.07187e-09 2379.74 3116.4 -0.0557807 0.482167 0.277427 0.253322 -0.59336 -0.169539 0.495396 -0.26693 -0.228476 2.119 1 0 297.507 0 2.15861 2.117 0.000299645 0.854564 0.676425 0.345375 0.42178 2.1588 135.077 83.9105 18.7203 60.8615 0.00402572 0 -40 10
1.218 3.52654e-08 2.53924e-06 0.125047 0.125046 0.0120338 1.60297e-05 0.0011542 0.156309 0.000658397 0.156963 0.90557 101.714 0.240506 0.786145 4.28579 0.059494 0.040432 0.959568 0.0196938 0.00438844 0.0189561 0.00420644 0.00530621 0.00604392 0.212248 0.241757 58.0155 -87.8971 126.252 15.9552 145.025 0.000141257 0.267213 192.815 0.310421 0.0673532 0.00409686 0.00056202 0.00138393 0.986974 0.991725 -2.98209e-06 -85.6621 0.0930385 31181.1 304.491 0.983508 0.319146 0.732771 0.732766 9.99958 2.98381e-06 1.19351e-05 0.132128 0.982997 0.931743 -0.0132924 4.91467e-06 0.506983 -1.9393e-20 7.17027e-24 -1.93858e-20 0.00139584 0.997816 8.59796e-05 0.15265 2.85229 0.00139584 0.997818 0.746762 0.0010583 0.00188059 0.000859796 0.455508 0.00188059 0.441272 0.000129835 1.02 0.888175 0.534542 0.286738 1.718e-07 3.07189e-09 2379.73 3116.42 -0.0557837 0.482167 0.277427 0.253324 -0.59336 -0.169539 0.495386 -0.266927 -0.228468 2.12 1 0 297.504 0 2.15875 2.118 0.000299644 0.854578 0.676471 0.345298 0.421804 2.15895 135.085 83.9102 18.7203 60.8613 0.00402573 0 -40 10
1.219 3.52943e-08 2.53924e-06 0.125098 0.125097 0.0120338 1.60429e-05 0.0011542 0.156372 0.000658398 0.157026 0.905649 101.714 0.240496 0.786264 4.28617 0.0595035 0.0404355 0.959564 0.0196934 0.00438876 0.0189557 0.00420671 0.0053066 0.00604431 0.212264 0.241773 58.0155 -87.8971 126.252 15.9551 145.025 0.000141258 0.267213 192.815 0.310421 0.0673531 0.00409686 0.000562021 0.00138393 0.986974 0.991725 -2.9821e-06 -85.6621 0.0930386 31181 304.5 0.983508 0.319146 0.732776 0.732772 9.99958 2.98381e-06 1.19351e-05 0.132131 0.982998 0.931743 -0.0132924 4.9147e-06 0.506997 -1.93941e-20 7.17074e-24 -1.93869e-20 0.00139584 0.997816 8.59797e-05 0.15265 2.8523 0.00139584 0.997818 0.74685 0.00105832 0.00188059 0.000859797 0.455508 0.00188059 0.441279 0.000129838 1.02 0.888176 0.534542 0.286739 1.71801e-07 3.07191e-09 2379.71 3116.44 -0.0557868 0.482167 0.277426 0.253325 -0.593359 -0.16954 0.495376 -0.266925 -0.22846 2.121 1 0 297.501 0 2.1589 2.119 0.000299644 0.854592 0.676516 0.345221 0.421828 2.1591 135.093 83.9099 18.7203 60.8612 0.00402574 0 -40 10
1.22 3.53232e-08 2.53924e-06 0.125149 0.125148 0.0120337 1.6056e-05 0.0011542 0.156436 0.000658399 0.15709 0.905728 101.713 0.240487 0.786383 4.28655 0.0595131 0.0404391 0.959561 0.019693 0.00438908 0.0189553 0.00420698 0.005307 0.00604471 0.21228 0.241788 58.0156 -87.8971 126.252 15.9551 145.025 0.000141259 0.267213 192.815 0.310421 0.0673531 0.00409686 0.000562021 0.00138394 0.986974 0.991725 -2.98212e-06 -85.662 0.0930387 31181 304.509 0.983508 0.319146 0.732782 0.732778 9.99958 2.98382e-06 1.19352e-05 0.132135 0.983 0.931743 -0.0132924 4.91473e-06 0.507011 -1.93953e-20 7.17121e-24 -1.93881e-20 0.00139585 0.997816 8.59798e-05 0.15265 2.8523 0.00139585 0.997817 0.746938 0.00105834 0.0018806 0.000859798 0.455507 0.00188059 0.441286 0.000129841 1.02 0.888177 0.534541 0.286741 1.71801e-07 3.07194e-09 2379.69 3116.47 -0.0557898 0.482167 0.277426 0.253327 -0.593359 -0.16954 0.495366 -0.266923 -0.228453 2.122 1 0 297.499 0 2.15904 2.12 0.000299643 0.854607 0.676562 0.345144 0.421852 2.15924 135.101 83.9097 18.7203 60.8611 0.00402575 0 -40 10
1.221 3.53521e-08 2.53924e-06 0.125199 0.125198 0.0120337 1.60691e-05 0.0011542 0.156499 0.000658401 0.157153 0.905808 101.713 0.240477 0.786502 4.28693 0.0595226 0.0404427 0.959557 0.0196926 0.0043894 0.0189549 0.00420725 0.00530739 0.00604511 0.212296 0.241804 58.0157 -87.8971 126.252 15.955 145.025 0.00014126 0.267213 192.815 0.31042 0.067353 0.00409687 0.000562022 0.00138394 0.986974 0.991725 -2.98213e-06 -85.662 0.0930388 31181 304.517 0.983508 0.319146 0.732788 0.732784 9.99958 2.98382e-06 1.19352e-05 0.132138 0.983001 0.931743 -0.0132924 4.91476e-06 0.507024 -1.93964e-20 7.17168e-24 -1.93892e-20 0.00139585 0.997816 8.59799e-05 0.15265 2.8523 0.00139585 0.997817 0.747026 0.00105835 0.0018806 0.000859799 0.455507 0.0018806 0.441293 0.000129843 1.02 0.888178 0.534541 0.286742 1.71801e-07 3.07196e-09 2379.68 3116.49 -0.0557929 0.482168 0.277426 0.253328 -0.593359 -0.16954 0.495356 -0.266921 -0.228445 2.123 1 0 297.496 0 2.15919 2.121 0.000299642 0.854621 0.676608 0.345068 0.421876 2.15939 135.109 83.9094 18.7202 60.8609 0.00402577 0 -40 10
1.222 3.5381e-08 2.53924e-06 0.12525 0.125249 0.0120337 1.60823e-05 0.0011542 0.156563 0.000658402 0.157216 0.905887 101.713 0.240468 0.786621 4.28731 0.0595321 0.0404463 0.959554 0.0196922 0.00438972 0.0189545 0.00420752 0.00530778 0.00604551 0.212311 0.24182 58.0157 -87.8972 126.252 15.955 145.025 0.000141261 0.267214 192.814 0.31042 0.067353 0.00409687 0.000562023 0.00138394 0.986974 0.991725 -2.98215e-06 -85.662 0.0930389 31181 304.526 0.983508 0.319146 0.732794 0.732789 9.99958 2.98383e-06 1.19352e-05 0.132141 0.983003 0.931742 -0.0132924 4.91479e-06 0.507038 -1.93976e-20 7.17215e-24 -1.93904e-20 0.00139585 0.997816 8.598e-05 0.15265 2.8523 0.00139585 0.997817 0.747114 0.00105837 0.0018806 0.0008598 0.455507 0.0018806 0.441299 0.000129846 1.02 0.888179 0.534541 0.286744 1.71801e-07 3.07198e-09 2379.66 3116.52 -0.055796 0.482168 0.277426 0.25333 -0.593358 -0.16954 0.495346 -0.266919 -0.228437 2.124 1 0 297.493 0 2.15934 2.122 0.000299641 0.854635 0.676653 0.344991 0.4219 2.15953 135.116 83.9091 18.7202 60.8608 0.00402578 0 -40 10
1.223 3.54099e-08 2.53925e-06 0.125301 0.1253 0.0120337 1.60954e-05 0.0011542 0.156626 0.000658403 0.15728 0.905966 101.712 0.240458 0.78674 4.2877 0.0595417 0.04045 0.95955 0.0196918 0.00439004 0.0189541 0.00420779 0.00530818 0.00604591 0.212327 0.241836 58.0158 -87.8972 126.252 15.955 145.025 0.000141263 0.267214 192.814 0.310419 0.0673529 0.00409687 0.000562023 0.00138394 0.986974 0.991725 -2.98216e-06 -85.662 0.093039 31180.9 304.535 0.983508 0.319146 0.732799 0.732795 9.99958 2.98383e-06 1.19352e-05 0.132144 0.983004 0.931742 -0.0132924 4.91482e-06 0.507052 -1.93987e-20 7.17262e-24 -1.93916e-20 0.00139585 0.997816 8.598e-05 0.15265 2.8523 0.00139585 0.997817 0.747201 0.00105839 0.0018806 0.0008598 0.455507 0.0018806 0.441306 0.000129849 1.02 0.88818 0.53454 0.286745 1.71802e-07 3.07201e-09 2379.64 3116.54 -0.055799 0.482168 0.277425 0.253331 -0.593358 -0.16954 0.495336 -0.266917 -0.228429 2.125 1 0 297.491 0 2.15948 2.123 0.000299641 0.85465 0.676699 0.344915 0.421924 2.15968 135.124 83.9088 18.7202 60.8606 0.00402579 0 -40 10
1.224 3.54388e-08 2.53925e-06 0.125351 0.12535 0.0120337 1.61085e-05 0.0011542 0.156689 0.000658404 0.157343 0.906045 101.712 0.240449 0.786859 4.28808 0.0595512 0.0404536 0.959546 0.0196914 0.00439036 0.0189537 0.00420807 0.00530857 0.00604631 0.212343 0.241852 58.0158 -87.8972 126.251 15.9549 145.025 0.000141264 0.267214 192.814 0.310419 0.0673529 0.00409688 0.000562024 0.00138395 0.986974 0.991725 -2.98218e-06 -85.662 0.0930391 31180.9 304.544 0.983508 0.319146 0.732805 0.732801 9.99958 2.98384e-06 1.19352e-05 0.132148 0.983006 0.931742 -0.0132924 4.91485e-06 0.507065 -1.93999e-20 7.1731e-24 -1.93927e-20 0.00139585 0.997816 8.59801e-05 0.15265 2.8523 0.00139585 0.997817 0.747289 0.00105841 0.0018806 0.000859801 0.455506 0.0018806 0.441313 0.000129852 1.02 0.888181 0.53454 0.286747 1.71802e-07 3.07203e-09 2379.63 3116.56 -0.0558021 0.482168 0.277425 0.253333 -0.593358 -0.16954 0.495326 -0.266915 -0.22842 2.126 1 0 297.488 0 2.15963 2.124 0.00029964 0.854664 0.676744 0.344838 0.421948 2.15982 135.132 83.9085 18.7202 60.8605 0.0040258 0 -40 10
1.225 3.54677e-08 2.53925e-06 0.125402 0.125401 0.0120337 1.61217e-05 0.0011542 0.156752 0.000658405 0.157406 0.906124 101.712 0.240439 0.786978 4.28846 0.0595608 0.0404572 0.959543 0.019691 0.00439068 0.0189533 0.00420834 0.00530897 0.0060467 0.212359 0.241868 58.0159 -87.8972 126.251 15.9549 145.025 0.000141265 0.267214 192.814 0.310418 0.0673528 0.00409688 0.000562025 0.00138395 0.986974 0.991725 -2.98219e-06 -85.662 0.0930391 31180.9 304.552 0.983508 0.319146 0.732811 0.732807 9.99958 2.98384e-06 1.19353e-05 0.132151 0.983008 0.931742 -0.0132924 4.91488e-06 0.507079 -1.9401e-20 7.17357e-24 -1.93939e-20 0.00139585 0.997816 8.59802e-05 0.152651 2.8523 0.00139585 0.997817 0.747377 0.00105843 0.0018806 0.000859802 0.455506 0.0018806 0.44132 0.000129855 1.02 0.888182 0.53454 0.286749 1.71802e-07 3.07205e-09 2379.61 3116.59 -0.0558052 0.482168 0.277425 0.253335 -0.593357 -0.16954 0.495316 -0.266913 -0.228412 2.127 1 0 297.485 0 2.15977 2.125 0.000299639 0.854679 0.67679 0.344762 0.421972 2.15997 135.14 83.9082 18.7202 60.8604 0.00402581 0 -40 10
1.226 3.54966e-08 2.53925e-06 0.125452 0.125451 0.0120337 1.61348e-05 0.0011542 0.156816 0.000658406 0.157469 0.906204 101.711 0.24043 0.787097 4.28885 0.0595703 0.0404608 0.959539 0.0196906 0.004391 0.0189529 0.00420861 0.00530936 0.0060471 0.212375 0.241884 58.016 -87.8972 126.251 15.9549 145.025 0.000141266 0.267214 192.814 0.310418 0.0673528 0.00409688 0.000562025 0.00138395 0.986974 0.991725 -2.98221e-06 -85.662 0.0930392 31180.9 304.561 0.983508 0.319146 0.732817 0.732813 9.99958 2.98385e-06 1.19353e-05 0.132154 0.983009 0.931742 -0.0132924 4.9149e-06 0.507093 -1.94022e-20 7.17404e-24 -1.9395e-20 0.00139585 0.997816 8.59803e-05 0.152651 2.8523 0.00139585 0.997817 0.747465 0.00105844 0.0018806 0.000859803 0.455506 0.0018806 0.441326 0.000129858 1.02 0.888183 0.53454 0.28675 1.71802e-07 3.07207e-09 2379.59 3116.61 -0.0558083 0.482168 0.277424 0.253336 -0.593357 -0.16954 0.495305 -0.266911 -0.228404 2.128 1 0 297.483 0 2.15992 2.126 0.000299639 0.854694 0.676836 0.344686 0.421996 2.16011 135.148 83.9079 18.7202 60.8602 0.00402583 0 -40 10
1.227 3.55255e-08 2.53925e-06 0.125503 0.125502 0.0120336 1.61479e-05 0.0011542 0.156879 0.000658407 0.157532 0.906283 101.711 0.24042 0.787216 4.28923 0.0595799 0.0404644 0.959536 0.0196902 0.00439132 0.0189525 0.00420888 0.00530976 0.0060475 0.21239 0.2419 58.016 -87.8972 126.251 15.9548 145.025 0.000141267 0.267215 192.814 0.310418 0.0673527 0.00409689 0.000562026 0.00138395 0.986974 0.991725 -2.98222e-06 -85.662 0.0930393 31180.9 304.57 0.983508 0.319146 0.732823 0.732818 9.99958 2.98385e-06 1.19353e-05 0.132158 0.983011 0.931741 -0.0132924 4.91493e-06 0.507106 -1.94034e-20 7.17451e-24 -1.93962e-20 0.00139585 0.997816 8.59804e-05 0.152651 2.8523 0.00139585 0.997817 0.747553 0.00105846 0.00188061 0.000859804 0.455506 0.0018806 0.441333 0.000129861 1.02 0.888184 0.534539 0.286752 1.71803e-07 3.0721e-09 2379.58 3116.64 -0.0558114 0.482168 0.277424 0.253338 -0.593357 -0.16954 0.495295 -0.266908 -0.228396 2.129 1 0 297.48 0 2.16006 2.127 0.000299638 0.854708 0.676881 0.34461 0.42202 2.16026 135.155 83.9076 18.7201 60.8601 0.00402584 0 -40 10
1.228 3.55544e-08 2.53925e-06 0.125553 0.125552 0.0120336 1.61611e-05 0.0011542 0.156942 0.000658408 0.157596 0.906362 101.71 0.240411 0.787335 4.28961 0.0595894 0.0404681 0.959532 0.0196898 0.00439165 0.0189521 0.00420916 0.00531015 0.00604791 0.212406 0.241916 58.0161 -87.8972 126.251 15.9548 145.025 0.000141268 0.267215 192.813 0.310417 0.0673527 0.00409689 0.000562027 0.00138395 0.986974 0.991725 -2.98224e-06 -85.662 0.0930394 31180.8 304.578 0.983508 0.319146 0.732829 0.732824 9.99958 2.98386e-06 1.19353e-05 0.132161 0.983012 0.931741 -0.0132924 4.91496e-06 0.50712 -1.94045e-20 7.17499e-24 -1.93973e-20 0.00139585 0.997816 8.59804e-05 0.152651 2.8523 0.00139585 0.997817 0.74764 0.00105848 0.00188061 0.000859804 0.455506 0.00188061 0.44134 0.000129863 1.02 0.888186 0.534539 0.286753 1.71803e-07 3.07212e-09 2379.56 3116.66 -0.0558145 0.482168 0.277424 0.253339 -0.593356 -0.16954 0.495285 -0.266906 -0.228388 2.13 1 0 297.477 0 2.16021 2.128 0.000299637 0.854723 0.676927 0.344534 0.422044 2.1604 135.163 83.9073 18.7201 60.8599 0.00402585 0 -40 10
1.229 3.55833e-08 2.53925e-06 0.125604 0.125603 0.0120336 1.61742e-05 0.00115421 0.157005 0.000658409 0.157659 0.906442 101.71 0.240401 0.787454 4.29 0.059599 0.0404717 0.959528 0.0196894 0.00439197 0.0189517 0.00420943 0.00531055 0.00604831 0.212422 0.241932 58.0162 -87.8972 126.251 15.9547 145.025 0.000141269 0.267215 192.813 0.310417 0.0673526 0.00409689 0.000562027 0.00138396 0.986974 0.991725 -2.98225e-06 -85.662 0.0930395 31180.8 304.587 0.983508 0.319146 0.732835 0.73283 9.99958 2.98386e-06 1.19353e-05 0.132164 0.983014 0.931741 -0.0132924 4.91499e-06 0.507134 -1.94057e-20 7.17546e-24 -1.93985e-20 0.00139586 0.997816 8.59805e-05 0.152651 2.8523 0.00139586 0.997817 0.747728 0.0010585 0.00188061 0.000859805 0.455505 0.00188061 0.441347 0.000129866 1.02 0.888187 0.534539 0.286755 1.71803e-07 3.07214e-09 2379.54 3116.68 -0.0558177 0.482168 0.277424 0.253341 -0.593356 -0.16954 0.495275 -0.266904 -0.22838 2.131 1 0 297.475 0 2.16035 2.129 0.000299636 0.854738 0.676972 0.344459 0.422068 2.16055 135.171 83.9071 18.7201 60.8598 0.00402586 0 -40 10
1.23 3.56122e-08 2.53925e-06 0.125654 0.125653 0.0120336 1.61873e-05 0.00115421 0.157068 0.000658411 0.157722 0.906521 101.71 0.240391 0.787574 4.29039 0.0596086 0.0404753 0.959525 0.0196891 0.00439229 0.0189513 0.0042097 0.00531095 0.00604871 0.212438 0.241948 58.0162 -87.8972 126.251 15.9547 145.025 0.00014127 0.267215 192.813 0.310416 0.0673526 0.00409689 0.000562028 0.00138396 0.986974 0.991725 -2.98227e-06 -85.6619 0.0930396 31180.8 304.596 0.983508 0.319146 0.732841 0.732836 9.99958 2.98387e-06 1.19354e-05 0.132167 0.983015 0.931741 -0.0132924 4.91502e-06 0.507148 -1.94068e-20 7.17593e-24 -1.93997e-20 0.00139586 0.997816 8.59806e-05 0.152651 2.85231 0.00139586 0.997817 0.747816 0.00105852 0.00188061 0.000859806 0.455505 0.00188061 0.441353 0.000129869 1.02 0.888188 0.534538 0.286756 1.71803e-07 3.07217e-09 2379.53 3116.71 -0.0558208 0.482168 0.277423 0.253342 -0.593356 -0.16954 0.495264 -0.266902 -0.228372 2.132 1 0 297.472 0 2.1605 2.13 0.000299636 0.854753 0.677018 0.344383 0.422092 2.1607 135.179 83.9068 18.7201 60.8597 0.00402587 0 -40 10
1.231 3.5641e-08 2.53925e-06 0.125705 0.125703 0.0120336 1.62005e-05 0.00115421 0.157131 0.000658412 0.157784 0.906601 101.709 0.240382 0.787693 4.29077 0.0596181 0.040479 0.959521 0.0196887 0.00439261 0.0189509 0.00420998 0.00531134 0.00604911 0.212454 0.241964 58.0163 -87.8972 126.251 15.9547 145.025 0.000141272 0.267215 192.813 0.310416 0.0673525 0.0040969 0.000562029 0.00138396 0.986974 0.991725 -2.98228e-06 -85.6619 0.0930397 31180.8 304.605 0.983508 0.319146 0.732847 0.732842 9.99958 2.98387e-06 1.19354e-05 0.132171 0.983017 0.93174 -0.0132924 4.91505e-06 0.507161 -1.9408e-20 7.17641e-24 -1.94008e-20 0.00139586 0.997816 8.59807e-05 0.152652 2.85231 0.00139586 0.997817 0.747903 0.00105853 0.00188061 0.000859807 0.455505 0.00188061 0.44136 0.000129872 1.02 0.888189 0.534538 0.286758 1.71804e-07 3.07219e-09 2379.51 3116.73 -0.0558239 0.482168 0.277423 0.253344 -0.593355 -0.16954 0.495254 -0.2669 -0.228363 2.133 1 0 297.469 0 2.16064 2.131 0.000299635 0.854768 0.677063 0.344308 0.422116 2.16084 135.187 83.9065 18.7201 60.8595 0.00402589 0 -40 10
1.232 3.56699e-08 2.53925e-06 0.125755 0.125754 0.0120336 1.62136e-05 0.00115421 0.157194 0.000658413 0.157847 0.90668 101.709 0.240372 0.787812 4.29116 0.0596277 0.0404826 0.959517 0.0196883 0.00439294 0.0189505 0.00421025 0.00531174 0.00604951 0.21247 0.24198 58.0163 -87.8972 126.251 15.9546 145.025 0.000141273 0.267215 192.813 0.310415 0.0673525 0.0040969 0.000562029 0.00138396 0.986974 0.991725 -2.9823e-06 -85.6619 0.0930398 31180.7 304.613 0.983508 0.319146 0.732853 0.732848 9.99958 2.98388e-06 1.19354e-05 0.132174 0.983018 0.93174 -0.0132924 4.91508e-06 0.507175 -1.94092e-20 7.17688e-24 -1.9402e-20 0.00139586 0.997816 8.59808e-05 0.152652 2.85231 0.00139586 0.997817 0.747991 0.00105855 0.00188061 0.000859808 0.455505 0.00188061 0.441367 0.000129875 1.02 0.88819 0.534538 0.286759 1.71804e-07 3.07221e-09 2379.5 3116.76 -0.0558271 0.482168 0.277423 0.253346 -0.593355 -0.16954 0.495244 -0.266898 -0.228355 2.134 1 0 297.467 0 2.16079 2.132 0.000299634 0.854783 0.677109 0.344232 0.42214 2.16099 135.194 83.9062 18.7201 60.8594 0.0040259 0 -40 10
1.233 3.56988e-08 2.53925e-06 0.125805 0.125804 0.0120336 1.62267e-05 0.00115421 0.157256 0.000658414 0.15791 0.90676 101.708 0.240363 0.787932 4.29155 0.0596373 0.0404863 0.959514 0.0196879 0.00439326 0.0189501 0.00421053 0.00531214 0.00604991 0.212486 0.241997 58.0164 -87.8972 126.25 15.9546 145.025 0.000141274 0.267216 192.813 0.310415 0.0673524 0.0040969 0.00056203 0.00138397 0.986974 0.991725 -2.98231e-06 -85.6619 0.0930398 31180.7 304.622 0.983508 0.319146 0.732859 0.732854 9.99958 2.98388e-06 1.19354e-05 0.132177 0.98302 0.93174 -0.0132924 4.91511e-06 0.507189 -1.94103e-20 7.17736e-24 -1.94031e-20 0.00139586 0.997816 8.59808e-05 0.152652 2.85231 0.00139586 0.997817 0.748078 0.00105857 0.00188061 0.000859808 0.455504 0.00188061 0.441374 0.000129878 1.02 0.888191 0.534537 0.286761 1.71804e-07 3.07223e-09 2379.48 3116.78 -0.0558302 0.482168 0.277422 0.253347 -0.593355 -0.16954 0.495233 -0.266896 -0.228347 2.135 1 0 297.464 0 2.16093 2.133 0.000299633 0.854798 0.677154 0.344157 0.422164 2.16113 135.202 83.9059 18.72 60.8592 0.00402591 0 -40 10
1.234 3.57277e-08 2.53926e-06 0.125855 0.125854 0.0120336 1.62399e-05 0.00115421 0.157319 0.000658415 0.157973 0.906839 101.708 0.240353 0.788051 4.29193 0.0596468 0.0404899 0.95951 0.0196875 0.00439358 0.0189497 0.0042108 0.00531254 0.00605032 0.212501 0.242013 58.0165 -87.8972 126.25 15.9546 145.025 0.000141275 0.267216 192.812 0.310415 0.0673523 0.00409691 0.000562031 0.00138397 0.986974 0.991725 -2.98233e-06 -85.6619 0.0930399 31180.7 304.631 0.983508 0.319146 0.732865 0.73286 9.99958 2.98389e-06 1.19354e-05 0.132181 0.983022 0.93174 -0.0132924 4.91514e-06 0.507203 -1.94115e-20 7.17783e-24 -1.94043e-20 0.00139586 0.997816 8.59809e-05 0.152652 2.85231 0.00139586 0.997817 0.748166 0.00105859 0.00188062 0.000859809 0.455504 0.00188062 0.44138 0.00012988 1.02 0.888192 0.534537 0.286762 1.71805e-07 3.07226e-09 2379.46 3116.81 -0.0558334 0.482169 0.277422 0.253349 -0.593354 -0.16954 0.495223 -0.266894 -0.228339 2.136 1 0 297.461 0 2.16108 2.134 0.000299633 0.854813 0.6772 0.344082 0.422188 2.16128 135.21 83.9056 18.72 60.8591 0.00402592 0 -40 10
1.235 3.57566e-08 2.53926e-06 0.125905 0.125904 0.0120335 1.6253e-05 0.00115421 0.157382 0.000658416 0.158036 0.906919 101.708 0.240344 0.78817 4.29232 0.0596564 0.0404936 0.959506 0.0196871 0.00439391 0.0189493 0.00421108 0.00531294 0.00605072 0.212517 0.242029 58.0165 -87.8972 126.25 15.9545 145.025 0.000141276 0.267216 192.812 0.310414 0.0673523 0.00409691 0.000562031 0.00138397 0.986974 0.991725 -2.98234e-06 -85.6619 0.09304 31180.7 304.64 0.983508 0.319146 0.732871 0.732866 9.99958 2.98389e-06 1.19355e-05 0.132184 0.983023 0.931739 -0.0132923 4.91517e-06 0.507216 -1.94127e-20 7.17831e-24 -1.94055e-20 0.00139586 0.997816 8.5981e-05 0.152652 2.85231 0.00139586 0.997817 0.748254 0.00105861 0.00188062 0.00085981 0.455504 0.00188062 0.441387 0.000129883 1.02 0.888193 0.534537 0.286764 1.71805e-07 3.07228e-09 2379.45 3116.83 -0.0558365 0.482169 0.277422 0.253351 -0.593354 -0.169541 0.495213 -0.266892 -0.22833 2.137 1 0 297.458 0 2.16123 2.135 0.000299632 0.854828 0.677245 0.344007 0.422212 2.16142 135.218 83.9053 18.72 60.8589 0.00402594 0 -40 10
1.236 3.57855e-08 2.53926e-06 0.125956 0.125954 0.0120335 1.62661e-05 0.00115421 0.157444 0.000658417 0.158098 0.906998 101.707 0.240334 0.78829 4.29271 0.059666 0.0404973 0.959503 0.0196867 0.00439423 0.0189489 0.00421135 0.00531333 0.00605112 0.212533 0.242045 58.0166 -87.8972 126.25 15.9545 145.025 0.000141277 0.267216 192.812 0.310414 0.0673522 0.00409691 0.000562032 0.00138397 0.986974 0.991725 -2.98236e-06 -85.6619 0.0930401 31180.7 304.648 0.983508 0.319146 0.732877 0.732872 9.99958 2.9839e-06 1.19355e-05 0.132187 0.983025 0.931739 -0.0132923 4.9152e-06 0.50723 -1.94138e-20 7.17878e-24 -1.94066e-20 0.00139586 0.997816 8.59811e-05 0.152652 2.85231 0.00139586 0.997817 0.748341 0.00105862 0.00188062 0.000859811 0.455504 0.00188062 0.441394 0.000129886 1.02 0.888194 0.534536 0.286765 1.71805e-07 3.0723e-09 2379.43 3116.86 -0.0558397 0.482169 0.277422 0.253352 -0.593354 -0.169541 0.495202 -0.266889 -0.228322 2.138 1 0 297.456 0 2.16137 2.136 0.000299631 0.854843 0.677291 0.343932 0.422236 2.16157 135.225 83.905 18.72 60.8588 0.00402595 0 -40 10
1.237 3.58144e-08 2.53926e-06 0.126006 0.126005 0.0120335 1.62793e-05 0.00115421 0.157507 0.000658418 0.158161 0.907078 101.707 0.240324 0.788409 4.2931 0.0596756 0.0405009 0.959499 0.0196863 0.00439455 0.0189485 0.00421163 0.00531373 0.00605153 0.212549 0.242061 58.0167 -87.8972 126.25 15.9544 145.025 0.000141279 0.267216 192.812 0.310413 0.0673522 0.00409692 0.000562033 0.00138397 0.986974 0.991725 -2.98237e-06 -85.6619 0.0930402 31180.6 304.657 0.983508 0.319146 0.732883 0.732879 9.99958 2.9839e-06 1.19355e-05 0.132191 0.983026 0.931739 -0.0132923 4.91523e-06 0.507244 -1.9415e-20 7.17926e-24 -1.94078e-20 0.00139586 0.997816 8.59812e-05 0.152652 2.85231 0.00139586 0.997817 0.748428 0.00105864 0.00188062 0.000859812 0.455504 0.00188062 0.441401 0.000129889 1.02 0.888195 0.534536 0.286767 1.71805e-07 3.07233e-09 2379.41 3116.88 -0.0558429 0.482169 0.277421 0.253354 -0.593353 -0.169541 0.495192 -0.266887 -0.228314 2.139 1 0 297.453 0 2.16152 2.137 0.00029963 0.854858 0.677336 0.343857 0.42226 2.16171 135.233 83.9047 18.72 60.8587 0.00402596 0 -40 10
1.238 3.58433e-08 2.53926e-06 0.126056 0.126055 0.0120335 1.62924e-05 0.00115421 0.15757 0.000658419 0.158223 0.907157 101.707 0.240315 0.788529 4.29349 0.0596852 0.0405046 0.959495 0.0196859 0.00439488 0.0189481 0.0042119 0.00531413 0.00605193 0.212565 0.242077 58.0167 -87.8972 126.25 15.9544 145.025 0.00014128 0.267217 192.812 0.310413 0.0673521 0.00409692 0.000562033 0.00138398 0.986974 0.991725 -2.98239e-06 -85.6619 0.0930403 31180.6 304.666 0.983508 0.319146 0.732889 0.732885 9.99958 2.98391e-06 1.19355e-05 0.132194 0.983028 0.931739 -0.0132923 4.91526e-06 0.507258 -1.94162e-20 7.17973e-24 -1.9409e-20 0.00139587 0.997816 8.59812e-05 0.152653 2.85231 0.00139587 0.997817 0.748516 0.00105866 0.00188062 0.000859812 0.455503 0.00188062 0.441407 0.000129892 1.02 0.888197 0.534536 0.286768 1.71806e-07 3.07235e-09 2379.4 3116.91 -0.0558461 0.482169 0.277421 0.253356 -0.593353 -0.169541 0.495181 -0.266885 -0.228305 2.14 1 0 297.45 0 2.16166 2.138 0.00029963 0.854873 0.677382 0.343783 0.422284 2.16186 135.241 83.9044 18.72 60.8585 0.00402597 0 -40 10
1.239 3.58722e-08 2.53926e-06 0.126106 0.126105 0.0120335 1.63055e-05 0.00115421 0.157632 0.00065842 0.158286 0.907237 101.706 0.240305 0.788649 4.29388 0.0596948 0.0405083 0.959492 0.0196855 0.0043952 0.0189477 0.00421218 0.00531453 0.00605234 0.212581 0.242093 58.0168 -87.8972 126.25 15.9544 145.025 0.000141281 0.267217 192.812 0.310412 0.0673521 0.00409692 0.000562034 0.00138398 0.986974 0.991725 -2.9824e-06 -85.6619 0.0930404 31180.6 304.675 0.983508 0.319146 0.732895 0.732891 9.99958 2.98391e-06 1.19355e-05 0.132197 0.983029 0.931738 -0.0132923 4.91529e-06 0.507272 -1.94173e-20 7.18021e-24 -1.94101e-20 0.00139587 0.997816 8.59813e-05 0.152653 2.85231 0.00139587 0.997817 0.748603 0.00105868 0.00188062 0.000859813 0.455503 0.00188062 0.441414 0.000129895 1.02 0.888198 0.534536 0.28677 1.71806e-07 3.07237e-09 2379.38 3116.94 -0.0558493 0.482169 0.277421 0.253357 -0.593353 -0.169541 0.495171 -0.266883 -0.228297 2.141 1 0 297.447 0 2.16181 2.139 0.000299629 0.854889 0.677427 0.343708 0.422307 2.162 135.249 83.9041 18.7199 60.8584 0.00402598 0 -40 10
1.24 3.59011e-08 2.53926e-06 0.126156 0.126155 0.0120335 1.63187e-05 0.00115421 0.157695 0.000658421 0.158348 0.907317 101.706 0.240296 0.788768 4.29427 0.0597044 0.040512 0.959488 0.0196851 0.00439553 0.0189473 0.00421246 0.00531493 0.00605274 0.212597 0.24211 58.0169 -87.8972 126.25 15.9543 145.025 0.000141282 0.267217 192.811 0.310412 0.067352 0.00409692 0.000562035 0.00138398 0.986974 0.991725 -2.98242e-06 -85.6619 0.0930405 31180.6 304.684 0.983508 0.319146 0.732901 0.732897 9.99958 2.98392e-06 1.19356e-05 0.132201 0.983031 0.931738 -0.0132923 4.91532e-06 0.507286 -1.94185e-20 7.18069e-24 -1.94113e-20 0.00139587 0.997816 8.59814e-05 0.152653 2.85231 0.00139587 0.997817 0.748691 0.0010587 0.00188063 0.000859814 0.455503 0.00188062 0.441421 0.000129898 1.02 0.888199 0.534535 0.286771 1.71806e-07 3.07239e-09 2379.36 3116.96 -0.0558525 0.482169 0.27742 0.253359 -0.593352 -0.169541 0.49516 -0.266881 -0.228288 2.142 1 0 297.445 0 2.16195 2.14 0.000299628 0.854904 0.677473 0.343634 0.422331 2.16215 135.257 83.9038 18.7199 60.8582 0.004026 0 -40 10
1.241 3.593e-08 2.53926e-06 0.126206 0.126205 0.0120335 1.63318e-05 0.00115421 0.157757 0.000658423 0.158411 0.907396 101.705 0.240286 0.788888 4.29466 0.059714 0.0405156 0.959484 0.0196847 0.00439585 0.0189469 0.00421273 0.00531533 0.00605315 0.212613 0.242126 58.0169 -87.8972 126.25 15.9543 145.025 0.000141283 0.267217 192.811 0.310412 0.067352 0.00409693 0.000562035 0.00138398 0.986974 0.991725 -2.98243e-06 -85.6618 0.0930405 31180.5 304.693 0.983508 0.319146 0.732908 0.732903 9.99958 2.98392e-06 1.19356e-05 0.132204 0.983032 0.931738 -0.0132923 4.91535e-06 0.5073 -1.94197e-20 7.18116e-24 -1.94125e-20 0.00139587 0.997816 8.59815e-05 0.152653 2.85232 0.00139587 0.997817 0.748778 0.00105871 0.00188063 0.000859815 0.455503 0.00188063 0.441427 0.0001299 1.02 0.8882 0.534535 0.286773 1.71806e-07 3.07242e-09 2379.35 3116.99 -0.0558557 0.482169 0.27742 0.253361 -0.593352 -0.169541 0.49515 -0.266879 -0.22828 2.143 1 0 297.442 0 2.1621 2.141 0.000299627 0.854919 0.677518 0.34356 0.422355 2.16229 135.264 83.9034 18.7199 60.8581 0.00402601 0 -40 10
1.242 3.59589e-08 2.53926e-06 0.126255 0.126254 0.0120334 1.63449e-05 0.00115421 0.157819 0.000658424 0.158473 0.907476 101.705 0.240276 0.789008 4.29505 0.0597236 0.0405193 0.959481 0.0196843 0.00439618 0.0189464 0.00421301 0.00531573 0.00605355 0.212629 0.242142 58.017 -87.8972 126.249 15.9543 145.025 0.000141285 0.267217 192.811 0.310411 0.0673519 0.00409693 0.000562036 0.00138398 0.986974 0.991725 -2.98245e-06 -85.6618 0.0930406 31180.5 304.701 0.983508 0.319146 0.732914 0.73291 9.99958 2.98393e-06 1.19356e-05 0.132207 0.983034 0.931737 -0.0132923 4.91538e-06 0.507313 -1.94208e-20 7.18164e-24 -1.94137e-20 0.00139587 0.997816 8.59816e-05 0.152653 2.85232 0.00139587 0.997817 0.748865 0.00105873 0.00188063 0.000859816 0.455502 0.00188063 0.441434 0.000129903 1.02 0.888201 0.534535 0.286774 1.71807e-07 3.07244e-09 2379.33 3117.01 -0.0558589 0.482169 0.27742 0.253362 -0.593352 -0.169541 0.495139 -0.266877 -0.228272 2.144 1 0 297.439 0 2.16224 2.142 0.000299626 0.854935 0.677564 0.343486 0.422379 2.16244 135.272 83.9031 18.7199 60.8579 0.00402602 0 -40 10
1.243 3.59878e-08 2.53926e-06 0.126305 0.126304 0.0120334 1.63581e-05 0.00115421 0.157882 0.000658425 0.158536 0.907556 101.705 0.240267 0.789127 4.29544 0.0597332 0.040523 0.959477 0.0196839 0.00439651 0.018946 0.00421329 0.00531614 0.00605396 0.212645 0.242158 58.017 -87.8972 126.249 15.9542 145.025 0.000141286 0.267218 192.811 0.310411 0.0673519 0.00409693 0.000562037 0.00138399 0.986974 0.991725 -2.98246e-06 -85.6618 0.0930407 31180.5 304.71 0.983508 0.319146 0.73292 0.732916 9.99958 2.98393e-06 1.19356e-05 0.132211 0.983035 0.931737 -0.0132923 4.91541e-06 0.507327 -1.9422e-20 7.18212e-24 -1.94148e-20 0.00139587 0.997816 8.59816e-05 0.152653 2.85232 0.00139587 0.997817 0.748953 0.00105875 0.00188063 0.000859816 0.455502 0.00188063 0.441441 0.000129906 1.02 0.888202 0.534534 0.286776 1.71807e-07 3.07246e-09 2379.31 3117.04 -0.0558622 0.482169 0.27742 0.253364 -0.593351 -0.169541 0.495128 -0.266875 -0.228263 2.145 1 0 297.436 0 2.16239 2.143 0.000299626 0.85495 0.677609 0.343412 0.422403 2.16258 135.28 83.9028 18.7199 60.8578 0.00402604 0 -40 10
1.244 3.60167e-08 2.53927e-06 0.126355 0.126354 0.0120334 1.63712e-05 0.00115421 0.157944 0.000658426 0.158598 0.907636 101.704 0.240257 0.789247 4.29583 0.0597428 0.0405267 0.959473 0.0196835 0.00439683 0.0189456 0.00421357 0.00531654 0.00605437 0.212661 0.242175 58.0171 -87.8972 126.249 15.9542 145.025 0.000141287 0.267218 192.811 0.31041 0.0673518 0.00409694 0.000562037 0.00138399 0.986974 0.991724 -2.98248e-06 -85.6618 0.0930408 31180.5 304.719 0.983508 0.319146 0.732926 0.732922 9.99958 2.98394e-06 1.19356e-05 0.132214 0.983037 0.931737 -0.0132923 4.91544e-06 0.507341 -1.94232e-20 7.1826e-24 -1.9416e-20 0.00139587 0.997816 8.59817e-05 0.152654 2.85232 0.00139587 0.997817 0.74904 0.00105877 0.00188063 0.000859817 0.455502 0.00188063 0.441447 0.000129909 1.02 0.888203 0.534534 0.286777 1.71807e-07 3.07249e-09 2379.3 3117.06 -0.0558654 0.482169 0.277419 0.253366 -0.593351 -0.169541 0.495118 -0.266873 -0.228255 2.146 1 0 297.434 0 2.16253 2.144 0.000299625 0.854966 0.677655 0.343338 0.422427 2.16273 135.288 83.9025 18.7199 60.8576 0.00402605 0 -40 10
1.245 3.60456e-08 2.53927e-06 0.126405 0.126404 0.0120334 1.63843e-05 0.00115421 0.158006 0.000658427 0.15866 0.907716 101.704 0.240248 0.789367 4.29622 0.0597524 0.0405304 0.95947 0.0196831 0.00439716 0.0189452 0.00421384 0.00531694 0.00605477 0.212678 0.242191 58.0172 -87.8972 126.249 15.9541 145.026 0.000141288 0.267218 192.811 0.31041 0.0673518 0.00409694 0.000562038 0.00138399 0.986974 0.991724 -2.98249e-06 -85.6618 0.0930409 31180.5 304.728 0.983508 0.319146 0.732933 0.732928 9.99958 2.98394e-06 1.19357e-05 0.132217 0.983038 0.931737 -0.0132923 4.91547e-06 0.507355 -1.94244e-20 7.18307e-24 -1.94172e-20 0.00139587 0.997816 8.59818e-05 0.152654 2.85232 0.00139587 0.997817 0.749127 0.00105879 0.00188063 0.000859818 0.455502 0.00188063 0.441454 0.000129912 1.02 0.888204 0.534534 0.286779 1.71808e-07 3.07251e-09 2379.28 3117.09 -0.0558686 0.482169 0.277419 0.253367 -0.593351 -0.169541 0.495107 -0.26687 -0.228246 2.147 1 0 297.431 0 2.16268 2.145 0.000299624 0.854981 0.6777 0.343264 0.422451 2.16287 135.296 83.9022 18.7198 60.8575 0.00402606 0 -40 10
1.246 3.60744e-08 2.53927e-06 0.126455 0.126454 0.0120334 1.63975e-05 0.00115421 0.158068 0.000658428 0.158722 0.907795 101.703 0.240238 0.789487 4.29662 0.059762 0.0405341 0.959466 0.0196827 0.00439749 0.0189448 0.00421412 0.00531734 0.00605518 0.212694 0.242207 58.0172 -87.8972 126.249 15.9541 145.026 0.000141289 0.267218 192.81 0.310409 0.0673517 0.00409694 0.000562039 0.00138399 0.986974 0.991724 -2.98251e-06 -85.6618 0.093041 31180.4 304.737 0.983508 0.319146 0.732939 0.732935 9.99958 2.98395e-06 1.19357e-05 0.132221 0.983039 0.931736 -0.0132923 4.9155e-06 0.507369 -1.94255e-20 7.18355e-24 -1.94183e-20 0.00139588 0.997816 8.59819e-05 0.152654 2.85232 0.00139587 0.997817 0.749214 0.0010588 0.00188063 0.000859819 0.455501 0.00188063 0.441461 0.000129915 1.02 0.888205 0.534533 0.28678 1.71808e-07 3.07253e-09 2379.26 3117.12 -0.0558719 0.482169 0.277419 0.253369 -0.59335 -0.169541 0.495096 -0.266868 -0.228238 2.148 1 0 297.428 0 2.16282 2.146 0.000299623 0.854997 0.677745 0.34319 0.422475 2.16302 135.303 83.9019 18.7198 60.8573 0.00402607 0 -40 10
1.247 3.61033e-08 2.53927e-06 0.126504 0.126503 0.0120334 1.64106e-05 0.00115421 0.15813 0.000658429 0.158784 0.907875 101.703 0.240228 0.789607 4.29701 0.0597716 0.0405378 0.959462 0.0196823 0.00439781 0.0189444 0.0042144 0.00531774 0.00605559 0.21271 0.242224 58.0173 -87.8972 126.249 15.9541 145.026 0.000141291 0.267218 192.81 0.310409 0.0673517 0.00409695 0.000562039 0.001384 0.986973 0.991724 -2.98252e-06 -85.6618 0.0930411 31180.4 304.746 0.983508 0.319146 0.732945 0.732941 9.99958 2.98395e-06 1.19357e-05 0.132224 0.983041 0.931736 -0.0132923 4.91553e-06 0.507383 -1.94267e-20 7.18403e-24 -1.94195e-20 0.00139588 0.997816 8.5982e-05 0.152654 2.85232 0.00139588 0.997817 0.749301 0.00105882 0.00188064 0.00085982 0.455501 0.00188063 0.441468 0.000129917 1.02 0.888206 0.534533 0.286782 1.71808e-07 3.07255e-09 2379.25 3117.14 -0.0558751 0.482169 0.277418 0.253371 -0.59335 -0.169541 0.495086 -0.266866 -0.228229 2.149 1 0 297.425 0 2.16297 2.147 0.000299623 0.855013 0.677791 0.343117 0.422499 2.16316 135.311 83.9016 18.7198 60.8572 0.00402609 0 -40 10
1.248 3.61322e-08 2.53927e-06 0.126554 0.126553 0.0120334 1.64237e-05 0.00115421 0.158192 0.00065843 0.158846 0.907955 101.703 0.240219 0.789727 4.2974 0.0597812 0.0405416 0.959458 0.0196819 0.00439814 0.018944 0.00421468 0.00531815 0.006056 0.212726 0.24224 58.0174 -87.8972 126.249 15.954 145.026 0.000141292 0.267219 192.81 0.310409 0.0673516 0.00409695 0.00056204 0.001384 0.986973 0.991724 -2.98254e-06 -85.6618 0.0930412 31180.4 304.755 0.983508 0.319146 0.732952 0.732947 9.99958 2.98396e-06 1.19357e-05 0.132227 0.983042 0.931736 -0.0132923 4.91556e-06 0.507397 -1.94279e-20 7.18451e-24 -1.94207e-20 0.00139588 0.997816 8.5982e-05 0.152654 2.85232 0.00139588 0.997817 0.749388 0.00105884 0.00188064 0.00085982 0.455501 0.00188064 0.441474 0.00012992 1.02 0.888208 0.534533 0.286784 1.71808e-07 3.07258e-09 2379.23 3117.17 -0.0558784 0.48217 0.277418 0.253372 -0.59335 -0.169541 0.495075 -0.266864 -0.22822 2.15 1 0 297.422 0 2.16311 2.148 0.000299622 0.855028 0.677836 0.343043 0.422522 2.16331 135.319 83.9013 18.7198 60.857 0.0040261 0 -40 10
1.249 3.61611e-08 2.53927e-06 0.126604 0.126603 0.0120333 1.64369e-05 0.00115421 0.158255 0.000658431 0.158908 0.908035 101.702 0.240209 0.789847 4.2978 0.0597909 0.0405453 0.959455 0.0196814 0.00439847 0.0189436 0.00421496 0.00531855 0.0060564 0.212742 0.242256 58.0174 -87.8973 126.249 15.954 145.026 0.000141293 0.267219 192.81 0.310408 0.0673516 0.00409695 0.000562041 0.001384 0.986973 0.991724 -2.98255e-06 -85.6618 0.0930412 31180.4 304.763 0.983508 0.319146 0.732958 0.732954 9.99958 2.98396e-06 1.19357e-05 0.132231 0.983044 0.931735 -0.0132923 4.91559e-06 0.507411 -1.94291e-20 7.18499e-24 -1.94219e-20 0.00139588 0.997816 8.59821e-05 0.152654 2.85232 0.00139588 0.997817 0.749475 0.00105886 0.00188064 0.000859821 0.455501 0.00188064 0.441481 0.000129923 1.02 0.888209 0.534532 0.286785 1.71809e-07 3.0726e-09 2379.21 3117.2 -0.0558817 0.48217 0.277418 0.253374 -0.593349 -0.169541 0.495064 -0.266862 -0.228212 2.151 1 0 297.419 0 2.16326 2.149 0.000299621 0.855044 0.677882 0.34297 0.422546 2.16345 135.327 83.9009 18.7198 60.8569 0.00402611 0 -40 10
1.25 3.619e-08 2.53927e-06 0.126653 0.126652 0.0120333 1.645e-05 0.00115421 0.158316 0.000658432 0.15897 0.908115 101.702 0.2402 0.789967 4.29819 0.0598005 0.040549 0.959451 0.019681 0.0043988 0.0189432 0.00421523 0.00531895 0.00605681 0.212758 0.242273 58.0175 -87.8973 126.249 15.9539 145.026 0.000141294 0.267219 192.81 0.310408 0.0673515 0.00409695 0.000562041 0.001384 0.986973 0.991724 -2.98257e-06 -85.6618 0.0930413 31180.3 304.772 0.983508 0.319146 0.732965 0.73296 9.99958 2.98397e-06 1.19358e-05 0.132234 0.983045 0.931735 -0.0132923 4.91562e-06 0.507425 -1.94302e-20 7.18547e-24 -1.94231e-20 0.00139588 0.997816 8.59822e-05 0.152654 2.85232 0.00139588 0.997817 0.749563 0.00105888 0.00188064 0.000859822 0.455501 0.00188064 0.441488 0.000129926 1.02 0.88821 0.534532 0.286787 1.71809e-07 3.07262e-09 2379.2 3117.22 -0.0558849 0.48217 0.277418 0.253376 -0.593349 -0.169542 0.495054 -0.26686 -0.228203 2.152 1 0 297.417 0 2.1634 2.15 0.00029962 0.85506 0.677927 0.342897 0.42257 2.1636 135.334 83.9006 18.7197 60.8567 0.00402613 0 -40 10
1.251 3.62189e-08 2.53927e-06 0.126703 0.126702 0.0120333 1.64631e-05 0.00115421 0.158378 0.000658433 0.159032 0.908195 101.701 0.24019 0.790087 4.29859 0.0598101 0.0405527 0.959447 0.0196806 0.00439913 0.0189428 0.00421551 0.00531936 0.00605722 0.212774 0.242289 58.0176 -87.8973 126.248 15.9539 145.026 0.000141296 0.267219 192.81 0.310407 0.0673515 0.00409696 0.000562042 0.001384 0.986973 0.991724 -2.98258e-06 -85.6618 0.0930414 31180.3 304.781 0.983508 0.319146 0.732971 0.732967 9.99958 2.98397e-06 1.19358e-05 0.132237 0.983047 0.931735 -0.0132923 4.91565e-06 0.507439 -1.94314e-20 7.18595e-24 -1.94242e-20 0.00139588 0.997816 8.59823e-05 0.152655 2.85233 0.00139588 0.997817 0.74965 0.00105889 0.00188064 0.000859823 0.4555 0.00188064 0.441494 0.000129929 1.02 0.888211 0.534532 0.286788 1.71809e-07 3.07265e-09 2379.18 3117.25 -0.0558882 0.48217 0.277417 0.253378 -0.593349 -0.169542 0.495043 -0.266858 -0.228194 2.153 1 0 297.414 0 2.16355 2.151 0.00029962 0.855076 0.677972 0.342824 0.422594 2.16374 135.342 83.9003 18.7197 60.8566 0.00402614 0 -40 10
1.252 3.62478e-08 2.53927e-06 0.126752 0.126751 0.0120333 1.64763e-05 0.00115422 0.15844 0.000658434 0.159094 0.908275 101.701 0.24018 0.790207 4.29898 0.0598198 0.0405565 0.959444 0.0196802 0.00439945 0.0189424 0.00421579 0.00531976 0.00605763 0.212791 0.242305 58.0176 -87.8973 126.248 15.9539 145.026 0.000141297 0.267219 192.809 0.310407 0.0673514 0.00409696 0.000562043 0.00138401 0.986973 0.991724 -2.9826e-06 -85.6617 0.0930415 31180.3 304.79 0.983508 0.319146 0.732977 0.732973 9.99958 2.98398e-06 1.19358e-05 0.132241 0.983048 0.931734 -0.0132923 4.91568e-06 0.507453 -1.94326e-20 7.18643e-24 -1.94254e-20 0.00139588 0.997816 8.59824e-05 0.152655 2.85233 0.00139588 0.997817 0.749737 0.00105891 0.00188064 0.000859824 0.4555 0.00188064 0.441501 0.000129932 1.02 0.888212 0.534532 0.28679 1.71809e-07 3.07267e-09 2379.16 3117.28 -0.0558915 0.48217 0.277417 0.253379 -0.593348 -0.169542 0.495032 -0.266856 -0.228186 2.154 1 0 297.411 0 2.16369 2.152 0.000299619 0.855092 0.678018 0.342751 0.422618 2.16389 135.35 83.9 18.7197 60.8564 0.00402615 0 -40 10
1.253 3.62767e-08 2.53927e-06 0.126802 0.126801 0.0120333 1.64894e-05 0.00115422 0.158502 0.000658435 0.159156 0.908355 101.701 0.240171 0.790327 4.29938 0.0598294 0.0405602 0.95944 0.0196798 0.00439978 0.018942 0.00421607 0.00532017 0.00605804 0.212807 0.242322 58.0177 -87.8973 126.248 15.9538 145.026 0.000141298 0.26722 192.809 0.310406 0.0673513 0.00409696 0.000562043 0.00138401 0.986973 0.991724 -2.98261e-06 -85.6617 0.0930416 31180.3 304.799 0.983508 0.319146 0.732984 0.73298 9.99958 2.98398e-06 1.19358e-05 0.132244 0.98305 0.931734 -0.0132923 4.91571e-06 0.507467 -1.94338e-20 7.18691e-24 -1.94266e-20 0.00139588 0.997816 8.59824e-05 0.152655 2.85233 0.00139588 0.997817 0.749823 0.00105893 0.00188064 0.000859824 0.4555 0.00188064 0.441508 0.000129934 1.02 0.888213 0.534531 0.286791 1.7181e-07 3.07269e-09 2379.15 3117.3 -0.0558948 0.48217 0.277417 0.253381 -0.593348 -0.169542 0.495021 -0.266854 -0.228177 2.155 1 0 297.408 0 2.16384 2.153 0.000299618 0.855108 0.678063 0.342678 0.422642 2.16403 135.358 83.8997 18.7197 60.8562 0.00402617 0 -40 10
1.254 3.63056e-08 2.53928e-06 0.126851 0.12685 0.0120333 1.65025e-05 0.00115422 0.158564 0.000658436 0.159218 0.908435 101.7 0.240161 0.790447 4.29978 0.059839 0.0405639 0.959436 0.0196794 0.00440011 0.0189415 0.00421635 0.00532057 0.00605845 0.212823 0.242338 58.0177 -87.8973 126.248 15.9538 145.026 0.000141299 0.26722 192.809 0.310406 0.0673513 0.00409697 0.000562044 0.00138401 0.986973 0.991724 -2.98263e-06 -85.6617 0.0930417 31180.2 304.808 0.983508 0.319146 0.73299 0.732986 9.99958 2.98399e-06 1.19358e-05 0.132247 0.983051 0.931734 -0.0132923 4.91574e-06 0.507481 -1.9435e-20 7.18739e-24 -1.94278e-20 0.00139588 0.997816 8.59825e-05 0.152655 2.85233 0.00139588 0.997817 0.74991 0.00105895 0.00188065 0.000859825 0.4555 0.00188064 0.441514 0.000129937 1.02 0.888214 0.534531 0.286793 1.7181e-07 3.07272e-09 2379.13 3117.33 -0.0558981 0.48217 0.277416 0.253383 -0.593347 -0.169542 0.49501 -0.266851 -0.228168 2.156 1 0 297.405 0 2.16398 2.154 0.000299617 0.855124 0.678108 0.342605 0.422666 2.16418 135.365 83.8994 18.7197 60.8561 0.00402618 0 -40 10
1.255 3.63345e-08 2.53928e-06 0.1269 0.126899 0.0120333 1.65157e-05 0.00115422 0.158626 0.000658438 0.159279 0.908515 101.7 0.240151 0.790567 4.30017 0.0598487 0.0405677 0.959432 0.019679 0.00440044 0.0189411 0.00421663 0.00532098 0.00605886 0.212839 0.242355 58.0178 -87.8973 126.248 15.9538 145.026 0.000141301 0.26722 192.809 0.310406 0.0673512 0.00409697 0.000562045 0.00138401 0.986973 0.991724 -2.98264e-06 -85.6617 0.0930418 31180.2 304.817 0.983508 0.319146 0.732997 0.732993 9.99958 2.98399e-06 1.19359e-05 0.132251 0.983053 0.931734 -0.0132923 4.91577e-06 0.507495 -1.94361e-20 7.18787e-24 -1.9429e-20 0.00139589 0.997816 8.59826e-05 0.152655 2.85233 0.00139589 0.997817 0.749997 0.00105896 0.00188065 0.000859826 0.455499 0.00188065 0.441521 0.00012994 1.02 0.888215 0.534531 0.286794 1.7181e-07 3.07274e-09 2379.11 3117.36 -0.0559014 0.48217 0.277416 0.253385 -0.593347 -0.169542 0.495 -0.266849 -0.22816 2.157 1 0 297.402 0 2.16413 2.155 0.000299617 0.85514 0.678154 0.342532 0.422689 2.16432 135.373 83.899 18.7196 60.8559 0.00402619 0 -40 10
1.256 3.63634e-08 2.53928e-06 0.12695 0.126949 0.0120333 1.65288e-05 0.00115422 0.158687 0.000658439 0.159341 0.908595 101.699 0.240142 0.790687 4.30057 0.0598583 0.0405714 0.959429 0.0196786 0.00440077 0.0189407 0.00421691 0.00532138 0.00605927 0.212855 0.242371 58.0179 -87.8973 126.248 15.9537 145.026 0.000141302 0.26722 192.809 0.310405 0.0673512 0.00409697 0.000562045 0.00138401 0.986973 0.991724 -2.98266e-06 -85.6617 0.0930419 31180.2 304.826 0.983508 0.319146 0.733004 0.732999 9.99958 2.984e-06 1.19359e-05 0.132254 0.983054 0.931733 -0.0132923 4.91579e-06 0.507509 -1.94373e-20 7.18835e-24 -1.94301e-20 0.00139589 0.997816 8.59827e-05 0.152655 2.85233 0.00139589 0.997817 0.750084 0.00105898 0.00188065 0.000859827 0.455499 0.00188065 0.441528 0.000129943 1.02 0.888216 0.53453 0.286796 1.71811e-07 3.07276e-09 2379.1 3117.38 -0.0559048 0.48217 0.277416 0.253386 -0.593347 -0.169542 0.494989 -0.266847 -0.228151 2.158 1 0 297.399 0 2.16427 2.156 0.000299616 0.855156 0.678199 0.34246 0.422713 2.16447 135.381 83.8987 18.7196 60.8558 0.00402621 0 -40 10
1.257 3.63923e-08 2.53928e-06 0.126999 0.126998 0.0120332 1.65419e-05 0.00115422 0.158749 0.00065844 0.159403 0.908675 101.699 0.240132 0.790808 4.30097 0.059868 0.0405752 0.959425 0.0196782 0.0044011 0.0189403 0.00421719 0.00532179 0.00605969 0.212872 0.242387 58.0179 -87.8973 126.248 15.9537 145.026 0.000141303 0.26722 192.809 0.310405 0.0673511 0.00409698 0.000562046 0.00138402 0.986973 0.991724 -2.98267e-06 -85.6617 0.0930419 31180.2 304.835 0.983508 0.319146 0.73301 0.733006 9.99958 2.984e-06 1.19359e-05 0.132257 0.983055 0.931733 -0.0132923 4.91582e-06 0.507524 -1.94385e-20 7.18884e-24 -1.94313e-20 0.00139589 0.997816 8.59828e-05 0.152656 2.85233 0.00139589 0.997817 0.750171 0.001059 0.00188065 0.000859828 0.455499 0.00188065 0.441534 0.000129946 1.02 0.888217 0.53453 0.286797 1.71811e-07 3.07278e-09 2379.08 3117.41 -0.0559081 0.48217 0.277416 0.253388 -0.593346 -0.169542 0.494978 -0.266845 -0.228142 2.159 1 0 297.397 0 2.16442 2.157 0.000299615 0.855172 0.678245 0.342387 0.422737 2.16461 135.389 83.8984 18.7196 60.8556 0.00402622 0 -40 10
1.258 3.64211e-08 2.53928e-06 0.127048 0.127047 0.0120332 1.65551e-05 0.00115422 0.15881 0.000658441 0.159464 0.908755 101.699 0.240122 0.790928 4.30137 0.0598776 0.0405789 0.959421 0.0196778 0.00440143 0.0189399 0.00421748 0.0053222 0.0060601 0.212888 0.242404 58.018 -87.8973 126.248 15.9536 145.026 0.000141304 0.26722 192.808 0.310404 0.0673511 0.00409698 0.000562047 0.00138402 0.986973 0.991724 -2.98269e-06 -85.6617 0.093042 31180.2 304.844 0.983508 0.319146 0.733017 0.733012 9.99958 2.984e-06 1.19359e-05 0.132261 0.983057 0.931733 -0.0132923 4.91585e-06 0.507538 -1.94397e-20 7.18932e-24 -1.94325e-20 0.00139589 0.997816 8.59829e-05 0.152656 2.85233 0.00139589 0.997817 0.750258 0.00105902 0.00188065 0.000859829 0.455499 0.00188065 0.441541 0.000129949 1.02 0.888218 0.53453 0.286799 1.71811e-07 3.07281e-09 2379.06 3117.44 -0.0559114 0.48217 0.277415 0.25339 -0.593346 -0.169542 0.494967 -0.266843 -0.228133 2.16 1 0 297.394 0 2.16456 2.158 0.000299614 0.855188 0.67829 0.342315 0.422761 2.16475 135.396 83.8981 18.7196 60.8555 0.00402623 0 -40 10
1.259 3.645e-08 2.53928e-06 0.127098 0.127096 0.0120332 1.65682e-05 0.00115422 0.158872 0.000658442 0.159526 0.908836 101.698 0.240113 0.791048 4.30177 0.0598873 0.0405827 0.959417 0.0196774 0.00440176 0.0189395 0.00421776 0.0053226 0.00606051 0.212904 0.24242 58.0181 -87.8973 126.247 15.9536 145.026 0.000141306 0.267221 192.808 0.310404 0.067351 0.00409698 0.000562047 0.00138402 0.986973 0.991724 -2.9827e-06 -85.6617 0.0930421 31180.1 304.853 0.983508 0.319146 0.733023 0.733019 9.99958 2.98401e-06 1.19359e-05 0.132264 0.983058 0.931732 -0.0132923 4.91588e-06 0.507552 -1.94409e-20 7.1898e-24 -1.94337e-20 0.00139589 0.997816 8.59829e-05 0.152656 2.85233 0.00139589 0.997817 0.750345 0.00105904 0.00188065 0.000859829 0.455499 0.00188065 0.441547 0.000129951 1.02 0.88822 0.534529 0.2868 1.71811e-07 3.07283e-09 2379.05 3117.47 -0.0559148 0.48217 0.277415 0.253392 -0.593346 -0.169542 0.494956 -0.266841 -0.228124 2.161 1 0 297.391 0 2.1647 2.159 0.000299613 0.855204 0.678335 0.342243 0.422785 2.1649 135.404 83.8977 18.7196 60.8553 0.00402625 0 -40 10
1.26 3.64789e-08 2.53928e-06 0.127147 0.127146 0.0120332 1.65813e-05 0.00115422 0.158933 0.000658443 0.159587 0.908916 101.698 0.240103 0.791169 4.30216 0.059897 0.0405865 0.959414 0.019677 0.00440209 0.0189391 0.00421804 0.00532301 0.00606092 0.21292 0.242437 58.0181 -87.8973 126.247 15.9536 145.026 0.000141307 0.267221 192.808 0.310403 0.067351 0.00409699 0.000562048 0.00138402 0.986973 0.991724 -2.98272e-06 -85.6617 0.0930422 31180.1 304.862 0.983508 0.319146 0.73303 0.733026 9.99958 2.98401e-06 1.1936e-05 0.132268 0.98306 0.931732 -0.0132923 4.91591e-06 0.507566 -1.94421e-20 7.19028e-24 -1.94349e-20 0.00139589 0.997816 8.5983e-05 0.152656 2.85233 0.00139589 0.997817 0.750431 0.00105905 0.00188066 0.00085983 0.455498 0.00188065 0.441554 0.000129954 1.02 0.888221 0.534529 0.286802 1.71812e-07 3.07285e-09 2379.03 3117.49 -0.0559181 0.48217 0.277415 0.253394 -0.593345 -0.169542 0.494945 -0.266839 -0.228116 2.162 1 0 297.388 0 2.16485 2.16 0.000299613 0.855221 0.678381 0.342171 0.422809 2.16504 135.412 83.8974 18.7196 60.8552 0.00402626 0 -40 10
1.261 3.65078e-08 2.53928e-06 0.127196 0.127195 0.0120332 1.65945e-05 0.00115422 0.158995 0.000658444 0.159649 0.908996 101.697 0.240093 0.791289 4.30256 0.0599066 0.0405902 0.95941 0.0196766 0.00440243 0.0189387 0.00421832 0.00532342 0.00606134 0.212937 0.242453 58.0182 -87.8973 126.247 15.9535 145.026 0.000141308 0.267221 192.808 0.310403 0.0673509 0.00409699 0.000562049 0.00138403 0.986973 0.991724 -2.98273e-06 -85.6617 0.0930423 31180.1 304.871 0.983508 0.319146 0.733037 0.733032 9.99958 2.98402e-06 1.1936e-05 0.132271 0.983061 0.931732 -0.0132923 4.91594e-06 0.50758 -1.94433e-20 7.19077e-24 -1.94361e-20 0.00139589 0.997816 8.59831e-05 0.152656 2.85233 0.00139589 0.997817 0.750518 0.00105907 0.00188066 0.000859831 0.455498 0.00188066 0.441561 0.000129957 1.02 0.888222 0.534529 0.286803 1.71812e-07 3.07288e-09 2379.01 3117.52 -0.0559215 0.482171 0.277415 0.253395 -0.593345 -0.169542 0.494934 -0.266837 -0.228107 2.163 1 0 297.385 0 2.16499 2.161 0.000299612 0.855237 0.678426 0.342099 0.422832 2.16519 135.42 83.8971 18.7195 60.855 0.00402627 0 -40 10
1.262 3.65367e-08 2.53928e-06 0.127245 0.127244 0.0120332 1.66076e-05 0.00115422 0.159056 0.000658445 0.15971 0.909076 101.697 0.240084 0.79141 4.30296 0.0599163 0.040594 0.959406 0.0196762 0.00440276 0.0189383 0.0042186 0.00532383 0.00606175 0.212953 0.24247 58.0183 -87.8973 126.247 15.9535 145.026 0.00014131 0.267221 192.808 0.310403 0.0673509 0.00409699 0.000562049 0.00138403 0.986973 0.991724 -2.98275e-06 -85.6616 0.0930424 31180.1 304.88 0.983508 0.319146 0.733043 0.733039 9.99958 2.98402e-06 1.1936e-05 0.132274 0.983062 0.931731 -0.0132923 4.91597e-06 0.507594 -1.94444e-20 7.19125e-24 -1.94372e-20 0.00139589 0.997816 8.59832e-05 0.152656 2.85234 0.00139589 0.997817 0.750605 0.00105909 0.00188066 0.000859832 0.455498 0.00188066 0.441567 0.00012996 1.02 0.888223 0.534528 0.286805 1.71812e-07 3.0729e-09 2379 3117.55 -0.0559248 0.482171 0.277414 0.253397 -0.593345 -0.169542 0.494923 -0.266835 -0.228098 2.164 1 0 297.382 0 2.16514 2.162 0.000299611 0.855253 0.678471 0.342027 0.422856 2.16533 135.428 83.8967 18.7195 60.8548 0.00402629 0 -40 10
1.263 3.65656e-08 2.53928e-06 0.127294 0.127293 0.0120332 1.66207e-05 0.00115422 0.159117 0.000658446 0.159771 0.909157 101.697 0.240074 0.79153 4.30337 0.059926 0.0405978 0.959402 0.0196758 0.00440309 0.0189378 0.00421888 0.00532424 0.00606216 0.212969 0.242487 58.0183 -87.8973 126.247 15.9535 145.026 0.000141311 0.267221 192.808 0.310402 0.0673508 0.00409699 0.00056205 0.00138403 0.986973 0.991724 -2.98276e-06 -85.6616 0.0930425 31180 304.889 0.983507 0.319146 0.73305 0.733046 9.99958 2.98403e-06 1.1936e-05 0.132278 0.983064 0.931731 -0.0132923 4.916e-06 0.507608 -1.94456e-20 7.19173e-24 -1.94384e-20 0.00139589 0.997816 8.59833e-05 0.152656 2.85234 0.00139589 0.997817 0.750691 0.00105911 0.00188066 0.000859833 0.455498 0.00188066 0.441574 0.000129963 1.02 0.888224 0.534528 0.286806 1.71812e-07 3.07292e-09 2378.98 3117.58 -0.0559282 0.482171 0.277414 0.253399 -0.593344 -0.169542 0.494912 -0.266832 -0.228089 2.165 1 0 297.379 0 2.16528 2.163 0.00029961 0.85527 0.678516 0.341955 0.42288 2.16548 135.435 83.8964 18.7195 60.8547 0.0040263 0 -40 10
1.264 3.65945e-08 2.53929e-06 0.127343 0.127342 0.0120331 1.66339e-05 0.00115422 0.159179 0.000658447 0.159833 0.909237 101.696 0.240064 0.791651 4.30377 0.0599356 0.0406016 0.959398 0.0196754 0.00440342 0.0189374 0.00421917 0.00532464 0.00606258 0.212986 0.242503 58.0184 -87.8973 126.247 15.9534 145.026 0.000141312 0.267222 192.807 0.310402 0.0673508 0.004097 0.000562051 0.00138403 0.986973 0.991724 -2.98278e-06 -85.6616 0.0930426 31180 304.898 0.983507 0.319146 0.733057 0.733052 9.99958 2.98403e-06 1.1936e-05 0.132281 0.983065 0.931731 -0.0132923 4.91603e-06 0.507623 -1.94468e-20 7.19222e-24 -1.94396e-20 0.0013959 0.997816 8.59833e-05 0.152657 2.85234 0.0013959 0.997817 0.750778 0.00105913 0.00188066 0.000859833 0.455497 0.00188066 0.441581 0.000129965 1.02 0.888225 0.534528 0.286808 1.71813e-07 3.07294e-09 2378.96 3117.6 -0.0559316 0.482171 0.277414 0.253401 -0.593344 -0.169542 0.494901 -0.26683 -0.22808 2.166 1 0 297.376 0 2.16543 2.164 0.00029961 0.855286 0.678562 0.341884 0.422904 2.16562 135.443 83.8961 18.7195 60.8545 0.00402631 0 -40 10
1.265 3.66234e-08 2.53929e-06 0.127392 0.127391 0.0120331 1.6647e-05 0.00115422 0.15924 0.000658448 0.159894 0.909317 101.696 0.240055 0.791771 4.30417 0.0599453 0.0406054 0.959395 0.0196749 0.00440375 0.018937 0.00421945 0.00532505 0.00606299 0.213002 0.24252 58.0184 -87.8973 126.247 15.9534 145.026 0.000141313 0.267222 192.807 0.310401 0.0673507 0.004097 0.000562051 0.00138403 0.986973 0.991724 -2.98279e-06 -85.6616 0.0930426 31180 304.907 0.983507 0.319146 0.733063 0.733059 9.99958 2.98404e-06 1.19361e-05 0.132285 0.983067 0.93173 -0.0132923 4.91606e-06 0.507637 -1.9448e-20 7.1927e-24 -1.94408e-20 0.0013959 0.997816 8.59834e-05 0.152657 2.85234 0.0013959 0.997817 0.750865 0.00105914 0.00188066 0.000859834 0.455497 0.00188066 0.441587 0.000129968 1.02 0.888226 0.534528 0.286809 1.71813e-07 3.07297e-09 2378.95 3117.63 -0.055935 0.482171 0.277413 0.253403 -0.593343 -0.169542 0.49489 -0.266828 -0.228071 2.167 1 0 297.373 0 2.16557 2.165 0.000299609 0.855303 0.678607 0.341812 0.422928 2.16577 135.451 83.8957 18.7195 60.8544 0.00402633 0 -40 10
1.266 3.66523e-08 2.53929e-06 0.127441 0.12744 0.0120331 1.66601e-05 0.00115422 0.159301 0.000658449 0.159955 0.909398 101.695 0.240045 0.791892 4.30457 0.059955 0.0406091 0.959391 0.0196745 0.00440409 0.0189366 0.00421973 0.00532546 0.00606341 0.213019 0.242536 58.0185 -87.8973 126.247 15.9533 145.026 0.000141315 0.267222 192.807 0.310401 0.0673507 0.004097 0.000562052 0.00138404 0.986973 0.991724 -2.98281e-06 -85.6616 0.0930427 31180 304.916 0.983507 0.319146 0.73307 0.733066 9.99958 2.98404e-06 1.19361e-05 0.132288 0.983068 0.93173 -0.0132923 4.91609e-06 0.507651 -1.94492e-20 7.19319e-24 -1.9442e-20 0.0013959 0.997816 8.59835e-05 0.152657 2.85234 0.0013959 0.997817 0.750951 0.00105916 0.00188066 0.000859835 0.455497 0.00188066 0.441594 0.000129971 1.02 0.888227 0.534527 0.286811 1.71813e-07 3.07299e-09 2378.93 3117.66 -0.0559383 0.482171 0.277413 0.253404 -0.593343 -0.169543 0.494879 -0.266826 -0.228062 2.168 1 0 297.37 0 2.16572 2.166 0.000299608 0.855319 0.678652 0.341741 0.422951 2.16591 135.459 83.8954 18.7194 60.8542 0.00402634 0 -40 10
1.267 3.66812e-08 2.53929e-06 0.12749 0.127489 0.0120331 1.66733e-05 0.00115422 0.159362 0.00065845 0.160016 0.909478 101.695 0.240035 0.792012 4.30497 0.0599647 0.0406129 0.959387 0.0196741 0.00440442 0.0189362 0.00422002 0.00532587 0.00606382 0.213035 0.242553 58.0186 -87.8973 126.246 15.9533 145.026 0.000141316 0.267222 192.807 0.3104 0.0673506 0.00409701 0.000562053 0.00138404 0.986973 0.991724 -2.98282e-06 -85.6616 0.0930428 31180 304.925 0.983507 0.319146 0.733077 0.733073 9.99958 2.98405e-06 1.19361e-05 0.132291 0.983069 0.93173 -0.0132923 4.91612e-06 0.507665 -1.94504e-20 7.19367e-24 -1.94432e-20 0.0013959 0.997816 8.59836e-05 0.152657 2.85234 0.0013959 0.997817 0.751038 0.00105918 0.00188067 0.000859836 0.455497 0.00188066 0.441601 0.000129974 1.02 0.888228 0.534527 0.286812 1.71813e-07 3.07301e-09 2378.91 3117.69 -0.0559417 0.482171 0.277413 0.253406 -0.593343 -0.169543 0.494868 -0.266824 -0.228053 2.169 1 0 297.367 0 2.16586 2.167 0.000299607 0.855336 0.678698 0.341669 0.422975 2.16606 135.466 83.8951 18.7194 60.854 0.00402636 0 -40 10
1.268 3.67101e-08 2.53929e-06 0.127539 0.127538 0.0120331 1.66864e-05 0.00115422 0.159423 0.000658451 0.160077 0.909558 101.695 0.240026 0.792133 4.30537 0.0599743 0.0406167 0.959383 0.0196737 0.00440475 0.0189358 0.0042203 0.00532628 0.00606424 0.213051 0.24257 58.0186 -87.8973 126.246 15.9533 145.026 0.000141317 0.267222 192.807 0.3104 0.0673506 0.00409701 0.000562053 0.00138404 0.986973 0.991724 -2.98284e-06 -85.6616 0.0930429 31179.9 304.934 0.983507 0.319146 0.733084 0.733079 9.99958 2.98405e-06 1.19361e-05 0.132295 0.983071 0.931729 -0.0132923 4.91615e-06 0.507679 -1.94516e-20 7.19416e-24 -1.94444e-20 0.0013959 0.997816 8.59837e-05 0.152657 2.85234 0.0013959 0.997817 0.751124 0.0010592 0.00188067 0.000859837 0.455497 0.00188067 0.441607 0.000129977 1.02 0.888229 0.534527 0.286814 1.71814e-07 3.07304e-09 2378.9 3117.72 -0.0559451 0.482171 0.277413 0.253408 -0.593342 -0.169543 0.494856 -0.266822 -0.228044 2.17 1 0 297.364 0 2.16601 2.168 0.000299606 0.855352 0.678743 0.341598 0.422999 2.1662 135.474 83.8947 18.7194 60.8539 0.00402637 0 -40 10
1.269 3.67389e-08 2.53929e-06 0.127587 0.127586 0.0120331 1.66995e-05 0.00115422 0.159484 0.000658452 0.160138 0.909639 101.694 0.240016 0.792254 4.30578 0.059984 0.0406205 0.959379 0.0196733 0.00440509 0.0189353 0.00422058 0.00532669 0.00606465 0.213068 0.242586 58.0187 -87.8973 126.246 15.9532 145.026 0.000141319 0.267223 192.807 0.3104 0.0673505 0.00409701 0.000562054 0.00138404 0.986973 0.991724 -2.98285e-06 -85.6616 0.093043 31179.9 304.943 0.983507 0.319146 0.733091 0.733086 9.99958 2.98406e-06 1.19361e-05 0.132298 0.983072 0.931729 -0.0132923 4.91618e-06 0.507694 -1.94528e-20 7.19464e-24 -1.94456e-20 0.0013959 0.997816 8.59837e-05 0.152657 2.85234 0.0013959 0.997817 0.751211 0.00105922 0.00188067 0.000859837 0.455496 0.00188067 0.441614 0.00012998 1.02 0.888231 0.534526 0.286815 1.71814e-07 3.07306e-09 2378.88 3117.74 -0.0559486 0.482171 0.277412 0.25341 -0.593342 -0.169543 0.494845 -0.26682 -0.228035 2.171 1 0 297.361 0 2.16615 2.169 0.000299606 0.855369 0.678788 0.341527 0.423023 2.16634 135.482 83.8944 18.7194 60.8537 0.00402638 0 -40 10
1.27 3.67678e-08 2.53929e-06 0.127636 0.127635 0.0120331 1.67127e-05 0.00115422 0.159545 0.000658453 0.160199 0.909719 101.694 0.240006 0.792375 4.30618 0.0599937 0.0406244 0.959376 0.0196729 0.00440542 0.0189349 0.00422087 0.0053271 0.00606507 0.213084 0.242603 58.0188 -87.8973 126.246 15.9532 145.026 0.00014132 0.267223 192.806 0.310399 0.0673505 0.00409702 0.000562055 0.00138405 0.986973 0.991724 -2.98287e-06 -85.6616 0.0930431 31179.9 304.952 0.983507 0.319146 0.733098 0.733093 9.99958 2.98406e-06 1.19362e-05 0.132302 0.983073 0.931728 -0.0132923 4.91621e-06 0.507708 -1.9454e-20 7.19513e-24 -1.94468e-20 0.0013959 0.997816 8.59838e-05 0.152658 2.85234 0.0013959 0.997817 0.751297 0.00105923 0.00188067 0.000859838 0.455496 0.00188067 0.44162 0.000129982 1.02 0.888232 0.534526 0.286817 1.71814e-07 3.07308e-09 2378.86 3117.77 -0.055952 0.482171 0.277412 0.253412 -0.593342 -0.169543 0.494834 -0.266818 -0.228026 2.172 1 0 297.358 0 2.16629 2.17 0.000299605 0.855386 0.678833 0.341456 0.423047 2.16649 135.49 83.8941 18.7194 60.8535 0.0040264 0 -40 10
1.271 3.67967e-08 2.53929e-06 0.127685 0.127684 0.0120331 1.67258e-05 0.00115422 0.159606 0.000658454 0.16026 0.9098 101.693 0.239997 0.792495 4.30659 0.0600034 0.0406282 0.959372 0.0196725 0.00440575 0.0189345 0.00422115 0.00532752 0.00606549 0.213101 0.242619 58.0188 -87.8973 126.246 15.9532 145.026 0.000141321 0.267223 192.806 0.310399 0.0673504 0.00409702 0.000562056 0.00138405 0.986973 0.991724 -2.98288e-06 -85.6616 0.0930432 31179.9 304.961 0.983507 0.319146 0.733104 0.7331 9.99958 2.98407e-06 1.19362e-05 0.132305 0.983075 0.931728 -0.0132923 4.91624e-06 0.507722 -1.94552e-20 7.19562e-24 -1.9448e-20 0.0013959 0.997816 8.59839e-05 0.152658 2.85234 0.0013959 0.997817 0.751384 0.00105925 0.00188067 0.000859839 0.455496 0.00188067 0.441627 0.000129985 1.02 0.888233 0.534526 0.286819 1.71815e-07 3.0731e-09 2378.85 3117.8 -0.0559554 0.482171 0.277412 0.253414 -0.593341 -0.169543 0.494823 -0.266816 -0.228017 2.173 1 0 297.355 0 2.16644 2.171 0.000299604 0.855403 0.678879 0.341385 0.42307 2.16663 135.497 83.8937 18.7193 60.8534 0.00402641 0 -40 10
1.272 3.68256e-08 2.53929e-06 0.127734 0.127733 0.012033 1.67389e-05 0.00115422 0.159667 0.000658455 0.160321 0.90988 101.693 0.239987 0.792616 4.30699 0.0600131 0.040632 0.959368 0.0196721 0.00440609 0.0189341 0.00422144 0.00532793 0.0060659 0.213117 0.242636 58.0189 -87.8973 126.246 15.9531 145.026 0.000141323 0.267223 192.806 0.310398 0.0673503 0.00409702 0.000562056 0.00138405 0.986973 0.991724 -2.9829e-06 -85.6616 0.0930433 31179.8 304.97 0.983507 0.319146 0.733111 0.733107 9.99958 2.98407e-06 1.19362e-05 0.132308 0.983076 0.931728 -0.0132923 4.91627e-06 0.507736 -1.94564e-20 7.1961e-24 -1.94492e-20 0.0013959 0.997816 8.5984e-05 0.152658 2.85234 0.0013959 0.997817 0.75147 0.00105927 0.00188067 0.00085984 0.455496 0.00188067 0.441634 0.000129988 1.02 0.888234 0.534525 0.28682 1.71815e-07 3.07313e-09 2378.83 3117.83 -0.0559588 0.482171 0.277411 0.253415 -0.593341 -0.169543 0.494812 -0.266813 -0.228008 2.174 1 0 297.352 0 2.16658 2.172 0.000299603 0.85542 0.678924 0.341315 0.423094 2.16678 135.505 83.8934 18.7193 60.8532 0.00402642 0 -40 10
1.273 3.68545e-08 2.53929e-06 0.127782 0.127781 0.012033 1.6752e-05 0.00115422 0.159728 0.000658456 0.160382 0.909961 101.693 0.239977 0.792737 4.3074 0.0600228 0.0406358 0.959364 0.0196717 0.00440642 0.0189337 0.00422172 0.00532834 0.00606632 0.213134 0.242653 58.0189 -87.8973 126.246 15.9531 145.026 0.000141324 0.267223 192.806 0.310398 0.0673503 0.00409702 0.000562057 0.00138405 0.986973 0.991724 -2.98291e-06 -85.6615 0.0930433 31179.8 304.979 0.983507 0.319146 0.733118 0.733114 9.99958 2.98408e-06 1.19362e-05 0.132312 0.983077 0.931727 -0.0132923 4.9163e-06 0.507751 -1.94576e-20 7.19659e-24 -1.94504e-20 0.00139591 0.997816 8.59841e-05 0.152658 2.85235 0.00139591 0.997817 0.751556 0.00105929 0.00188067 0.000859841 0.455495 0.00188067 0.44164 0.000129991 1.02 0.888235 0.534525 0.286822 1.71815e-07 3.07315e-09 2378.81 3117.86 -0.0559623 0.482171 0.277411 0.253417 -0.59334 -0.169543 0.494801 -0.266811 -0.227999 2.175 1 0 297.349 0 2.16673 2.173 0.000299603 0.855436 0.678969 0.341244 0.423118 2.16692 135.513 83.893 18.7193 60.8531 0.00402644 0 -40 10
1.274 3.68834e-08 2.53929e-06 0.127831 0.12783 0.012033 1.67652e-05 0.00115422 0.159789 0.000658457 0.160443 0.910042 101.692 0.239967 0.792858 4.3078 0.0600325 0.0406396 0.95936 0.0196712 0.00440676 0.0189333 0.00422201 0.00532875 0.00606674 0.21315 0.24267 58.019 -87.8973 126.246 15.953 145.026 0.000141325 0.267224 192.806 0.310397 0.0673502 0.00409703 0.000562058 0.00138405 0.986973 0.991724 -2.98293e-06 -85.6615 0.0930434 31179.8 304.988 0.983507 0.319146 0.733125 0.733121 9.99958 2.98408e-06 1.19362e-05 0.132315 0.983079 0.931727 -0.0132923 4.91633e-06 0.507765 -1.94588e-20 7.19708e-24 -1.94516e-20 0.00139591 0.997816 8.59841e-05 0.152658 2.85235 0.00139591 0.997817 0.751643 0.0010593 0.00188068 0.000859841 0.455495 0.00188067 0.441647 0.000129994 1.02 0.888236 0.534525 0.286823 1.71815e-07 3.07317e-09 2378.8 3117.89 -0.0559657 0.482172 0.277411 0.253419 -0.59334 -0.169543 0.494789 -0.266809 -0.227989 2.176 1 0 297.346 0 2.16687 2.174 0.000299602 0.855453 0.679014 0.341173 0.423142 2.16707 135.52 83.8927 18.7193 60.8529 0.00402645 0 -40 10
1.275 3.69123e-08 2.5393e-06 0.12788 0.127879 0.012033 1.67783e-05 0.00115423 0.159849 0.000658458 0.160503 0.910122 101.692 0.239958 0.792979 4.30821 0.0600422 0.0406435 0.959357 0.0196708 0.00440709 0.0189328 0.00422229 0.00532916 0.00606716 0.213167 0.242686 58.0191 -87.8973 126.245 15.953 145.026 0.000141327 0.267224 192.806 0.310397 0.0673502 0.00409703 0.000562058 0.00138406 0.986973 0.991724 -2.98294e-06 -85.6615 0.0930435 31179.8 304.998 0.983507 0.319146 0.733132 0.733128 9.99958 2.98409e-06 1.19362e-05 0.132319 0.98308 0.931727 -0.0132923 4.91636e-06 0.507779 -1.946e-20 7.19756e-24 -1.94528e-20 0.00139591 0.997816 8.59842e-05 0.152658 2.85235 0.00139591 0.997817 0.751729 0.00105932 0.00188068 0.000859842 0.455495 0.00188068 0.441653 0.000129996 1.02 0.888237 0.534524 0.286825 1.71816e-07 3.0732e-09 2378.78 3117.92 -0.0559692 0.482172 0.277411 0.253421 -0.59334 -0.169543 0.494778 -0.266807 -0.22798 2.177 1 0 297.343 0 2.16702 2.175 0.000299601 0.85547 0.67906 0.341103 0.423165 2.16721 135.528 83.8923 18.7193 60.8527 0.00402647 0 -40 10
1.276 3.69412e-08 2.5393e-06 0.127928 0.127927 0.012033 1.67914e-05 0.00115423 0.15991 0.000658459 0.160564 0.910203 101.691 0.239948 0.7931 4.30861 0.0600519 0.0406473 0.959353 0.0196704 0.00440743 0.0189324 0.00422258 0.00532958 0.00606758 0.213183 0.242703 58.0191 -87.8974 126.245 15.953 145.026 0.000141328 0.267224 192.805 0.310397 0.0673501 0.00409703 0.000562059 0.00138406 0.986973 0.991724 -2.98296e-06 -85.6615 0.0930436 31179.8 305.007 0.983507 0.319146 0.733139 0.733135 9.99958 2.98409e-06 1.19363e-05 0.132322 0.983081 0.931726 -0.0132923 4.91639e-06 0.507794 -1.94612e-20 7.19805e-24 -1.9454e-20 0.00139591 0.997816 8.59843e-05 0.152658 2.85235 0.00139591 0.997817 0.751815 0.00105934 0.00188068 0.000859843 0.455495 0.00188068 0.44166 0.000129999 1.02 0.888238 0.534524 0.286826 1.71816e-07 3.07322e-09 2378.76 3117.95 -0.0559726 0.482172 0.27741 0.253423 -0.593339 -0.169543 0.494767 -0.266805 -0.227971 2.178 1 0 297.34 0 2.16716 2.176 0.0002996 0.855487 0.679105 0.341033 0.423189 2.16736 135.536 83.892 18.7192 60.8526 0.00402648 0 -40 10
1.277 3.69701e-08 2.5393e-06 0.127977 0.127976 0.012033 1.68046e-05 0.00115423 0.159971 0.00065846 0.160625 0.910283 101.691 0.239938 0.793221 4.30902 0.0600616 0.0406511 0.959349 0.01967 0.00440776 0.018932 0.00422286 0.00532999 0.006068 0.2132 0.24272 58.0192 -87.8974 126.245 15.9529 145.026 0.000141329 0.267224 192.805 0.310396 0.0673501 0.00409704 0.00056206 0.00138406 0.986973 0.991724 -2.98297e-06 -85.6615 0.0930437 31179.7 305.016 0.983507 0.319146 0.733146 0.733142 9.99958 2.9841e-06 1.19363e-05 0.132325 0.983083 0.931726 -0.0132923 4.91642e-06 0.507808 -1.94624e-20 7.19854e-24 -1.94552e-20 0.00139591 0.997816 8.59844e-05 0.152659 2.85235 0.00139591 0.997817 0.751901 0.00105936 0.00188068 0.000859844 0.455494 0.00188068 0.441667 0.000130002 1.02 0.888239 0.534524 0.286828 1.71816e-07 3.07324e-09 2378.75 3117.97 -0.0559761 0.482172 0.27741 0.253425 -0.593339 -0.169543 0.494755 -0.266803 -0.227962 2.179 1 0 297.337 0 2.16731 2.177 0.000299599 0.855504 0.67915 0.340962 0.423213 2.1675 135.544 83.8917 18.7192 60.8524 0.0040265 0 -40 10
1.278 3.6999e-08 2.5393e-06 0.128025 0.128024 0.012033 1.68177e-05 0.00115423 0.160031 0.000658461 0.160685 0.910364 101.691 0.239929 0.793342 4.30943 0.0600714 0.040655 0.959345 0.0196696 0.0044081 0.0189316 0.00422315 0.0053304 0.00606841 0.213216 0.242737 58.0193 -87.8974 126.245 15.9529 145.026 0.000141331 0.267224 192.805 0.310396 0.06735 0.00409704 0.00056206 0.00138406 0.986973 0.991724 -2.98299e-06 -85.6615 0.0930438 31179.7 305.025 0.983507 0.319146 0.733153 0.733149 9.99958 2.9841e-06 1.19363e-05 0.132329 0.983084 0.931726 -0.0132923 4.91645e-06 0.507822 -1.94636e-20 7.19903e-24 -1.94564e-20 0.00139591 0.997816 8.59845e-05 0.152659 2.85235 0.00139591 0.997817 0.751988 0.00105938 0.00188068 0.000859845 0.455494 0.00188068 0.441673 0.000130005 1.02 0.88824 0.534524 0.286829 1.71816e-07 3.07326e-09 2378.73 3118 -0.0559796 0.482172 0.27741 0.253427 -0.593339 -0.169543 0.494744 -0.266801 -0.227953 2.18 1 0 297.334 0 2.16745 2.178 0.000299599 0.855521 0.679195 0.340892 0.423237 2.16764 135.551 83.8913 18.7192 60.8522 0.00402651 0 -40 10
1.279 3.70278e-08 2.5393e-06 0.128073 0.128072 0.0120329 1.68308e-05 0.00115423 0.160092 0.000658462 0.160746 0.910445 101.69 0.239919 0.793463 4.30983 0.0600811 0.0406588 0.959341 0.0196692 0.00440844 0.0189312 0.00422343 0.00533082 0.00606883 0.213233 0.242753 58.0193 -87.8974 126.245 15.9529 145.026 0.000141332 0.267224 192.805 0.310395 0.06735 0.00409704 0.000562061 0.00138406 0.986973 0.991724 -2.983e-06 -85.6615 0.0930439 31179.7 305.034 0.983507 0.319146 0.73316 0.733156 9.99958 2.98411e-06 1.19363e-05 0.132332 0.983085 0.931725 -0.0132923 4.91648e-06 0.507837 -1.94648e-20 7.19952e-24 -1.94576e-20 0.00139591 0.997816 8.59845e-05 0.152659 2.85235 0.00139591 0.997817 0.752074 0.00105939 0.00188068 0.000859845 0.455494 0.00188068 0.44168 0.000130008 1.02 0.888242 0.534523 0.286831 1.71817e-07 3.07329e-09 2378.71 3118.03 -0.055983 0.482172 0.277409 0.253429 -0.593338 -0.169543 0.494733 -0.266799 -0.227943 2.181 1 0 297.331 0 2.16759 2.179 0.000299598 0.855538 0.67924 0.340822 0.42326 2.16779 135.559 83.891 18.7192 60.8521 0.00402652 0 -40 10
1.28 3.70567e-08 2.5393e-06 0.128122 0.128121 0.0120329 1.6844e-05 0.00115423 0.160152 0.000658463 0.160806 0.910526 101.69 0.239909 0.793584 4.31024 0.0600908 0.0406627 0.959337 0.0196688 0.00440877 0.0189307 0.00422372 0.00533123 0.00606925 0.213249 0.24277 58.0194 -87.8974 126.245 15.9528 145.026 0.000141333 0.267225 192.805 0.310395 0.0673499 0.00409705 0.000562062 0.00138407 0.986973 0.991724 -2.98302e-06 -85.6615 0.093044 31179.7 305.043 0.983507 0.319146 0.733167 0.733163 9.99958 2.98411e-06 1.19363e-05 0.132336 0.983087 0.931725 -0.0132923 4.91651e-06 0.507851 -1.9466e-20 7.20001e-24 -1.94588e-20 0.00139591 0.997816 8.59846e-05 0.152659 2.85235 0.00139591 0.997817 0.75216 0.00105941 0.00188069 0.000859846 0.455494 0.00188068 0.441686 0.00013001 1.02 0.888243 0.534523 0.286832 1.71817e-07 3.07331e-09 2378.7 3118.06 -0.0559865 0.482172 0.277409 0.25343 -0.593338 -0.169543 0.494721 -0.266797 -0.227934 2.182 1 0 297.328 0 2.16774 2.18 0.000299597 0.855556 0.679285 0.340752 0.423284 2.16793 135.567 83.8906 18.7192 60.8519 0.00402654 0 -40 10
1.281 3.70856e-08 2.5393e-06 0.12817 0.128169 0.0120329 1.68571e-05 0.00115423 0.160213 0.000658464 0.160867 0.910606 101.689 0.239899 0.793705 4.31065 0.0601005 0.0406665 0.959333 0.0196684 0.00440911 0.0189303 0.00422401 0.00533165 0.00606967 0.213266 0.242787 58.0195 -87.8974 126.245 15.9528 145.026 0.000141335 0.267225 192.805 0.310394 0.0673499 0.00409705 0.000562062 0.00138407 0.986973 0.991724 -2.98304e-06 -85.6615 0.093044 31179.6 305.052 0.983507 0.319146 0.733174 0.73317 9.99958 2.98412e-06 1.19364e-05 0.132339 0.983088 0.931724 -0.0132923 4.91654e-06 0.507866 -1.94672e-20 7.2005e-24 -1.946e-20 0.00139592 0.997816 8.59847e-05 0.152659 2.85235 0.00139592 0.997817 0.752246 0.00105943 0.00188069 0.000859847 0.455494 0.00188069 0.441693 0.000130013 1.02 0.888244 0.534523 0.286834 1.71817e-07 3.07333e-09 2378.68 3118.09 -0.05599 0.482172 0.277409 0.253432 -0.593337 -0.169543 0.49471 -0.266794 -0.227925 2.183 1 0 297.325 0 2.16788 2.181 0.000299596 0.855573 0.679331 0.340683 0.423308 2.16808 135.575 83.8903 18.7191 60.8517 0.00402655 0 -40 10
1.282 3.71145e-08 2.5393e-06 0.128219 0.128218 0.0120329 1.68702e-05 0.00115423 0.160273 0.000658465 0.160927 0.910687 101.689 0.23989 0.793827 4.31106 0.0601103 0.0406704 0.95933 0.0196679 0.00440945 0.0189299 0.00422429 0.00533206 0.0060701 0.213283 0.242804 58.0195 -87.8974 126.245 15.9527 145.026 0.000141336 0.267225 192.805 0.310394 0.0673498 0.00409705 0.000562063 0.00138407 0.986973 0.991724 -2.98305e-06 -85.6615 0.0930441 31179.6 305.061 0.983507 0.319146 0.733181 0.733177 9.99958 2.98412e-06 1.19364e-05 0.132343 0.983089 0.931724 -0.0132923 4.91657e-06 0.50788 -1.94684e-20 7.20099e-24 -1.94612e-20 0.00139592 0.997816 8.59848e-05 0.152659 2.85235 0.00139592 0.997817 0.752332 0.00105945 0.00188069 0.000859848 0.455493 0.00188069 0.441699 0.000130016 1.02 0.888245 0.534522 0.286835 1.71818e-07 3.07336e-09 2378.66 3118.12 -0.0559935 0.482172 0.277409 0.253434 -0.593337 -0.169544 0.494699 -0.266792 -0.227916 2.184 1 0 297.322 0 2.16803 2.182 0.000299595 0.85559 0.679376 0.340613 0.423331 2.16822 135.582 83.8899 18.7191 60.8515 0.00402657 0 -40 10
1.283 3.71434e-08 2.5393e-06 0.128267 0.128266 0.0120329 1.68834e-05 0.00115423 0.160334 0.000658466 0.160987 0.910768 101.689 0.23988 0.793948 4.31147 0.06012 0.0406742 0.959326 0.0196675 0.00440979 0.0189295 0.00422458 0.00533248 0.00607052 0.213299 0.242821 58.0196 -87.8974 126.244 15.9527 145.026 0.000141338 0.267225 192.804 0.310394 0.0673498 0.00409706 0.000562064 0.00138407 0.986972 0.991724 -2.98307e-06 -85.6615 0.0930442 31179.6 305.071 0.983507 0.319146 0.733188 0.733184 9.99958 2.98413e-06 1.19364e-05 0.132346 0.983091 0.931724 -0.0132923 4.9166e-06 0.507894 -1.94696e-20 7.20148e-24 -1.94624e-20 0.00139592 0.997816 8.59849e-05 0.15266 2.85235 0.00139592 0.997817 0.752418 0.00105947 0.00188069 0.000859849 0.455493 0.00188069 0.441706 0.000130019 1.02 0.888246 0.534522 0.286837 1.71818e-07 3.07338e-09 2378.65 3118.15 -0.055997 0.482172 0.277408 0.253436 -0.593337 -0.169544 0.494687 -0.26679 -0.227906 2.185 1 0 297.319 0 2.16817 2.183 0.000299595 0.855607 0.679421 0.340543 0.423355 2.16836 135.59 83.8896 18.7191 60.8514 0.00402658 0 -40 10
1.284 3.71723e-08 2.53931e-06 0.128315 0.128314 0.0120329 1.68965e-05 0.00115423 0.160394 0.000658467 0.161048 0.910849 101.688 0.23987 0.794069 4.31188 0.0601297 0.0406781 0.959322 0.0196671 0.00441012 0.0189291 0.00422487 0.00533289 0.00607094 0.213316 0.242838 58.0196 -87.8974 126.244 15.9527 145.026 0.000141339 0.267225 192.804 0.310393 0.0673497 0.00409706 0.000562064 0.00138408 0.986972 0.991724 -2.98308e-06 -85.6614 0.0930443 31179.6 305.08 0.983507 0.319146 0.733196 0.733191 9.99958 2.98413e-06 1.19364e-05 0.13235 0.983092 0.931723 -0.0132923 4.91663e-06 0.507909 -1.94708e-20 7.20197e-24 -1.94636e-20 0.00139592 0.997816 8.59849e-05 0.15266 2.85236 0.00139592 0.997817 0.752504 0.00105948 0.00188069 0.000859849 0.455493 0.00188069 0.441713 0.000130022 1.02 0.888247 0.534522 0.286838 1.71818e-07 3.0734e-09 2378.63 3118.18 -0.0560005 0.482172 0.277408 0.253438 -0.593336 -0.169544 0.494676 -0.266788 -0.227897 2.186 1 0 297.316 0 2.16831 2.184 0.000299594 0.855625 0.679466 0.340474 0.423379 2.16851 135.598 83.8892 18.7191 60.8512 0.0040266 0 -40 10
1.285 3.72012e-08 2.53931e-06 0.128363 0.128362 0.0120329 1.69096e-05 0.00115423 0.160454 0.000658468 0.161108 0.91093 101.688 0.239861 0.79419 4.31229 0.0601395 0.040682 0.959318 0.0196667 0.00441046 0.0189286 0.00422516 0.00533331 0.00607136 0.213332 0.242854 58.0197 -87.8974 126.244 15.9526 145.026 0.00014134 0.267226 192.804 0.310393 0.0673497 0.00409706 0.000562065 0.00138408 0.986972 0.991724 -2.9831e-06 -85.6614 0.0930444 31179.6 305.089 0.983507 0.319146 0.733203 0.733198 9.99958 2.98414e-06 1.19364e-05 0.132353 0.983093 0.931723 -0.0132923 4.91666e-06 0.507923 -1.9472e-20 7.20246e-24 -1.94648e-20 0.00139592 0.997816 8.5985e-05 0.15266 2.85236 0.00139592 0.997817 0.75259 0.0010595 0.00188069 0.00085985 0.455493 0.00188069 0.441719 0.000130024 1.02 0.888248 0.534521 0.28684 1.71818e-07 3.07343e-09 2378.61 3118.21 -0.056004 0.482172 0.277408 0.25344 -0.593336 -0.169544 0.494664 -0.266786 -0.227888 2.187 1 0 297.313 0 2.16846 2.185 0.000299593 0.855642 0.679511 0.340405 0.423403 2.16865 135.606 83.8889 18.7191 60.851 0.00402661 0 -40 10
1.286 3.72301e-08 2.53931e-06 0.128411 0.12841 0.0120328 1.69228e-05 0.00115423 0.160514 0.00065847 0.161168 0.91101 101.687 0.239851 0.794312 4.3127 0.0601492 0.0406859 0.959314 0.0196663 0.0044108 0.0189282 0.00422545 0.00533373 0.00607178 0.213349 0.242871 58.0198 -87.8974 126.244 15.9526 145.026 0.000141342 0.267226 192.804 0.310392 0.0673496 0.00409706 0.000562066 0.00138408 0.986972 0.991724 -2.98311e-06 -85.6614 0.0930445 31179.5 305.098 0.983507 0.319146 0.73321 0.733206 9.99958 2.98414e-06 1.19365e-05 0.132356 0.983095 0.931722 -0.0132923 4.91669e-06 0.507938 -1.94732e-20 7.20295e-24 -1.9466e-20 0.00139592 0.997816 8.59851e-05 0.15266 2.85236 0.00139592 0.997817 0.752676 0.00105952 0.00188069 0.000859851 0.455492 0.00188069 0.441726 0.000130027 1.02 0.888249 0.534521 0.286841 1.71819e-07 3.07345e-09 2378.6 3118.24 -0.0560076 0.482172 0.277407 0.253442 -0.593335 -0.169544 0.494653 -0.266784 -0.227878 2.188 1 0 297.31 0 2.1686 2.186 0.000299592 0.85566 0.679556 0.340335 0.423426 2.1688 135.613 83.8885 18.719 60.8509 0.00402663 0 -40 10
1.287 3.7259e-08 2.53931e-06 0.12846 0.128459 0.0120328 1.69359e-05 0.00115423 0.160574 0.000658471 0.161228 0.911091 101.687 0.239841 0.794433 4.31311 0.0601589 0.0406897 0.95931 0.0196659 0.00441114 0.0189278 0.00422573 0.00533414 0.00607221 0.213366 0.242888 58.0198 -87.8974 126.244 15.9526 145.026 0.000141343 0.267226 192.804 0.310392 0.0673496 0.00409707 0.000562066 0.00138408 0.986972 0.991724 -2.98313e-06 -85.6614 0.0930446 31179.5 305.107 0.983507 0.319146 0.733217 0.733213 9.99958 2.98415e-06 1.19365e-05 0.13236 0.983096 0.931722 -0.0132923 4.91671e-06 0.507952 -1.94744e-20 7.20344e-24 -1.94672e-20 0.00139592 0.997816 8.59852e-05 0.15266 2.85236 0.00139592 0.997817 0.752762 0.00105954 0.0018807 0.000859852 0.455492 0.00188069 0.441732 0.00013003 1.02 0.88825 0.534521 0.286843 1.71819e-07 3.07347e-09 2378.58 3118.27 -0.0560111 0.482172 0.277407 0.253444 -0.593335 -0.169544 0.494641 -0.266782 -0.227869 2.189 1 0 297.307 0 2.16875 2.187 0.000299592 0.855677 0.679602 0.340266 0.42345 2.16894 135.621 83.8881 18.719 60.8507 0.00402664 0 -40 10
1.288 3.72878e-08 2.53931e-06 0.128508 0.128507 0.0120328 1.6949e-05 0.00115423 0.160634 0.000658472 0.161288 0.911172 101.686 0.239831 0.794554 4.31352 0.0601687 0.0406936 0.959306 0.0196654 0.00441148 0.0189274 0.00422602 0.00533456 0.00607263 0.213382 0.242905 58.0199 -87.8974 126.244 15.9525 145.026 0.000141344 0.267226 192.804 0.310391 0.0673495 0.00409707 0.000562067 0.00138408 0.986972 0.991724 -2.98314e-06 -85.6614 0.0930447 31179.5 305.116 0.983507 0.319146 0.733224 0.73322 9.99958 2.98415e-06 1.19365e-05 0.132363 0.983097 0.931722 -0.0132923 4.91674e-06 0.507967 -1.94756e-20 7.20393e-24 -1.94684e-20 0.00139592 0.997816 8.59853e-05 0.15266 2.85236 0.00139592 0.997817 0.752848 0.00105955 0.0018807 0.000859853 0.455492 0.0018807 0.441739 0.000130033 1.02 0.888251 0.53452 0.286844 1.71819e-07 3.07349e-09 2378.56 3118.3 -0.0560146 0.482173 0.277407 0.253446 -0.593335 -0.169544 0.49463 -0.26678 -0.227859 2.19 1 0 297.304 0 2.16889 2.188 0.000299591 0.855695 0.679647 0.340197 0.423474 2.16909 135.629 83.8878 18.719 60.8505 0.00402665 0 -40 10
1.289 3.73167e-08 2.53931e-06 0.128556 0.128555 0.0120328 1.69622e-05 0.00115423 0.160695 0.000658473 0.161348 0.911253 101.686 0.239822 0.794676 4.31394 0.0601784 0.0406975 0.959302 0.019665 0.00441182 0.0189269 0.00422631 0.00533498 0.00607305 0.213399 0.242922 58.02 -87.8974 126.244 15.9525 145.026 0.000141346 0.267226 192.803 0.310391 0.0673494 0.00409707 0.000562068 0.00138409 0.986972 0.991724 -2.98316e-06 -85.6614 0.0930447 31179.5 305.126 0.983507 0.319146 0.733232 0.733227 9.99958 2.98416e-06 1.19365e-05 0.132367 0.983098 0.931721 -0.0132923 4.91677e-06 0.507981 -1.94768e-20 7.20442e-24 -1.94696e-20 0.00139592 0.997816 8.59854e-05 0.15266 2.85236 0.00139592 0.997817 0.752934 0.00105957 0.0018807 0.000859854 0.455492 0.0018807 0.441745 0.000130036 1.02 0.888253 0.53452 0.286846 1.71819e-07 3.07352e-09 2378.55 3118.33 -0.0560182 0.482173 0.277407 0.253448 -0.593334 -0.169544 0.494618 -0.266778 -0.22785 2.191 1 0 297.301 0 2.16904 2.189 0.00029959 0.855712 0.679692 0.340128 0.423497 2.16923 135.636 83.8874 18.719 60.8504 0.00402667 0 -40 10
1.29 3.73456e-08 2.53931e-06 0.128604 0.128603 0.0120328 1.69753e-05 0.00115423 0.160755 0.000658474 0.161408 0.911334 101.686 0.239812 0.794797 4.31435 0.0601882 0.0407014 0.959299 0.0196646 0.00441216 0.0189265 0.0042266 0.0053354 0.00607348 0.213416 0.242939 58.02 -87.8974 126.244 15.9524 145.026 0.000141347 0.267227 192.803 0.310391 0.0673494 0.00409708 0.000562068 0.00138409 0.986972 0.991724 -2.98317e-06 -85.6614 0.0930448 31179.4 305.135 0.983507 0.319146 0.733239 0.733235 9.99958 2.98416e-06 1.19365e-05 0.13237 0.9831 0.931721 -0.0132923 4.9168e-06 0.507996 -1.9478e-20 7.20491e-24 -1.94708e-20 0.00139593 0.997816 8.59854e-05 0.152661 2.85236 0.00139593 0.997817 0.75302 0.00105959 0.0018807 0.000859854 0.455492 0.0018807 0.441752 0.000130038 1.02 0.888254 0.53452 0.286847 1.7182e-07 3.07354e-09 2378.53 3118.36 -0.0560217 0.482173 0.277406 0.25345 -0.593334 -0.169544 0.494607 -0.266775 -0.227841 2.192 1 0 297.297 0 2.16918 2.19 0.000299589 0.85573 0.679737 0.340059 0.423521 2.16937 135.644 83.8871 18.719 60.8502 0.00402668 0 -40 10
1.291 3.73745e-08 2.53931e-06 0.128652 0.128651 0.0120328 1.69884e-05 0.00115423 0.160814 0.000658475 0.161468 0.911415 101.685 0.239802 0.794919 4.31476 0.060198 0.0407053 0.959295 0.0196642 0.0044125 0.0189261 0.00422689 0.00533582 0.0060739 0.213433 0.242956 58.0201 -87.8974 126.243 15.9524 145.026 0.000141349 0.267227 192.803 0.31039 0.0673493 0.00409708 0.000562069 0.00138409 0.986972 0.991724 -2.98319e-06 -85.6614 0.0930449 31179.4 305.144 0.983507 0.319146 0.733246 0.733242 9.99958 2.98417e-06 1.19366e-05 0.132374 0.983101 0.93172 -0.0132923 4.91683e-06 0.50801 -1.94792e-20 7.20541e-24 -1.9472e-20 0.00139593 0.997816 8.59855e-05 0.152661 2.85236 0.00139593 0.997817 0.753105 0.00105961 0.0018807 0.000859855 0.455491 0.0018807 0.441758 0.000130041 1.02 0.888255 0.53452 0.286849 1.7182e-07 3.07356e-09 2378.51 3118.39 -0.0560253 0.482173 0.277406 0.253452 -0.593333 -0.169544 0.494595 -0.266773 -0.227831 2.193 1 0 297.294 0 2.16932 2.191 0.000299588 0.855747 0.679782 0.339991 0.423545 2.16952 135.652 83.8867 18.7189 60.85 0.0040267 0 -40 10
1.292 3.74034e-08 2.53931e-06 0.1287 0.128699 0.0120328 1.70015e-05 0.00115423 0.160874 0.000658476 0.161528 0.911496 101.685 0.239792 0.79504 4.31518 0.0602077 0.0407092 0.959291 0.0196638 0.00441284 0.0189257 0.00422718 0.00533623 0.00607432 0.213449 0.242973 58.0201 -87.8974 126.243 15.9524 145.026 0.00014135 0.267227 192.803 0.31039 0.0673493 0.00409708 0.00056207 0.00138409 0.986972 0.991724 -2.9832e-06 -85.6614 0.093045 31179.4 305.153 0.983507 0.319146 0.733253 0.733249 9.99958 2.98417e-06 1.19366e-05 0.132377 0.983102 0.93172 -0.0132923 4.91686e-06 0.508025 -1.94805e-20 7.2059e-24 -1.94732e-20 0.00139593 0.997816 8.59856e-05 0.152661 2.85236 0.00139593 0.997817 0.753191 0.00105963 0.0018807 0.000859856 0.455491 0.0018807 0.441765 0.000130044 1.02 0.888256 0.534519 0.28685 1.7182e-07 3.07359e-09 2378.5 3118.42 -0.0560288 0.482173 0.277406 0.253454 -0.593333 -0.169544 0.494583 -0.266771 -0.227822 2.194 1 0 297.291 0 2.16947 2.192 0.000299588 0.855765 0.679827 0.339922 0.423568 2.16966 135.66 83.8863 18.7189 60.8498 0.00402671 0 -40 10
1.293 3.74323e-08 2.53931e-06 0.128747 0.128746 0.0120328 1.70147e-05 0.00115423 0.160934 0.000658477 0.161588 0.911577 101.684 0.239783 0.795162 4.31559 0.0602175 0.0407131 0.959287 0.0196633 0.00441318 0.0189253 0.00422747 0.00533665 0.00607475 0.213466 0.24299 58.0202 -87.8974 126.243 15.9523 145.026 0.000141351 0.267227 192.803 0.310389 0.0673492 0.00409709 0.00056207 0.0013841 0.986972 0.991724 -2.98322e-06 -85.6614 0.0930451 31179.4 305.163 0.983507 0.319146 0.733261 0.733256 9.99958 2.98418e-06 1.19366e-05 0.132381 0.983104 0.93172 -0.0132923 4.91689e-06 0.508039 -1.94817e-20 7.20639e-24 -1.94745e-20 0.00139593 0.997816 8.59857e-05 0.152661 2.85236 0.00139593 0.997817 0.753277 0.00105964 0.0018807 0.000859857 0.455491 0.0018807 0.441771 0.000130047 1.02 0.888257 0.534519 0.286852 1.7182e-07 3.07361e-09 2378.48 3118.45 -0.0560324 0.482173 0.277405 0.253456 -0.593333 -0.169544 0.494572 -0.266769 -0.227812 2.195 1 0 297.288 0 2.16961 2.193 0.000299587 0.855783 0.679872 0.339853 0.423592 2.16981 135.667 83.886 18.7189 60.8497 0.00402673 0 -40 10
1.294 3.74612e-08 2.53932e-06 0.128795 0.128794 0.0120327 1.70278e-05 0.00115423 0.160994 0.000658478 0.161648 0.911658 101.684 0.239773 0.795284 4.31601 0.0602272 0.040717 0.959283 0.0196629 0.00441352 0.0189248 0.00422776 0.00533707 0.00607517 0.213483 0.243007 58.0203 -87.8974 126.243 15.9523 145.027 0.000141353 0.267227 192.803 0.310389 0.0673492 0.00409709 0.000562071 0.0013841 0.986972 0.991724 -2.98323e-06 -85.6613 0.0930452 31179.3 305.172 0.983507 0.319146 0.733268 0.733264 9.99958 2.98418e-06 1.19366e-05 0.132384 0.983105 0.931719 -0.0132923 4.91692e-06 0.508054 -1.94829e-20 7.20689e-24 -1.94757e-20 0.00139593 0.997816 8.59858e-05 0.152661 2.85236 0.00139593 0.997817 0.753363 0.00105966 0.00188071 0.000859858 0.455491 0.0018807 0.441778 0.00013005 1.02 0.888258 0.534519 0.286854 1.71821e-07 3.07363e-09 2378.46 3118.48 -0.056036 0.482173 0.277405 0.253458 -0.593332 -0.169544 0.49456 -0.266767 -0.227803 2.196 1 0 297.285 0 2.16976 2.194 0.000299586 0.8558 0.679917 0.339785 0.423616 2.16995 135.675 83.8856 18.7189 60.8495 0.00402674 0 -40 10
1.295 3.74901e-08 2.53932e-06 0.128843 0.128842 0.0120327 1.70409e-05 0.00115423 0.161054 0.000658479 0.161708 0.91174 101.684 0.239763 0.795405 4.31642 0.060237 0.0407209 0.959279 0.0196625 0.00441386 0.0189244 0.00422805 0.00533749 0.0060756 0.2135 0.243024 58.0203 -87.8974 126.243 15.9522 145.027 0.000141354 0.267228 192.802 0.310388 0.0673491 0.00409709 0.000562072 0.0013841 0.986972 0.991724 -2.98325e-06 -85.6613 0.0930453 31179.3 305.181 0.983507 0.319146 0.733275 0.733271 9.99958 2.98419e-06 1.19366e-05 0.132388 0.983106 0.931719 -0.0132923 4.91695e-06 0.508068 -1.94841e-20 7.20738e-24 -1.94769e-20 0.00139593 0.997816 8.59858e-05 0.152661 2.85237 0.00139593 0.997817 0.753448 0.00105968 0.00188071 0.000859858 0.45549 0.00188071 0.441785 0.000130052 1.02 0.888259 0.534518 0.286855 1.71821e-07 3.07365e-09 2378.45 3118.51 -0.0560395 0.482173 0.277405 0.25346 -0.593332 -0.169544 0.494549 -0.266765 -0.227793 2.197 1 0 297.282 0 2.1699 2.195 0.000299585 0.855818 0.679962 0.339717 0.423639 2.17009 135.683 83.8853 18.7189 60.8493 0.00402676 0 -40 10
1.296 3.75189e-08 2.53932e-06 0.128891 0.12889 0.0120327 1.70541e-05 0.00115424 0.161114 0.000658479 0.161767 0.911821 101.683 0.239753 0.795527 4.31684 0.0602468 0.0407249 0.959275 0.0196621 0.0044142 0.018924 0.00422834 0.00533791 0.00607603 0.213516 0.243041 58.0204 -87.8974 126.243 15.9522 145.027 0.000141356 0.267228 192.802 0.310388 0.0673491 0.00409709 0.000562072 0.0013841 0.986972 0.991724 -2.98326e-06 -85.6613 0.0930454 31179.3 305.19 0.983507 0.319146 0.733283 0.733278 9.99958 2.98419e-06 1.19367e-05 0.132391 0.983107 0.931718 -0.0132923 4.91698e-06 0.508083 -1.94853e-20 7.20787e-24 -1.94781e-20 0.00139593 0.997816 8.59859e-05 0.152662 2.85237 0.00139593 0.997817 0.753534 0.0010597 0.00188071 0.000859859 0.45549 0.00188071 0.441791 0.000130055 1.02 0.88826 0.534518 0.286857 1.71821e-07 3.07368e-09 2378.43 3118.54 -0.0560431 0.482173 0.277405 0.253462 -0.593331 -0.169544 0.494537 -0.266763 -0.227783 2.198 1 0 297.279 0 2.17004 2.196 0.000299584 0.855836 0.680008 0.339648 0.423663 2.17024 135.691 83.8849 18.7188 60.8491 0.00402677 0 -40 10
1.297 3.75478e-08 2.53932e-06 0.128939 0.128938 0.0120327 1.70672e-05 0.00115424 0.161173 0.00065848 0.161827 0.911902 101.683 0.239743 0.795649 4.31725 0.0602565 0.0407288 0.959271 0.0196617 0.00441454 0.0189235 0.00422863 0.00533833 0.00607645 0.213533 0.243058 58.0205 -87.8974 126.243 15.9522 145.027 0.000141357 0.267228 192.802 0.310388 0.067349 0.0040971 0.000562073 0.0013841 0.986972 0.991724 -2.98328e-06 -85.6613 0.0930454 31179.3 305.2 0.983507 0.319146 0.73329 0.733286 9.99958 2.9842e-06 1.19367e-05 0.132395 0.983109 0.931718 -0.0132923 4.91701e-06 0.508098 -1.94865e-20 7.20837e-24 -1.94793e-20 0.00139593 0.997816 8.5986e-05 0.152662 2.85237 0.00139593 0.997817 0.75362 0.00105971 0.00188071 0.00085986 0.45549 0.00188071 0.441798 0.000130058 1.02 0.888261 0.534518 0.286858 1.71822e-07 3.0737e-09 2378.41 3118.57 -0.0560467 0.482173 0.277404 0.253464 -0.593331 -0.169545 0.494525 -0.266761 -0.227774 2.199 1 0 297.276 0 2.17019 2.197 0.000299583 0.855854 0.680053 0.33958 0.423687 2.17038 135.698 83.8845 18.7188 60.849 0.00402679 0 -40 10
1.298 3.75767e-08 2.53932e-06 0.128986 0.128985 0.0120327 1.70803e-05 0.00115424 0.161233 0.000658481 0.161887 0.911983 101.682 0.239734 0.79577 4.31767 0.0602663 0.0407327 0.959267 0.0196612 0.00441488 0.0189231 0.00422892 0.00533875 0.00607688 0.21355 0.243075 58.0205 -87.8974 126.242 15.9521 145.027 0.000141359 0.267228 192.802 0.310387 0.067349 0.0040971 0.000562074 0.00138411 0.986972 0.991724 -2.98329e-06 -85.6613 0.0930455 31179.3 305.209 0.983507 0.319146 0.733298 0.733293 9.99958 2.9842e-06 1.19367e-05 0.132398 0.98311 0.931717 -0.0132923 4.91704e-06 0.508112 -1.94877e-20 7.20886e-24 -1.94805e-20 0.00139593 0.997816 8.59861e-05 0.152662 2.85237 0.00139593 0.997817 0.753705 0.00105973 0.00188071 0.000859861 0.45549 0.00188071 0.441804 0.000130061 1.02 0.888262 0.534517 0.28686 1.71822e-07 3.07372e-09 2378.4 3118.6 -0.0560503 0.482173 0.277404 0.253466 -0.593331 -0.169545 0.494513 -0.266759 -0.227764 2.2 1 0 297.272 0 2.17033 2.198 0.000299583 0.855872 0.680098 0.339512 0.42371 2.17052 135.706 83.8842 18.7188 60.8488 0.0040268 0 -40 10
1.299 3.76056e-08 2.53932e-06 0.129034 0.129033 0.0120327 1.70935e-05 0.00115424 0.161292 0.000658482 0.161946 0.912064 101.682 0.239724 0.795892 4.31808 0.0602761 0.0407366 0.959263 0.0196608 0.00441523 0.0189227 0.00422921 0.00533917 0.00607731 0.213567 0.243092 58.0206 -87.8974 126.242 15.9521 145.027 0.00014136 0.267228 192.802 0.310387 0.0673489 0.0040971 0.000562074 0.00138411 0.986972 0.991724 -2.98331e-06 -85.6613 0.0930456 31179.2 305.218 0.983507 0.319146 0.733305 0.733301 9.99958 2.98421e-06 1.19367e-05 0.132402 0.983111 0.931717 -0.0132923 4.91707e-06 0.508127 -1.9489e-20 7.20936e-24 -1.94818e-20 0.00139594 0.997816 8.59862e-05 0.152662 2.85237 0.00139594 0.997817 0.753791 0.00105975 0.00188071 0.000859862 0.455489 0.00188071 0.441811 0.000130064 1.02 0.888264 0.534517 0.286861 1.71822e-07 3.07375e-09 2378.38 3118.64 -0.0560539 0.482173 0.277404 0.253468 -0.59333 -0.169545 0.494502 -0.266756 -0.227755 2.201 1 0 297.269 0 2.17047 2.199 0.000299582 0.85589 0.680143 0.339444 0.423734 2.17067 135.714 83.8838 18.7188 60.8486 0.00402682 0 -40 10
1.3 3.76345e-08 2.53932e-06 0.129082 0.129081 0.0120327 1.71066e-05 0.00115424 0.161352 0.000658483 0.162006 0.912146 101.681 0.239714 0.796014 4.3185 0.0602859 0.0407406 0.959259 0.0196604 0.00441557 0.0189223 0.00422951 0.0053396 0.00607773 0.213584 0.243109 58.0207 -87.8974 126.242 15.9521 145.027 0.000141361 0.267229 192.802 0.310386 0.0673489 0.00409711 0.000562075 0.00138411 0.986972 0.991724 -2.98332e-06 -85.6613 0.0930457 31179.2 305.227 0.983507 0.319146 0.733313 0.733308 9.99958 2.98421e-06 1.19367e-05 0.132405 0.983112 0.931717 -0.0132923 4.9171e-06 0.508142 -1.94902e-20 7.20985e-24 -1.9483e-20 0.00139594 0.997816 8.59862e-05 0.152662 2.85237 0.00139594 0.997817 0.753876 0.00105977 0.00188071 0.000859862 0.455489 0.00188071 0.441817 0.000130066 1.02 0.888265 0.534517 0.286863 1.71822e-07 3.07377e-09 2378.36 3118.67 -0.0560575 0.482173 0.277403 0.25347 -0.59333 -0.169545 0.49449 -0.266754 -0.227745 2.202 1 0 297.266 0 2.17062 2.2 0.000299581 0.855908 0.680188 0.339376 0.423758 2.17081 135.721 83.8834 18.7187 60.8484 0.00402683 0 -40 10
1.301 3.76634e-08 2.53932e-06 0.129129 0.129128 0.0120326 1.71197e-05 0.00115424 0.161411 0.000658484 0.162065 0.912227 101.681 0.239704 0.796136 4.31892 0.0602957 0.0407445 0.959255 0.01966 0.00441591 0.0189218 0.0042298 0.00534002 0.00607816 0.213601 0.243126 58.0207 -87.8974 126.242 15.952 145.027 0.000141363 0.267229 192.801 0.310386 0.0673488 0.00409711 0.000562076 0.00138411 0.986972 0.991724 -2.98334e-06 -85.6613 0.0930458 31179.2 305.237 0.983507 0.319146 0.73332 0.733316 9.99958 2.98422e-06 1.19368e-05 0.132409 0.983114 0.931716 -0.0132923 4.91713e-06 0.508156 -1.94914e-20 7.21035e-24 -1.94842e-20 0.00139594 0.997816 8.59863e-05 0.152662 2.85237 0.00139594 0.997817 0.753962 0.00105979 0.00188072 0.000859863 0.455489 0.00188072 0.441824 0.000130069 1.02 0.888266 0.534516 0.286864 1.71823e-07 3.07379e-09 2378.35 3118.7 -0.0560612 0.482174 0.277403 0.253472 -0.593329 -0.169545 0.494478 -0.266752 -0.227735 2.203 1 0 297.263 0 2.17076 2.201 0.00029958 0.855926 0.680233 0.339309 0.423781 2.17096 135.729 83.8831 18.7187 60.8482 0.00402685 0 -40 10
1.302 3.76923e-08 2.53932e-06 0.129177 0.129176 0.0120326 1.71329e-05 0.00115424 0.161471 0.000658485 0.162125 0.912308 101.681 0.239695 0.796258 4.31934 0.0603055 0.0407485 0.959252 0.0196596 0.00441625 0.0189214 0.00423009 0.00534044 0.00607859 0.213618 0.243144 58.0208 -87.8975 126.242 15.952 145.027 0.000141364 0.267229 192.801 0.310385 0.0673488 0.00409711 0.000562076 0.00138411 0.986972 0.991724 -2.98335e-06 -85.6613 0.0930459 31179.2 305.246 0.983507 0.319146 0.733328 0.733323 9.99958 2.98422e-06 1.19368e-05 0.132412 0.983115 0.931716 -0.0132923 4.91716e-06 0.508171 -1.94926e-20 7.21084e-24 -1.94854e-20 0.00139594 0.997816 8.59864e-05 0.152662 2.85237 0.00139594 0.997817 0.754047 0.0010598 0.00188072 0.000859864 0.455489 0.00188072 0.44183 0.000130072 1.02 0.888267 0.534516 0.286866 1.71823e-07 3.07381e-09 2378.33 3118.73 -0.0560648 0.482174 0.277403 0.253474 -0.593329 -0.169545 0.494466 -0.26675 -0.227726 2.204 1 0 297.26 0 2.17091 2.202 0.000299579 0.855944 0.680278 0.339241 0.423805 2.1711 135.737 83.8827 18.7187 60.8481 0.00402686 0 -40 10
1.303 3.77212e-08 2.53932e-06 0.129224 0.129223 0.0120326 1.7146e-05 0.00115424 0.16153 0.000658486 0.162184 0.912389 101.68 0.239685 0.79638 4.31976 0.0603153 0.0407524 0.959248 0.0196591 0.0044166 0.018921 0.00423038 0.00534086 0.00607902 0.213634 0.243161 58.0208 -87.8975 126.242 15.9519 145.027 0.000141366 0.267229 192.801 0.310385 0.0673487 0.00409712 0.000562077 0.00138412 0.986972 0.991724 -2.98337e-06 -85.6613 0.093046 31179.1 305.255 0.983507 0.319146 0.733335 0.733331 9.99958 2.98423e-06 1.19368e-05 0.132416 0.983116 0.931715 -0.0132923 4.91719e-06 0.508186 -1.94938e-20 7.21134e-24 -1.94866e-20 0.00139594 0.997816 8.59865e-05 0.152663 2.85237 0.00139594 0.997817 0.754133 0.00105982 0.00188072 0.000859865 0.455489 0.00188072 0.441837 0.000130075 1.02 0.888268 0.534516 0.286867 1.71823e-07 3.07384e-09 2378.31 3118.76 -0.0560684 0.482174 0.277403 0.253476 -0.593329 -0.169545 0.494455 -0.266748 -0.227716 2.205 1 0 297.257 0 2.17105 2.203 0.000299579 0.855962 0.680323 0.339174 0.423829 2.17124 135.745 83.8823 18.7187 60.8479 0.00402688 0 -40 10
1.304 3.775e-08 2.53933e-06 0.129272 0.129271 0.0120326 1.71591e-05 0.00115424 0.16159 0.000658487 0.162243 0.912471 101.68 0.239675 0.796502 4.32018 0.060325 0.0407564 0.959244 0.0196587 0.00441694 0.0189206 0.00423067 0.00534128 0.00607945 0.213651 0.243178 58.0209 -87.8975 126.242 15.9519 145.027 0.000141367 0.267229 192.801 0.310385 0.0673487 0.00409712 0.000562078 0.00138412 0.986972 0.991724 -2.98338e-06 -85.6613 0.0930461 31179.1 305.265 0.983507 0.319146 0.733343 0.733338 9.99958 2.98423e-06 1.19368e-05 0.132419 0.983117 0.931715 -0.0132923 4.91722e-06 0.5082 -1.94951e-20 7.21184e-24 -1.94879e-20 0.00139594 0.997816 8.59866e-05 0.152663 2.85237 0.00139594 0.997817 0.754218 0.00105984 0.00188072 0.000859866 0.455488 0.00188072 0.441843 0.000130077 1.02 0.888269 0.534516 0.286869 1.71823e-07 3.07386e-09 2378.3 3118.79 -0.056072 0.482174 0.277402 0.253478 -0.593328 -0.169545 0.494443 -0.266746 -0.227706 2.206 1 0 297.253 0 2.17119 2.204 0.000299578 0.85598 0.680368 0.339106 0.423852 2.17139 135.752 83.8819 18.7187 60.8477 0.0040269 0 -40 10
1.305 3.77789e-08 2.53933e-06 0.129319 0.129318 0.0120326 1.71722e-05 0.00115424 0.161649 0.000658488 0.162303 0.912552 101.679 0.239665 0.796624 4.32059 0.0603348 0.0407603 0.95924 0.0196583 0.00441728 0.0189201 0.00423097 0.00534171 0.00607988 0.213668 0.243195 58.021 -87.8975 126.242 15.9519 145.027 0.000141369 0.267229 192.801 0.310384 0.0673486 0.00409712 0.000562078 0.00138412 0.986972 0.991724 -2.9834e-06 -85.6612 0.0930461 31179.1 305.274 0.983507 0.319146 0.73335 0.733346 9.99958 2.98424e-06 1.19368e-05 0.132423 0.983118 0.931714 -0.0132922 4.91725e-06 0.508215 -1.94963e-20 7.21233e-24 -1.94891e-20 0.00139594 0.997816 8.59866e-05 0.152663 2.85237 0.00139594 0.997817 0.754304 0.00105986 0.00188072 0.000859866 0.455488 0.00188072 0.44185 0.00013008 1.02 0.88827 0.534515 0.28687 1.71824e-07 3.07388e-09 2378.28 3118.82 -0.0560757 0.482174 0.277402 0.25348 -0.593328 -0.169545 0.494431 -0.266744 -0.227697 2.207 1 0 297.25 0 2.17134 2.205 0.000299577 0.855999 0.680413 0.339039 0.423876 2.17153 135.76 83.8816 18.7186 60.8475 0.00402691 0 -40 10
1.306 3.78078e-08 2.53933e-06 0.129366 0.129365 0.0120326 1.71854e-05 0.00115424 0.161708 0.000658489 0.162362 0.912633 101.679 0.239655 0.796746 4.32101 0.0603446 0.0407643 0.959236 0.0196579 0.00441763 0.0189197 0.00423126 0.00534213 0.00608031 0.213685 0.243212 58.021 -87.8975 126.241 15.9518 145.027 0.00014137 0.26723 192.801 0.310384 0.0673486 0.00409713 0.000562079 0.00138412 0.986972 0.991723 -2.98341e-06 -85.6612 0.0930462 31179.1 305.283 0.983507 0.319146 0.733358 0.733353 9.99958 2.98424e-06 1.19369e-05 0.132426 0.98312 0.931714 -0.0132922 4.91728e-06 0.50823 -1.94975e-20 7.21283e-24 -1.94903e-20 0.00139594 0.997816 8.59867e-05 0.152663 2.85238 0.00139594 0.997817 0.754389 0.00105987 0.00188072 0.000859867 0.455488 0.00188072 0.441856 0.000130083 1.02 0.888271 0.534515 0.286872 1.71824e-07 3.07391e-09 2378.26 3118.85 -0.0560793 0.482174 0.277402 0.253482 -0.593327 -0.169545 0.494419 -0.266742 -0.227687 2.208 1 0 297.247 0 2.17148 2.206 0.000299576 0.856017 0.680458 0.338972 0.4239 2.17167 135.768 83.8812 18.7186 60.8474 0.00402693 0 -40 10
1.307 3.78367e-08 2.53933e-06 0.129414 0.129413 0.0120326 1.71985e-05 0.00115424 0.161767 0.00065849 0.162421 0.912715 101.679 0.239646 0.796868 4.32144 0.0603545 0.0407683 0.959232 0.0196574 0.00441797 0.0189193 0.00423155 0.00534256 0.00608074 0.213702 0.243229 58.0211 -87.8975 126.241 15.9518 145.027 0.000141372 0.26723 192.8 0.310383 0.0673485 0.00409713 0.00056208 0.00138413 0.986972 0.991723 -2.98343e-06 -85.6612 0.0930463 31179.1 305.293 0.983507 0.319146 0.733365 0.733361 9.99958 2.98425e-06 1.19369e-05 0.13243 0.983121 0.931714 -0.0132922 4.91731e-06 0.508244 -1.94987e-20 7.21333e-24 -1.94915e-20 0.00139595 0.997816 8.59868e-05 0.152663 2.85238 0.00139594 0.997817 0.754474 0.00105989 0.00188073 0.000859868 0.455488 0.00188072 0.441863 0.000130086 1.02 0.888272 0.534515 0.286873 1.71824e-07 3.07393e-09 2378.25 3118.89 -0.056083 0.482174 0.277401 0.253484 -0.593327 -0.169545 0.494407 -0.26674 -0.227677 2.209 1 0 297.244 0 2.17162 2.207 0.000299575 0.856035 0.680503 0.338904 0.423923 2.17182 135.775 83.8808 18.7186 60.8472 0.00402694 0 -40 10
1.308 3.78656e-08 2.53933e-06 0.129461 0.12946 0.0120325 1.72116e-05 0.00115424 0.161826 0.000658491 0.16248 0.912796 101.678 0.239636 0.79699 4.32186 0.0603643 0.0407722 0.959228 0.019657 0.00441832 0.0189188 0.00423185 0.00534298 0.00608117 0.213719 0.243247 58.0212 -87.8975 126.241 15.9518 145.027 0.000141373 0.26723 192.8 0.310383 0.0673484 0.00409713 0.00056208 0.00138413 0.986972 0.991723 -2.98344e-06 -85.6612 0.0930464 31179 305.302 0.983507 0.319146 0.733373 0.733369 9.99958 2.98425e-06 1.19369e-05 0.132433 0.983122 0.931713 -0.0132922 4.91734e-06 0.508259 -1.95e-20 7.21383e-24 -1.94928e-20 0.00139595 0.997816 8.59869e-05 0.152663 2.85238 0.00139595 0.997817 0.75456 0.00105991 0.00188073 0.000859869 0.455487 0.00188073 0.441869 0.000130089 1.02 0.888273 0.534514 0.286875 1.71825e-07 3.07395e-09 2378.23 3118.92 -0.0560866 0.482174 0.277401 0.253486 -0.593327 -0.169545 0.494395 -0.266737 -0.227667 2.21 1 0 297.241 0 2.17177 2.208 0.000299575 0.856053 0.680548 0.338837 0.423947 2.17196 135.783 83.8804 18.7186 60.847 0.00402696 0 -40 10
1.309 3.78945e-08 2.53933e-06 0.129508 0.129507 0.0120325 1.72248e-05 0.00115424 0.161885 0.000658492 0.162539 0.912878 101.678 0.239626 0.797112 4.32228 0.0603741 0.0407762 0.959224 0.0196566 0.00441866 0.0189184 0.00423214 0.0053434 0.0060816 0.213736 0.243264 58.0212 -87.8975 126.241 15.9517 145.027 0.000141375 0.26723 192.8 0.310382 0.0673484 0.00409713 0.000562081 0.00138413 0.986972 0.991723 -2.98346e-06 -85.6612 0.0930465 31179 305.311 0.983507 0.319146 0.733381 0.733376 9.99958 2.98426e-06 1.19369e-05 0.132437 0.983123 0.931713 -0.0132922 4.91737e-06 0.508274 -1.95012e-20 7.21432e-24 -1.9494e-20 0.00139595 0.997816 8.5987e-05 0.152664 2.85238 0.00139595 0.997817 0.754645 0.00105993 0.00188073 0.00085987 0.455487 0.00188073 0.441876 0.000130091 1.02 0.888275 0.534514 0.286876 1.71825e-07 3.07397e-09 2378.21 3118.95 -0.0560903 0.482174 0.277401 0.253488 -0.593326 -0.169545 0.494383 -0.266735 -0.227658 2.211 1 0 297.237 0 2.17191 2.209 0.000299574 0.856072 0.680593 0.338771 0.42397 2.17211 135.791 83.8801 18.7186 60.8468 0.00402697 0 -40 10
1.31 3.79234e-08 2.53933e-06 0.129556 0.129555 0.0120325 1.72379e-05 0.00115424 0.161945 0.000658493 0.162598 0.912959 101.677 0.239616 0.797234 4.3227 0.0603839 0.0407802 0.95922 0.0196562 0.00441901 0.018918 0.00423243 0.00534383 0.00608203 0.213753 0.243281 58.0213 -87.8975 126.241 15.9517 145.027 0.000141376 0.26723 192.8 0.310382 0.0673483 0.00409714 0.000562082 0.00138413 0.986972 0.991723 -2.98347e-06 -85.6612 0.0930466 31179 305.321 0.983507 0.319146 0.733388 0.733384 9.99958 2.98426e-06 1.19369e-05 0.13244 0.983124 0.931712 -0.0132922 4.9174e-06 0.508289 -1.95024e-20 7.21482e-24 -1.94952e-20 0.00139595 0.997816 8.5987e-05 0.152664 2.85238 0.00139595 0.997817 0.75473 0.00105994 0.00188073 0.00085987 0.455487 0.00188073 0.441882 0.000130094 1.02 0.888276 0.534514 0.286878 1.71825e-07 3.074e-09 2378.2 3118.98 -0.056094 0.482174 0.277401 0.25349 -0.593326 -0.169545 0.494372 -0.266733 -0.227648 2.212 1 0 297.234 0 2.17206 2.21 0.000299573 0.85609 0.680638 0.338704 0.423994 2.17225 135.798 83.8797 18.7185 60.8466 0.00402699 0 -40 10
1.311 3.79523e-08 2.53933e-06 0.129603 0.129602 0.0120325 1.7251e-05 0.00115424 0.162004 0.000658494 0.162657 0.913041 101.677 0.239606 0.797356 4.32312 0.0603937 0.0407842 0.959216 0.0196557 0.00441935 0.0189175 0.00423273 0.00534425 0.00608246 0.21377 0.243298 58.0214 -87.8975 126.241 15.9516 145.027 0.000141378 0.267231 192.8 0.310382 0.0673483 0.00409714 0.000562082 0.00138413 0.986972 0.991723 -2.98349e-06 -85.6612 0.0930467 31179 305.33 0.983507 0.319146 0.733396 0.733391 9.99958 2.98427e-06 1.1937e-05 0.132444 0.983126 0.931712 -0.0132922 4.91743e-06 0.508303 -1.95037e-20 7.21532e-24 -1.94964e-20 0.00139595 0.997816 8.59871e-05 0.152664 2.85238 0.00139595 0.997817 0.754815 0.00105996 0.00188073 0.000859871 0.455487 0.00188073 0.441889 0.000130097 1.02 0.888277 0.534513 0.286879 1.71825e-07 3.07402e-09 2378.18 3119.01 -0.0560977 0.482174 0.2774 0.253492 -0.593325 -0.169545 0.49436 -0.266731 -0.227638 2.213 1 0 297.231 0 2.1722 2.211 0.000299572 0.856109 0.680683 0.338637 0.424018 2.17239 135.806 83.8793 18.7185 60.8464 0.004027 0 -40 10
1.312 3.79811e-08 2.53933e-06 0.12965 0.129649 0.0120325 1.72642e-05 0.00115424 0.162062 0.000658495 0.162716 0.913122 101.676 0.239596 0.797479 4.32354 0.0604035 0.0407882 0.959212 0.0196553 0.0044197 0.0189171 0.00423302 0.00534468 0.00608289 0.213787 0.243316 58.0214 -87.8975 126.241 15.9516 145.027 0.000141379 0.267231 192.8 0.310381 0.0673482 0.00409714 0.000562083 0.00138414 0.986972 0.991723 -2.9835e-06 -85.6612 0.0930468 31178.9 305.34 0.983506 0.319146 0.733403 0.733399 9.99958 2.98427e-06 1.1937e-05 0.132447 0.983127 0.931711 -0.0132922 4.91746e-06 0.508318 -1.95049e-20 7.21582e-24 -1.94977e-20 0.00139595 0.997816 8.59872e-05 0.152664 2.85238 0.00139595 0.997817 0.7549 0.00105998 0.00188073 0.000859872 0.455487 0.00188073 0.441895 0.0001301 1.02 0.888278 0.534513 0.286881 1.71826e-07 3.07404e-09 2378.16 3119.04 -0.0561013 0.482174 0.2774 0.253494 -0.593325 -0.169545 0.494348 -0.266729 -0.227628 2.214 1 0 297.228 0 2.17234 2.212 0.000299571 0.856127 0.680728 0.33857 0.424041 2.17254 135.814 83.8789 18.7185 60.8463 0.00402702 0 -40 10
1.313 3.801e-08 2.53933e-06 0.129697 0.129696 0.0120325 1.72773e-05 0.00115424 0.162121 0.000658496 0.162775 0.913204 101.676 0.239587 0.797601 4.32397 0.0604133 0.0407921 0.959208 0.0196549 0.00442005 0.0189167 0.00423332 0.00534511 0.00608332 0.213804 0.243333 58.0215 -87.8975 126.24 15.9516 145.027 0.00014138 0.267231 192.799 0.310381 0.0673482 0.00409715 0.000562084 0.00138414 0.986972 0.991723 -2.98352e-06 -85.6612 0.0930468 31178.9 305.349 0.983506 0.319146 0.733411 0.733407 9.99958 2.98428e-06 1.1937e-05 0.132451 0.983128 0.931711 -0.0132922 4.91749e-06 0.508333 -1.95061e-20 7.21632e-24 -1.94989e-20 0.00139595 0.997816 8.59873e-05 0.152664 2.85238 0.00139595 0.997817 0.754986 0.00106 0.00188073 0.000859873 0.455486 0.00188073 0.441901 0.000130102 1.02 0.888279 0.534513 0.286882 1.71826e-07 3.07407e-09 2378.15 3119.08 -0.056105 0.482174 0.2774 0.253496 -0.593324 -0.169546 0.494336 -0.266727 -0.227618 2.215 1 0 297.224 0 2.17249 2.213 0.00029957 0.856146 0.680773 0.338504 0.424065 2.17268 135.822 83.8785 18.7185 60.8461 0.00402704 0 -40 10
1.314 3.80389e-08 2.53934e-06 0.129744 0.129743 0.0120325 1.72904e-05 0.00115424 0.16218 0.000658497 0.162834 0.913286 101.676 0.239577 0.797723 4.32439 0.0604232 0.0407961 0.959204 0.0196545 0.00442039 0.0189162 0.00423361 0.00534553 0.00608376 0.213821 0.24335 58.0215 -87.8975 126.24 15.9515 145.027 0.000141382 0.267231 192.799 0.31038 0.0673481 0.00409715 0.000562084 0.00138414 0.986972 0.991723 -2.98353e-06 -85.6612 0.0930469 31178.9 305.358 0.983506 0.319146 0.733419 0.733415 9.99958 2.98428e-06 1.1937e-05 0.132454 0.983129 0.93171 -0.0132922 4.91752e-06 0.508348 -1.95073e-20 7.21682e-24 -1.95001e-20 0.00139595 0.997816 8.59874e-05 0.152664 2.85238 0.00139595 0.997817 0.755071 0.00106002 0.00188074 0.000859874 0.455486 0.00188073 0.441908 0.000130105 1.02 0.88828 0.534512 0.286884 1.71826e-07 3.07409e-09 2378.13 3119.11 -0.0561087 0.482175 0.277399 0.253498 -0.593324 -0.169546 0.494324 -0.266725 -0.227608 2.216 1 0 297.221 0 2.17263 2.214 0.00029957 0.856164 0.680818 0.338437 0.424088 2.17282 135.829 83.8782 18.7184 60.8459 0.00402705 0 -40 10
1.315 3.80678e-08 2.53934e-06 0.129791 0.12979 0.0120325 1.73035e-05 0.00115424 0.162239 0.000658498 0.162893 0.913367 101.675 0.239567 0.797846 4.32481 0.060433 0.0408001 0.9592 0.019654 0.00442074 0.0189158 0.00423391 0.00534596 0.00608419 0.213838 0.243368 58.0216 -87.8975 126.24 15.9515 145.027 0.000141383 0.267231 192.799 0.31038 0.0673481 0.00409715 0.000562085 0.00138414 0.986972 0.991723 -2.98355e-06 -85.6611 0.093047 31178.9 305.368 0.983506 0.319146 0.733427 0.733422 9.99958 2.98429e-06 1.1937e-05 0.132458 0.98313 0.93171 -0.0132922 4.91755e-06 0.508363 -1.95086e-20 7.21732e-24 -1.95014e-20 0.00139595 0.997816 8.59875e-05 0.152664 2.85238 0.00139595 0.997817 0.755156 0.00106003 0.00188074 0.000859875 0.455486 0.00188074 0.441914 0.000130108 1.02 0.888281 0.534512 0.286886 1.71826e-07 3.07411e-09 2378.12 3119.14 -0.0561124 0.482175 0.277399 0.2535 -0.593324 -0.169546 0.494312 -0.266723 -0.227598 2.217 1 0 297.218 0 2.17277 2.215 0.000299569 0.856183 0.680863 0.338371 0.424112 2.17297 135.837 83.8778 18.7184 60.8457 0.00402707 0 -40 10
1.316 3.80967e-08 2.53934e-06 0.129838 0.129837 0.0120324 1.73167e-05 0.00115424 0.162298 0.000658499 0.162952 0.913449 101.675 0.239557 0.797968 4.32524 0.0604428 0.0408041 0.959196 0.0196536 0.00442108 0.0189154 0.0042342 0.00534639 0.00608462 0.213855 0.243385 58.0217 -87.8975 126.24 15.9515 145.027 0.000141385 0.267232 192.799 0.310379 0.067348 0.00409716 0.000562086 0.00138415 0.986972 0.991723 -2.98356e-06 -85.6611 0.0930471 31178.9 305.377 0.983506 0.319146 0.733434 0.73343 9.99958 2.98429e-06 1.19371e-05 0.132461 0.983132 0.931709 -0.0132922 4.91758e-06 0.508378 -1.95098e-20 7.21782e-24 -1.95026e-20 0.00139596 0.997816 8.59875e-05 0.152665 2.85238 0.00139596 0.997817 0.755241 0.00106005 0.00188074 0.000859875 0.455486 0.00188074 0.441921 0.000130111 1.02 0.888282 0.534512 0.286887 1.71827e-07 3.07414e-09 2378.1 3119.17 -0.0561161 0.482175 0.277399 0.253502 -0.593323 -0.169546 0.4943 -0.266721 -0.227588 2.218 1 0 297.215 0 2.17292 2.216 0.000299568 0.856202 0.680908 0.338305 0.424136 2.17311 135.845 83.8774 18.7184 60.8455 0.00402708 0 -40 10
1.317 3.81256e-08 2.53934e-06 0.129885 0.129884 0.0120324 1.73298e-05 0.00115425 0.162356 0.0006585 0.16301 0.91353 101.674 0.239547 0.79809 4.32566 0.0604526 0.0408082 0.959192 0.0196532 0.00442143 0.0189149 0.0042345 0.00534681 0.00608506 0.213873 0.243402 58.0217 -87.8975 126.24 15.9514 145.027 0.000141386 0.267232 192.799 0.310379 0.067348 0.00409716 0.000562086 0.00138415 0.986972 0.991723 -2.98358e-06 -85.6611 0.0930472 31178.8 305.387 0.983506 0.319146 0.733442 0.733438 9.99958 2.9843e-06 1.19371e-05 0.132465 0.983133 0.931709 -0.0132922 4.91761e-06 0.508392 -1.9511e-20 7.21832e-24 -1.95038e-20 0.00139596 0.997816 8.59876e-05 0.152665 2.85239 0.00139596 0.997817 0.755326 0.00106007 0.00188074 0.000859876 0.455485 0.00188074 0.441927 0.000130113 1.02 0.888283 0.534512 0.286889 1.71827e-07 3.07416e-09 2378.08 3119.21 -0.0561198 0.482175 0.277399 0.253505 -0.593323 -0.169546 0.494288 -0.266718 -0.227578 2.219 1 0 297.211 0 2.17306 2.217 0.000299567 0.85622 0.680953 0.338239 0.424159 2.17325 135.852 83.877 18.7184 60.8453 0.0040271 0 -40 10
1.318 3.81545e-08 2.53934e-06 0.129932 0.129931 0.0120324 1.73429e-05 0.00115425 0.162415 0.000658501 0.163069 0.913612 101.674 0.239538 0.798213 4.32609 0.0604625 0.0408122 0.959188 0.0196528 0.00442178 0.0189145 0.0042348 0.00534724 0.00608549 0.21389 0.24342 58.0218 -87.8975 126.24 15.9514 145.027 0.000141388 0.267232 192.799 0.310379 0.0673479 0.00409716 0.000562087 0.00138415 0.986972 0.991723 -2.98359e-06 -85.6611 0.0930473 31178.8 305.396 0.983506 0.319146 0.73345 0.733446 9.99958 2.9843e-06 1.19371e-05 0.132469 0.983134 0.931709 -0.0132922 4.91764e-06 0.508407 -1.95123e-20 7.21882e-24 -1.95051e-20 0.00139596 0.997816 8.59877e-05 0.152665 2.85239 0.00139596 0.997817 0.755411 0.00106009 0.00188074 0.000859877 0.455485 0.00188074 0.441934 0.000130116 1.02 0.888284 0.534511 0.28689 1.71827e-07 3.07418e-09 2378.07 3119.24 -0.0561236 0.482175 0.277398 0.253507 -0.593322 -0.169546 0.494275 -0.266716 -0.227569 2.22 1 0 297.208 0 2.1732 2.218 0.000299566 0.856239 0.680998 0.338173 0.424183 2.1734 135.86 83.8766 18.7184 60.8452 0.00402711 0 -40 10
1.319 3.81833e-08 2.53934e-06 0.129979 0.129978 0.0120324 1.73561e-05 0.00115425 0.162474 0.000658502 0.163128 0.913694 101.673 0.239528 0.798335 4.32652 0.0604723 0.0408162 0.959184 0.0196523 0.00442213 0.0189141 0.00423509 0.00534767 0.00608593 0.213907 0.243437 58.0219 -87.8975 126.24 15.9513 145.027 0.000141389 0.267232 192.798 0.310378 0.0673479 0.00409716 0.000562088 0.00138415 0.986972 0.991723 -2.98361e-06 -85.6611 0.0930474 31178.8 305.405 0.983506 0.319146 0.733458 0.733453 9.99958 2.98431e-06 1.19371e-05 0.132472 0.983135 0.931708 -0.0132922 4.91766e-06 0.508422 -1.95135e-20 7.21932e-24 -1.95063e-20 0.00139596 0.997816 8.59878e-05 0.152665 2.85239 0.00139596 0.997817 0.755496 0.0010601 0.00188074 0.000859878 0.455485 0.00188074 0.44194 0.000130119 1.02 0.888286 0.534511 0.286892 1.71828e-07 3.0742e-09 2378.05 3119.27 -0.0561273 0.482175 0.277398 0.253509 -0.593322 -0.169546 0.494263 -0.266714 -0.227559 2.221 1 0 297.205 0 2.17335 2.219 0.000299566 0.856258 0.681043 0.338107 0.424206 2.17354 135.868 83.8762 18.7183 60.845 0.00402713 0 -40 10
1.32 3.82122e-08 2.53934e-06 0.130026 0.130025 0.0120324 1.73692e-05 0.00115425 0.162532 0.000658503 0.163186 0.913776 101.673 0.239518 0.798458 4.32694 0.0604822 0.0408202 0.95918 0.0196519 0.00442248 0.0189136 0.00423539 0.0053481 0.00608636 0.213924 0.243454 58.0219 -87.8975 126.239 15.9513 145.027 0.000141391 0.267232 192.798 0.310378 0.0673478 0.00409717 0.000562088 0.00138415 0.986971 0.991723 -2.98362e-06 -85.6611 0.0930475 31178.8 305.415 0.983506 0.319146 0.733466 0.733461 9.99958 2.98431e-06 1.19371e-05 0.132476 0.983136 0.931708 -0.0132922 4.91769e-06 0.508437 -1.95147e-20 7.21982e-24 -1.95075e-20 0.00139596 0.997816 8.59879e-05 0.152665 2.85239 0.00139596 0.997817 0.755581 0.00106012 0.00188074 0.000859879 0.455485 0.00188074 0.441947 0.000130122 1.02 0.888287 0.534511 0.286893 1.71828e-07 3.07423e-09 2378.03 3119.3 -0.056131 0.482175 0.277398 0.253511 -0.593321 -0.169546 0.494251 -0.266712 -0.227549 2.222 1 0 297.201 0 2.17349 2.22 0.000299565 0.856277 0.681088 0.338041 0.42423 2.17368 135.875 83.8759 18.7183 60.8448 0.00402715 0 -40 10
1.321 3.82411e-08 2.53934e-06 0.130073 0.130072 0.0120324 1.73823e-05 0.00115425 0.162591 0.000658504 0.163245 0.913857 101.673 0.239508 0.79858 4.32737 0.060492 0.0408242 0.959176 0.0196515 0.00442282 0.0189132 0.00423569 0.00534853 0.0060868 0.213941 0.243472 58.022 -87.8975 126.239 15.9513 145.027 0.000141392 0.267233 192.798 0.310377 0.0673478 0.00409717 0.000562089 0.00138416 0.986971 0.991723 -2.98364e-06 -85.6611 0.0930475 31178.7 305.424 0.983506 0.319146 0.733473 0.733469 9.99958 2.98432e-06 1.19372e-05 0.132479 0.983137 0.931707 -0.0132922 4.91772e-06 0.508452 -1.9516e-20 7.22033e-24 -1.95088e-20 0.00139596 0.997816 8.59879e-05 0.152665 2.85239 0.00139596 0.997817 0.755666 0.00106014 0.00188075 0.000859879 0.455485 0.00188074 0.441953 0.000130125 1.02 0.888288 0.53451 0.286895 1.71828e-07 3.07425e-09 2378.02 3119.34 -0.0561347 0.482175 0.277397 0.253513 -0.593321 -0.169546 0.494239 -0.26671 -0.227539 2.223 1 0 297.198 0 2.17363 2.221 0.000299564 0.856295 0.681132 0.337975 0.424253 2.17383 135.883 83.8755 18.7183 60.8446 0.00402716 0 -40 10
1.322 3.827e-08 2.53934e-06 0.130119 0.130119 0.0120324 1.73955e-05 0.00115425 0.162649 0.000658505 0.163303 0.913939 101.672 0.239498 0.798703 4.3278 0.0605019 0.0408283 0.959172 0.019651 0.00442317 0.0189128 0.00423598 0.00534895 0.00608723 0.213958 0.243489 58.022 -87.8975 126.239 15.9512 145.027 0.000141394 0.267233 192.798 0.310377 0.0673477 0.00409717 0.00056209 0.00138416 0.986971 0.991723 -2.98365e-06 -85.6611 0.0930476 31178.7 305.434 0.983506 0.319146 0.733481 0.733477 9.99958 2.98432e-06 1.19372e-05 0.132483 0.983139 0.931707 -0.0132922 4.91775e-06 0.508467 -1.95172e-20 7.22083e-24 -1.951e-20 0.00139596 0.997816 8.5988e-05 0.152666 2.85239 0.00139596 0.997817 0.755751 0.00106016 0.00188075 0.00085988 0.455484 0.00188075 0.44196 0.000130127 1.02 0.888289 0.53451 0.286896 1.71828e-07 3.07427e-09 2378 3119.37 -0.0561385 0.482175 0.277397 0.253515 -0.593321 -0.169546 0.494227 -0.266708 -0.227529 2.224 1 0 297.195 0 2.17378 2.222 0.000299563 0.856314 0.681177 0.337909 0.424277 2.17397 135.891 83.8751 18.7183 60.8444 0.00402718 0 -40 10
1.323 3.82989e-08 2.53935e-06 0.130166 0.130165 0.0120323 1.74086e-05 0.00115425 0.162708 0.000658506 0.163362 0.914021 101.672 0.239488 0.798826 4.32822 0.0605117 0.0408323 0.959168 0.0196506 0.00442352 0.0189123 0.00423628 0.00534938 0.00608767 0.213975 0.243507 58.0221 -87.8975 126.239 15.9512 145.027 0.000141396 0.267233 192.798 0.310376 0.0673477 0.00409718 0.00056209 0.00138416 0.986971 0.991723 -2.98367e-06 -85.6611 0.0930477 31178.7 305.443 0.983506 0.319146 0.733489 0.733485 9.99958 2.98433e-06 1.19372e-05 0.132486 0.98314 0.931706 -0.0132922 4.91778e-06 0.508482 -1.95185e-20 7.22133e-24 -1.95112e-20 0.00139596 0.997816 8.59881e-05 0.152666 2.85239 0.00139596 0.997817 0.755835 0.00106017 0.00188075 0.000859881 0.455484 0.00188075 0.441966 0.00013013 1.02 0.88829 0.53451 0.286898 1.71829e-07 3.0743e-09 2377.98 3119.4 -0.0561422 0.482175 0.277397 0.253517 -0.59332 -0.169546 0.494215 -0.266706 -0.227518 2.225 1 0 297.192 0 2.17392 2.223 0.000299562 0.856333 0.681222 0.337844 0.4243 2.17411 135.898 83.8747 18.7182 60.8442 0.00402719 0 -40 10
1.324 3.83278e-08 2.53935e-06 0.130213 0.130212 0.0120323 1.74217e-05 0.00115425 0.162766 0.000658507 0.16342 0.914103 101.671 0.239478 0.798948 4.32865 0.0605216 0.0408363 0.959164 0.0196502 0.00442387 0.0189119 0.00423658 0.00534981 0.0060881 0.213993 0.243524 58.0222 -87.8975 126.239 15.9512 145.027 0.000141397 0.267233 192.798 0.310376 0.0673476 0.00409718 0.000562091 0.00138416 0.986971 0.991723 -2.98368e-06 -85.6611 0.0930478 31178.7 305.453 0.983506 0.319146 0.733497 0.733493 9.99958 2.98433e-06 1.19372e-05 0.13249 0.983141 0.931706 -0.0132922 4.91781e-06 0.508497 -1.95197e-20 7.22183e-24 -1.95125e-20 0.00139596 0.997816 8.59882e-05 0.152666 2.85239 0.00139596 0.997817 0.75592 0.00106019 0.00188075 0.000859882 0.455484 0.00188075 0.441972 0.000130133 1.02 0.888291 0.534509 0.286899 1.71829e-07 3.07432e-09 2377.97 3119.43 -0.056146 0.482175 0.277397 0.253519 -0.59332 -0.169546 0.494203 -0.266704 -0.227508 2.226 1 0 297.188 0 2.17406 2.224 0.000299561 0.856352 0.681267 0.337778 0.424324 2.17426 135.906 83.8743 18.7182 60.844 0.00402721 0 -40 10
1.325 3.83566e-08 2.53935e-06 0.13026 0.130259 0.0120323 1.74348e-05 0.00115425 0.162825 0.000658508 0.163478 0.914185 101.671 0.239469 0.799071 4.32908 0.0605314 0.0408404 0.95916 0.0196498 0.00442422 0.0189115 0.00423688 0.00535024 0.00608854 0.21401 0.243542 58.0222 -87.8975 126.239 15.9511 145.027 0.000141399 0.267233 192.797 0.310376 0.0673476 0.00409718 0.000562092 0.00138416 0.986971 0.991723 -2.9837e-06 -85.6611 0.0930479 31178.6 305.462 0.983506 0.319146 0.733505 0.733501 9.99958 2.98434e-06 1.19372e-05 0.132493 0.983142 0.931705 -0.0132922 4.91784e-06 0.508512 -1.95209e-20 7.22234e-24 -1.95137e-20 0.00139597 0.997816 8.59883e-05 0.152666 2.85239 0.00139597 0.997817 0.756005 0.00106021 0.00188075 0.000859883 0.455484 0.00188075 0.441979 0.000130136 1.02 0.888292 0.534509 0.286901 1.71829e-07 3.07434e-09 2377.95 3119.47 -0.0561497 0.482175 0.277396 0.253522 -0.593319 -0.169546 0.494191 -0.266702 -0.227498 2.227 1 0 297.185 0 2.17421 2.225 0.000299561 0.856371 0.681312 0.337713 0.424348 2.1744 135.914 83.8739 18.7182 60.8438 0.00402723 0 -40 10
1.326 3.83855e-08 2.53935e-06 0.130306 0.130305 0.0120323 1.7448e-05 0.00115425 0.162883 0.000658509 0.163537 0.914267 101.67 0.239459 0.799194 4.32951 0.0605413 0.0408444 0.959156 0.0196493 0.00442457 0.018911 0.00423717 0.00535067 0.00608898 0.214027 0.243559 58.0223 -87.8975 126.239 15.9511 145.027 0.0001414 0.267233 192.797 0.310375 0.0673475 0.00409719 0.000562092 0.00138417 0.986971 0.991723 -2.98371e-06 -85.661 0.093048 31178.6 305.472 0.983506 0.319146 0.733513 0.733509 9.99958 2.98434e-06 1.19373e-05 0.132497 0.983143 0.931705 -0.0132922 4.91787e-06 0.508527 -1.95222e-20 7.22284e-24 -1.95149e-20 0.00139597 0.997816 8.59883e-05 0.152666 2.85239 0.00139597 0.997817 0.75609 0.00106023 0.00188075 0.000859883 0.455483 0.00188075 0.441985 0.000130138 1.02 0.888293 0.534509 0.286902 1.71829e-07 3.07436e-09 2377.93 3119.5 -0.0561535 0.482175 0.277396 0.253524 -0.593319 -0.169546 0.494178 -0.2667 -0.227488 2.228 1 0 297.182 0 2.17435 2.226 0.00029956 0.85639 0.681357 0.337648 0.424371 2.17454 135.922 83.8735 18.7182 60.8437 0.00402724 0 -40 10
1.327 3.84144e-08 2.53935e-06 0.130353 0.130352 0.0120323 1.74611e-05 0.00115425 0.162941 0.00065851 0.163595 0.914348 101.67 0.239449 0.799316 4.32994 0.0605511 0.0408485 0.959152 0.0196489 0.00442492 0.0189106 0.00423747 0.0053511 0.00608941 0.214044 0.243577 58.0224 -87.8975 126.238 15.951 145.027 0.000141402 0.267234 192.797 0.310375 0.0673474 0.00409719 0.000562093 0.00138417 0.986971 0.991723 -2.98373e-06 -85.661 0.0930481 31178.6 305.481 0.983506 0.319146 0.733521 0.733516 9.99958 2.98435e-06 1.19373e-05 0.132501 0.983144 0.931704 -0.0132922 4.9179e-06 0.508542 -1.95234e-20 7.22334e-24 -1.95162e-20 0.00139597 0.997816 8.59884e-05 0.152666 2.8524 0.00139597 0.997817 0.756175 0.00106025 0.00188076 0.000859884 0.455483 0.00188075 0.441992 0.000130141 1.02 0.888294 0.534508 0.286904 1.7183e-07 3.07439e-09 2377.92 3119.53 -0.0561573 0.482176 0.277396 0.253526 -0.593318 -0.169546 0.494166 -0.266697 -0.227478 2.229 1 0 297.178 0 2.17449 2.227 0.000299559 0.856409 0.681402 0.337582 0.424395 2.17469 135.929 83.8731 18.7181 60.8435 0.00402726 0 -40 10
1.328 3.84433e-08 2.53935e-06 0.130399 0.130398 0.0120323 1.74742e-05 0.00115425 0.162999 0.00065851 0.163653 0.91443 101.67 0.239439 0.799439 4.33037 0.060561 0.0408525 0.959147 0.0196485 0.00442527 0.0189101 0.00423777 0.00535154 0.00608985 0.214061 0.243594 58.0224 -87.8975 126.238 15.951 145.027 0.000141403 0.267234 192.797 0.310374 0.0673474 0.00409719 0.000562094 0.00138417 0.986971 0.991723 -2.98374e-06 -85.661 0.0930482 31178.6 305.491 0.983506 0.319146 0.733529 0.733524 9.99958 2.98435e-06 1.19373e-05 0.132504 0.983145 0.931704 -0.0132922 4.91793e-06 0.508557 -1.95247e-20 7.22385e-24 -1.95174e-20 0.00139597 0.997816 8.59885e-05 0.152666 2.8524 0.00139597 0.997817 0.756259 0.00106026 0.00188076 0.000859885 0.455483 0.00188076 0.441998 0.000130144 1.02 0.888295 0.534508 0.286905 1.7183e-07 3.07441e-09 2377.9 3119.57 -0.056161 0.482176 0.277395 0.253528 -0.593318 -0.169546 0.494154 -0.266695 -0.227468 2.23 1 0 297.175 0 2.17464 2.228 0.000299558 0.856428 0.681447 0.337517 0.424418 2.17483 135.937 83.8727 18.7181 60.8433 0.00402727 0 -40 10
1.329 3.84722e-08 2.53935e-06 0.130446 0.130445 0.0120323 1.74874e-05 0.00115425 0.163057 0.000658511 0.163711 0.914512 101.669 0.239429 0.799562 4.3308 0.0605709 0.0408566 0.959143 0.019648 0.00442562 0.0189097 0.00423807 0.00535197 0.00609029 0.214079 0.243612 58.0225 -87.8976 126.238 15.951 145.027 0.000141405 0.267234 192.797 0.310374 0.0673473 0.0040972 0.000562094 0.00138417 0.986971 0.991723 -2.98376e-06 -85.661 0.0930482 31178.6 305.5 0.983506 0.319146 0.733537 0.733532 9.99958 2.98436e-06 1.19373e-05 0.132508 0.983147 0.931703 -0.0132922 4.91796e-06 0.508572 -1.95259e-20 7.22435e-24 -1.95187e-20 0.00139597 0.997816 8.59886e-05 0.152667 2.8524 0.00139597 0.997817 0.756344 0.00106028 0.00188076 0.000859886 0.455483 0.00188076 0.442005 0.000130147 1.02 0.888297 0.534508 0.286907 1.7183e-07 3.07443e-09 2377.88 3119.6 -0.0561648 0.482176 0.277395 0.25353 -0.593318 -0.169547 0.494142 -0.266693 -0.227458 2.231 1 0 297.172 0 2.17478 2.229 0.000299557 0.856448 0.681492 0.337452 0.424442 2.17497 135.945 83.8723 18.7181 60.8431 0.00402729 0 -40 10
1.33 3.85011e-08 2.53935e-06 0.130492 0.130491 0.0120322 1.75005e-05 0.00115425 0.163116 0.000658512 0.163769 0.914594 101.669 0.239419 0.799685 4.33123 0.0605807 0.0408607 0.959139 0.0196476 0.00442597 0.0189093 0.00423837 0.0053524 0.00609073 0.214096 0.243629 58.0226 -87.8976 126.238 15.9509 145.027 0.000141406 0.267234 192.797 0.310373 0.0673473 0.0040972 0.000562095 0.00138418 0.986971 0.991723 -2.98377e-06 -85.661 0.0930483 31178.5 305.51 0.983506 0.319146 0.733545 0.73354 9.99958 2.98436e-06 1.19373e-05 0.132511 0.983148 0.931703 -0.0132922 4.91799e-06 0.508587 -1.95271e-20 7.22486e-24 -1.95199e-20 0.00139597 0.997816 8.59887e-05 0.152667 2.8524 0.00139597 0.997817 0.756429 0.0010603 0.00188076 0.000859887 0.455482 0.00188076 0.442011 0.000130149 1.02 0.888298 0.534508 0.286908 1.7183e-07 3.07446e-09 2377.87 3119.63 -0.0561686 0.482176 0.277395 0.253532 -0.593317 -0.169547 0.494129 -0.266691 -0.227448 2.232 1 0 297.168 0 2.17492 2.23 0.000299556 0.856467 0.681536 0.337387 0.424465 2.17512 135.952 83.8719 18.7181 60.8429 0.00402731 0 -40 10
1.331 3.853e-08 2.53935e-06 0.130539 0.130538 0.0120322 1.75136e-05 0.00115425 0.163174 0.000658513 0.163827 0.914676 101.668 0.239409 0.799808 4.33166 0.0605906 0.0408647 0.959135 0.0196472 0.00442632 0.0189088 0.00423867 0.00535283 0.00609117 0.214113 0.243647 58.0226 -87.8976 126.238 15.9509 145.027 0.000141408 0.267234 192.796 0.310373 0.0673472 0.0040972 0.000562096 0.00138418 0.986971 0.991723 -2.98379e-06 -85.661 0.0930484 31178.5 305.519 0.983506 0.319146 0.733553 0.733548 9.99958 2.98437e-06 1.19374e-05 0.132515 0.983149 0.931702 -0.0132922 4.91802e-06 0.508602 -1.95284e-20 7.22536e-24 -1.95212e-20 0.00139597 0.997816 8.59887e-05 0.152667 2.8524 0.00139597 0.997817 0.756513 0.00106032 0.00188076 0.000859887 0.455482 0.00188076 0.442017 0.000130152 1.02 0.888299 0.534507 0.28691 1.71831e-07 3.07448e-09 2377.85 3119.67 -0.0561724 0.482176 0.277395 0.253534 -0.593317 -0.169547 0.494117 -0.266689 -0.227437 2.233 1 0 297.165 0 2.17507 2.231 0.000299556 0.856486 0.681581 0.337322 0.424489 2.17526 135.96 83.8715 18.7181 60.8427 0.00402732 0 -40 10
1.332 3.85588e-08 2.53936e-06 0.130585 0.130584 0.0120322 1.75267e-05 0.00115425 0.163232 0.000658514 0.163885 0.914758 101.668 0.2394 0.799931 4.33209 0.0606005 0.0408688 0.959131 0.0196467 0.00442667 0.0189084 0.00423897 0.00535326 0.00609161 0.214131 0.243664 58.0227 -87.8976 126.238 15.9508 145.027 0.000141409 0.267235 192.796 0.310373 0.0673472 0.0040972 0.000562096 0.00138418 0.986971 0.991723 -2.9838e-06 -85.661 0.0930485 31178.5 305.529 0.983506 0.319146 0.733561 0.733557 9.99958 2.98437e-06 1.19374e-05 0.132519 0.98315 0.931702 -0.0132922 4.91805e-06 0.508617 -1.95296e-20 7.22587e-24 -1.95224e-20 0.00139597 0.997816 8.59888e-05 0.152667 2.8524 0.00139597 0.997817 0.756598 0.00106033 0.00188076 0.000859888 0.455482 0.00188076 0.442024 0.000130155 1.02 0.8883 0.534507 0.286911 1.71831e-07 3.0745e-09 2377.83 3119.7 -0.0561762 0.482176 0.277394 0.253537 -0.593316 -0.169547 0.494105 -0.266687 -0.227427 2.234 1 0 297.162 0 2.17521 2.232 0.000299555 0.856505 0.681626 0.337258 0.424512 2.1754 135.968 83.8711 18.718 60.8425 0.00402734 0 -40 10
1.333 3.85877e-08 2.53936e-06 0.130632 0.130631 0.0120322 1.75399e-05 0.00115425 0.16329 0.000658515 0.163943 0.91484 101.667 0.23939 0.800054 4.33252 0.0606104 0.0408729 0.959127 0.0196463 0.00442702 0.018908 0.00423927 0.0053537 0.00609205 0.214148 0.243682 58.0227 -87.8976 126.238 15.9508 145.027 0.000141411 0.267235 192.796 0.310372 0.0673471 0.00409721 0.000562097 0.00138418 0.986971 0.991723 -2.98382e-06 -85.661 0.0930486 31178.5 305.538 0.983506 0.319146 0.733569 0.733565 9.99958 2.98438e-06 1.19374e-05 0.132522 0.983151 0.931701 -0.0132922 4.91808e-06 0.508632 -1.95309e-20 7.22637e-24 -1.95237e-20 0.00139597 0.997816 8.59889e-05 0.152667 2.8524 0.00139597 0.997817 0.756682 0.00106035 0.00188076 0.000859889 0.455482 0.00188076 0.44203 0.000130158 1.02 0.888301 0.534507 0.286913 1.71831e-07 3.07452e-09 2377.82 3119.73 -0.05618 0.482176 0.277394 0.253539 -0.593316 -0.169547 0.494092 -0.266685 -0.227417 2.235 1 0 297.158 0 2.17535 2.233 0.000299554 0.856524 0.681671 0.337193 0.424536 2.17555 135.975 83.8708 18.718 60.8423 0.00402736 0 -40 10
1.334 3.86166e-08 2.53936e-06 0.130678 0.130677 0.0120322 1.7553e-05 0.00115425 0.163347 0.000658516 0.164001 0.914922 101.667 0.23938 0.800177 4.33296 0.0606202 0.040877 0.959123 0.0196459 0.00442738 0.0189075 0.00423957 0.00535413 0.00609249 0.214165 0.243699 58.0228 -87.8976 126.237 15.9508 145.027 0.000141412 0.267235 192.796 0.310372 0.0673471 0.00409721 0.000562098 0.00138418 0.986971 0.991723 -2.98383e-06 -85.661 0.0930487 31178.4 305.548 0.983506 0.319146 0.733577 0.733573 9.99958 2.98438e-06 1.19374e-05 0.132526 0.983152 0.931701 -0.0132922 4.91811e-06 0.508647 -1.95321e-20 7.22688e-24 -1.95249e-20 0.00139598 0.997816 8.5989e-05 0.152667 2.8524 0.00139598 0.997817 0.756767 0.00106037 0.00188077 0.00085989 0.455482 0.00188076 0.442037 0.00013016 1.02 0.888302 0.534506 0.286914 1.71832e-07 3.07455e-09 2377.8 3119.77 -0.0561838 0.482176 0.277394 0.253541 -0.593315 -0.169547 0.49408 -0.266683 -0.227407 2.236 1 0 297.155 0 2.1755 2.234 0.000299553 0.856544 0.681716 0.337128 0.424559 2.17569 135.983 83.8704 18.718 60.8421 0.00402737 0 -40 10
1.335 3.86455e-08 2.53936e-06 0.130724 0.130723 0.0120322 1.75661e-05 0.00115425 0.163405 0.000658517 0.164059 0.915005 101.667 0.23937 0.8003 4.33339 0.0606301 0.040881 0.959119 0.0196454 0.00442773 0.0189071 0.00423987 0.00535456 0.00609293 0.214183 0.243717 58.0229 -87.8976 126.237 15.9507 145.027 0.000141414 0.267235 192.796 0.310371 0.067347 0.00409721 0.000562098 0.00138419 0.986971 0.991723 -2.98385e-06 -85.661 0.0930488 31178.4 305.557 0.983506 0.319146 0.733585 0.733581 9.99958 2.98439e-06 1.19374e-05 0.132529 0.983153 0.9317 -0.0132922 4.91814e-06 0.508662 -1.95334e-20 7.22738e-24 -1.95261e-20 0.00139598 0.997816 8.59891e-05 0.152668 2.8524 0.00139598 0.997817 0.756851 0.00106039 0.00188077 0.000859891 0.455481 0.00188077 0.442043 0.000130163 1.02 0.888303 0.534506 0.286916 1.71832e-07 3.07457e-09 2377.78 3119.8 -0.0561876 0.482176 0.277394 0.253543 -0.593315 -0.169547 0.494068 -0.266681 -0.227397 2.237 1 0 297.152 0 2.17564 2.235 0.000299552 0.856563 0.681761 0.337064 0.424583 2.17583 135.991 83.87 18.718 60.8419 0.00402739 0 -40 10
1.336 3.86744e-08 2.53936e-06 0.130771 0.13077 0.0120322 1.75793e-05 0.00115425 0.163463 0.000658518 0.164117 0.915087 101.666 0.23936 0.800423 4.33382 0.06064 0.0408851 0.959115 0.019645 0.00442808 0.0189066 0.00424017 0.005355 0.00609337 0.2142 0.243735 58.0229 -87.8976 126.237 15.9507 145.027 0.000141416 0.267235 192.796 0.310371 0.067347 0.00409722 0.000562099 0.00138419 0.986971 0.991723 -2.98386e-06 -85.661 0.0930489 31178.4 305.567 0.983506 0.319146 0.733593 0.733589 9.99958 2.98439e-06 1.19375e-05 0.132533 0.983154 0.9317 -0.0132922 4.91817e-06 0.508677 -1.95346e-20 7.22789e-24 -1.95274e-20 0.00139598 0.997816 8.59891e-05 0.152668 2.8524 0.00139598 0.997817 0.756936 0.0010604 0.00188077 0.000859891 0.455481 0.00188077 0.442049 0.000130166 1.02 0.888304 0.534506 0.286917 1.71832e-07 3.07459e-09 2377.77 3119.83 -0.0561914 0.482176 0.277393 0.253545 -0.593315 -0.169547 0.494055 -0.266678 -0.227386 2.238 1 0 297.148 0 2.17578 2.236 0.000299551 0.856583 0.681805 0.337 0.424606 2.17597 135.998 83.8696 18.7179 60.8417 0.00402741 0 -40 10
1.337 3.87033e-08 2.53936e-06 0.130817 0.130816 0.0120322 1.75924e-05 0.00115425 0.163521 0.000658519 0.164175 0.915169 101.666 0.23935 0.800546 4.33426 0.0606499 0.0408892 0.959111 0.0196446 0.00442843 0.0189062 0.00424047 0.00535543 0.00609381 0.214217 0.243752 58.023 -87.8976 126.237 15.9507 145.027 0.000141417 0.267236 192.795 0.31037 0.0673469 0.00409722 0.0005621 0.00138419 0.986971 0.991723 -2.98388e-06 -85.6609 0.0930489 31178.4 305.577 0.983506 0.319146 0.733601 0.733597 9.99958 2.9844e-06 1.19375e-05 0.132536 0.983155 0.931699 -0.0132922 4.9182e-06 0.508692 -1.95359e-20 7.2284e-24 -1.95286e-20 0.00139598 0.997816 8.59892e-05 0.152668 2.8524 0.00139598 0.997817 0.75702 0.00106042 0.00188077 0.000859892 0.455481 0.00188077 0.442056 0.000130169 1.02 0.888305 0.534505 0.286919 1.71832e-07 3.07462e-09 2377.75 3119.87 -0.0561953 0.482176 0.277393 0.253547 -0.593314 -0.169547 0.494043 -0.266676 -0.227376 2.239 1 0 297.145 0 2.17593 2.237 0.000299551 0.856602 0.68185 0.336935 0.42463 2.17612 136.006 83.8691 18.7179 60.8416 0.00402742 0 -40 10
1.338 3.87321e-08 2.53936e-06 0.130863 0.130862 0.0120321 1.76055e-05 0.00115426 0.163579 0.00065852 0.164233 0.915251 101.665 0.23934 0.800669 4.33469 0.0606598 0.0408933 0.959107 0.0196441 0.00442879 0.0189058 0.00424077 0.00535587 0.00609425 0.214235 0.24377 58.0231 -87.8976 126.237 15.9506 145.027 0.000141419 0.267236 192.795 0.31037 0.0673469 0.00409722 0.0005621 0.00138419 0.986971 0.991723 -2.98389e-06 -85.6609 0.093049 31178.4 305.586 0.983506 0.319146 0.733609 0.733605 9.99958 2.9844e-06 1.19375e-05 0.13254 0.983157 0.931699 -0.0132922 4.91823e-06 0.508707 -1.95371e-20 7.2289e-24 -1.95299e-20 0.00139598 0.997816 8.59893e-05 0.152668 2.85241 0.00139598 0.997817 0.757105 0.00106044 0.00188077 0.000859893 0.455481 0.00188077 0.442062 0.000130171 1.02 0.888306 0.534505 0.286921 1.71833e-07 3.07464e-09 2377.73 3119.9 -0.0561991 0.482176 0.277393 0.25355 -0.593314 -0.169547 0.494031 -0.266674 -0.227366 2.24 1 0 297.141 0 2.17607 2.238 0.00029955 0.856622 0.681895 0.336871 0.424653 2.17626 136.014 83.8687 18.7179 60.8414 0.00402744 0 -40 10
1.339 3.8761e-08 2.53936e-06 0.130909 0.130908 0.0120321 1.76186e-05 0.00115426 0.163636 0.000658521 0.16429 0.915333 101.665 0.23933 0.800792 4.33513 0.0606697 0.0408974 0.959103 0.0196437 0.00442914 0.0189053 0.00424107 0.0053563 0.00609469 0.214252 0.243788 58.0231 -87.8976 126.237 15.9506 145.027 0.00014142 0.267236 192.795 0.31037 0.0673468 0.00409723 0.000562101 0.0013842 0.986971 0.991723 -2.98391e-06 -85.6609 0.0930491 31178.3 305.596 0.983506 0.319146 0.733618 0.733613 9.99958 2.98441e-06 1.19375e-05 0.132544 0.983158 0.931698 -0.0132922 4.91826e-06 0.508722 -1.95384e-20 7.22941e-24 -1.95311e-20 0.00139598 0.997816 8.59894e-05 0.152668 2.85241 0.00139598 0.997817 0.757189 0.00106046 0.00188077 0.000859894 0.45548 0.00188077 0.442069 0.000130174 1.02 0.888308 0.534505 0.286922 1.71833e-07 3.07466e-09 2377.72 3119.94 -0.0562029 0.482176 0.277392 0.253552 -0.593313 -0.169547 0.494018 -0.266672 -0.227355 2.241 1 0 297.138 0 2.17621 2.239 0.000299549 0.856641 0.68194 0.336807 0.424677 2.1764 136.021 83.8683 18.7179 60.8412 0.00402746 0 -40 10
1.34 3.87899e-08 2.53936e-06 0.130955 0.130954 0.0120321 1.76318e-05 0.00115426 0.163694 0.000658522 0.164348 0.915415 101.664 0.23932 0.800915 4.33556 0.0606796 0.0409015 0.959098 0.0196433 0.00442949 0.0189049 0.00424137 0.00535674 0.00609513 0.214269 0.243805 58.0232 -87.8976 126.237 15.9505 145.027 0.000141422 0.267236 192.795 0.310369 0.0673468 0.00409723 0.000562102 0.0013842 0.986971 0.991723 -2.98392e-06 -85.6609 0.0930492 31178.3 305.605 0.983506 0.319146 0.733626 0.733621 9.99958 2.98441e-06 1.19375e-05 0.132547 0.983159 0.931698 -0.0132922 4.91829e-06 0.508737 -1.95396e-20 7.22992e-24 -1.95324e-20 0.00139598 0.997816 8.59895e-05 0.152668 2.85241 0.00139598 0.997817 0.757273 0.00106047 0.00188077 0.000859895 0.45548 0.00188077 0.442075 0.000130177 1.02 0.888309 0.534504 0.286924 1.71833e-07 3.07469e-09 2377.7 3119.97 -0.0562068 0.482176 0.277392 0.253554 -0.593313 -0.169547 0.494006 -0.26667 -0.227345 2.242 1 0 297.135 0 2.17636 2.24 0.000299548 0.856661 0.681985 0.336743 0.4247 2.17655 136.029 83.8679 18.7178 60.841 0.00402747 0 -40 10
1.341 3.88188e-08 2.53936e-06 0.131001 0.131 0.0120321 1.76449e-05 0.00115426 0.163752 0.000658523 0.164405 0.915498 101.664 0.239311 0.801038 4.336 0.0606895 0.0409056 0.959094 0.0196428 0.00442985 0.0189044 0.00424167 0.00535717 0.00609558 0.214287 0.243823 58.0232 -87.8976 126.236 15.9505 145.027 0.000141423 0.267236 192.795 0.310369 0.0673467 0.00409723 0.000562102 0.0013842 0.986971 0.991723 -2.98394e-06 -85.6609 0.0930493 31178.3 305.615 0.983506 0.319146 0.733634 0.73363 9.99958 2.98442e-06 1.19376e-05 0.132551 0.98316 0.931697 -0.0132922 4.91832e-06 0.508753 -1.95409e-20 7.23043e-24 -1.95337e-20 0.00139598 0.997816 8.59895e-05 0.152668 2.85241 0.00139598 0.997817 0.757358 0.00106049 0.00188078 0.000859895 0.45548 0.00188077 0.442081 0.00013018 1.02 0.88831 0.534504 0.286925 1.71833e-07 3.07471e-09 2377.68 3120 -0.0562106 0.482177 0.277392 0.253556 -0.593312 -0.169547 0.493993 -0.266668 -0.227335 2.243 1 0 297.131 0 2.1765 2.241 0.000299547 0.85668 0.68203 0.336679 0.424724 2.17669 136.037 83.8675 18.7178 60.8408 0.00402749 0 -40 10
1.342 3.88477e-08 2.53937e-06 0.131047 0.131046 0.0120321 1.7658e-05 0.00115426 0.163809 0.000658524 0.164463 0.91558 101.664 0.239301 0.801162 4.33643 0.0606994 0.0409098 0.95909 0.0196424 0.0044302 0.018904 0.00424198 0.00535761 0.00609602 0.214304 0.243841 58.0233 -87.8976 126.236 15.9505 145.027 0.000141425 0.267237 192.795 0.310368 0.0673467 0.00409723 0.000562103 0.0013842 0.986971 0.991723 -2.98395e-06 -85.6609 0.0930494 31178.3 305.625 0.983506 0.319146 0.733642 0.733638 9.99958 2.98442e-06 1.19376e-05 0.132555 0.983161 0.931697 -0.0132922 4.91835e-06 0.508768 -1.95421e-20 7.23094e-24 -1.95349e-20 0.00139599 0.997816 8.59896e-05 0.152669 2.85241 0.00139599 0.997817 0.757442 0.00106051 0.00188078 0.000859896 0.45548 0.00188078 0.442088 0.000130182 1.02 0.888311 0.534504 0.286927 1.71834e-07 3.07473e-09 2377.67 3120.04 -0.0562145 0.482177 0.277392 0.253558 -0.593312 -0.169547 0.493981 -0.266666 -0.227324 2.244 1 0 297.128 0 2.17664 2.242 0.000299546 0.8567 0.682074 0.336615 0.424747 2.17683 136.044 83.8671 18.7178 60.8406 0.00402751 0 -40 10
1.343 3.88766e-08 2.53937e-06 0.131093 0.131092 0.0120321 1.76712e-05 0.00115426 0.163867 0.000658524 0.164521 0.915662 101.663 0.239291 0.801285 4.33687 0.0607093 0.0409139 0.959086 0.019642 0.00443056 0.0189035 0.00424228 0.00535804 0.00609646 0.214322 0.243858 58.0234 -87.8976 126.236 15.9504 145.028 0.000141427 0.267237 192.794 0.310368 0.0673466 0.00409724 0.000562104 0.0013842 0.986971 0.991723 -2.98397e-06 -85.6609 0.0930495 31178.2 305.634 0.983506 0.319146 0.73365 0.733646 9.99958 2.98443e-06 1.19376e-05 0.132558 0.983162 0.931696 -0.0132922 4.91838e-06 0.508783 -1.95434e-20 7.23144e-24 -1.95362e-20 0.00139599 0.997816 8.59897e-05 0.152669 2.85241 0.00139599 0.997817 0.757526 0.00106053 0.00188078 0.000859897 0.45548 0.00188078 0.442094 0.000130185 1.02 0.888312 0.534504 0.286928 1.71834e-07 3.07475e-09 2377.65 3120.07 -0.0562183 0.482177 0.277391 0.253561 -0.593311 -0.169547 0.493968 -0.266664 -0.227314 2.245 1 0 297.124 0 2.17678 2.243 0.000299545 0.856719 0.682119 0.336552 0.424771 2.17698 136.052 83.8667 18.7178 60.8404 0.00402752 0 -40 10
1.344 3.89054e-08 2.53937e-06 0.131139 0.131138 0.0120321 1.76843e-05 0.00115426 0.163924 0.000658525 0.164578 0.915745 101.663 0.239281 0.801408 4.33731 0.0607192 0.040918 0.959082 0.0196415 0.00443091 0.0189031 0.00424258 0.00535848 0.00609691 0.214339 0.243876 58.0234 -87.8976 126.236 15.9504 145.028 0.000141428 0.267237 192.794 0.310367 0.0673465 0.00409724 0.000562104 0.00138421 0.986971 0.991723 -2.98398e-06 -85.6609 0.0930495 31178.2 305.644 0.983506 0.319146 0.733659 0.733654 9.99958 2.98443e-06 1.19376e-05 0.132562 0.983163 0.931696 -0.0132922 4.91841e-06 0.508798 -1.95446e-20 7.23195e-24 -1.95374e-20 0.00139599 0.997816 8.59898e-05 0.152669 2.85241 0.00139599 0.997817 0.75761 0.00106054 0.00188078 0.000859898 0.455479 0.00188078 0.442101 0.000130188 1.02 0.888313 0.534503 0.28693 1.71834e-07 3.07478e-09 2377.63 3120.11 -0.0562222 0.482177 0.277391 0.253563 -0.593311 -0.169547 0.493956 -0.266662 -0.227304 2.246 1 0 297.121 0 2.17693 2.244 0.000299545 0.856739 0.682164 0.336488 0.424794 2.17712 136.06 83.8663 18.7178 60.8402 0.00402754 0 -40 10
1.345 3.89343e-08 2.53937e-06 0.131185 0.131184 0.012032 1.76974e-05 0.00115426 0.163981 0.000658526 0.164635 0.915827 101.662 0.239271 0.801531 4.33775 0.0607291 0.0409221 0.959078 0.0196411 0.00443127 0.0189027 0.00424288 0.00535892 0.00609735 0.214357 0.243894 58.0235 -87.8976 126.236 15.9504 145.028 0.00014143 0.267237 192.794 0.310367 0.0673465 0.00409724 0.000562105 0.00138421 0.986971 0.991723 -2.984e-06 -85.6609 0.0930496 31178.2 305.653 0.983506 0.319146 0.733667 0.733663 9.99958 2.98444e-06 1.19376e-05 0.132565 0.983164 0.931695 -0.0132922 4.91844e-06 0.508813 -1.95459e-20 7.23246e-24 -1.95387e-20 0.00139599 0.997816 8.59899e-05 0.152669 2.85241 0.00139599 0.997817 0.757695 0.00106056 0.00188078 0.000859899 0.455479 0.00188078 0.442107 0.000130191 1.02 0.888314 0.534503 0.286931 1.71835e-07 3.0748e-09 2377.62 3120.14 -0.0562261 0.482177 0.277391 0.253565 -0.593311 -0.169548 0.493943 -0.266659 -0.227293 2.247 1 0 297.118 0 2.17707 2.245 0.000299544 0.856759 0.682209 0.336424 0.424818 2.17726 136.067 83.8659 18.7177 60.84 0.00402756 0 -40 10
1.346 3.89632e-08 2.53937e-06 0.131231 0.13123 0.012032 1.77105e-05 0.00115426 0.164039 0.000658527 0.164693 0.915909 101.662 0.239261 0.801655 4.33818 0.060739 0.0409263 0.959074 0.0196406 0.00443162 0.0189022 0.00424319 0.00535935 0.00609779 0.214374 0.243912 58.0236 -87.8976 126.236 15.9503 145.028 0.000141431 0.267237 192.794 0.310367 0.0673464 0.00409725 0.000562106 0.00138421 0.986971 0.991723 -2.98401e-06 -85.6609 0.0930497 31178.2 305.663 0.983506 0.319146 0.733675 0.733671 9.99958 2.98444e-06 1.19377e-05 0.132569 0.983165 0.931694 -0.0132922 4.91847e-06 0.508829 -1.95472e-20 7.23297e-24 -1.95399e-20 0.00139599 0.997816 8.599e-05 0.152669 2.85241 0.00139599 0.997817 0.757779 0.00106058 0.00188078 0.0008599 0.455479 0.00188078 0.442113 0.000130193 1.02 0.888315 0.534503 0.286933 1.71835e-07 3.07482e-09 2377.6 3120.18 -0.0562299 0.482177 0.27739 0.253567 -0.59331 -0.169548 0.493931 -0.266657 -0.227283 2.248 1 0 297.114 0 2.17721 2.246 0.000299543 0.856779 0.682253 0.336361 0.424841 2.1774 136.075 83.8655 18.7177 60.8398 0.00402757 0 -40 10
1.347 3.89921e-08 2.53937e-06 0.131277 0.131276 0.012032 1.77237e-05 0.00115426 0.164096 0.000658528 0.16475 0.915992 101.661 0.239251 0.801778 4.33862 0.060749 0.0409304 0.95907 0.0196402 0.00443198 0.0189018 0.00424349 0.00535979 0.00609824 0.214392 0.24393 58.0236 -87.8976 126.235 15.9503 145.028 0.000141433 0.267237 192.794 0.310366 0.0673464 0.00409725 0.000562106 0.00138421 0.986971 0.991723 -2.98403e-06 -85.6608 0.0930498 31178.2 305.673 0.983506 0.319146 0.733683 0.733679 9.99958 2.98445e-06 1.19377e-05 0.132573 0.983166 0.931694 -0.0132922 4.9185e-06 0.508844 -1.95484e-20 7.23348e-24 -1.95412e-20 0.00139599 0.997816 8.599e-05 0.152669 2.85241 0.00139599 0.997817 0.757863 0.0010606 0.00188079 0.0008599 0.455479 0.00188078 0.44212 0.000130196 1.02 0.888316 0.534502 0.286934 1.71835e-07 3.07485e-09 2377.58 3120.21 -0.0562338 0.482177 0.27739 0.25357 -0.59331 -0.169548 0.493918 -0.266655 -0.227272 2.249 1 0 297.111 0 2.17736 2.247 0.000299542 0.856798 0.682298 0.336298 0.424864 2.17755 136.083 83.8651 18.7177 60.8396 0.00402759 0 -40 10
1.348 3.9021e-08 2.53937e-06 0.131323 0.131322 0.012032 1.77368e-05 0.00115426 0.164153 0.000658529 0.164807 0.916074 101.661 0.239241 0.801902 4.33906 0.0607589 0.0409345 0.959065 0.0196398 0.00443233 0.0189013 0.00424379 0.00536023 0.00609868 0.214409 0.243947 58.0237 -87.8976 126.235 15.9502 145.028 0.000141435 0.267238 192.794 0.310366 0.0673463 0.00409725 0.000562107 0.00138421 0.986971 0.991723 -2.98404e-06 -85.6608 0.0930499 31178.1 305.682 0.983506 0.319146 0.733692 0.733687 9.99958 2.98445e-06 1.19377e-05 0.132576 0.983167 0.931693 -0.0132922 4.91853e-06 0.508859 -1.95497e-20 7.23399e-24 -1.95424e-20 0.00139599 0.997816 8.59901e-05 0.15267 2.85241 0.00139599 0.997817 0.757947 0.00106062 0.00188079 0.000859901 0.455478 0.00188079 0.442126 0.000130199 1.02 0.888317 0.534502 0.286936 1.71835e-07 3.07487e-09 2377.57 3120.25 -0.0562377 0.482177 0.27739 0.253572 -0.593309 -0.169548 0.493906 -0.266653 -0.227262 2.25 1 0 297.107 0 2.1775 2.248 0.000299541 0.856818 0.682343 0.336234 0.424888 2.17769 136.09 83.8647 18.7177 60.8394 0.00402761 0 -40 10
1.349 3.90499e-08 2.53937e-06 0.131369 0.131368 0.012032 1.77499e-05 0.00115426 0.164211 0.00065853 0.164865 0.916157 101.66 0.239231 0.802025 4.3395 0.0607688 0.0409387 0.959061 0.0196393 0.00443269 0.0189009 0.0042441 0.00536067 0.00609913 0.214427 0.243965 58.0238 -87.8976 126.235 15.9502 145.028 0.000141436 0.267238 192.793 0.310365 0.0673463 0.00409726 0.000562108 0.00138422 0.986971 0.991723 -2.98406e-06 -85.6608 0.09305 31178.1 305.692 0.983506 0.319146 0.7337 0.733696 9.99958 2.98446e-06 1.19377e-05 0.13258 0.983168 0.931693 -0.0132922 4.91856e-06 0.508874 -1.95509e-20 7.2345e-24 -1.95437e-20 0.00139599 0.997816 8.59902e-05 0.15267 2.85242 0.00139599 0.997817 0.758031 0.00106063 0.00188079 0.000859902 0.455478 0.00188079 0.442132 0.000130202 1.02 0.888318 0.534502 0.286937 1.71836e-07 3.07489e-09 2377.55 3120.28 -0.0562416 0.482177 0.27739 0.253574 -0.593309 -0.169548 0.493893 -0.266651 -0.227251 2.251 1 0 297.104 0 2.17764 2.249 0.00029954 0.856838 0.682388 0.336171 0.424911 2.17783 136.098 83.8643 18.7176 60.8392 0.00402762 0 -40 10
1.35 3.90787e-08 2.53937e-06 0.131414 0.131413 0.012032 1.77631e-05 0.00115426 0.164268 0.000658531 0.164922 0.916239 101.66 0.239221 0.802149 4.33994 0.0607787 0.0409428 0.959057 0.0196389 0.00443304 0.0189004 0.0042444 0.00536111 0.00609957 0.214444 0.243983 58.0238 -87.8976 126.235 15.9502 145.028 0.000141438 0.267238 192.793 0.310365 0.0673462 0.00409726 0.000562109 0.00138422 0.986971 0.991723 -2.98407e-06 -85.6608 0.0930501 31178.1 305.702 0.983506 0.319146 0.733708 0.733704 9.99958 2.98446e-06 1.19377e-05 0.132584 0.983169 0.931692 -0.0132922 4.91858e-06 0.50889 -1.95522e-20 7.23501e-24 -1.9545e-20 0.00139599 0.997816 8.59903e-05 0.15267 2.85242 0.00139599 0.997817 0.758115 0.00106065 0.00188079 0.000859903 0.455478 0.00188079 0.442139 0.000130204 1.02 0.88832 0.534501 0.286939 1.71836e-07 3.07491e-09 2377.53 3120.31 -0.0562455 0.482177 0.277389 0.253576 -0.593308 -0.169548 0.49388 -0.266649 -0.227241 2.252 1 0 297.1 0 2.17778 2.25 0.00029954 0.856858 0.682432 0.336108 0.424935 2.17798 136.106 83.8639 18.7176 60.839 0.00402764 0 -40 10
1.351 3.91076e-08 2.53938e-06 0.13146 0.131459 0.012032 1.77762e-05 0.00115426 0.164325 0.000658532 0.164979 0.916321 101.66 0.239211 0.802272 4.34038 0.0607887 0.040947 0.959053 0.0196385 0.0044334 0.0189 0.00424471 0.00536155 0.00610002 0.214462 0.244001 58.0239 -87.8976 126.235 15.9501 145.028 0.000141439 0.267238 192.793 0.310364 0.0673462 0.00409726 0.000562109 0.00138422 0.986971 0.991723 -2.98409e-06 -85.6608 0.0930502 31178.1 305.711 0.983506 0.319146 0.733717 0.733712 9.99958 2.98447e-06 1.19378e-05 0.132587 0.98317 0.931692 -0.0132922 4.91861e-06 0.508905 -1.95535e-20 7.23552e-24 -1.95462e-20 0.001396 0.997816 8.59904e-05 0.15267 2.85242 0.001396 0.997817 0.758199 0.00106067 0.00188079 0.000859904 0.455478 0.00188079 0.442145 0.000130207 1.02 0.888321 0.534501 0.28694 1.71836e-07 3.07494e-09 2377.52 3120.35 -0.0562494 0.482177 0.277389 0.253579 -0.593308 -0.169548 0.493868 -0.266647 -0.227231 2.253 1 0 297.097 0 2.17793 2.251 0.000299539 0.856878 0.682477 0.336045 0.424958 2.17812 136.113 83.8634 18.7176 60.8388 0.00402766 0 -40 10
1.352 3.91365e-08 2.53938e-06 0.131506 0.131505 0.0120319 1.77893e-05 0.00115426 0.164382 0.000658533 0.165036 0.916404 101.659 0.239201 0.802396 4.34082 0.0607986 0.0409512 0.959049 0.019638 0.00443376 0.0188995 0.00424501 0.00536199 0.00610047 0.214479 0.244019 58.0239 -87.8976 126.235 15.9501 145.028 0.000141441 0.267238 192.793 0.310364 0.0673461 0.00409727 0.00056211 0.00138422 0.986971 0.991723 -2.9841e-06 -85.6608 0.0930502 31178 305.721 0.983506 0.319146 0.733725 0.733721 9.99958 2.98447e-06 1.19378e-05 0.132591 0.983172 0.931691 -0.0132922 4.91864e-06 0.50892 -1.95547e-20 7.23604e-24 -1.95475e-20 0.001396 0.997816 8.59904e-05 0.15267 2.85242 0.001396 0.997817 0.758283 0.00106069 0.00188079 0.000859904 0.455477 0.00188079 0.442151 0.00013021 1.02 0.888322 0.534501 0.286942 1.71836e-07 3.07496e-09 2377.5 3120.38 -0.0562533 0.482177 0.277389 0.253581 -0.593307 -0.169548 0.493855 -0.266645 -0.22722 2.254 1 0 297.094 0 2.17807 2.252 0.000299538 0.856898 0.682522 0.335982 0.424982 2.17826 136.121 83.863 18.7176 60.8386 0.00402767 0 -40 10
1.353 3.91654e-08 2.53938e-06 0.131551 0.13155 0.0120319 1.78024e-05 0.00115426 0.164439 0.000658534 0.165093 0.916487 101.659 0.239191 0.802519 4.34126 0.0608085 0.0409553 0.959045 0.0196376 0.00443412 0.0188991 0.00424531 0.00536242 0.00610091 0.214497 0.244037 58.024 -87.8976 126.235 15.9501 145.028 0.000141443 0.267239 192.793 0.310364 0.0673461 0.00409727 0.000562111 0.00138423 0.986971 0.991723 -2.98412e-06 -85.6608 0.0930503 31178 305.731 0.983506 0.319146 0.733734 0.733729 9.99958 2.98448e-06 1.19378e-05 0.132594 0.983173 0.931691 -0.0132922 4.91867e-06 0.508935 -1.9556e-20 7.23655e-24 -1.95487e-20 0.001396 0.997816 8.59905e-05 0.15267 2.85242 0.001396 0.997817 0.758367 0.0010607 0.00188079 0.000859905 0.455477 0.00188079 0.442158 0.000130213 1.02 0.888323 0.5345 0.286943 1.71837e-07 3.07498e-09 2377.48 3120.42 -0.0562572 0.482177 0.277388 0.253583 -0.593307 -0.169548 0.493843 -0.266643 -0.227209 2.255 1 0 297.09 0 2.17821 2.253 0.000299537 0.856918 0.682567 0.335919 0.425005 2.1784 136.129 83.8626 18.7175 60.8384 0.00402769 0 -40 10
1.354 3.91943e-08 2.53938e-06 0.131597 0.131596 0.0120319 1.78156e-05 0.00115426 0.164496 0.000658535 0.16515 0.916569 101.658 0.239182 0.802643 4.34171 0.0608185 0.0409595 0.959041 0.0196371 0.00443447 0.0188986 0.00424562 0.00536286 0.00610136 0.214515 0.244054 58.0241 -87.8976 126.234 15.95 145.028 0.000141444 0.267239 192.793 0.310363 0.067346 0.00409727 0.000562111 0.00138423 0.986971 0.991723 -2.98413e-06 -85.6608 0.0930504 31178 305.741 0.983506 0.319146 0.733742 0.733738 9.99958 2.98448e-06 1.19378e-05 0.132598 0.983174 0.93169 -0.0132922 4.9187e-06 0.508951 -1.95572e-20 7.23706e-24 -1.955e-20 0.001396 0.997816 8.59906e-05 0.15267 2.85242 0.001396 0.997817 0.758451 0.00106072 0.0018808 0.000859906 0.455477 0.00188079 0.442164 0.000130215 1.02 0.888324 0.5345 0.286945 1.71837e-07 3.07501e-09 2377.47 3120.45 -0.0562611 0.482178 0.277388 0.253585 -0.593306 -0.169548 0.49383 -0.26664 -0.227199 2.256 1 0 297.087 0 2.17836 2.254 0.000299536 0.856938 0.682611 0.335856 0.425029 2.17855 136.136 83.8622 18.7175 60.8382 0.00402771 0 -40 10
1.355 3.92232e-08 2.53938e-06 0.131642 0.131642 0.0120319 1.78287e-05 0.00115426 0.164553 0.000658535 0.165207 0.916652 101.658 0.239172 0.802767 4.34215 0.0608284 0.0409637 0.959036 0.0196367 0.00443483 0.0188982 0.00424592 0.0053633 0.00610181 0.214532 0.244072 58.0241 -87.8976 126.234 15.95 145.028 0.000141446 0.267239 192.792 0.310363 0.067346 0.00409727 0.000562112 0.00138423 0.986971 0.991723 -2.98415e-06 -85.6608 0.0930505 31178 305.75 0.983506 0.319146 0.73375 0.733746 9.99958 2.98449e-06 1.19378e-05 0.132602 0.983175 0.93169 -0.0132922 4.91873e-06 0.508966 -1.95585e-20 7.23757e-24 -1.95513e-20 0.001396 0.997816 8.59907e-05 0.152671 2.85242 0.001396 0.997817 0.758535 0.00106074 0.0018808 0.000859907 0.455477 0.0018808 0.44217 0.000130218 1.02 0.888325 0.5345 0.286946 1.71837e-07 3.07503e-09 2377.45 3120.49 -0.056265 0.482178 0.277388 0.253588 -0.593306 -0.169548 0.493817 -0.266638 -0.227188 2.257 1 0 297.083 0 2.1785 2.255 0.000299535 0.856958 0.682656 0.335794 0.425052 2.17869 136.144 83.8618 18.7175 60.838 0.00402773 0 -40 10
1.356 3.9252e-08 2.53938e-06 0.131688 0.131687 0.0120319 1.78418e-05 0.00115426 0.16461 0.000658536 0.165264 0.916734 101.657 0.239162 0.80289 4.34259 0.0608383 0.0409678 0.959032 0.0196363 0.00443519 0.0188977 0.00424623 0.00536375 0.00610226 0.21455 0.24409 58.0242 -87.8977 126.234 15.9499 145.028 0.000141447 0.267239 192.792 0.310362 0.0673459 0.00409728 0.000562113 0.00138423 0.986971 0.991723 -2.98416e-06 -85.6608 0.0930506 31177.9 305.76 0.983506 0.319146 0.733759 0.733754 9.99958 2.98449e-06 1.19379e-05 0.132605 0.983176 0.931689 -0.0132922 4.91876e-06 0.508981 -1.95598e-20 7.23808e-24 -1.95525e-20 0.001396 0.997816 8.59908e-05 0.152671 2.85242 0.001396 0.997817 0.758619 0.00106076 0.0018808 0.000859908 0.455477 0.0018808 0.442177 0.000130221 1.02 0.888326 0.5345 0.286948 1.71838e-07 3.07505e-09 2377.43 3120.52 -0.0562689 0.482178 0.277388 0.25359 -0.593306 -0.169548 0.493805 -0.266636 -0.227178 2.258 1 0 297.08 0 2.17864 2.256 0.000299534 0.856978 0.682701 0.335731 0.425075 2.17883 136.152 83.8614 18.7175 60.8378 0.00402774 0 -40 10
1.357 3.92809e-08 2.53938e-06 0.131733 0.131733 0.0120319 1.7855e-05 0.00115426 0.164667 0.000658537 0.165321 0.916817 101.657 0.239152 0.803014 4.34303 0.0608483 0.040972 0.959028 0.0196358 0.00443555 0.0188973 0.00424654 0.00536419 0.0061027 0.214567 0.244108 58.0243 -87.8977 126.234 15.9499 145.028 0.000141449 0.267239 192.792 0.310362 0.0673459 0.00409728 0.000562113 0.00138423 0.98697 0.991723 -2.98418e-06 -85.6608 0.0930507 31177.9 305.77 0.983506 0.319146 0.733767 0.733763 9.99958 2.9845e-06 1.19379e-05 0.132609 0.983177 0.931689 -0.0132922 4.91879e-06 0.508997 -1.9561e-20 7.2386e-24 -1.95538e-20 0.001396 0.997816 8.59908e-05 0.152671 2.85242 0.001396 0.997817 0.758703 0.00106077 0.0018808 0.000859908 0.455476 0.0018808 0.442183 0.000130224 1.02 0.888327 0.534499 0.286949 1.71838e-07 3.07507e-09 2377.42 3120.56 -0.0562729 0.482178 0.277387 0.253592 -0.593305 -0.169548 0.493792 -0.266634 -0.227167 2.259 1 0 297.076 0 2.17878 2.257 0.000299534 0.856998 0.682745 0.335669 0.425099 2.17897 136.159 83.8609 18.7174 60.8376 0.00402776 0 -40 10
1.358 3.93098e-08 2.53938e-06 0.131779 0.131778 0.0120319 1.78681e-05 0.00115427 0.164724 0.000658538 0.165378 0.9169 101.657 0.239142 0.803138 4.34348 0.0608582 0.0409762 0.959024 0.0196354 0.00443591 0.0188968 0.00424684 0.00536463 0.00610315 0.214585 0.244126 58.0243 -87.8977 126.234 15.9499 145.028 0.000141451 0.26724 192.792 0.310361 0.0673458 0.00409728 0.000562114 0.00138424 0.98697 0.991723 -2.98419e-06 -85.6607 0.0930508 31177.9 305.779 0.983506 0.319146 0.733776 0.733771 9.99958 2.9845e-06 1.19379e-05 0.132613 0.983178 0.931688 -0.0132922 4.91882e-06 0.509012 -1.95623e-20 7.23911e-24 -1.95551e-20 0.001396 0.997816 8.59909e-05 0.152671 2.85242 0.001396 0.997817 0.758786 0.00106079 0.0018808 0.000859909 0.455476 0.0018808 0.442189 0.000130226 1.02 0.888328 0.534499 0.286951 1.71838e-07 3.0751e-09 2377.4 3120.6 -0.0562768 0.482178 0.277387 0.253594 -0.593305 -0.169548 0.493779 -0.266632 -0.227157 2.26 1 0 297.073 0 2.17893 2.258 0.000299533 0.857019 0.68279 0.335606 0.425122 2.17912 136.167 83.8605 18.7174 60.8374 0.00402778 0 -40 10
1.359 3.93387e-08 2.53938e-06 0.131824 0.131823 0.0120319 1.78812e-05 0.00115427 0.16478 0.000658539 0.165434 0.916982 101.656 0.239132 0.803262 4.34392 0.0608682 0.0409804 0.95902 0.0196349 0.00443626 0.0188964 0.00424715 0.00536507 0.0061036 0.214603 0.244144 58.0244 -87.8977 126.234 15.9498 145.028 0.000141452 0.26724 192.792 0.310361 0.0673458 0.00409729 0.000562115 0.00138424 0.98697 0.991723 -2.98421e-06 -85.6607 0.0930509 31177.9 305.789 0.983506 0.319146 0.733784 0.73378 9.99958 2.98451e-06 1.19379e-05 0.132616 0.983179 0.931687 -0.0132922 4.91885e-06 0.509027 -1.95636e-20 7.23962e-24 -1.95563e-20 0.001396 0.997816 8.5991e-05 0.152671 2.85242 0.001396 0.997817 0.75887 0.00106081 0.0018808 0.00085991 0.455476 0.0018808 0.442196 0.000130229 1.02 0.888329 0.534499 0.286952 1.71838e-07 3.07512e-09 2377.38 3120.63 -0.0562807 0.482178 0.277387 0.253597 -0.593304 -0.169548 0.493766 -0.26663 -0.227146 2.261 1 0 297.069 0 2.17907 2.259 0.000299532 0.857039 0.682835 0.335544 0.425146 2.17926 136.175 83.8601 18.7174 60.8372 0.00402779 0 -40 10
1.36 3.93676e-08 2.53939e-06 0.13187 0.131869 0.0120318 1.78943e-05 0.00115427 0.164837 0.00065854 0.165491 0.917065 101.656 0.239122 0.803385 4.34437 0.0608781 0.0409846 0.959015 0.0196345 0.00443662 0.0188959 0.00424745 0.00536551 0.00610405 0.21462 0.244162 58.0245 -87.8977 126.233 15.9498 145.028 0.000141454 0.26724 192.792 0.310361 0.0673457 0.00409729 0.000562115 0.00138424 0.98697 0.991723 -2.98422e-06 -85.6607 0.0930509 31177.9 305.799 0.983506 0.319146 0.733793 0.733788 9.99958 2.98451e-06 1.19379e-05 0.13262 0.98318 0.931687 -0.0132922 4.91888e-06 0.509043 -1.95648e-20 7.24014e-24 -1.95576e-20 0.00139601 0.997816 8.59911e-05 0.152671 2.85243 0.00139601 0.997817 0.758954 0.00106083 0.0018808 0.000859911 0.455476 0.0018808 0.442202 0.000130232 1.02 0.888331 0.534498 0.286954 1.71839e-07 3.07514e-09 2377.37 3120.67 -0.0562847 0.482178 0.277386 0.253599 -0.593304 -0.169549 0.493754 -0.266628 -0.227135 2.262 1 0 297.066 0 2.17921 2.26 0.000299531 0.857059 0.68288 0.335482 0.425169 2.1794 136.182 83.8597 18.7174 60.837 0.00402781 0 -40 10
1.361 3.93964e-08 2.53939e-06 0.131915 0.131914 0.0120318 1.79075e-05 0.00115427 0.164894 0.000658541 0.165548 0.917148 101.655 0.239112 0.803509 4.34481 0.0608881 0.0409888 0.959011 0.019634 0.00443698 0.0188955 0.00424776 0.00536595 0.0061045 0.214638 0.24418 58.0245 -87.8977 126.233 15.9498 145.028 0.000141456 0.26724 192.791 0.31036 0.0673457 0.00409729 0.000562116 0.00138424 0.98697 0.991723 -2.98424e-06 -85.6607 0.093051 31177.8 305.809 0.983505 0.319146 0.733801 0.733797 9.99958 2.98452e-06 1.1938e-05 0.132624 0.983181 0.931686 -0.0132922 4.91891e-06 0.509058 -1.95661e-20 7.24065e-24 -1.95589e-20 0.00139601 0.997816 8.59912e-05 0.152672 2.85243 0.00139601 0.997817 0.759038 0.00106084 0.00188081 0.000859912 0.455475 0.0018808 0.442208 0.000130234 1.02 0.888332 0.534498 0.286956 1.71839e-07 3.07517e-09 2377.35 3120.7 -0.0562886 0.482178 0.277386 0.253601 -0.593303 -0.169549 0.493741 -0.266626 -0.227125 2.263 1 0 297.062 0 2.17935 2.261 0.00029953 0.857079 0.682924 0.335419 0.425192 2.17955 136.19 83.8593 18.7173 60.8368 0.00402783 0 -40 10
1.362 3.94253e-08 2.53939e-06 0.13196 0.131959 0.0120318 1.79206e-05 0.00115427 0.16495 0.000658542 0.165604 0.91723 101.655 0.239102 0.803633 4.34526 0.0608981 0.040993 0.959007 0.0196336 0.00443734 0.018895 0.00424807 0.0053664 0.00610495 0.214656 0.244198 58.0246 -87.8977 126.233 15.9497 145.028 0.000141457 0.26724 192.791 0.31036 0.0673456 0.0040973 0.000562117 0.00138425 0.98697 0.991723 -2.98425e-06 -85.6607 0.0930511 31177.8 305.818 0.983505 0.319146 0.73381 0.733805 9.99958 2.98452e-06 1.1938e-05 0.132627 0.983182 0.931686 -0.0132922 4.91894e-06 0.509074 -1.95674e-20 7.24117e-24 -1.95601e-20 0.00139601 0.997816 8.59912e-05 0.152672 2.85243 0.00139601 0.997817 0.759121 0.00106086 0.00188081 0.000859912 0.455475 0.00188081 0.442215 0.000130237 1.02 0.888333 0.534498 0.286957 1.71839e-07 3.07519e-09 2377.34 3120.74 -0.0562926 0.482178 0.277386 0.253604 -0.593303 -0.169549 0.493728 -0.266624 -0.227114 2.264 1 0 297.059 0 2.1795 2.262 0.000299529 0.8571 0.682969 0.335357 0.425216 2.17969 136.197 83.8588 18.7173 60.8366 0.00402785 0 -40 10
1.363 3.94542e-08 2.53939e-06 0.132006 0.132005 0.0120318 1.79337e-05 0.00115427 0.165007 0.000658543 0.165661 0.917313 101.654 0.239092 0.803757 4.3457 0.060908 0.0409972 0.959003 0.0196332 0.0044377 0.0188946 0.00424837 0.00536684 0.0061054 0.214674 0.244216 58.0246 -87.8977 126.233 15.9497 145.028 0.000141459 0.267241 192.791 0.310359 0.0673455 0.0040973 0.000562117 0.00138425 0.98697 0.991723 -2.98427e-06 -85.6607 0.0930512 31177.8 305.828 0.983505 0.319146 0.733818 0.733814 9.99958 2.98453e-06 1.1938e-05 0.132631 0.983183 0.931685 -0.0132922 4.91897e-06 0.509089 -1.95687e-20 7.24168e-24 -1.95614e-20 0.00139601 0.997816 8.59913e-05 0.152672 2.85243 0.00139601 0.997817 0.759205 0.00106088 0.00188081 0.000859913 0.455475 0.00188081 0.442221 0.00013024 1.02 0.888334 0.534497 0.286959 1.71839e-07 3.07521e-09 2377.32 3120.77 -0.0562966 0.482178 0.277386 0.253606 -0.593302 -0.169549 0.493715 -0.266621 -0.227103 2.265 1 0 297.055 0 2.17964 2.263 0.000299528 0.85712 0.683014 0.335295 0.425239 2.17983 136.205 83.8584 18.7173 60.8364 0.00402786 0 -40 10
1.364 3.94831e-08 2.53939e-06 0.132051 0.13205 0.0120318 1.79469e-05 0.00115427 0.165063 0.000658544 0.165717 0.917396 101.654 0.239082 0.803881 4.34615 0.060918 0.0410014 0.958999 0.0196327 0.00443806 0.0188941 0.00424868 0.00536728 0.00610585 0.214691 0.244234 58.0247 -87.8977 126.233 15.9496 145.028 0.000141461 0.267241 192.791 0.310359 0.0673455 0.0040973 0.000562118 0.00138425 0.98697 0.991723 -2.98428e-06 -85.6607 0.0930513 31177.8 305.838 0.983505 0.319146 0.733827 0.733823 9.99958 2.98453e-06 1.1938e-05 0.132635 0.983184 0.931685 -0.0132922 4.919e-06 0.509105 -1.95699e-20 7.2422e-24 -1.95627e-20 0.00139601 0.997816 8.59914e-05 0.152672 2.85243 0.00139601 0.997817 0.759289 0.0010609 0.00188081 0.000859914 0.455475 0.00188081 0.442227 0.000130243 1.02 0.888335 0.534497 0.28696 1.7184e-07 3.07524e-09 2377.3 3120.81 -0.0563005 0.482178 0.277385 0.253608 -0.593302 -0.169549 0.493703 -0.266619 -0.227093 2.266 1 0 297.052 0 2.17978 2.264 0.000299528 0.857141 0.683058 0.335233 0.425263 2.17997 136.213 83.858 18.7173 60.8362 0.00402788 0 -40 10
1.365 3.9512e-08 2.53939e-06 0.132096 0.132095 0.0120318 1.796e-05 0.00115427 0.16512 0.000658544 0.165774 0.917479 101.653 0.239072 0.804005 4.34659 0.060928 0.0410056 0.958994 0.0196323 0.00443842 0.0188937 0.00424899 0.00536773 0.0061063 0.214709 0.244252 58.0248 -87.8977 126.233 15.9496 145.028 0.000141462 0.267241 192.791 0.310358 0.0673454 0.0040973 0.000562119 0.00138425 0.98697 0.991723 -2.9843e-06 -85.6607 0.0930514 31177.7 305.848 0.983505 0.319146 0.733835 0.733831 9.99958 2.98454e-06 1.1938e-05 0.132638 0.983185 0.931684 -0.0132922 4.91903e-06 0.50912 -1.95712e-20 7.24271e-24 -1.9564e-20 0.00139601 0.997816 8.59915e-05 0.152672 2.85243 0.00139601 0.997817 0.759372 0.00106091 0.00188081 0.000859915 0.455475 0.00188081 0.442234 0.000130245 1.02 0.888336 0.534497 0.286962 1.7184e-07 3.07526e-09 2377.29 3120.84 -0.0563045 0.482178 0.277385 0.253611 -0.593301 -0.169549 0.49369 -0.266617 -0.227082 2.267 1 0 297.048 0 2.17992 2.265 0.000299527 0.857161 0.683103 0.335172 0.425286 2.18012 136.22 83.8576 18.7172 60.836 0.0040279 0 -40 10
1.366 3.95408e-08 2.53939e-06 0.132141 0.13214 0.0120318 1.79731e-05 0.00115427 0.165176 0.000658545 0.16583 0.917562 101.653 0.239062 0.804129 4.34704 0.0609379 0.0410098 0.95899 0.0196318 0.00443878 0.0188932 0.0042493 0.00536817 0.00610675 0.214727 0.24427 58.0248 -87.8977 126.233 15.9496 145.028 0.000141464 0.267241 192.791 0.310358 0.0673454 0.00409731 0.000562119 0.00138425 0.98697 0.991723 -2.98431e-06 -85.6607 0.0930515 31177.7 305.858 0.983505 0.319146 0.733844 0.73384 9.99958 2.98454e-06 1.19381e-05 0.132642 0.983186 0.931683 -0.0132922 4.91906e-06 0.509135 -1.95725e-20 7.24323e-24 -1.95652e-20 0.00139601 0.997816 8.59916e-05 0.152672 2.85243 0.00139601 0.997817 0.759456 0.00106093 0.00188081 0.000859916 0.455474 0.00188081 0.44224 0.000130248 1.02 0.888337 0.534496 0.286963 1.7184e-07 3.07528e-09 2377.27 3120.88 -0.0563085 0.482178 0.277385 0.253613 -0.593301 -0.169549 0.493677 -0.266615 -0.227071 2.268 1 0 297.045 0 2.18007 2.266 0.000299526 0.857181 0.683148 0.33511 0.425309 2.18026 136.228 83.8572 18.7172 60.8358 0.00402792 0 -40 10
1.367 3.95697e-08 2.53939e-06 0.132186 0.132185 0.0120317 1.79862e-05 0.00115427 0.165233 0.000658546 0.165887 0.917644 101.653 0.239052 0.804253 4.34749 0.0609479 0.041014 0.958986 0.0196314 0.00443914 0.0188928 0.00424961 0.00536861 0.00610721 0.214745 0.244288 58.0249 -87.8977 126.232 15.9495 145.028 0.000141466 0.267241 192.791 0.310358 0.0673453 0.00409731 0.00056212 0.00138426 0.98697 0.991723 -2.98433e-06 -85.6607 0.0930516 31177.7 305.867 0.983505 0.319146 0.733853 0.733848 9.99958 2.98455e-06 1.19381e-05 0.132646 0.983187 0.931683 -0.0132922 4.91909e-06 0.509151 -1.95737e-20 7.24375e-24 -1.95665e-20 0.00139601 0.997816 8.59916e-05 0.152672 2.85243 0.00139601 0.997817 0.759539 0.00106095 0.00188081 0.000859916 0.455474 0.00188081 0.442246 0.000130251 1.02 0.888338 0.534496 0.286965 1.7184e-07 3.0753e-09 2377.25 3120.92 -0.0563124 0.482179 0.277384 0.253615 -0.5933 -0.169549 0.493664 -0.266613 -0.22706 2.269 1 0 297.041 0 2.18021 2.267 0.000299525 0.857202 0.683192 0.335048 0.425333 2.1804 136.236 83.8567 18.7172 60.8356 0.00402793 0 -40 10
1.368 3.95986e-08 2.53939e-06 0.132231 0.13223 0.0120317 1.79994e-05 0.00115427 0.165289 0.000658547 0.165943 0.917727 101.652 0.239042 0.804377 4.34794 0.0609579 0.0410183 0.958982 0.0196309 0.00443951 0.0188923 0.00424991 0.00536906 0.00610766 0.214762 0.244306 58.025 -87.8977 126.232 15.9495 145.028 0.000141467 0.267242 192.79 0.310357 0.0673453 0.00409731 0.000562121 0.00138426 0.98697 0.991722 -2.98434e-06 -85.6607 0.0930516 31177.7 305.877 0.983505 0.319146 0.733861 0.733857 9.99958 2.98455e-06 1.19381e-05 0.132649 0.983188 0.931682 -0.0132922 4.91912e-06 0.509166 -1.9575e-20 7.24426e-24 -1.95678e-20 0.00139602 0.997816 8.59917e-05 0.152673 2.85243 0.00139601 0.997817 0.759623 0.00106097 0.00188082 0.000859917 0.455474 0.00188082 0.442253 0.000130254 1.02 0.888339 0.534496 0.286966 1.71841e-07 3.07533e-09 2377.24 3120.95 -0.0563164 0.482179 0.277384 0.253618 -0.5933 -0.169549 0.493651 -0.266611 -0.22705 2.27 1 0 297.038 0 2.18035 2.268 0.000299524 0.857223 0.683237 0.334987 0.425356 2.18054 136.243 83.8563 18.7172 60.8354 0.00402795 0 -40 10
1.369 3.96275e-08 2.5394e-06 0.132276 0.132276 0.0120317 1.80125e-05 0.00115427 0.165346 0.000658548 0.165999 0.91781 101.652 0.239032 0.804501 4.34839 0.0609678 0.0410225 0.958977 0.0196305 0.00443987 0.0188919 0.00425022 0.0053695 0.00610811 0.21478 0.244324 58.025 -87.8977 126.232 15.9495 145.028 0.000141469 0.267242 192.79 0.310357 0.0673452 0.00409732 0.000562121 0.00138426 0.98697 0.991722 -2.98436e-06 -85.6606 0.0930517 31177.7 305.887 0.983505 0.319146 0.73387 0.733866 9.99958 2.98456e-06 1.19381e-05 0.132653 0.983189 0.931682 -0.0132922 4.91915e-06 0.509182 -1.95763e-20 7.24478e-24 -1.95691e-20 0.00139602 0.997816 8.59918e-05 0.152673 2.85243 0.00139602 0.997817 0.759706 0.00106098 0.00188082 0.000859918 0.455474 0.00188082 0.442259 0.000130256 1.02 0.88834 0.534496 0.286968 1.71841e-07 3.07535e-09 2377.22 3120.99 -0.0563204 0.482179 0.277384 0.25362 -0.5933 -0.169549 0.493638 -0.266609 -0.227039 2.271 1 0 297.034 0 2.18049 2.269 0.000299523 0.857243 0.683281 0.334925 0.425379 2.18069 136.251 83.8559 18.7172 60.8352 0.00402797 0 -40 10
1.37 3.96564e-08 2.5394e-06 0.132321 0.132321 0.0120317 1.80256e-05 0.00115427 0.165402 0.000658549 0.166056 0.917893 101.651 0.239022 0.804625 4.34883 0.0609778 0.0410267 0.958973 0.0196301 0.00444023 0.0188914 0.00425053 0.00536995 0.00610856 0.214798 0.244343 58.0251 -87.8977 126.232 15.9494 145.028 0.000141471 0.267242 192.79 0.310356 0.0673452 0.00409732 0.000562122 0.00138426 0.98697 0.991722 -2.98437e-06 -85.6606 0.0930518 31177.6 305.897 0.983505 0.319146 0.733879 0.733874 9.99958 2.98456e-06 1.19381e-05 0.132657 0.98319 0.931681 -0.0132922 4.91918e-06 0.509197 -1.95776e-20 7.2453e-24 -1.95703e-20 0.00139602 0.997816 8.59919e-05 0.152673 2.85243 0.00139602 0.997817 0.75979 0.001061 0.00188082 0.000859919 0.455473 0.00188082 0.442265 0.000130259 1.02 0.888342 0.534495 0.286969 1.71841e-07 3.07537e-09 2377.2 3121.02 -0.0563244 0.482179 0.277384 0.253622 -0.593299 -0.169549 0.493625 -0.266607 -0.227028 2.272 1 0 297.031 0 2.18064 2.27 0.000299522 0.857264 0.683326 0.334864 0.425403 2.18083 136.259 83.8554 18.7171 60.835 0.00402799 0 -40 10
1.371 3.96853e-08 2.5394e-06 0.132366 0.132366 0.0120317 1.80388e-05 0.00115427 0.165458 0.00065855 0.166112 0.917976 101.651 0.239012 0.804749 4.34928 0.0609878 0.041031 0.958969 0.0196296 0.00444059 0.018891 0.00425084 0.0053704 0.00610902 0.214816 0.244361 58.0251 -87.8977 126.232 15.9494 145.028 0.000141472 0.267242 192.79 0.310356 0.0673451 0.00409732 0.000562123 0.00138426 0.98697 0.991722 -2.98439e-06 -85.6606 0.0930519 31177.6 305.907 0.983505 0.319146 0.733887 0.733883 9.99958 2.98457e-06 1.19382e-05 0.132661 0.983191 0.931681 -0.0132922 4.91921e-06 0.509213 -1.95789e-20 7.24581e-24 -1.95716e-20 0.00139602 0.997816 8.5992e-05 0.152673 2.85244 0.00139602 0.997817 0.759873 0.00106102 0.00188082 0.00085992 0.455473 0.00188082 0.442271 0.000130262 1.02 0.888343 0.534495 0.286971 1.71842e-07 3.0754e-09 2377.19 3121.06 -0.0563284 0.482179 0.277383 0.253625 -0.593299 -0.169549 0.493612 -0.266605 -0.227017 2.273 1 0 297.027 0 2.18078 2.271 0.000299521 0.857284 0.683371 0.334803 0.425426 2.18097 136.266 83.855 18.7171 60.8347 0.004028 0 -40 10
1.372 3.97141e-08 2.5394e-06 0.132411 0.13241 0.0120317 1.80519e-05 0.00115427 0.165514 0.000658551 0.166168 0.918059 101.65 0.239002 0.804874 4.34973 0.0609978 0.0410352 0.958965 0.0196292 0.00444095 0.0188905 0.00425115 0.00537084 0.00610947 0.214834 0.244379 58.0252 -87.8977 126.232 15.9493 145.028 0.000141474 0.267242 192.79 0.310355 0.0673451 0.00409733 0.000562123 0.00138427 0.98697 0.991722 -2.9844e-06 -85.6606 0.093052 31177.6 305.916 0.983505 0.319146 0.733896 0.733892 9.99958 2.98457e-06 1.19382e-05 0.132664 0.983192 0.93168 -0.0132922 4.91924e-06 0.509228 -1.95801e-20 7.24633e-24 -1.95729e-20 0.00139602 0.997816 8.59921e-05 0.152673 2.85244 0.00139602 0.997817 0.759957 0.00106104 0.00188082 0.000859921 0.455473 0.00188082 0.442278 0.000130264 1.02 0.888344 0.534495 0.286972 1.71842e-07 3.07542e-09 2377.17 3121.1 -0.0563324 0.482179 0.277383 0.253627 -0.593298 -0.169549 0.4936 -0.266602 -0.227006 2.274 1 0 297.023 0 2.18092 2.272 0.000299521 0.857305 0.683415 0.334741 0.42545 2.18111 136.274 83.8546 18.7171 60.8345 0.00402802 0 -40 10
1.373 3.9743e-08 2.5394e-06 0.132456 0.132455 0.0120317 1.8065e-05 0.00115427 0.16557 0.000658552 0.166224 0.918142 101.65 0.238992 0.804998 4.35018 0.0610078 0.0410395 0.958961 0.0196287 0.00444132 0.0188901 0.00425146 0.00537129 0.00610992 0.214852 0.244397 58.0253 -87.8977 126.231 15.9493 145.028 0.000141476 0.267242 192.79 0.310355 0.067345 0.00409733 0.000562124 0.00138427 0.98697 0.991722 -2.98442e-06 -85.6606 0.0930521 31177.6 305.926 0.983505 0.319146 0.733905 0.7339 9.99958 2.98458e-06 1.19382e-05 0.132668 0.983193 0.931679 -0.0132922 4.91927e-06 0.509244 -1.95814e-20 7.24685e-24 -1.95742e-20 0.00139602 0.997816 8.59921e-05 0.152673 2.85244 0.00139602 0.997817 0.76004 0.00106105 0.00188082 0.000859921 0.455473 0.00188082 0.442284 0.000130267 1.02 0.888345 0.534494 0.286974 1.71842e-07 3.07544e-09 2377.15 3121.13 -0.0563364 0.482179 0.277383 0.253629 -0.593298 -0.169549 0.493587 -0.2666 -0.226996 2.275 1 0 297.02 0 2.18106 2.273 0.00029952 0.857326 0.68346 0.33468 0.425473 2.18126 136.282 83.8542 18.7171 60.8343 0.00402804 0 -40 10
1.374 3.97719e-08 2.5394e-06 0.132501 0.1325 0.0120316 1.80781e-05 0.00115427 0.165626 0.000658552 0.16628 0.918225 101.649 0.238982 0.805122 4.35064 0.0610178 0.0410437 0.958956 0.0196283 0.00444168 0.0188896 0.00425177 0.00537173 0.00611038 0.214869 0.244415 58.0253 -87.8977 126.231 15.9493 145.028 0.000141477 0.267243 192.789 0.310355 0.067345 0.00409733 0.000562125 0.00138427 0.98697 0.991722 -2.98443e-06 -85.6606 0.0930522 31177.5 305.936 0.983505 0.319146 0.733913 0.733909 9.99958 2.98458e-06 1.19382e-05 0.132672 0.983194 0.931679 -0.0132921 4.9193e-06 0.50926 -1.95827e-20 7.24737e-24 -1.95754e-20 0.00139602 0.997816 8.59922e-05 0.152674 2.85244 0.00139602 0.997817 0.760123 0.00106107 0.00188083 0.000859922 0.455473 0.00188082 0.44229 0.00013027 1.02 0.888346 0.534494 0.286975 1.71842e-07 3.07546e-09 2377.14 3121.17 -0.0563404 0.482179 0.277382 0.253632 -0.593297 -0.169549 0.493574 -0.266598 -0.226985 2.276 1 0 297.016 0 2.18121 2.274 0.000299519 0.857346 0.683505 0.334619 0.425496 2.1814 136.289 83.8537 18.717 60.8341 0.00402806 0 -40 10
1.375 3.98008e-08 2.5394e-06 0.132546 0.132545 0.0120316 1.80913e-05 0.00115427 0.165682 0.000658553 0.166336 0.918308 101.649 0.238972 0.805246 4.35109 0.0610278 0.041048 0.958952 0.0196278 0.00444204 0.0188892 0.00425208 0.00537218 0.00611083 0.214887 0.244433 58.0254 -87.8977 126.231 15.9492 145.028 0.000141479 0.267243 192.789 0.310354 0.0673449 0.00409734 0.000562125 0.00138427 0.98697 0.991722 -2.98445e-06 -85.6606 0.0930523 31177.5 305.946 0.983505 0.319146 0.733922 0.733918 9.99958 2.98459e-06 1.19382e-05 0.132675 0.983195 0.931678 -0.0132921 4.91933e-06 0.509275 -1.9584e-20 7.24789e-24 -1.95767e-20 0.00139602 0.997816 8.59923e-05 0.152674 2.85244 0.00139602 0.997817 0.760207 0.00106109 0.00188083 0.000859923 0.455472 0.00188083 0.442297 0.000130273 1.02 0.888347 0.534494 0.286977 1.71843e-07 3.07549e-09 2377.12 3121.21 -0.0563445 0.482179 0.277382 0.253634 -0.593297 -0.169549 0.493561 -0.266596 -0.226974 2.277 1 0 297.013 0 2.18135 2.275 0.000299518 0.857367 0.683549 0.334558 0.42552 2.18154 136.297 83.8533 18.717 60.8339 0.00402808 0 -40 10
1.376 3.98297e-08 2.5394e-06 0.132591 0.13259 0.0120316 1.81044e-05 0.00115427 0.165738 0.000658554 0.166392 0.918391 101.648 0.238962 0.805371 4.35154 0.0610378 0.0410522 0.958948 0.0196274 0.0044424 0.0188887 0.00425239 0.00537263 0.00611129 0.214905 0.244452 58.0255 -87.8977 126.231 15.9492 145.028 0.000141481 0.267243 192.789 0.310354 0.0673449 0.00409734 0.000562126 0.00138428 0.98697 0.991722 -2.98446e-06 -85.6606 0.0930523 31177.5 305.956 0.983505 0.319146 0.733931 0.733926 9.99958 2.98459e-06 1.19383e-05 0.132679 0.983196 0.931678 -0.0132921 4.91936e-06 0.509291 -1.95853e-20 7.2484e-24 -1.9578e-20 0.00139602 0.997816 8.59924e-05 0.152674 2.85244 0.00139602 0.997817 0.76029 0.00106111 0.00188083 0.000859924 0.455472 0.00188083 0.442303 0.000130275 1.02 0.888348 0.534493 0.286978 1.71843e-07 3.07551e-09 2377.1 3121.24 -0.0563485 0.482179 0.277382 0.253636 -0.593296 -0.16955 0.493548 -0.266594 -0.226963 2.278 1 0 297.009 0 2.18149 2.276 0.000299517 0.857388 0.683594 0.334497 0.425543 2.18168 136.304 83.8529 18.717 60.8337 0.00402809 0 -40 10
1.377 3.98585e-08 2.5394e-06 0.132635 0.132635 0.0120316 1.81175e-05 0.00115427 0.165794 0.000658555 0.166448 0.918474 101.648 0.238952 0.805495 4.35199 0.0610478 0.0410565 0.958943 0.0196269 0.00444277 0.0188883 0.0042527 0.00537308 0.00611174 0.214923 0.24447 58.0255 -87.8977 126.231 15.9492 145.028 0.000141482 0.267243 192.789 0.310353 0.0673448 0.00409734 0.000562127 0.00138428 0.98697 0.991722 -2.98448e-06 -85.6606 0.0930524 31177.5 305.966 0.983505 0.319146 0.73394 0.733935 9.99958 2.9846e-06 1.19383e-05 0.132683 0.983197 0.931677 -0.0132921 4.91939e-06 0.509306 -1.95865e-20 7.24892e-24 -1.95793e-20 0.00139603 0.997816 8.59925e-05 0.152674 2.85244 0.00139603 0.997817 0.760373 0.00106112 0.00188083 0.000859925 0.455472 0.00188083 0.442309 0.000130278 1.02 0.888349 0.534493 0.28698 1.71843e-07 3.07553e-09 2377.09 3121.28 -0.0563525 0.482179 0.277382 0.253639 -0.593296 -0.16955 0.493535 -0.266592 -0.226952 2.279 1 0 297.006 0 2.18163 2.277 0.000299516 0.857409 0.683638 0.334436 0.425566 2.18182 136.312 83.8524 18.717 60.8335 0.00402811 0 -40 10
1.378 3.98874e-08 2.53941e-06 0.13268 0.132679 0.0120316 1.81306e-05 0.00115428 0.16585 0.000658556 0.166504 0.918557 101.648 0.238942 0.805619 4.35244 0.0610578 0.0410608 0.958939 0.0196265 0.00444313 0.0188878 0.00425301 0.00537352 0.0061122 0.214941 0.244488 58.0256 -87.8977 126.231 15.9491 145.028 0.000141484 0.267243 192.789 0.310353 0.0673448 0.00409734 0.000562127 0.00138428 0.98697 0.991722 -2.98449e-06 -85.6606 0.0930525 31177.5 305.976 0.983505 0.319146 0.733948 0.733944 9.99958 2.9846e-06 1.19383e-05 0.132687 0.983198 0.931677 -0.0132921 4.91942e-06 0.509322 -1.95878e-20 7.24944e-24 -1.95806e-20 0.00139603 0.997816 8.59925e-05 0.152674 2.85244 0.00139603 0.997817 0.760457 0.00106114 0.00188083 0.000859925 0.455472 0.00188083 0.442315 0.000130281 1.02 0.88835 0.534493 0.286981 1.71843e-07 3.07556e-09 2377.07 3121.32 -0.0563565 0.482179 0.277381 0.253641 -0.593295 -0.16955 0.493522 -0.26659 -0.226941 2.28 1 0 297.002 0 2.18178 2.278 0.000299515 0.85743 0.683683 0.334376 0.42559 2.18197 136.32 83.852 18.7169 60.8333 0.00402813 0 -40 10
1.379 3.99163e-08 2.53941e-06 0.132725 0.132724 0.0120316 1.81438e-05 0.00115428 0.165906 0.000658557 0.16656 0.918641 101.647 0.238932 0.805744 4.3529 0.0610678 0.0410651 0.958935 0.019626 0.0044435 0.0188873 0.00425332 0.00537397 0.00611265 0.214959 0.244506 58.0257 -87.8977 126.23 15.9491 145.028 0.000141486 0.267244 192.789 0.310352 0.0673447 0.00409735 0.000562128 0.00138428 0.98697 0.991722 -2.98451e-06 -85.6605 0.0930526 31177.4 305.985 0.983505 0.319146 0.733957 0.733953 9.99958 2.98461e-06 1.19383e-05 0.13269 0.983199 0.931676 -0.0132921 4.91945e-06 0.509337 -1.95891e-20 7.24996e-24 -1.95819e-20 0.00139603 0.997816 8.59926e-05 0.152674 2.85244 0.00139603 0.997817 0.76054 0.00106116 0.00188083 0.000859926 0.455471 0.00188083 0.442322 0.000130283 1.02 0.888351 0.534492 0.286983 1.71844e-07 3.07558e-09 2377.05 3121.35 -0.0563606 0.482179 0.277381 0.253643 -0.593295 -0.16955 0.493509 -0.266588 -0.22693 2.281 1 0 296.998 0 2.18192 2.279 0.000299514 0.857451 0.683727 0.334315 0.425613 2.18211 136.327 83.8516 18.7169 60.8331 0.00402815 0 -40 10
1.38 3.99452e-08 2.53941e-06 0.13277 0.132769 0.0120316 1.81569e-05 0.00115428 0.165962 0.000658558 0.166616 0.918724 101.647 0.238922 0.805868 4.35335 0.0610778 0.0410693 0.958931 0.0196256 0.00444386 0.0188869 0.00425363 0.00537442 0.00611311 0.214977 0.244524 58.0257 -87.8977 126.23 15.949 145.028 0.000141487 0.267244 192.788 0.310352 0.0673447 0.00409735 0.000562129 0.00138428 0.98697 0.991722 -2.98452e-06 -85.6605 0.0930527 31177.4 305.995 0.983505 0.319146 0.733966 0.733962 9.99958 2.98461e-06 1.19383e-05 0.132694 0.9832 0.931675 -0.0132921 4.91948e-06 0.509353 -1.95904e-20 7.25048e-24 -1.95831e-20 0.00139603 0.997816 8.59927e-05 0.152674 2.85244 0.00139603 0.997817 0.760623 0.00106118 0.00188083 0.000859927 0.455471 0.00188083 0.442328 0.000130286 1.02 0.888353 0.534492 0.286984 1.71844e-07 3.0756e-09 2377.04 3121.39 -0.0563646 0.482179 0.277381 0.253646 -0.593294 -0.16955 0.493496 -0.266586 -0.226919 2.282 1 0 296.995 0 2.18206 2.28 0.000299514 0.857472 0.683772 0.334254 0.425636 2.18225 136.335 83.8511 18.7169 60.8329 0.00402816 0 -40 10
1.381 3.9974e-08 2.53941e-06 0.132814 0.132813 0.0120316 1.817e-05 0.00115428 0.166018 0.000658559 0.166672 0.918807 101.646 0.238912 0.805993 4.3538 0.0610878 0.0410736 0.958926 0.0196251 0.00444423 0.0188864 0.00425394 0.00537487 0.00611357 0.214995 0.244543 58.0258 -87.8977 126.23 15.949 145.028 0.000141489 0.267244 192.788 0.310351 0.0673446 0.00409735 0.000562129 0.00138429 0.98697 0.991722 -2.98454e-06 -85.6605 0.0930528 31177.4 306.005 0.983505 0.319146 0.733975 0.73397 9.99958 2.98462e-06 1.19384e-05 0.132698 0.983201 0.931675 -0.0132921 4.91951e-06 0.509369 -1.95917e-20 7.251e-24 -1.95844e-20 0.00139603 0.997816 8.59928e-05 0.152675 2.85244 0.00139603 0.997817 0.760706 0.00106119 0.00188084 0.000859928 0.455471 0.00188083 0.442334 0.000130289 1.02 0.888354 0.534492 0.286986 1.71844e-07 3.07562e-09 2377.02 3121.43 -0.0563687 0.48218 0.27738 0.253648 -0.593294 -0.16955 0.493483 -0.266584 -0.226908 2.283 1 0 296.991 0 2.1822 2.281 0.000299513 0.857493 0.683817 0.334194 0.42566 2.18239 136.343 83.8507 18.7169 60.8327 0.00402818 0 -40 10
1.382 4.00029e-08 2.53941e-06 0.132859 0.132858 0.0120315 1.81831e-05 0.00115428 0.166073 0.000658559 0.166727 0.91889 101.646 0.238902 0.806117 4.35426 0.0610978 0.0410779 0.958922 0.0196247 0.00444459 0.018886 0.00425426 0.00537532 0.00611403 0.215013 0.244561 58.0258 -87.8978 126.23 15.949 145.028 0.000141491 0.267244 192.788 0.310351 0.0673445 0.00409736 0.00056213 0.00138429 0.98697 0.991722 -2.98455e-06 -85.6605 0.0930529 31177.4 306.015 0.983505 0.319146 0.733984 0.733979 9.99958 2.98462e-06 1.19384e-05 0.132701 0.983201 0.931674 -0.0132921 4.91953e-06 0.509384 -1.9593e-20 7.25152e-24 -1.95857e-20 0.00139603 0.997816 8.59929e-05 0.152675 2.85245 0.00139603 0.997817 0.760789 0.00106121 0.00188084 0.000859929 0.455471 0.00188084 0.44234 0.000130292 1.02 0.888355 0.534492 0.286987 1.71845e-07 3.07565e-09 2377 3121.46 -0.0563727 0.48218 0.27738 0.25365 -0.593293 -0.16955 0.49347 -0.266581 -0.226898 2.284 1 0 296.988 0 2.18235 2.282 0.000299512 0.857514 0.683861 0.334134 0.425683 2.18254 136.35 83.8503 18.7168 60.8325 0.0040282 0 -40 10
1.383 4.00318e-08 2.53941e-06 0.132903 0.132902 0.0120315 1.81963e-05 0.00115428 0.166129 0.00065856 0.166783 0.918973 101.645 0.238892 0.806242 4.35471 0.0611078 0.0410822 0.958918 0.0196242 0.00444496 0.0188855 0.00425457 0.00537577 0.00611448 0.215031 0.244579 58.0259 -87.8978 126.23 15.9489 145.028 0.000141493 0.267244 192.788 0.310351 0.0673445 0.00409736 0.000562131 0.00138429 0.98697 0.991722 -2.98457e-06 -85.6605 0.093053 31177.3 306.025 0.983505 0.319146 0.733993 0.733988 9.99958 2.98463e-06 1.19384e-05 0.132705 0.983202 0.931674 -0.0132921 4.91956e-06 0.5094 -1.95942e-20 7.25205e-24 -1.9587e-20 0.00139603 0.997816 8.59929e-05 0.152675 2.85245 0.00139603 0.997817 0.760872 0.00106123 0.00188084 0.000859929 0.45547 0.00188084 0.442347 0.000130294 1.02 0.888356 0.534491 0.286989 1.71845e-07 3.07567e-09 2376.99 3121.5 -0.0563768 0.48218 0.27738 0.253653 -0.593293 -0.16955 0.493456 -0.266579 -0.226887 2.285 1 0 296.984 0 2.18249 2.283 0.000299511 0.857535 0.683906 0.334073 0.425706 2.18268 136.358 83.8498 18.7168 60.8322 0.00402822 0 -40 10
1.384 4.00607e-08 2.53941e-06 0.132948 0.132947 0.0120315 1.82094e-05 0.00115428 0.166185 0.000658561 0.166839 0.919057 101.645 0.238882 0.806366 4.35517 0.0611178 0.0410865 0.958914 0.0196238 0.00444532 0.0188851 0.00425488 0.00537622 0.00611494 0.215049 0.244598 58.026 -87.8978 126.23 15.9489 145.028 0.000141494 0.267245 192.788 0.31035 0.0673444 0.00409736 0.000562131 0.00138429 0.98697 0.991722 -2.98458e-06 -85.6605 0.093053 31177.3 306.035 0.983505 0.319146 0.734001 0.733997 9.99958 2.98463e-06 1.19384e-05 0.132709 0.983203 0.931673 -0.0132921 4.91959e-06 0.509416 -1.95955e-20 7.25257e-24 -1.95883e-20 0.00139603 0.997816 8.5993e-05 0.152675 2.85245 0.00139603 0.997817 0.760955 0.00106125 0.00188084 0.00085993 0.45547 0.00188084 0.442353 0.000130297 1.02 0.888357 0.534491 0.286991 1.71845e-07 3.07569e-09 2376.97 3121.54 -0.0563808 0.48218 0.27738 0.253655 -0.593292 -0.16955 0.493443 -0.266577 -0.226876 2.286 1 0 296.98 0 2.18263 2.284 0.00029951 0.857556 0.68395 0.334013 0.42573 2.18282 136.366 83.8494 18.7168 60.832 0.00402824 0 -40 10
1.385 4.00896e-08 2.53941e-06 0.132992 0.132991 0.0120315 1.82225e-05 0.00115428 0.16624 0.000658562 0.166894 0.91914 101.644 0.238872 0.806491 4.35562 0.0611279 0.0410908 0.958909 0.0196233 0.00444569 0.0188846 0.00425519 0.00537667 0.0061154 0.215067 0.244616 58.026 -87.8978 126.23 15.9488 145.028 0.000141496 0.267245 192.788 0.31035 0.0673444 0.00409737 0.000562132 0.00138429 0.98697 0.991722 -2.9846e-06 -85.6605 0.0930531 31177.3 306.045 0.983505 0.319146 0.73401 0.734006 9.99958 2.98464e-06 1.19384e-05 0.132713 0.983204 0.931672 -0.0132921 4.91962e-06 0.509431 -1.95968e-20 7.25309e-24 -1.95896e-20 0.00139603 0.997816 8.59931e-05 0.152675 2.85245 0.00139603 0.997817 0.761038 0.00106126 0.00188084 0.000859931 0.45547 0.00188084 0.442359 0.0001303 1.02 0.888358 0.534491 0.286992 1.71845e-07 3.07572e-09 2376.95 3121.57 -0.0563849 0.48218 0.277379 0.253658 -0.593292 -0.16955 0.49343 -0.266575 -0.226865 2.287 1 0 296.977 0 2.18277 2.285 0.000299509 0.857577 0.683995 0.333953 0.425753 2.18296 136.373 83.8489 18.7167 60.8318 0.00402825 0 -40 10
1.386 4.01184e-08 2.53941e-06 0.133037 0.133036 0.0120315 1.82357e-05 0.00115428 0.166296 0.000658563 0.16695 0.919223 101.644 0.238862 0.806616 4.35608 0.0611379 0.0410951 0.958905 0.0196229 0.00444605 0.0188841 0.00425551 0.00537712 0.00611586 0.215085 0.244634 58.0261 -87.8978 126.229 15.9488 145.028 0.000141498 0.267245 192.787 0.310349 0.0673443 0.00409737 0.000562133 0.0013843 0.98697 0.991722 -2.98461e-06 -85.6605 0.0930532 31177.3 306.055 0.983505 0.319146 0.734019 0.734015 9.99958 2.98464e-06 1.19385e-05 0.132716 0.983205 0.931672 -0.0132921 4.91965e-06 0.509447 -1.95981e-20 7.25361e-24 -1.95909e-20 0.00139604 0.997816 8.59932e-05 0.152675 2.85245 0.00139604 0.997817 0.761121 0.00106128 0.00188084 0.000859932 0.45547 0.00188084 0.442365 0.000130302 1.02 0.888359 0.53449 0.286994 1.71846e-07 3.07574e-09 2376.94 3121.61 -0.056389 0.48218 0.277379 0.25366 -0.593292 -0.16955 0.493417 -0.266573 -0.226854 2.288 1 0 296.973 0 2.18291 2.286 0.000299508 0.857598 0.684039 0.333893 0.425776 2.1831 136.381 83.8485 18.7167 60.8316 0.00402827 0 -40 10
1.387 4.01473e-08 2.53942e-06 0.133081 0.13308 0.0120315 1.82488e-05 0.00115428 0.166351 0.000658564 0.167005 0.919307 101.643 0.238852 0.80674 4.35654 0.0611479 0.0410994 0.958901 0.0196224 0.00444642 0.0188837 0.00425582 0.00537757 0.00611632 0.215103 0.244653 58.0262 -87.8978 126.229 15.9488 145.028 0.000141499 0.267245 192.787 0.310349 0.0673443 0.00409737 0.000562133 0.0013843 0.98697 0.991722 -2.98463e-06 -85.6605 0.0930533 31177.3 306.065 0.983505 0.319146 0.734028 0.734024 9.99958 2.98465e-06 1.19385e-05 0.13272 0.983206 0.931671 -0.0132921 4.91968e-06 0.509463 -1.95994e-20 7.25413e-24 -1.95922e-20 0.00139604 0.997816 8.59933e-05 0.152676 2.85245 0.00139604 0.997817 0.761204 0.0010613 0.00188084 0.000859933 0.45547 0.00188084 0.442372 0.000130305 1.02 0.88836 0.53449 0.286995 1.71846e-07 3.07576e-09 2376.92 3121.65 -0.0563931 0.48218 0.277379 0.253662 -0.593291 -0.16955 0.493404 -0.266571 -0.226842 2.289 1 0 296.97 0 2.18306 2.287 0.000299507 0.857619 0.684084 0.333833 0.425799 2.18325 136.388 83.8481 18.7167 60.8314 0.00402829 0 -40 10
1.388 4.01762e-08 2.53942e-06 0.133125 0.133125 0.0120315 1.82619e-05 0.00115428 0.166407 0.000658565 0.167061 0.91939 101.643 0.238842 0.806865 4.35699 0.0611579 0.0411037 0.958896 0.019622 0.00444679 0.0188832 0.00425613 0.00537802 0.00611678 0.215121 0.244671 58.0262 -87.8978 126.229 15.9487 145.028 0.000141501 0.267245 192.787 0.310348 0.0673442 0.00409737 0.000562134 0.0013843 0.98697 0.991722 -2.98464e-06 -85.6605 0.0930534 31177.2 306.075 0.983505 0.319146 0.734037 0.734033 9.99958 2.98465e-06 1.19385e-05 0.132724 0.983207 0.93167 -0.0132921 4.91971e-06 0.509479 -1.96007e-20 7.25466e-24 -1.95934e-20 0.00139604 0.997816 8.59933e-05 0.152676 2.85245 0.00139604 0.997817 0.761287 0.00106132 0.00188085 0.000859933 0.455469 0.00188084 0.442378 0.000130308 1.02 0.888361 0.53449 0.286997 1.71846e-07 3.07579e-09 2376.9 3121.68 -0.0563971 0.48218 0.277378 0.253665 -0.593291 -0.16955 0.493391 -0.266569 -0.226831 2.29 1 0 296.966 0 2.1832 2.288 0.000299507 0.85764 0.684128 0.333773 0.425823 2.18339 136.396 83.8476 18.7167 60.8312 0.00402831 0 -40 10
1.389 4.02051e-08 2.53942e-06 0.13317 0.133169 0.0120314 1.8275e-05 0.00115428 0.166462 0.000658565 0.167116 0.919473 101.643 0.238832 0.80699 4.35745 0.061168 0.041108 0.958892 0.0196215 0.00444715 0.0188828 0.00425644 0.00537848 0.00611723 0.215139 0.244689 58.0263 -87.8978 126.229 15.9487 145.028 0.000141503 0.267246 192.787 0.310348 0.0673442 0.00409738 0.000562135 0.0013843 0.98697 0.991722 -2.98466e-06 -85.6605 0.0930535 31177.2 306.085 0.983505 0.319146 0.734046 0.734042 9.99958 2.98465e-06 1.19385e-05 0.132728 0.983208 0.93167 -0.0132921 4.91974e-06 0.509494 -1.9602e-20 7.25518e-24 -1.95947e-20 0.00139604 0.997816 8.59934e-05 0.152676 2.85245 0.00139604 0.997817 0.76137 0.00106133 0.00188085 0.000859934 0.455469 0.00188085 0.442384 0.000130311 1.02 0.888362 0.534489 0.286998 1.71846e-07 3.07581e-09 2376.89 3121.72 -0.0564012 0.48218 0.277378 0.253667 -0.59329 -0.16955 0.493378 -0.266567 -0.22682 2.291 1 0 296.962 0 2.18334 2.289 0.000299506 0.857661 0.684173 0.333713 0.425846 2.18353 136.404 83.8472 18.7166 60.831 0.00402833 0 -40 10
1.39 4.0234e-08 2.53942e-06 0.133214 0.133213 0.0120314 1.82882e-05 0.00115428 0.166518 0.000658566 0.167172 0.919557 101.642 0.238822 0.807114 4.35791 0.061178 0.0411124 0.958888 0.0196211 0.00444752 0.0188823 0.00425676 0.00537893 0.00611769 0.215157 0.244708 58.0263 -87.8978 126.229 15.9487 145.028 0.000141505 0.267246 192.787 0.310348 0.0673441 0.00409738 0.000562135 0.00138431 0.98697 0.991722 -2.98467e-06 -85.6604 0.0930536 31177.2 306.095 0.983505 0.319146 0.734055 0.73405 9.99958 2.98466e-06 1.19385e-05 0.132731 0.983209 0.931669 -0.0132921 4.91977e-06 0.50951 -1.96033e-20 7.2557e-24 -1.9596e-20 0.00139604 0.997816 8.59935e-05 0.152676 2.85245 0.00139604 0.997816 0.761453 0.00106135 0.00188085 0.000859935 0.455469 0.00188085 0.44239 0.000130313 1.02 0.888364 0.534489 0.287 1.71847e-07 3.07583e-09 2376.87 3121.76 -0.0564053 0.48218 0.277378 0.25367 -0.59329 -0.16955 0.493364 -0.266565 -0.226809 2.292 1 0 296.959 0 2.18348 2.29 0.000299505 0.857683 0.684217 0.333653 0.425869 2.18367 136.411 83.8467 18.7166 60.8308 0.00402835 0 -40 10
1.391 4.02628e-08 2.53942e-06 0.133258 0.133258 0.0120314 1.83013e-05 0.00115428 0.166573 0.000658567 0.167227 0.91964 101.642 0.238812 0.807239 4.35837 0.061188 0.0411167 0.958883 0.0196206 0.00444789 0.0188818 0.00425707 0.00537938 0.00611816 0.215175 0.244726 58.0264 -87.8978 126.229 15.9486 145.028 0.000141506 0.267246 192.787 0.310347 0.0673441 0.00409738 0.000562136 0.00138431 0.98697 0.991722 -2.98469e-06 -85.6604 0.0930537 31177.2 306.105 0.983505 0.319146 0.734064 0.734059 9.99958 2.98466e-06 1.19386e-05 0.132735 0.98321 0.931669 -0.0132921 4.9198e-06 0.509526 -1.96046e-20 7.25622e-24 -1.95973e-20 0.00139604 0.997816 8.59936e-05 0.152676 2.85245 0.00139604 0.997816 0.761536 0.00106137 0.00188085 0.000859936 0.455469 0.00188085 0.442396 0.000130316 1.02 0.888365 0.534489 0.287001 1.71847e-07 3.07585e-09 2376.85 3121.8 -0.0564094 0.48218 0.277378 0.253672 -0.593289 -0.16955 0.493351 -0.266562 -0.226798 2.293 1 0 296.955 0 2.18362 2.291 0.000299504 0.857704 0.684262 0.333593 0.425893 2.18381 136.419 83.8463 18.7166 60.8305 0.00402836 0 -40 10
1.392 4.02917e-08 2.53942e-06 0.133303 0.133302 0.0120314 1.83144e-05 0.00115428 0.166628 0.000658568 0.167282 0.919723 101.641 0.238802 0.807364 4.35883 0.0611981 0.041121 0.958879 0.0196202 0.00444826 0.0188814 0.00425739 0.00537983 0.00611862 0.215193 0.244745 58.0265 -87.8978 126.228 15.9486 145.029 0.000141508 0.267246 192.786 0.310347 0.067344 0.00409739 0.000562137 0.00138431 0.98697 0.991722 -2.9847e-06 -85.6604 0.0930537 31177.1 306.115 0.983505 0.319146 0.734073 0.734068 9.99958 2.98467e-06 1.19386e-05 0.132739 0.983211 0.931668 -0.0132921 4.91983e-06 0.509542 -1.96059e-20 7.25675e-24 -1.95986e-20 0.00139604 0.997816 8.59937e-05 0.152676 2.85246 0.00139604 0.997816 0.761619 0.00106139 0.00188085 0.000859937 0.455468 0.00188085 0.442403 0.000130319 1.02 0.888366 0.534488 0.287003 1.71847e-07 3.07588e-09 2376.84 3121.83 -0.0564135 0.48218 0.277377 0.253674 -0.593289 -0.169551 0.493338 -0.26656 -0.226787 2.294 1 0 296.951 0 2.18377 2.292 0.000299503 0.857725 0.684306 0.333534 0.425916 2.18396 136.427 83.8459 18.7166 60.8303 0.00402838 0 -40 10
1.393 4.03206e-08 2.53942e-06 0.133347 0.133346 0.0120314 1.83275e-05 0.00115428 0.166683 0.000658569 0.167337 0.919807 101.641 0.238792 0.807489 4.35929 0.0612081 0.0411254 0.958875 0.0196197 0.00444862 0.0188809 0.0042577 0.00538029 0.00611908 0.215211 0.244763 58.0265 -87.8978 126.228 15.9485 145.029 0.00014151 0.267246 192.786 0.310346 0.067344 0.00409739 0.000562137 0.00138431 0.986969 0.991722 -2.98472e-06 -85.6604 0.0930538 31177.1 306.125 0.983505 0.319146 0.734082 0.734077 9.99958 2.98467e-06 1.19386e-05 0.132743 0.983212 0.931667 -0.0132921 4.91986e-06 0.509557 -1.96072e-20 7.25727e-24 -1.95999e-20 0.00139604 0.997816 8.59937e-05 0.152676 2.85246 0.00139604 0.997816 0.761701 0.0010614 0.00188085 0.000859937 0.455468 0.00188085 0.442409 0.000130321 1.02 0.888367 0.534488 0.287004 1.71847e-07 3.0759e-09 2376.82 3121.87 -0.0564176 0.48218 0.277377 0.253677 -0.593288 -0.169551 0.493325 -0.266558 -0.226776 2.295 1 0 296.948 0 2.18391 2.293 0.000299502 0.857747 0.684351 0.333474 0.425939 2.1841 136.434 83.8454 18.7165 60.8301 0.0040284 0 -40 10
1.394 4.03495e-08 2.53942e-06 0.133391 0.13339 0.0120314 1.83407e-05 0.00115428 0.166739 0.00065857 0.167393 0.91989 101.64 0.238782 0.807614 4.35975 0.0612182 0.0411297 0.95887 0.0196193 0.00444899 0.0188805 0.00425802 0.00538074 0.00611954 0.21523 0.244782 58.0266 -87.8978 126.228 15.9485 145.029 0.000141511 0.267246 192.786 0.310346 0.0673439 0.00409739 0.000562138 0.00138431 0.986969 0.991722 -2.98473e-06 -85.6604 0.0930539 31177.1 306.135 0.983505 0.319146 0.734091 0.734086 9.99958 2.98468e-06 1.19386e-05 0.132746 0.983213 0.931667 -0.0132921 4.91989e-06 0.509573 -1.96085e-20 7.2578e-24 -1.96012e-20 0.00139604 0.997816 8.59938e-05 0.152677 2.85246 0.00139604 0.997816 0.761784 0.00106142 0.00188086 0.000859938 0.455468 0.00188085 0.442415 0.000130324 1.02 0.888368 0.534488 0.287006 1.71848e-07 3.07592e-09 2376.8 3121.91 -0.0564217 0.482181 0.277377 0.253679 -0.593288 -0.169551 0.493312 -0.266556 -0.226765 2.296 1 0 296.944 0 2.18405 2.294 0.000299501 0.857768 0.684395 0.333415 0.425963 2.18424 136.442 83.845 18.7165 60.8299 0.00402842 0 -40 10
1.395 4.03784e-08 2.53943e-06 0.133435 0.133434 0.0120314 1.83538e-05 0.00115428 0.166794 0.000658571 0.167448 0.919974 101.64 0.238772 0.807739 4.36021 0.0612282 0.041134 0.958866 0.0196188 0.00444936 0.01888 0.00425833 0.00538119 0.00612 0.215248 0.2448 58.0267 -87.8978 126.228 15.9485 145.029 0.000141513 0.267247 192.786 0.310345 0.0673439 0.0040974 0.000562139 0.00138432 0.986969 0.991722 -2.98475e-06 -85.6604 0.093054 31177.1 306.145 0.983505 0.319146 0.7341 0.734095 9.99958 2.98468e-06 1.19386e-05 0.13275 0.983214 0.931666 -0.0132921 4.91992e-06 0.509589 -1.96098e-20 7.25832e-24 -1.96025e-20 0.00139605 0.997816 8.59939e-05 0.152677 2.85246 0.00139605 0.997816 0.761867 0.00106144 0.00188086 0.000859939 0.455468 0.00188086 0.442421 0.000130327 1.02 0.888369 0.534487 0.287007 1.71848e-07 3.07595e-09 2376.79 3121.95 -0.0564258 0.482181 0.277377 0.253682 -0.593287 -0.169551 0.493298 -0.266554 -0.226754 2.297 1 0 296.94 0 2.18419 2.295 0.0002995 0.857789 0.68444 0.333356 0.425986 2.18438 136.449 83.8445 18.7165 60.8297 0.00402844 0 -40 10
1.396 4.04072e-08 2.53943e-06 0.133479 0.133478 0.0120313 1.83669e-05 0.00115428 0.166849 0.000658572 0.167503 0.920057 101.639 0.238762 0.807863 4.36067 0.0612383 0.0411384 0.958862 0.0196184 0.00444973 0.0188795 0.00425864 0.00538165 0.00612046 0.215266 0.244818 58.0267 -87.8978 126.228 15.9484 145.029 0.000141515 0.267247 192.786 0.310345 0.0673438 0.0040974 0.000562139 0.00138432 0.986969 0.991722 -2.98476e-06 -85.6604 0.0930541 31177 306.155 0.983505 0.319146 0.734109 0.734104 9.99958 2.98469e-06 1.19387e-05 0.132754 0.983214 0.931666 -0.0132921 4.91995e-06 0.509605 -1.96111e-20 7.25885e-24 -1.96038e-20 0.00139605 0.997816 8.5994e-05 0.152677 2.85246 0.00139605 0.997816 0.76195 0.00106146 0.00188086 0.00085994 0.455468 0.00188086 0.442428 0.000130329 1.02 0.88837 0.534487 0.287009 1.71848e-07 3.07597e-09 2376.77 3121.98 -0.0564299 0.482181 0.277376 0.253684 -0.593287 -0.169551 0.493285 -0.266552 -0.226743 2.298 1 0 296.937 0 2.18433 2.296 0.000299499 0.857811 0.684484 0.333296 0.426009 2.18452 136.457 83.8441 18.7165 60.8295 0.00402846 0 -40 10
1.397 4.04361e-08 2.53943e-06 0.133523 0.133522 0.0120313 1.838e-05 0.00115429 0.166904 0.000658572 0.167558 0.920141 101.639 0.238752 0.807988 4.36113 0.0612483 0.0411427 0.958857 0.0196179 0.0044501 0.0188791 0.00425896 0.0053821 0.00612092 0.215284 0.244837 58.0268 -87.8978 126.228 15.9484 145.029 0.000141517 0.267247 192.786 0.310345 0.0673438 0.0040974 0.00056214 0.00138432 0.986969 0.991722 -2.98478e-06 -85.6604 0.0930542 31177 306.165 0.983505 0.319146 0.734118 0.734114 9.99958 2.98469e-06 1.19387e-05 0.132758 0.983215 0.931665 -0.0132921 4.91998e-06 0.509621 -1.96124e-20 7.25937e-24 -1.96051e-20 0.00139605 0.997816 8.59941e-05 0.152677 2.85246 0.00139605 0.997816 0.762032 0.00106147 0.00188086 0.000859941 0.455467 0.00188086 0.442434 0.000130332 1.02 0.888371 0.534487 0.28701 1.71849e-07 3.07599e-09 2376.76 3122.02 -0.0564341 0.482181 0.277376 0.253687 -0.593286 -0.169551 0.493272 -0.26655 -0.226731 2.299 1 0 296.933 0 2.18448 2.297 0.000299499 0.857832 0.684529 0.333237 0.426032 2.18467 136.465 83.8436 18.7164 60.8293 0.00402847 0 -40 10
1.398 4.0465e-08 2.53943e-06 0.133567 0.133566 0.0120313 1.83932e-05 0.00115429 0.166959 0.000658573 0.167613 0.920225 101.638 0.238742 0.808113 4.36159 0.0612584 0.0411471 0.958853 0.0196174 0.00445047 0.0188786 0.00425928 0.00538256 0.00612139 0.215302 0.244855 58.0269 -87.8978 126.227 15.9484 145.029 0.000141518 0.267247 192.785 0.310344 0.0673437 0.00409741 0.000562141 0.00138432 0.986969 0.991722 -2.98479e-06 -85.6604 0.0930543 31177 306.175 0.983505 0.319146 0.734127 0.734123 9.99958 2.9847e-06 1.19387e-05 0.132761 0.983216 0.931664 -0.0132921 4.92001e-06 0.509637 -1.96137e-20 7.2599e-24 -1.96064e-20 0.00139605 0.997816 8.59941e-05 0.152677 2.85246 0.00139605 0.997816 0.762115 0.00106149 0.00188086 0.000859941 0.455467 0.00188086 0.44244 0.000130335 1.02 0.888372 0.534487 0.287012 1.71849e-07 3.07601e-09 2376.74 3122.06 -0.0564382 0.482181 0.277376 0.253689 -0.593286 -0.169551 0.493259 -0.266548 -0.22672 2.3 1 0 296.929 0 2.18462 2.298 0.000299498 0.857854 0.684573 0.333178 0.426056 2.18481 136.472 83.8432 18.7164 60.829 0.00402849 0 -40 10
1.399 4.04939e-08 2.53943e-06 0.133611 0.13361 0.0120313 1.84063e-05 0.00115429 0.167014 0.000658574 0.167668 0.920308 101.638 0.238732 0.808238 4.36205 0.0612684 0.0411514 0.958849 0.019617 0.00445084 0.0188781 0.00425959 0.00538301 0.00612185 0.21532 0.244874 58.0269 -87.8978 126.227 15.9483 145.029 0.00014152 0.267247 192.785 0.310344 0.0673436 0.00409741 0.000562141 0.00138433 0.986969 0.991722 -2.98481e-06 -85.6604 0.0930544 31177 306.185 0.983505 0.319146 0.734136 0.734132 9.99958 2.9847e-06 1.19387e-05 0.132765 0.983217 0.931664 -0.0132921 4.92004e-06 0.509652 -1.9615e-20 7.26042e-24 -1.96077e-20 0.00139605 0.997816 8.59942e-05 0.152677 2.85246 0.00139605 0.997816 0.762198 0.00106151 0.00188086 0.000859942 0.455467 0.00188086 0.442446 0.000130338 1.02 0.888373 0.534486 0.287013 1.71849e-07 3.07604e-09 2376.72 3122.1 -0.0564423 0.482181 0.277375 0.253692 -0.593285 -0.169551 0.493245 -0.266546 -0.226709 2.301 1 0 296.926 0 2.18476 2.299 0.000299497 0.857875 0.684618 0.333119 0.426079 2.18495 136.48 83.8427 18.7164 60.8288 0.00402851 0 -40 10
1.4 4.05227e-08 2.53943e-06 0.133655 0.133654 0.0120313 1.84194e-05 0.00115429 0.167069 0.000658575 0.167723 0.920392 101.637 0.238722 0.808363 4.36252 0.0612785 0.0411558 0.958844 0.0196165 0.00445121 0.0188777 0.00425991 0.00538347 0.00612231 0.215339 0.244893 58.027 -87.8978 126.227 15.9483 145.029 0.000141522 0.267248 192.785 0.310343 0.0673436 0.00409741 0.000562142 0.00138433 0.986969 0.991722 -2.98482e-06 -85.6604 0.0930544 31177 306.195 0.983505 0.319146 0.734145 0.734141 9.99958 2.98471e-06 1.19387e-05 0.132769 0.983218 0.931663 -0.0132921 4.92007e-06 0.509668 -1.96163e-20 7.26095e-24 -1.9609e-20 0.00139605 0.997816 8.59943e-05 0.152678 2.85246 0.00139605 0.997816 0.76228 0.00106152 0.00188086 0.000859943 0.455467 0.00188086 0.442452 0.00013034 1.02 0.888375 0.534486 0.287015 1.71849e-07 3.07606e-09 2376.71 3122.14 -0.0564464 0.482181 0.277375 0.253694 -0.593285 -0.169551 0.493232 -0.266543 -0.226698 2.302 1 0 296.922 0 2.1849 2.3 0.000299496 0.857897 0.684662 0.33306 0.426102 2.18509 136.487 83.8423 18.7164 60.8286 0.00402853 0 -40 10
1.401 4.05516e-08 2.53943e-06 0.133699 0.133698 0.0120313 1.84326e-05 0.00115429 0.167124 0.000658576 0.167778 0.920475 101.637 0.238711 0.808488 4.36298 0.0612885 0.0411602 0.95884 0.0196161 0.00445158 0.0188772 0.00426022 0.00538392 0.00612278 0.215357 0.244911 58.027 -87.8978 126.227 15.9482 145.029 0.000141524 0.267248 192.785 0.310343 0.0673435 0.00409741 0.000562143 0.00138433 0.986969 0.991722 -2.98484e-06 -85.6603 0.0930545 31176.9 306.205 0.983505 0.319146 0.734154 0.73415 9.99958 2.98471e-06 1.19388e-05 0.132773 0.983219 0.931662 -0.0132921 4.9201e-06 0.509684 -1.96176e-20 7.26148e-24 -1.96103e-20 0.00139605 0.997816 8.59944e-05 0.152678 2.85246 0.00139605 0.997816 0.762363 0.00106154 0.00188087 0.000859944 0.455466 0.00188086 0.442459 0.000130343 1.02 0.888376 0.534486 0.287016 1.7185e-07 3.07608e-09 2376.69 3122.17 -0.0564506 0.482181 0.277375 0.253696 -0.593284 -0.169551 0.493219 -0.266541 -0.226687 2.303 1 0 296.918 0 2.18504 2.301 0.000299495 0.857919 0.684707 0.333001 0.426125 2.18523 136.495 83.8418 18.7163 60.8284 0.00402855 0 -40 10
1.402 4.05805e-08 2.53943e-06 0.133743 0.133742 0.0120313 1.84457e-05 0.00115429 0.167179 0.000658577 0.167833 0.920559 101.637 0.238701 0.808614 4.36344 0.0612986 0.0411646 0.958835 0.0196156 0.00445195 0.0188768 0.00426054 0.00538438 0.00612324 0.215375 0.24493 58.0271 -87.8978 126.227 15.9482 145.029 0.000141525 0.267248 192.785 0.310342 0.0673435 0.00409742 0.000562143 0.00138433 0.986969 0.991722 -2.98485e-06 -85.6603 0.0930546 31176.9 306.215 0.983505 0.319146 0.734163 0.734159 9.99958 2.98472e-06 1.19388e-05 0.132776 0.98322 0.931662 -0.0132921 4.92013e-06 0.5097 -1.96189e-20 7.262e-24 -1.96116e-20 0.00139605 0.997816 8.59945e-05 0.152678 2.85246 0.00139605 0.997816 0.762445 0.00106156 0.00188087 0.000859945 0.455466 0.00188087 0.442465 0.000130346 1.02 0.888377 0.534485 0.287018 1.7185e-07 3.07611e-09 2376.67 3122.21 -0.0564547 0.482181 0.277375 0.253699 -0.593284 -0.169551 0.493205 -0.266539 -0.226675 2.304 1 0 296.915 0 2.18519 2.302 0.000299494 0.85794 0.684751 0.332942 0.426149 2.18538 136.503 83.8414 18.7163 60.8282 0.00402857 0 -40 10
1.403 4.06094e-08 2.53943e-06 0.133787 0.133786 0.0120313 1.84588e-05 0.00115429 0.167233 0.000658577 0.167887 0.920643 101.636 0.238691 0.808739 4.36391 0.0613087 0.0411689 0.958831 0.0196152 0.00445232 0.0188763 0.00426086 0.00538483 0.00612371 0.215393 0.244948 58.0272 -87.8978 126.227 15.9482 145.029 0.000141527 0.267248 192.785 0.310342 0.0673434 0.00409742 0.000562144 0.00138433 0.986969 0.991722 -2.98487e-06 -85.6603 0.0930547 31176.9 306.225 0.983505 0.319146 0.734173 0.734168 9.99958 2.98472e-06 1.19388e-05 0.13278 0.983221 0.931661 -0.0132921 4.92016e-06 0.509716 -1.96202e-20 7.26253e-24 -1.96129e-20 0.00139606 0.997816 8.59946e-05 0.152678 2.85247 0.00139606 0.997816 0.762528 0.00106158 0.00188087 0.000859946 0.455466 0.00188087 0.442471 0.000130348 1.02 0.888378 0.534485 0.287019 1.7185e-07 3.07613e-09 2376.66 3122.25 -0.0564589 0.482181 0.277374 0.253701 -0.593283 -0.169551 0.493192 -0.266537 -0.226664 2.305 1 0 296.911 0 2.18533 2.303 0.000299493 0.857962 0.684796 0.332883 0.426172 2.18552 136.51 83.8409 18.7163 60.828 0.00402859 0 -40 10
1.404 4.06383e-08 2.53944e-06 0.133831 0.13383 0.0120312 1.84719e-05 0.00115429 0.167288 0.000658578 0.167942 0.920726 101.636 0.238681 0.808864 4.36437 0.0613187 0.0411733 0.958827 0.0196147 0.00445269 0.0188758 0.00426117 0.00538529 0.00612417 0.215412 0.244967 58.0272 -87.8978 126.226 15.9481 145.029 0.000141529 0.267248 192.784 0.310342 0.0673434 0.00409742 0.000562145 0.00138434 0.986969 0.991722 -2.98488e-06 -85.6603 0.0930548 31176.9 306.235 0.983505 0.319146 0.734182 0.734177 9.99958 2.98473e-06 1.19388e-05 0.132784 0.983222 0.931661 -0.0132921 4.92019e-06 0.509732 -1.96215e-20 7.26306e-24 -1.96142e-20 0.00139606 0.997816 8.59946e-05 0.152678 2.85247 0.00139606 0.997816 0.76261 0.00106159 0.00188087 0.000859946 0.455466 0.00188087 0.442477 0.000130351 1.02 0.888379 0.534485 0.287021 1.7185e-07 3.07615e-09 2376.64 3122.29 -0.056463 0.482181 0.277374 0.253704 -0.593283 -0.169551 0.493179 -0.266535 -0.226653 2.306 1 0 296.907 0 2.18547 2.304 0.000299492 0.857983 0.68484 0.332825 0.426195 2.18566 136.518 83.8405 18.7163 60.8277 0.0040286 0 -40 10
1.405 4.06671e-08 2.53944e-06 0.133874 0.133873 0.0120312 1.84851e-05 0.00115429 0.167343 0.000658579 0.167997 0.92081 101.635 0.238671 0.808989 4.36484 0.0613288 0.0411777 0.958822 0.0196143 0.00445306 0.0188754 0.00426149 0.00538575 0.00612464 0.21543 0.244985 58.0273 -87.8978 126.226 15.9481 145.029 0.000141531 0.267249 192.784 0.310341 0.0673433 0.00409743 0.000562145 0.00138434 0.986969 0.991722 -2.9849e-06 -85.6603 0.0930549 31176.8 306.245 0.983505 0.319146 0.734191 0.734186 9.99958 2.98473e-06 1.19388e-05 0.132788 0.983223 0.93166 -0.0132921 4.92022e-06 0.509748 -1.96228e-20 7.26359e-24 -1.96155e-20 0.00139606 0.997816 8.59947e-05 0.152678 2.85247 0.00139606 0.997816 0.762693 0.00106161 0.00188087 0.000859947 0.455466 0.00188087 0.442483 0.000130354 1.02 0.88838 0.534484 0.287022 1.71851e-07 3.07617e-09 2376.62 3122.33 -0.0564672 0.482181 0.277374 0.253706 -0.593282 -0.169551 0.493165 -0.266533 -0.226642 2.307 1 0 296.904 0 2.18561 2.305 0.000299491 0.858005 0.684884 0.332766 0.426218 2.1858 136.525 83.84 18.7162 60.8275 0.00402862 0 -40 10
1.406 4.0696e-08 2.53944e-06 0.133918 0.133917 0.0120312 1.84982e-05 0.00115429 0.167397 0.00065858 0.168051 0.920894 101.635 0.238661 0.809114 4.3653 0.0613389 0.0411821 0.958818 0.0196138 0.00445343 0.0188749 0.00426181 0.0053862 0.0061251 0.215448 0.245004 58.0274 -87.8978 126.226 15.9481 145.029 0.000141533 0.267249 192.784 0.310341 0.0673433 0.00409743 0.000562146 0.00138434 0.986969 0.991722 -2.98491e-06 -85.6603 0.093055 31176.8 306.255 0.983505 0.319146 0.7342 0.734196 9.99958 2.98474e-06 1.19388e-05 0.132792 0.983223 0.931659 -0.0132921 4.92025e-06 0.509764 -1.96241e-20 7.26412e-24 -1.96168e-20 0.00139606 0.997816 8.59948e-05 0.152678 2.85247 0.00139606 0.997816 0.762775 0.00106163 0.00188087 0.000859948 0.455465 0.00188087 0.44249 0.000130356 1.02 0.888381 0.534484 0.287024 1.71851e-07 3.0762e-09 2376.61 3122.36 -0.0564713 0.482181 0.277373 0.253709 -0.593282 -0.169551 0.493152 -0.266531 -0.22663 2.308 1 0 296.9 0 2.18575 2.306 0.00029949 0.858027 0.684929 0.332708 0.426242 2.18594 136.533 83.8396 18.7162 60.8273 0.00402864 0 -40 10
1.407 4.07249e-08 2.53944e-06 0.133962 0.133961 0.0120312 1.85113e-05 0.00115429 0.167452 0.000658581 0.168106 0.920978 101.634 0.238651 0.809239 4.36577 0.061349 0.0411865 0.958814 0.0196133 0.0044538 0.0188744 0.00426213 0.00538666 0.00612557 0.215466 0.245023 58.0274 -87.8978 126.226 15.948 145.029 0.000141534 0.267249 192.784 0.31034 0.0673432 0.00409743 0.000562147 0.00138434 0.986969 0.991722 -2.98493e-06 -85.6603 0.0930551 31176.8 306.265 0.983505 0.319146 0.734209 0.734205 9.99958 2.98474e-06 1.19389e-05 0.132795 0.983224 0.931659 -0.0132921 4.92028e-06 0.50978 -1.96254e-20 7.26464e-24 -1.96181e-20 0.00139606 0.997816 8.59949e-05 0.152679 2.85247 0.00139606 0.997816 0.762858 0.00106165 0.00188087 0.000859949 0.455465 0.00188087 0.442496 0.000130359 1.02 0.888382 0.534484 0.287026 1.71851e-07 3.07622e-09 2376.59 3122.4 -0.0564755 0.482182 0.277373 0.253711 -0.593281 -0.169551 0.493138 -0.266529 -0.226619 2.309 1 0 296.896 0 2.1859 2.307 0.00029949 0.858049 0.684973 0.332649 0.426265 2.18609 136.541 83.8391 18.7162 60.8271 0.00402866 0 -40 10
1.408 4.07538e-08 2.53944e-06 0.134005 0.134005 0.0120312 1.85244e-05 0.00115429 0.167507 0.000658582 0.168161 0.921061 101.634 0.238641 0.809365 4.36623 0.061359 0.0411909 0.958809 0.0196129 0.00445418 0.018874 0.00426244 0.00538712 0.00612603 0.215485 0.245041 58.0275 -87.8978 126.226 15.948 145.029 0.000141536 0.267249 192.784 0.31034 0.0673432 0.00409744 0.000562147 0.00138434 0.986969 0.991722 -2.98494e-06 -85.6603 0.0930551 31176.8 306.275 0.983505 0.319146 0.734218 0.734214 9.99958 2.98475e-06 1.19389e-05 0.132799 0.983225 0.931658 -0.0132921 4.92031e-06 0.509796 -1.96267e-20 7.26517e-24 -1.96194e-20 0.00139606 0.997816 8.5995e-05 0.152679 2.85247 0.00139606 0.997816 0.76294 0.00106166 0.00188088 0.00085995 0.455465 0.00188087 0.442502 0.000130362 1.02 0.888383 0.534483 0.287027 1.71852e-07 3.07624e-09 2376.57 3122.44 -0.0564797 0.482182 0.277373 0.253714 -0.593281 -0.169552 0.493125 -0.266527 -0.226608 2.31 1 0 296.893 0 2.18604 2.308 0.000299489 0.858071 0.685018 0.332591 0.426288 2.18623 136.548 83.8387 18.7162 60.8269 0.00402868 0 -40 10
1.409 4.07826e-08 2.53944e-06 0.134049 0.134048 0.0120312 1.85376e-05 0.00115429 0.167561 0.000658582 0.168215 0.921145 101.633 0.238631 0.80949 4.3667 0.0613691 0.0411953 0.958805 0.0196124 0.00445455 0.0188735 0.00426276 0.00538758 0.0061265 0.215503 0.24506 58.0275 -87.8979 126.226 15.9479 145.029 0.000141538 0.267249 192.784 0.310339 0.0673431 0.00409744 0.000562148 0.00138435 0.986969 0.991722 -2.98496e-06 -85.6603 0.0930552 31176.8 306.285 0.983505 0.319146 0.734228 0.734223 9.99958 2.98475e-06 1.19389e-05 0.132803 0.983226 0.931657 -0.0132921 4.92034e-06 0.509812 -1.9628e-20 7.2657e-24 -1.96207e-20 0.00139606 0.997816 8.5995e-05 0.152679 2.85247 0.00139606 0.997816 0.763022 0.00106168 0.00188088 0.00085995 0.455465 0.00188088 0.442508 0.000130364 1.02 0.888384 0.534483 0.287029 1.71852e-07 3.07627e-09 2376.56 3122.48 -0.0564838 0.482182 0.277373 0.253716 -0.59328 -0.169552 0.493112 -0.266524 -0.226596 2.311 1 0 296.889 0 2.18618 2.309 0.000299488 0.858092 0.685062 0.332532 0.426311 2.18637 136.556 83.8382 18.7161 60.8266 0.0040287 0 -40 10
1.41 4.08115e-08 2.53944e-06 0.134093 0.134092 0.0120312 1.85507e-05 0.00115429 0.167616 0.000658583 0.16827 0.921229 101.633 0.238621 0.809615 4.36717 0.0613792 0.0411997 0.9588 0.019612 0.00445492 0.018873 0.00426308 0.00538804 0.00612697 0.215521 0.245079 58.0276 -87.8979 126.225 15.9479 145.029 0.00014154 0.26725 192.783 0.310339 0.0673431 0.00409744 0.000562149 0.00138435 0.986969 0.991722 -2.98497e-06 -85.6603 0.0930553 31176.7 306.296 0.983504 0.319146 0.734237 0.734232 9.99958 2.98476e-06 1.19389e-05 0.132807 0.983227 0.931657 -0.0132921 4.92037e-06 0.509828 -1.96293e-20 7.26623e-24 -1.96221e-20 0.00139606 0.997816 8.59951e-05 0.152679 2.85247 0.00139606 0.997816 0.763104 0.0010617 0.00188088 0.000859951 0.455464 0.00188088 0.442514 0.000130367 1.02 0.888386 0.534483 0.28703 1.71852e-07 3.07629e-09 2376.54 3122.52 -0.056488 0.482182 0.277372 0.253719 -0.59328 -0.169552 0.493098 -0.266522 -0.226585 2.312 1 0 296.885 0 2.18632 2.31 0.000299487 0.858114 0.685107 0.332474 0.426334 2.18651 136.564 83.8377 18.7161 60.8264 0.00402872 0 -40 10
1.411 4.08404e-08 2.53944e-06 0.134136 0.134135 0.0120311 1.85638e-05 0.00115429 0.16767 0.000658584 0.168324 0.921313 101.632 0.238611 0.809741 4.36764 0.0613893 0.0412041 0.958796 0.0196115 0.00445529 0.0188726 0.0042634 0.0053885 0.00612743 0.21554 0.245097 58.0277 -87.8979 126.225 15.9479 145.029 0.000141541 0.26725 192.783 0.310339 0.067343 0.00409744 0.000562149 0.00138435 0.986969 0.991722 -2.98499e-06 -85.6602 0.0930554 31176.7 306.306 0.983504 0.319146 0.734246 0.734242 9.99958 2.98476e-06 1.19389e-05 0.132811 0.983228 0.931656 -0.0132921 4.9204e-06 0.509844 -1.96306e-20 7.26676e-24 -1.96234e-20 0.00139606 0.997816 8.59952e-05 0.152679 2.85247 0.00139606 0.997816 0.763187 0.00106172 0.00188088 0.000859952 0.455464 0.00188088 0.44252 0.00013037 1.02 0.888387 0.534483 0.287032 1.71852e-07 3.07631e-09 2376.52 3122.56 -0.0564922 0.482182 0.277372 0.253721 -0.593279 -0.169552 0.493085 -0.26652 -0.226574 2.313 1 0 296.881 0 2.18646 2.311 0.000299486 0.858136 0.685151 0.332416 0.426358 2.18665 136.571 83.8373 18.7161 60.8262 0.00402874 0 -40 10
1.412 4.08693e-08 2.53944e-06 0.13418 0.134179 0.0120311 1.85769e-05 0.00115429 0.167725 0.000658585 0.168379 0.921397 101.632 0.238601 0.809866 4.3681 0.0613994 0.0412085 0.958791 0.019611 0.00445567 0.0188721 0.00426372 0.00538896 0.0061279 0.215558 0.245116 58.0277 -87.8979 126.225 15.9478 145.029 0.000141543 0.26725 192.783 0.310338 0.067343 0.00409745 0.00056215 0.00138435 0.986969 0.991722 -2.985e-06 -85.6602 0.0930555 31176.7 306.316 0.983504 0.319146 0.734255 0.734251 9.99958 2.98477e-06 1.1939e-05 0.132814 0.983229 0.931655 -0.0132921 4.92043e-06 0.50986 -1.96319e-20 7.26729e-24 -1.96247e-20 0.00139607 0.997816 8.59953e-05 0.152679 2.85247 0.00139607 0.997816 0.763269 0.00106173 0.00188088 0.000859953 0.455464 0.00188088 0.442527 0.000130373 1.02 0.888388 0.534482 0.287033 1.71853e-07 3.07634e-09 2376.51 3122.6 -0.0564964 0.482182 0.277372 0.253724 -0.593279 -0.169552 0.493071 -0.266518 -0.226562 2.314 1 0 296.878 0 2.1866 2.312 0.000299485 0.858158 0.685195 0.332358 0.426381 2.18679 136.579 83.8368 18.716 60.826 0.00402875 0 -40 10
1.413 4.08981e-08 2.53945e-06 0.134223 0.134222 0.0120311 1.85901e-05 0.00115429 0.167779 0.000658586 0.168433 0.921481 101.631 0.238591 0.809992 4.36857 0.0614095 0.0412129 0.958787 0.0196106 0.00445604 0.0188716 0.00426404 0.00538941 0.00612837 0.215577 0.245135 58.0278 -87.8979 126.225 15.9478 145.029 0.000141545 0.26725 192.783 0.310338 0.0673429 0.00409745 0.000562151 0.00138436 0.986969 0.991722 -2.98502e-06 -85.6602 0.0930556 31176.7 306.326 0.983504 0.319146 0.734265 0.73426 9.99958 2.98477e-06 1.1939e-05 0.132818 0.98323 0.931655 -0.0132921 4.92045e-06 0.509876 -1.96333e-20 7.26782e-24 -1.9626e-20 0.00139607 0.997816 8.59954e-05 0.15268 2.85247 0.00139607 0.997816 0.763351 0.00106175 0.00188088 0.000859954 0.455464 0.00188088 0.442533 0.000130375 1.02 0.888389 0.534482 0.287035 1.71853e-07 3.07636e-09 2376.49 3122.63 -0.0565006 0.482182 0.277371 0.253726 -0.593278 -0.169552 0.493058 -0.266516 -0.226551 2.315 1 0 296.874 0 2.18675 2.313 0.000299484 0.85818 0.68524 0.3323 0.426404 2.18694 136.586 83.8364 18.716 60.8258 0.00402877 0 -40 10
1.414 4.0927e-08 2.53945e-06 0.134267 0.134266 0.0120311 1.86032e-05 0.00115429 0.167833 0.000658587 0.168487 0.921565 101.631 0.23858 0.810117 4.36904 0.0614196 0.0412174 0.958783 0.0196101 0.00445641 0.0188712 0.00426436 0.00538987 0.00612884 0.215595 0.245154 58.0279 -87.8979 126.225 15.9478 145.029 0.000141547 0.26725 192.783 0.310337 0.0673429 0.00409745 0.000562151 0.00138436 0.986969 0.991722 -2.98503e-06 -85.6602 0.0930557 31176.6 306.336 0.983504 0.319146 0.734274 0.734269 9.99958 2.98478e-06 1.1939e-05 0.132822 0.98323 0.931654 -0.0132921 4.92048e-06 0.509892 -1.96346e-20 7.26835e-24 -1.96273e-20 0.00139607 0.997816 8.59954e-05 0.15268 2.85248 0.00139607 0.997816 0.763433 0.00106177 0.00188089 0.000859954 0.455463 0.00188088 0.442539 0.000130378 1.02 0.88839 0.534482 0.287036 1.71853e-07 3.07638e-09 2376.47 3122.67 -0.0565048 0.482182 0.277371 0.253729 -0.593278 -0.169552 0.493044 -0.266514 -0.22654 2.316 1 0 296.87 0 2.18689 2.314 0.000299483 0.858202 0.685284 0.332242 0.426427 2.18708 136.594 83.8359 18.716 60.8255 0.00402879 0 -40 10
1.415 4.09559e-08 2.53945e-06 0.13431 0.134309 0.0120311 1.86163e-05 0.00115429 0.167887 0.000658587 0.168541 0.921649 101.63 0.23857 0.810242 4.36951 0.0614297 0.0412218 0.958778 0.0196097 0.00445679 0.0188707 0.00426468 0.00539033 0.00612931 0.215613 0.245172 58.0279 -87.8979 126.225 15.9477 145.029 0.000141549 0.267251 192.783 0.310337 0.0673428 0.00409746 0.000562152 0.00138436 0.986969 0.991722 -2.98505e-06 -85.6602 0.0930558 31176.6 306.346 0.983504 0.319146 0.734283 0.734279 9.99958 2.98478e-06 1.1939e-05 0.132826 0.983231 0.931653 -0.0132921 4.92051e-06 0.509908 -1.96359e-20 7.26888e-24 -1.96286e-20 0.00139607 0.997816 8.59955e-05 0.15268 2.85248 0.00139607 0.997816 0.763516 0.00106179 0.00188089 0.000859955 0.455463 0.00188089 0.442545 0.000130381 1.02 0.888391 0.534481 0.287038 1.71853e-07 3.0764e-09 2376.46 3122.71 -0.056509 0.482182 0.277371 0.253731 -0.593277 -0.169552 0.493031 -0.266512 -0.226528 2.317 1 0 296.866 0 2.18703 2.315 0.000299482 0.858224 0.685328 0.332184 0.42645 2.18722 136.602 83.8355 18.716 60.8253 0.00402881 0 -40 10
1.416 4.09848e-08 2.53945e-06 0.134353 0.134353 0.0120311 1.86294e-05 0.0011543 0.167942 0.000658588 0.168596 0.921733 101.63 0.23856 0.810368 4.36998 0.0614398 0.0412262 0.958774 0.0196092 0.00445716 0.0188702 0.004265 0.0053908 0.00612978 0.215632 0.245191 58.028 -87.8979 126.224 15.9477 145.029 0.00014155 0.267251 192.782 0.310336 0.0673428 0.00409746 0.000562153 0.00138436 0.986969 0.991722 -2.98506e-06 -85.6602 0.0930558 31176.6 306.356 0.983504 0.319146 0.734292 0.734288 9.99958 2.98479e-06 1.1939e-05 0.13283 0.983232 0.931653 -0.0132921 4.92054e-06 0.509924 -1.96372e-20 7.26941e-24 -1.96299e-20 0.00139607 0.997816 8.59956e-05 0.15268 2.85248 0.00139607 0.997816 0.763598 0.0010618 0.00188089 0.000859956 0.455463 0.00188089 0.442551 0.000130383 1.02 0.888392 0.534481 0.287039 1.71854e-07 3.07643e-09 2376.44 3122.75 -0.0565132 0.482182 0.277371 0.253734 -0.593277 -0.169552 0.493017 -0.26651 -0.226517 2.318 1 0 296.863 0 2.18717 2.316 0.000299481 0.858246 0.685373 0.332126 0.426474 2.18736 136.609 83.835 18.7159 60.8251 0.00402883 0 -40 10
1.417 4.10136e-08 2.53945e-06 0.134397 0.134396 0.0120311 1.86426e-05 0.0011543 0.167996 0.000658589 0.16865 0.921817 101.63 0.23855 0.810493 4.37045 0.0614499 0.0412307 0.958769 0.0196087 0.00445753 0.0188698 0.00426532 0.00539126 0.00613025 0.21565 0.24521 58.0281 -87.8979 126.224 15.9476 145.029 0.000141552 0.267251 192.782 0.310336 0.0673427 0.00409746 0.000562153 0.00138436 0.986969 0.991722 -2.98508e-06 -85.6602 0.0930559 31176.6 306.367 0.983504 0.319146 0.734302 0.734297 9.99958 2.98479e-06 1.19391e-05 0.132833 0.983233 0.931652 -0.0132921 4.92057e-06 0.50994 -1.96385e-20 7.26995e-24 -1.96312e-20 0.00139607 0.997816 8.59957e-05 0.15268 2.85248 0.00139607 0.997816 0.76368 0.00106182 0.00188089 0.000859957 0.455463 0.00188089 0.442557 0.000130386 1.02 0.888393 0.534481 0.287041 1.71854e-07 3.07645e-09 2376.42 3122.79 -0.0565174 0.482182 0.27737 0.253736 -0.593276 -0.169552 0.493004 -0.266508 -0.226505 2.319 1 0 296.859 0 2.18731 2.317 0.00029948 0.858268 0.685417 0.332069 0.426497 2.1875 136.617 83.8345 18.7159 60.8249 0.00402885 0 -40 10
1.418 4.10425e-08 2.53945e-06 0.13444 0.134439 0.012031 1.86557e-05 0.0011543 0.16805 0.00065859 0.168704 0.921901 101.629 0.23854 0.810619 4.37092 0.06146 0.0412351 0.958765 0.0196083 0.00445791 0.0188693 0.00426564 0.00539172 0.00613072 0.215669 0.245229 58.0281 -87.8979 126.224 15.9476 145.029 0.000141554 0.267251 192.782 0.310336 0.0673426 0.00409747 0.000562154 0.00138437 0.986969 0.991722 -2.98509e-06 -85.6602 0.093056 31176.6 306.377 0.983504 0.319146 0.734311 0.734307 9.99958 2.9848e-06 1.19391e-05 0.132837 0.983234 0.931651 -0.0132921 4.9206e-06 0.509956 -1.96398e-20 7.27048e-24 -1.96326e-20 0.00139607 0.997816 8.59958e-05 0.15268 2.85248 0.00139607 0.997816 0.763762 0.00106184 0.00188089 0.000859958 0.455463 0.00188089 0.442563 0.000130389 1.02 0.888394 0.53448 0.287042 1.71854e-07 3.07647e-09 2376.41 3122.83 -0.0565216 0.482182 0.27737 0.253739 -0.593276 -0.169552 0.49299 -0.266506 -0.226494 2.32 1 0 296.855 0 2.18745 2.318 0.00029948 0.85829 0.685462 0.332011 0.42652 2.18764 136.624 83.8341 18.7159 60.8247 0.00402887 0 -40 10
1.419 4.10714e-08 2.53945e-06 0.134483 0.134482 0.012031 1.86688e-05 0.0011543 0.168104 0.000658591 0.168758 0.921985 101.629 0.23853 0.810745 4.37139 0.0614701 0.0412396 0.95876 0.0196078 0.00445828 0.0188688 0.00426596 0.00539218 0.00613119 0.215687 0.245247 58.0282 -87.8979 126.224 15.9476 145.029 0.000141556 0.267251 192.782 0.310335 0.0673426 0.00409747 0.000562155 0.00138437 0.986969 0.991722 -2.98511e-06 -85.6602 0.0930561 31176.5 306.387 0.983504 0.319146 0.73432 0.734316 9.99958 2.9848e-06 1.19391e-05 0.132841 0.983235 0.931651 -0.0132921 4.92063e-06 0.509972 -1.96411e-20 7.27101e-24 -1.96339e-20 0.00139607 0.997816 8.59958e-05 0.15268 2.85248 0.00139607 0.997816 0.763844 0.00106185 0.00188089 0.000859958 0.455462 0.00188089 0.44257 0.000130391 1.02 0.888395 0.53448 0.287044 1.71855e-07 3.0765e-09 2376.39 3122.87 -0.0565258 0.482182 0.27737 0.253741 -0.593275 -0.169552 0.492977 -0.266503 -0.226483 2.321 1 0 296.851 0 2.1876 2.319 0.000299479 0.858312 0.685506 0.331954 0.426543 2.18778 136.632 83.8336 18.7159 60.8244 0.00402889 0 -40 10
1.42 4.11003e-08 2.53945e-06 0.134527 0.134526 0.012031 1.86819e-05 0.0011543 0.168158 0.000658592 0.168812 0.922069 101.628 0.23852 0.81087 4.37186 0.0614802 0.041244 0.958756 0.0196074 0.00445866 0.0188683 0.00426628 0.00539264 0.00613166 0.215706 0.245266 58.0282 -87.8979 126.224 15.9475 145.029 0.000141558 0.267251 192.782 0.310335 0.0673425 0.00409747 0.000562155 0.00138437 0.986969 0.991722 -2.98512e-06 -85.6602 0.0930562 31176.5 306.397 0.983504 0.319146 0.73433 0.734325 9.99958 2.98481e-06 1.19391e-05 0.132845 0.983236 0.93165 -0.0132921 4.92066e-06 0.509988 -1.96425e-20 7.27154e-24 -1.96352e-20 0.00139607 0.997816 8.59959e-05 0.152681 2.85248 0.00139607 0.997816 0.763926 0.00106187 0.00188089 0.000859959 0.455462 0.00188089 0.442576 0.000130394 1.02 0.888397 0.53448 0.287045 1.71855e-07 3.07652e-09 2376.37 3122.91 -0.05653 0.482182 0.277369 0.253744 -0.593275 -0.169552 0.492963 -0.266501 -0.226471 2.322 1 0 296.848 0 2.18774 2.32 0.000299478 0.858335 0.68555 0.331896 0.426566 2.18793 136.639 83.8332 18.7158 60.8242 0.00402891 0 -40 10
1.421 4.11292e-08 2.53946e-06 0.13457 0.134569 0.012031 1.86951e-05 0.0011543 0.168212 0.000658592 0.168866 0.922153 101.628 0.23851 0.810996 4.37234 0.0614903 0.0412485 0.958752 0.0196069 0.00445903 0.0188679 0.0042666 0.0053931 0.00613213 0.215724 0.245285 58.0283 -87.8979 126.224 15.9475 145.029 0.000141559 0.267252 192.782 0.310334 0.0673425 0.00409748 0.000562156 0.00138437 0.986969 0.991722 -2.98514e-06 -85.6602 0.0930563 31176.5 306.407 0.983504 0.319146 0.734339 0.734335 9.99958 2.98481e-06 1.19391e-05 0.132849 0.983236 0.931649 -0.0132921 4.92069e-06 0.510004 -1.96438e-20 7.27207e-24 -1.96365e-20 0.00139608 0.997816 8.5996e-05 0.152681 2.85248 0.00139608 0.997816 0.764008 0.00106189 0.0018809 0.00085996 0.455462 0.00188089 0.442582 0.000130397 1.02 0.888398 0.534479 0.287047 1.71855e-07 3.07654e-09 2376.36 3122.95 -0.0565342 0.482183 0.277369 0.253746 -0.593274 -0.169552 0.492949 -0.266499 -0.22646 2.323 1 0 296.844 0 2.18788 2.321 0.000299477 0.858357 0.685595 0.331839 0.42659 2.18807 136.647 83.8327 18.7158 60.824 0.00402892 0 -40 10
1.422 4.1158e-08 2.53946e-06 0.134613 0.134612 0.012031 1.87082e-05 0.0011543 0.168266 0.000658593 0.16892 0.922237 101.627 0.2385 0.811122 4.37281 0.0615004 0.0412529 0.958747 0.0196064 0.00445941 0.0188674 0.00426692 0.00539357 0.0061326 0.215743 0.245304 58.0284 -87.8979 126.223 15.9475 145.029 0.000141561 0.267252 192.781 0.310334 0.0673424 0.00409748 0.000562157 0.00138438 0.986969 0.991722 -2.98515e-06 -85.6601 0.0930564 31176.5 306.417 0.983504 0.319146 0.734349 0.734344 9.99958 2.98482e-06 1.19392e-05 0.132853 0.983237 0.931649 -0.0132921 4.92072e-06 0.51002 -1.96451e-20 7.27261e-24 -1.96378e-20 0.00139608 0.997816 8.59961e-05 0.152681 2.85248 0.00139608 0.997816 0.76409 0.00106191 0.0018809 0.000859961 0.455462 0.0018809 0.442588 0.000130399 1.02 0.888399 0.534479 0.287048 1.71855e-07 3.07656e-09 2376.34 3122.99 -0.0565385 0.482183 0.277369 0.253749 -0.593274 -0.169552 0.492936 -0.266497 -0.226448 2.324 1 0 296.84 0 2.18802 2.322 0.000299476 0.858379 0.685639 0.331781 0.426613 2.18821 136.655 83.8322 18.7158 60.8238 0.00402894 0 -40 10
1.423 4.11869e-08 2.53946e-06 0.134656 0.134655 0.012031 1.87213e-05 0.0011543 0.16832 0.000658594 0.168974 0.922321 101.627 0.238489 0.811247 4.37328 0.0615105 0.0412574 0.958743 0.019606 0.00445979 0.0188669 0.00426724 0.00539403 0.00613307 0.215761 0.245323 58.0284 -87.8979 126.223 15.9474 145.029 0.000141563 0.267252 192.781 0.310333 0.0673424 0.00409748 0.000562158 0.00138438 0.986969 0.991722 -2.98517e-06 -85.6601 0.0930565 31176.4 306.428 0.983504 0.319146 0.734358 0.734354 9.99958 2.98482e-06 1.19392e-05 0.132856 0.983238 0.931648 -0.0132921 4.92075e-06 0.510037 -1.96464e-20 7.27314e-24 -1.96391e-20 0.00139608 0.997816 8.59962e-05 0.152681 2.85248 0.00139608 0.997816 0.764172 0.00106192 0.0018809 0.000859962 0.455461 0.0018809 0.442594 0.000130402 1.02 0.8884 0.534479 0.28705 1.71856e-07 3.07659e-09 2376.32 3123.02 -0.0565427 0.482183 0.277369 0.253751 -0.593273 -0.169553 0.492922 -0.266495 -0.226437 2.325 1 0 296.836 0 2.18816 2.323 0.000299475 0.858401 0.685683 0.331724 0.426636 2.18835 136.662 83.8318 18.7158 60.8235 0.00402896 0 -40 10
1.424 4.12158e-08 2.53946e-06 0.134699 0.134698 0.012031 1.87344e-05 0.0011543 0.168374 0.000658595 0.169028 0.922405 101.626 0.238479 0.811373 4.37376 0.0615207 0.0412618 0.958738 0.0196055 0.00446016 0.0188665 0.00426756 0.00539449 0.00613354 0.21578 0.245342 58.0285 -87.8979 126.223 15.9474 145.029 0.000141565 0.267252 192.781 0.310333 0.0673423 0.00409748 0.000562158 0.00138438 0.986969 0.991722 -2.98518e-06 -85.6601 0.0930565 31176.4 306.438 0.983504 0.319146 0.734367 0.734363 9.99958 2.98483e-06 1.19392e-05 0.13286 0.983239 0.931647 -0.0132921 4.92078e-06 0.510053 -1.96477e-20 7.27368e-24 -1.96405e-20 0.00139608 0.997816 8.59962e-05 0.152681 2.85248 0.00139608 0.997816 0.764254 0.00106194 0.0018809 0.000859962 0.455461 0.0018809 0.4426 0.000130405 1.02 0.888401 0.534479 0.287051 1.71856e-07 3.07661e-09 2376.31 3123.06 -0.0565469 0.482183 0.277368 0.253754 -0.593273 -0.169553 0.492909 -0.266493 -0.226425 2.326 1 0 296.833 0 2.1883 2.324 0.000299474 0.858424 0.685728 0.331667 0.426659 2.18849 136.67 83.8313 18.7157 60.8233 0.00402898 0 -40 10
1.425 4.12447e-08 2.53946e-06 0.134742 0.134741 0.012031 1.87476e-05 0.0011543 0.168428 0.000658596 0.169082 0.922489 101.626 0.238469 0.811499 4.37423 0.0615308 0.0412663 0.958734 0.019605 0.00446054 0.018866 0.00426789 0.00539495 0.00613401 0.215798 0.245361 58.0286 -87.8979 126.223 15.9473 145.029 0.000141567 0.267252 192.781 0.310333 0.0673423 0.00409749 0.000562159 0.00138438 0.986969 0.991722 -2.9852e-06 -85.6601 0.0930566 31176.4 306.448 0.983504 0.319146 0.734377 0.734372 9.99958 2.98483e-06 1.19392e-05 0.132864 0.98324 0.931647 -0.0132921 4.92081e-06 0.510069 -1.96491e-20 7.27421e-24 -1.96418e-20 0.00139608 0.997816 8.59963e-05 0.152681 2.85249 0.00139608 0.997816 0.764335 0.00106196 0.0018809 0.000859963 0.455461 0.0018809 0.442606 0.000130407 1.02 0.888402 0.534478 0.287053 1.71856e-07 3.07663e-09 2376.29 3123.1 -0.0565512 0.482183 0.277368 0.253756 -0.593272 -0.169553 0.492895 -0.266491 -0.226414 2.327 1 0 296.829 0 2.18845 2.325 0.000299473 0.858446 0.685772 0.33161 0.426682 2.18863 136.677 83.8308 18.7157 60.8231 0.004029 0 -40 10
1.426 4.12735e-08 2.53946e-06 0.134785 0.134784 0.0120309 1.87607e-05 0.0011543 0.168482 0.000658597 0.169136 0.922573 101.625 0.238459 0.811625 4.3747 0.0615409 0.0412708 0.958729 0.0196046 0.00446092 0.0188655 0.00426821 0.00539542 0.00613449 0.215817 0.245379 58.0286 -87.8979 126.223 15.9473 145.029 0.000141568 0.267253 192.781 0.310332 0.0673422 0.00409749 0.00056216 0.00138438 0.986969 0.991722 -2.98521e-06 -85.6601 0.0930567 31176.4 306.458 0.983504 0.319146 0.734386 0.734382 9.99958 2.98484e-06 1.19392e-05 0.132868 0.983241 0.931646 -0.0132921 4.92084e-06 0.510085 -1.96504e-20 7.27474e-24 -1.96431e-20 0.00139608 0.997816 8.59964e-05 0.152682 2.85249 0.00139608 0.997816 0.764417 0.00106198 0.0018809 0.000859964 0.455461 0.0018809 0.442612 0.00013041 1.02 0.888403 0.534478 0.287054 1.71856e-07 3.07666e-09 2376.27 3123.14 -0.0565554 0.482183 0.277368 0.253759 -0.593272 -0.169553 0.492881 -0.266489 -0.226402 2.328 1 0 296.825 0 2.18859 2.326 0.000299472 0.858468 0.685816 0.331553 0.426705 2.18878 136.685 83.8304 18.7157 60.8229 0.00402902 0 -40 10
1.427 4.13024e-08 2.53946e-06 0.134828 0.134827 0.0120309 1.87738e-05 0.0011543 0.168535 0.000658597 0.169189 0.922658 101.625 0.238449 0.81175 4.37518 0.061551 0.0412753 0.958725 0.0196041 0.00446129 0.018865 0.00426853 0.00539588 0.00613496 0.215835 0.245398 58.0287 -87.8979 126.222 15.9473 145.029 0.00014157 0.267253 192.781 0.310332 0.0673422 0.00409749 0.00056216 0.00138439 0.986969 0.991722 -2.98523e-06 -85.6601 0.0930568 31176.3 306.469 0.983504 0.319146 0.734396 0.734391 9.99958 2.98484e-06 1.19393e-05 0.132872 0.983241 0.931645 -0.0132921 4.92087e-06 0.510101 -1.96517e-20 7.27528e-24 -1.96444e-20 0.00139608 0.997816 8.59965e-05 0.152682 2.85249 0.00139608 0.997816 0.764499 0.00106199 0.0018809 0.000859965 0.455461 0.0018809 0.442619 0.000130413 1.02 0.888404 0.534478 0.287056 1.71857e-07 3.07668e-09 2376.26 3123.18 -0.0565597 0.482183 0.277367 0.253761 -0.593271 -0.169553 0.492868 -0.266487 -0.22639 2.329 1 0 296.821 0 2.18873 2.327 0.000299471 0.858491 0.685861 0.331496 0.426729 2.18892 136.693 83.8299 18.7156 60.8226 0.00402904 0 -40 10
1.428 4.13313e-08 2.53946e-06 0.134871 0.13487 0.0120309 1.87869e-05 0.0011543 0.168589 0.000658598 0.169243 0.922742 101.624 0.238439 0.811876 4.37565 0.0615612 0.0412798 0.95872 0.0196037 0.00446167 0.0188646 0.00426885 0.00539635 0.00613543 0.215854 0.245417 58.0287 -87.8979 126.222 15.9472 145.029 0.000141572 0.267253 192.78 0.310331 0.0673421 0.0040975 0.000562161 0.00138439 0.986969 0.991722 -2.98524e-06 -85.6601 0.0930569 31176.3 306.479 0.983504 0.319146 0.734405 0.734401 9.99958 2.98485e-06 1.19393e-05 0.132876 0.983242 0.931645 -0.0132921 4.9209e-06 0.510118 -1.9653e-20 7.27581e-24 -1.96458e-20 0.00139608 0.997816 8.59966e-05 0.152682 2.85249 0.00139608 0.997816 0.764581 0.00106201 0.00188091 0.000859966 0.45546 0.0018809 0.442625 0.000130415 1.02 0.888405 0.534477 0.287057 1.71857e-07 3.0767e-09 2376.24 3123.22 -0.0565639 0.482183 0.277367 0.253764 -0.593271 -0.169553 0.492854 -0.266484 -0.226379 2.33 1 0 296.817 0 2.18887 2.328 0.00029947 0.858513 0.685905 0.331439 0.426752 2.18906 136.7 83.8294 18.7156 60.8224 0.00402906 0 -40 10
1.429 4.13602e-08 2.53947e-06 0.134914 0.134913 0.0120309 1.88001e-05 0.0011543 0.168643 0.000658599 0.169297 0.922826 101.624 0.238429 0.812002 4.37613 0.0615713 0.0412843 0.958716 0.0196032 0.00446205 0.0188641 0.00426918 0.00539681 0.00613591 0.215872 0.245436 58.0288 -87.8979 126.222 15.9472 145.029 0.000141574 0.267253 192.78 0.310331 0.0673421 0.0040975 0.000562162 0.00138439 0.986969 0.991721 -2.98526e-06 -85.6601 0.093057 31176.3 306.489 0.983504 0.319146 0.734415 0.73441 9.99958 2.98485e-06 1.19393e-05 0.13288 0.983243 0.931644 -0.0132921 4.92093e-06 0.510134 -1.96544e-20 7.27635e-24 -1.96471e-20 0.00139609 0.997816 8.59967e-05 0.152682 2.85249 0.00139608 0.997816 0.764663 0.00106203 0.00188091 0.000859967 0.45546 0.00188091 0.442631 0.000130418 1.02 0.888406 0.534477 0.287059 1.71857e-07 3.07672e-09 2376.23 3123.26 -0.0565682 0.482183 0.277367 0.253767 -0.59327 -0.169553 0.49284 -0.266482 -0.226367 2.331 1 0 296.814 0 2.18901 2.329 0.000299469 0.858535 0.685949 0.331382 0.426775 2.1892 136.708 83.829 18.7156 60.8222 0.00402908 0 -40 10
1.43 4.1389e-08 2.53947e-06 0.134957 0.134956 0.0120309 1.88132e-05 0.0011543 0.168696 0.0006586 0.16935 0.92291 101.623 0.238419 0.812128 4.37661 0.0615814 0.0412887 0.958711 0.0196027 0.00446243 0.0188636 0.0042695 0.00539728 0.00613638 0.215891 0.245455 58.0289 -87.8979 126.222 15.9472 145.029 0.000141576 0.267253 192.78 0.31033 0.067342 0.0040975 0.000562162 0.00138439 0.986968 0.991721 -2.98527e-06 -85.6601 0.0930571 31176.3 306.499 0.983504 0.319146 0.734424 0.73442 9.99958 2.98486e-06 1.19393e-05 0.132883 0.983244 0.931643 -0.0132921 4.92096e-06 0.51015 -1.96557e-20 7.27688e-24 -1.96484e-20 0.00139609 0.997816 8.59967e-05 0.152682 2.85249 0.00139609 0.997816 0.764744 0.00106205 0.00188091 0.000859967 0.45546 0.00188091 0.442637 0.000130421 1.02 0.888408 0.534477 0.287061 1.71857e-07 3.07675e-09 2376.21 3123.3 -0.0565724 0.482183 0.277367 0.253769 -0.59327 -0.169553 0.492827 -0.26648 -0.226356 2.332 1 0 296.81 0 2.18915 2.33 0.000299469 0.858558 0.685994 0.331325 0.426798 2.18934 136.715 83.8285 18.7156 60.822 0.0040291 0 -40 10
1.431 4.14179e-08 2.53947e-06 0.135 0.134999 0.0120309 1.88263e-05 0.0011543 0.16875 0.000658601 0.169404 0.922995 101.623 0.238408 0.812254 4.37708 0.0615916 0.0412932 0.958707 0.0196023 0.0044628 0.0188631 0.00426982 0.00539774 0.00613685 0.21591 0.245474 58.0289 -87.8979 126.222 15.9471 145.029 0.000141578 0.267254 192.78 0.31033 0.067342 0.00409751 0.000562163 0.00138439 0.986968 0.991721 -2.98529e-06 -85.6601 0.0930572 31176.3 306.51 0.983504 0.319146 0.734434 0.734429 9.99958 2.98486e-06 1.19393e-05 0.132887 0.983245 0.931643 -0.0132921 4.92099e-06 0.510166 -1.9657e-20 7.27742e-24 -1.96497e-20 0.00139609 0.997816 8.59968e-05 0.152682 2.85249 0.00139609 0.997816 0.764826 0.00106206 0.00188091 0.000859968 0.45546 0.00188091 0.442643 0.000130423 1.02 0.888409 0.534476 0.287062 1.71858e-07 3.07677e-09 2376.19 3123.34 -0.0565767 0.482183 0.277366 0.253772 -0.593269 -0.169553 0.492813 -0.266478 -0.226344 2.333 1 0 296.806 0 2.18929 2.331 0.000299468 0.85858 0.686038 0.331269 0.426821 2.18948 136.723 83.828 18.7155 60.8217 0.00402912 0 -40 10
1.432 4.14468e-08 2.53947e-06 0.135043 0.135042 0.0120309 1.88394e-05 0.0011543 0.168803 0.000658601 0.169457 0.923079 101.622 0.238398 0.81238 4.37756 0.0616017 0.0412977 0.958702 0.0196018 0.00446318 0.0188627 0.00427015 0.00539821 0.00613733 0.215928 0.245493 58.029 -87.8979 126.222 15.9471 145.029 0.000141579 0.267254 192.78 0.31033 0.0673419 0.00409751 0.000562164 0.0013844 0.986968 0.991721 -2.9853e-06 -85.66 0.0930572 31176.2 306.52 0.983504 0.319146 0.734443 0.734439 9.99958 2.98487e-06 1.19394e-05 0.132891 0.983245 0.931642 -0.0132921 4.92102e-06 0.510182 -1.96583e-20 7.27796e-24 -1.96511e-20 0.00139609 0.997816 8.59969e-05 0.152682 2.85249 0.00139609 0.997816 0.764908 0.00106208 0.00188091 0.000859969 0.455459 0.00188091 0.442649 0.000130426 1.02 0.88841 0.534476 0.287064 1.71858e-07 3.07679e-09 2376.18 3123.38 -0.056581 0.482183 0.277366 0.253774 -0.593269 -0.169553 0.492799 -0.266476 -0.226333 2.334 1 0 296.802 0 2.18944 2.332 0.000299467 0.858603 0.686082 0.331212 0.426844 2.18962 136.731 83.8276 18.7155 60.8215 0.00402914 0 -40 10
1.433 4.14757e-08 2.53947e-06 0.135085 0.135085 0.0120308 1.88526e-05 0.0011543 0.168857 0.000658602 0.169511 0.923163 101.622 0.238388 0.812506 4.37804 0.0616118 0.0413022 0.958698 0.0196013 0.00446356 0.0188622 0.00427047 0.00539867 0.0061378 0.215947 0.245512 58.0291 -87.8979 126.221 15.947 145.029 0.000141581 0.267254 192.78 0.310329 0.0673419 0.00409751 0.000562164 0.0013844 0.986968 0.991721 -2.98532e-06 -85.66 0.0930573 31176.2 306.53 0.983504 0.319146 0.734453 0.734448 9.99958 2.98487e-06 1.19394e-05 0.132895 0.983246 0.931641 -0.0132921 4.92105e-06 0.510199 -1.96597e-20 7.27849e-24 -1.96524e-20 0.00139609 0.997816 8.5997e-05 0.152683 2.85249 0.00139609 0.997816 0.764989 0.0010621 0.00188091 0.00085997 0.455459 0.00188091 0.442655 0.000130429 1.02 0.888411 0.534476 0.287065 1.71858e-07 3.07682e-09 2376.16 3123.42 -0.0565852 0.482183 0.277366 0.253777 -0.593268 -0.169553 0.492785 -0.266474 -0.226321 2.335 1 0 296.798 0 2.18958 2.333 0.000299466 0.858625 0.686126 0.331156 0.426868 2.18977 136.738 83.8271 18.7155 60.8213 0.00402916 0 -40 10
1.434 4.15045e-08 2.53947e-06 0.135128 0.135127 0.0120308 1.88657e-05 0.0011543 0.16891 0.000658603 0.169564 0.923248 101.621 0.238378 0.812632 4.37852 0.061622 0.0413068 0.958693 0.0196009 0.00446394 0.0188617 0.00427079 0.00539914 0.00613828 0.215966 0.245531 58.0291 -87.8979 126.221 15.947 145.029 0.000141583 0.267254 192.779 0.310329 0.0673418 0.00409751 0.000562165 0.0013844 0.986968 0.991721 -2.98533e-06 -85.66 0.0930574 31176.2 306.54 0.983504 0.319146 0.734462 0.734458 9.99958 2.98488e-06 1.19394e-05 0.132899 0.983247 0.931641 -0.0132921 4.92108e-06 0.510215 -1.9661e-20 7.27903e-24 -1.96537e-20 0.00139609 0.997816 8.59971e-05 0.152683 2.85249 0.00139609 0.997816 0.765071 0.00106211 0.00188091 0.000859971 0.455459 0.00188091 0.442661 0.000130431 1.02 0.888412 0.534475 0.287067 1.71859e-07 3.07684e-09 2376.14 3123.46 -0.0565895 0.482184 0.277365 0.253779 -0.593268 -0.169553 0.492772 -0.266472 -0.226309 2.336 1 0 296.795 0 2.18972 2.334 0.000299465 0.858648 0.686171 0.331099 0.426891 2.18991 136.746 83.8266 18.7155 60.8211 0.00402918 0 -40 10
1.435 4.15334e-08 2.53947e-06 0.135171 0.13517 0.0120308 1.88788e-05 0.00115431 0.168964 0.000658604 0.169618 0.923332 101.621 0.238368 0.812758 4.379 0.0616321 0.0413113 0.958689 0.0196004 0.00446432 0.0188612 0.00427112 0.00539961 0.00613875 0.215984 0.24555 58.0292 -87.8979 126.221 15.947 145.029 0.000141585 0.267254 192.779 0.310328 0.0673418 0.00409752 0.000562166 0.0013844 0.986968 0.991721 -2.98535e-06 -85.66 0.0930575 31176.2 306.551 0.983504 0.319146 0.734472 0.734467 9.99958 2.98488e-06 1.19394e-05 0.132903 0.983248 0.93164 -0.0132921 4.92111e-06 0.510231 -1.96623e-20 7.27957e-24 -1.9655e-20 0.00139609 0.997816 8.59971e-05 0.152683 2.85249 0.00139609 0.997816 0.765153 0.00106213 0.00188092 0.000859971 0.455459 0.00188092 0.442667 0.000130434 1.02 0.888413 0.534475 0.287068 1.71859e-07 3.07686e-09 2376.13 3123.5 -0.0565938 0.482184 0.277365 0.253782 -0.593267 -0.169553 0.492758 -0.26647 -0.226298 2.337 1 0 296.791 0 2.18986 2.335 0.000299464 0.85867 0.686215 0.331043 0.426914 2.19005 136.753 83.8261 18.7154 60.8208 0.00402919 0 -40 10
1.436 4.15623e-08 2.53947e-06 0.135214 0.135213 0.0120308 1.88919e-05 0.00115431 0.169017 0.000658605 0.169671 0.923417 101.621 0.238358 0.812884 4.37947 0.0616423 0.0413158 0.958684 0.0195999 0.0044647 0.0188608 0.00427144 0.00540007 0.00613923 0.216003 0.245569 58.0293 -87.898 126.221 15.9469 145.029 0.000141587 0.267255 192.779 0.310328 0.0673417 0.00409752 0.000562166 0.00138441 0.986968 0.991721 -2.98536e-06 -85.66 0.0930576 31176.1 306.561 0.983504 0.319146 0.734481 0.734477 9.99958 2.98489e-06 1.19394e-05 0.132907 0.983249 0.931639 -0.0132921 4.92114e-06 0.510248 -1.96637e-20 7.2801e-24 -1.96564e-20 0.00139609 0.997816 8.59972e-05 0.152683 2.8525 0.00139609 0.997816 0.765234 0.00106215 0.00188092 0.000859972 0.455458 0.00188092 0.442674 0.000130437 1.02 0.888414 0.534475 0.28707 1.71859e-07 3.07689e-09 2376.11 3123.54 -0.0565981 0.482184 0.277365 0.253784 -0.593267 -0.169553 0.492744 -0.266468 -0.226286 2.338 1 0 296.787 0 2.19 2.336 0.000299463 0.858693 0.686259 0.330986 0.426937 2.19019 136.761 83.8257 18.7154 60.8206 0.00402921 0 -40 10
1.437 4.15911e-08 2.53947e-06 0.135256 0.135255 0.0120308 1.89051e-05 0.00115431 0.16907 0.000658605 0.169724 0.923501 101.62 0.238348 0.81301 4.37995 0.0616524 0.0413203 0.95868 0.0195995 0.00446508 0.0188603 0.00427177 0.00540054 0.00613971 0.216022 0.245588 58.0293 -87.898 126.221 15.9469 145.029 0.000141589 0.267255 192.779 0.310327 0.0673416 0.00409752 0.000562167 0.00138441 0.986968 0.991721 -2.98538e-06 -85.66 0.0930577 31176.1 306.571 0.983504 0.319146 0.734491 0.734486 9.99958 2.98489e-06 1.19395e-05 0.13291 0.983249 0.931639 -0.0132921 4.92117e-06 0.510264 -1.9665e-20 7.28064e-24 -1.96577e-20 0.00139609 0.997816 8.59973e-05 0.152683 2.8525 0.00139609 0.997816 0.765316 0.00106217 0.00188092 0.000859973 0.455458 0.00188092 0.44268 0.000130439 1.02 0.888415 0.534475 0.287071 1.71859e-07 3.07691e-09 2376.09 3123.58 -0.0566024 0.482184 0.277365 0.253787 -0.593266 -0.169553 0.49273 -0.266465 -0.226274 2.339 1 0 296.783 0 2.19014 2.337 0.000299462 0.858716 0.686304 0.33093 0.42696 2.19033 136.768 83.8252 18.7154 60.8204 0.00402923 0 -40 10
1.438 4.162e-08 2.53948e-06 0.135299 0.135298 0.0120308 1.89182e-05 0.00115431 0.169124 0.000658606 0.169778 0.923585 101.62 0.238337 0.813136 4.38043 0.0616626 0.0413248 0.958675 0.019599 0.00446546 0.0188598 0.00427209 0.00540101 0.00614018 0.21604 0.245607 58.0294 -87.898 126.221 15.9469 145.029 0.00014159 0.267255 192.779 0.310327 0.0673416 0.00409753 0.000562168 0.00138441 0.986968 0.991721 -2.98539e-06 -85.66 0.0930578 31176.1 306.582 0.983504 0.319146 0.7345 0.734496 9.99958 2.9849e-06 1.19395e-05 0.132914 0.98325 0.931638 -0.0132921 4.9212e-06 0.51028 -1.96663e-20 7.28118e-24 -1.9659e-20 0.0013961 0.997816 8.59974e-05 0.152683 2.8525 0.0013961 0.997816 0.765397 0.00106218 0.00188092 0.000859974 0.455458 0.00188092 0.442686 0.000130442 1.02 0.888416 0.534474 0.287073 1.7186e-07 3.07693e-09 2376.08 3123.62 -0.0566067 0.482184 0.277364 0.25379 -0.593266 -0.169553 0.492717 -0.266463 -0.226263 2.34 1 0 296.779 0 2.19028 2.338 0.000299461 0.858738 0.686348 0.330874 0.426983 2.19047 136.776 83.8247 18.7153 60.8202 0.00402925 0 -40 10
1.439 4.16489e-08 2.53948e-06 0.135341 0.135341 0.0120308 1.89313e-05 0.00115431 0.169177 0.000658607 0.169831 0.92367 101.619 0.238327 0.813262 4.38091 0.0616727 0.0413294 0.958671 0.0195985 0.00446584 0.0188593 0.00427242 0.00540148 0.00614066 0.216059 0.245626 58.0294 -87.898 126.22 15.9468 145.029 0.000141592 0.267255 192.779 0.310327 0.0673415 0.00409753 0.000562168 0.00138441 0.986968 0.991721 -2.98541e-06 -85.66 0.0930579 31176.1 306.592 0.983504 0.319146 0.73451 0.734506 9.99958 2.9849e-06 1.19395e-05 0.132918 0.983251 0.931637 -0.0132921 4.92123e-06 0.510297 -1.96677e-20 7.28172e-24 -1.96604e-20 0.0013961 0.997816 8.59975e-05 0.152684 2.8525 0.0013961 0.997816 0.765479 0.0010622 0.00188092 0.000859975 0.455458 0.00188092 0.442692 0.000130445 1.02 0.888417 0.534474 0.287074 1.7186e-07 3.07695e-09 2376.06 3123.66 -0.0566109 0.482184 0.277364 0.253792 -0.593265 -0.169554 0.492703 -0.266461 -0.226251 2.341 1 0 296.775 0 2.19042 2.339 0.00029946 0.858761 0.686392 0.330818 0.427006 2.19061 136.784 83.8243 18.7153 60.8199 0.00402927 0 -40 10
1.44 4.16778e-08 2.53948e-06 0.135384 0.135383 0.0120307 1.89444e-05 0.00115431 0.16923 0.000658608 0.169884 0.923754 101.619 0.238317 0.813388 4.38139 0.0616829 0.0413339 0.958666 0.0195981 0.00446622 0.0188589 0.00427274 0.00540195 0.00614114 0.216078 0.245645 58.0295 -87.898 126.22 15.9468 145.029 0.000141594 0.267255 192.778 0.310326 0.0673415 0.00409753 0.000562169 0.00138441 0.986968 0.991721 -2.98542e-06 -85.66 0.0930579 31176.1 306.602 0.983504 0.319146 0.73452 0.734515 9.99958 2.98491e-06 1.19395e-05 0.132922 0.983252 0.931637 -0.0132921 4.92126e-06 0.510313 -1.9669e-20 7.28226e-24 -1.96617e-20 0.0013961 0.997816 8.59975e-05 0.152684 2.8525 0.0013961 0.997816 0.76556 0.00106222 0.00188092 0.000859975 0.455458 0.00188092 0.442698 0.000130447 1.02 0.888419 0.534474 0.287076 1.7186e-07 3.07698e-09 2376.04 3123.7 -0.0566152 0.482184 0.277364 0.253795 -0.593265 -0.169554 0.492689 -0.266459 -0.226239 2.342 1 0 296.772 0 2.19057 2.34 0.000299459 0.858784 0.686436 0.330762 0.427029 2.19075 136.791 83.8238 18.7153 60.8197 0.00402929 0 -40 10
1.441 4.17066e-08 2.53948e-06 0.135427 0.135426 0.0120307 1.89576e-05 0.00115431 0.169283 0.000658609 0.169937 0.923839 101.618 0.238307 0.813515 4.38188 0.0616931 0.0413385 0.958662 0.0195976 0.0044666 0.0188584 0.00427307 0.00540241 0.00614161 0.216097 0.245665 58.0296 -87.898 126.22 15.9467 145.03 0.000141596 0.267255 192.778 0.310326 0.0673414 0.00409754 0.00056217 0.00138442 0.986968 0.991721 -2.98544e-06 -85.66 0.093058 31176 306.613 0.983504 0.319146 0.734529 0.734525 9.99958 2.98491e-06 1.19395e-05 0.132926 0.983253 0.931636 -0.0132921 4.92129e-06 0.510329 -1.96703e-20 7.2828e-24 -1.9663e-20 0.0013961 0.997816 8.59976e-05 0.152684 2.8525 0.0013961 0.997816 0.765641 0.00106224 0.00188093 0.000859976 0.455457 0.00188092 0.442704 0.00013045 1.02 0.88842 0.534473 0.287077 1.7186e-07 3.077e-09 2376.03 3123.74 -0.0566195 0.482184 0.277363 0.253797 -0.593264 -0.169554 0.492675 -0.266457 -0.226228 2.343 1 0 296.768 0 2.19071 2.341 0.000299458 0.858807 0.686481 0.330706 0.427052 2.1909 136.799 83.8233 18.7153 60.8195 0.00402931 0 -40 10
1.442 4.17355e-08 2.53948e-06 0.135469 0.135468 0.0120307 1.89707e-05 0.00115431 0.169336 0.000658609 0.16999 0.923923 101.618 0.238297 0.813641 4.38236 0.0617032 0.041343 0.958657 0.0195971 0.00446698 0.0188579 0.00427339 0.00540288 0.00614209 0.216115 0.245684 58.0296 -87.898 126.22 15.9467 145.03 0.000141598 0.267256 192.778 0.310325 0.0673414 0.00409754 0.00056217 0.00138442 0.986968 0.991721 -2.98545e-06 -85.66 0.0930581 31176 306.623 0.983504 0.319146 0.734539 0.734535 9.99958 2.98492e-06 1.19396e-05 0.13293 0.983253 0.931635 -0.0132921 4.92132e-06 0.510346 -1.96717e-20 7.28334e-24 -1.96644e-20 0.0013961 0.997816 8.59977e-05 0.152684 2.8525 0.0013961 0.997816 0.765723 0.00106225 0.00188093 0.000859977 0.455457 0.00188093 0.44271 0.000130453 1.02 0.888421 0.534473 0.287079 1.71861e-07 3.07702e-09 2376.01 3123.78 -0.0566239 0.482184 0.277363 0.2538 -0.593264 -0.169554 0.492661 -0.266455 -0.226216 2.344 1 0 296.764 0 2.19085 2.342 0.000299457 0.858829 0.686525 0.33065 0.427076 2.19104 136.806 83.8228 18.7152 60.8192 0.00402933 0 -40 10
1.443 4.17644e-08 2.53948e-06 0.135511 0.135511 0.0120307 1.89838e-05 0.00115431 0.169389 0.00065861 0.170043 0.924008 101.617 0.238287 0.813767 4.38284 0.0617134 0.0413475 0.958652 0.0195966 0.00446736 0.0188574 0.00427372 0.00540335 0.00614257 0.216134 0.245703 58.0297 -87.898 126.22 15.9467 145.03 0.0001416 0.267256 192.778 0.310325 0.0673413 0.00409754 0.000562171 0.00138442 0.986968 0.991721 -2.98547e-06 -85.6599 0.0930582 31176 306.633 0.983504 0.319146 0.734549 0.734544 9.99958 2.98492e-06 1.19396e-05 0.132934 0.983254 0.931634 -0.013292 4.92135e-06 0.510362 -1.9673e-20 7.28387e-24 -1.96657e-20 0.0013961 0.997816 8.59978e-05 0.152684 2.8525 0.0013961 0.997816 0.765804 0.00106227 0.00188093 0.000859978 0.455457 0.00188093 0.442716 0.000130455 1.02 0.888422 0.534473 0.28708 1.71861e-07 3.07705e-09 2375.99 3123.82 -0.0566282 0.482184 0.277363 0.253803 -0.593263 -0.169554 0.492648 -0.266453 -0.226204 2.345 1 0 296.76 0 2.19099 2.343 0.000299456 0.858852 0.686569 0.330594 0.427099 2.19118 136.814 83.8224 18.7152 60.819 0.00402935 0 -40 10
1.444 4.17933e-08 2.53948e-06 0.135554 0.135553 0.0120307 1.89969e-05 0.00115431 0.169442 0.000658611 0.170096 0.924093 101.617 0.238276 0.813893 4.38332 0.0617236 0.0413521 0.958648 0.0195962 0.00446774 0.018857 0.00427405 0.00540382 0.00614305 0.216153 0.245722 58.0298 -87.898 126.22 15.9466 145.03 0.000141602 0.267256 192.778 0.310324 0.0673413 0.00409755 0.000562172 0.00138442 0.986968 0.991721 -2.98548e-06 -85.6599 0.0930583 31176 306.644 0.983504 0.319146 0.734558 0.734554 9.99958 2.98493e-06 1.19396e-05 0.132938 0.983255 0.931634 -0.013292 4.92138e-06 0.510378 -1.96743e-20 7.28441e-24 -1.96671e-20 0.0013961 0.997816 8.59979e-05 0.152684 2.8525 0.0013961 0.997816 0.765886 0.00106229 0.00188093 0.000859979 0.455457 0.00188093 0.442722 0.000130458 1.02 0.888423 0.534472 0.287082 1.71861e-07 3.07707e-09 2375.98 3123.86 -0.0566325 0.482184 0.277363 0.253805 -0.593263 -0.169554 0.492634 -0.266451 -0.226192 2.346 1 0 296.756 0 2.19113 2.344 0.000299456 0.858875 0.686613 0.330538 0.427122 2.19132 136.821 83.8219 18.7152 60.8188 0.00402937 0 -40 10
1.445 4.18221e-08 2.53948e-06 0.135596 0.135595 0.0120307 1.90101e-05 0.00115431 0.169495 0.000658612 0.170149 0.924177 101.616 0.238266 0.81402 4.38381 0.0617337 0.0413567 0.958643 0.0195957 0.00446812 0.0188565 0.00427437 0.00540429 0.00614353 0.216172 0.245741 58.0298 -87.898 126.219 15.9466 145.03 0.000141603 0.267256 192.778 0.310324 0.0673412 0.00409755 0.000562172 0.00138443 0.986968 0.991721 -2.9855e-06 -85.6599 0.0930584 31175.9 306.654 0.983504 0.319146 0.734568 0.734563 9.99958 2.98493e-06 1.19396e-05 0.132941 0.983256 0.931633 -0.013292 4.9214e-06 0.510395 -1.96757e-20 7.28495e-24 -1.96684e-20 0.0013961 0.997816 8.59979e-05 0.152684 2.8525 0.0013961 0.997816 0.765967 0.0010623 0.00188093 0.000859979 0.455456 0.00188093 0.442728 0.000130461 1.02 0.888424 0.534472 0.287083 1.71862e-07 3.07709e-09 2375.96 3123.9 -0.0566368 0.482184 0.277362 0.253808 -0.593262 -0.169554 0.49262 -0.266449 -0.226181 2.347 1 0 296.752 0 2.19127 2.345 0.000299455 0.858898 0.686657 0.330483 0.427145 2.19146 136.829 83.8214 18.7152 60.8185 0.00402939 0 -40 10
1.446 4.1851e-08 2.53949e-06 0.135639 0.135638 0.0120307 1.90232e-05 0.00115431 0.169548 0.000658613 0.170202 0.924262 101.616 0.238256 0.814146 4.38429 0.0617439 0.0413612 0.958639 0.0195952 0.0044685 0.018856 0.0042747 0.00540476 0.00614401 0.216191 0.24576 58.0299 -87.898 126.219 15.9466 145.03 0.000141605 0.267256 192.777 0.310324 0.0673412 0.00409755 0.000562173 0.00138443 0.986968 0.991721 -2.98551e-06 -85.6599 0.0930585 31175.9 306.664 0.983504 0.319146 0.734578 0.734573 9.99958 2.98494e-06 1.19396e-05 0.132945 0.983257 0.931632 -0.013292 4.92143e-06 0.510411 -1.9677e-20 7.2855e-24 -1.96697e-20 0.0013961 0.997816 8.5998e-05 0.152685 2.8525 0.0013961 0.997816 0.766048 0.00106232 0.00188093 0.00085998 0.455456 0.00188093 0.442734 0.000130463 1.02 0.888425 0.534472 0.287085 1.71862e-07 3.07711e-09 2375.94 3123.94 -0.0566411 0.482184 0.277362 0.25381 -0.593261 -0.169554 0.492606 -0.266447 -0.226169 2.348 1 0 296.748 0 2.19141 2.346 0.000299454 0.858921 0.686702 0.330427 0.427168 2.1916 136.837 83.8209 18.7151 60.8183 0.00402941 0 -40 10
1.447 4.18799e-08 2.53949e-06 0.135681 0.13568 0.0120307 1.90363e-05 0.00115431 0.169601 0.000658613 0.170255 0.924346 101.615 0.238246 0.814272 4.38477 0.0617541 0.0413658 0.958634 0.0195948 0.00446889 0.0188555 0.00427503 0.00540523 0.00614449 0.216209 0.24578 58.0299 -87.898 126.219 15.9465 145.03 0.000141607 0.267257 192.777 0.310323 0.0673411 0.00409755 0.000562174 0.00138443 0.986968 0.991721 -2.98553e-06 -85.6599 0.0930586 31175.9 306.675 0.983504 0.319146 0.734587 0.734583 9.99958 2.98494e-06 1.19397e-05 0.132949 0.983257 0.931632 -0.013292 4.92146e-06 0.510428 -1.96784e-20 7.28604e-24 -1.96711e-20 0.00139611 0.997816 8.59981e-05 0.152685 2.85251 0.00139611 0.997816 0.766129 0.00106234 0.00188093 0.000859981 0.455456 0.00188093 0.44274 0.000130466 1.02 0.888426 0.534471 0.287086 1.71862e-07 3.07714e-09 2375.93 3123.98 -0.0566454 0.482185 0.277362 0.253813 -0.593261 -0.169554 0.492592 -0.266444 -0.226157 2.349 1 0 296.745 0 2.19155 2.347 0.000299453 0.858944 0.686746 0.330371 0.427191 2.19174 136.844 83.8204 18.7151 60.8181 0.00402943 0 -40 10
1.448 4.19088e-08 2.53949e-06 0.135723 0.135722 0.0120306 1.90494e-05 0.00115431 0.169654 0.000658614 0.170308 0.924431 101.615 0.238236 0.814399 4.38526 0.0617643 0.0413704 0.95863 0.0195943 0.00446927 0.018855 0.00427535 0.0054057 0.00614497 0.216228 0.245799 58.03 -87.898 126.219 15.9465 145.03 0.000141609 0.267257 192.777 0.310323 0.0673411 0.00409756 0.000562174 0.00138443 0.986968 0.991721 -2.98554e-06 -85.6599 0.0930586 31175.9 306.685 0.983504 0.319146 0.734597 0.734593 9.99958 2.98495e-06 1.19397e-05 0.132953 0.983258 0.931631 -0.013292 4.92149e-06 0.510444 -1.96797e-20 7.28658e-24 -1.96724e-20 0.00139611 0.997816 8.59982e-05 0.152685 2.85251 0.00139611 0.997816 0.766211 0.00106236 0.00188094 0.000859982 0.455456 0.00188093 0.442746 0.000130469 1.02 0.888427 0.534471 0.287088 1.71862e-07 3.07716e-09 2375.91 3124.02 -0.0566498 0.482185 0.277362 0.253816 -0.59326 -0.169554 0.492578 -0.266442 -0.226145 2.35 1 0 296.741 0 2.19169 2.348 0.000299452 0.858967 0.68679 0.330316 0.427214 2.19188 136.852 83.82 18.7151 60.8179 0.00402945 0 -40 10
1.449 4.19376e-08 2.53949e-06 0.135765 0.135765 0.0120306 1.90626e-05 0.00115431 0.169707 0.000658615 0.170361 0.924516 101.614 0.238226 0.814525 4.38574 0.0617744 0.0413749 0.958625 0.0195938 0.00446965 0.0188546 0.00427568 0.00540618 0.00614545 0.216247 0.245818 58.0301 -87.898 126.219 15.9464 145.03 0.000141611 0.267257 192.777 0.310322 0.067341 0.00409756 0.000562175 0.00138443 0.986968 0.991721 -2.98556e-06 -85.6599 0.0930587 31175.9 306.695 0.983504 0.319146 0.734607 0.734602 9.99958 2.98495e-06 1.19397e-05 0.132957 0.983259 0.93163 -0.013292 4.92152e-06 0.510461 -1.9681e-20 7.28712e-24 -1.96737e-20 0.00139611 0.997816 8.59983e-05 0.152685 2.85251 0.00139611 0.997816 0.766292 0.00106237 0.00188094 0.000859983 0.455456 0.00188094 0.442752 0.000130471 1.02 0.888428 0.534471 0.287089 1.71863e-07 3.07718e-09 2375.89 3124.06 -0.0566541 0.482185 0.277361 0.253818 -0.59326 -0.169554 0.492564 -0.26644 -0.226133 2.351 1 0 296.737 0 2.19184 2.349 0.000299451 0.85899 0.686834 0.330261 0.427237 2.19202 136.859 83.8195 18.715 60.8176 0.00402947 0 -40 10
1.45 4.19665e-08 2.53949e-06 0.135808 0.135807 0.0120306 1.90757e-05 0.00115431 0.16976 0.000658616 0.170414 0.9246 101.614 0.238215 0.814652 4.38623 0.0617846 0.0413795 0.95862 0.0195934 0.00447003 0.0188541 0.00427601 0.00540665 0.00614593 0.216266 0.245837 58.0301 -87.898 126.218 15.9464 145.03 0.000141613 0.267257 192.777 0.310322 0.067341 0.00409756 0.000562176 0.00138444 0.986968 0.991721 -2.98557e-06 -85.6599 0.0930588 31175.8 306.706 0.983504 0.319146 0.734616 0.734612 9.99958 2.98496e-06 1.19397e-05 0.132961 0.98326 0.931629 -0.013292 4.92155e-06 0.510477 -1.96824e-20 7.28766e-24 -1.96751e-20 0.00139611 0.997816 8.59983e-05 0.152685 2.85251 0.00139611 0.997816 0.766373 0.00106239 0.00188094 0.000859983 0.455455 0.00188094 0.442758 0.000130474 1.02 0.88843 0.534471 0.287091 1.71863e-07 3.07721e-09 2375.88 3124.1 -0.0566584 0.482185 0.277361 0.253821 -0.593259 -0.169554 0.49255 -0.266438 -0.226122 2.352 1 0 296.733 0 2.19198 2.35 0.00029945 0.859013 0.686878 0.330205 0.42726 2.19217 136.867 83.819 18.715 60.8174 0.00402949 0 -40 10
1.451 4.19954e-08 2.53949e-06 0.13585 0.135849 0.0120306 1.90888e-05 0.00115431 0.169812 0.000658617 0.170466 0.924685 101.613 0.238205 0.814778 4.38671 0.0617948 0.0413841 0.958616 0.0195929 0.00447042 0.0188536 0.00427634 0.00540712 0.00614641 0.216285 0.245856 58.0302 -87.898 126.218 15.9464 145.03 0.000141615 0.267257 192.777 0.310321 0.0673409 0.00409757 0.000562176 0.00138444 0.986968 0.991721 -2.98559e-06 -85.6599 0.0930589 31175.8 306.716 0.983504 0.319146 0.734626 0.734622 9.99958 2.98496e-06 1.19397e-05 0.132965 0.98326 0.931629 -0.013292 4.92158e-06 0.510493 -1.96837e-20 7.2882e-24 -1.96764e-20 0.00139611 0.997816 8.59984e-05 0.152685 2.85251 0.00139611 0.997816 0.766454 0.00106241 0.00188094 0.000859984 0.455455 0.00188094 0.442765 0.000130477 1.02 0.888431 0.53447 0.287092 1.71863e-07 3.07723e-09 2375.86 3124.15 -0.0566628 0.482185 0.277361 0.253823 -0.593259 -0.169554 0.492536 -0.266436 -0.22611 2.353 1 0 296.729 0 2.19212 2.351 0.000299449 0.859036 0.686923 0.33015 0.427283 2.19231 136.874 83.8185 18.715 60.8172 0.00402951 0 -40 10
1.452 4.20242e-08 2.53949e-06 0.135892 0.135891 0.0120306 1.91019e-05 0.00115431 0.169865 0.000658617 0.170519 0.92477 101.613 0.238195 0.814905 4.3872 0.061805 0.0413887 0.958611 0.0195924 0.0044708 0.0188531 0.00427667 0.00540759 0.00614689 0.216304 0.245876 58.0303 -87.898 126.218 15.9463 145.03 0.000141617 0.267258 192.777 0.310321 0.0673409 0.00409757 0.000562177 0.00138444 0.986968 0.991721 -2.98561e-06 -85.6599 0.093059 31175.8 306.727 0.983504 0.319146 0.734636 0.734631 9.99958 2.98497e-06 1.19398e-05 0.132969 0.983261 0.931628 -0.013292 4.92161e-06 0.51051 -1.96851e-20 7.28874e-24 -1.96778e-20 0.00139611 0.997816 8.59985e-05 0.152686 2.85251 0.00139611 0.997816 0.766535 0.00106242 0.00188094 0.000859985 0.455455 0.00188094 0.442771 0.000130479 1.02 0.888432 0.53447 0.287094 1.71863e-07 3.07725e-09 2375.84 3124.19 -0.0566671 0.482185 0.27736 0.253826 -0.593258 -0.169554 0.492522 -0.266434 -0.226098 2.354 1 0 296.725 0 2.19226 2.352 0.000299448 0.859059 0.686967 0.330095 0.427306 2.19245 136.882 83.818 18.715 60.8169 0.00402953 0 -40 10
1.453 4.20531e-08 2.53949e-06 0.135934 0.135933 0.0120306 1.91151e-05 0.00115432 0.169918 0.000658618 0.170572 0.924855 101.612 0.238185 0.815031 4.38769 0.0618152 0.0413933 0.958607 0.0195919 0.00447119 0.0188526 0.00427699 0.00540806 0.00614737 0.216323 0.245895 58.0303 -87.898 126.218 15.9463 145.03 0.000141618 0.267258 192.776 0.310321 0.0673408 0.00409757 0.000562178 0.00138444 0.986968 0.991721 -2.98562e-06 -85.6599 0.0930591 31175.8 306.737 0.983504 0.319146 0.734646 0.734641 9.99958 2.98497e-06 1.19398e-05 0.132973 0.983262 0.931627 -0.013292 4.92164e-06 0.510526 -1.96864e-20 7.28929e-24 -1.96791e-20 0.00139611 0.997816 8.59986e-05 0.152686 2.85251 0.00139611 0.997816 0.766616 0.00106244 0.00188094 0.000859986 0.455455 0.00188094 0.442777 0.000130482 1.02 0.888433 0.53447 0.287096 1.71864e-07 3.07727e-09 2375.83 3124.23 -0.0566715 0.482185 0.27736 0.253829 -0.593258 -0.169554 0.492509 -0.266432 -0.226086 2.355 1 0 296.721 0 2.1924 2.353 0.000299447 0.859082 0.687011 0.33004 0.42733 2.19259 136.89 83.8176 18.7149 60.8167 0.00402955 0 -40 10
1.454 4.2082e-08 2.5395e-06 0.135976 0.135975 0.0120306 1.91282e-05 0.00115432 0.16997 0.000658619 0.170624 0.924939 101.612 0.238175 0.815158 4.38817 0.0618254 0.0413979 0.958602 0.0195915 0.00447157 0.0188521 0.00427732 0.00540854 0.00614786 0.216341 0.245914 58.0304 -87.898 126.218 15.9462 145.03 0.00014162 0.267258 192.776 0.31032 0.0673407 0.00409758 0.000562178 0.00138444 0.986968 0.991721 -2.98564e-06 -85.6598 0.0930592 31175.7 306.747 0.983504 0.319146 0.734655 0.734651 9.99958 2.98498e-06 1.19398e-05 0.132977 0.983263 0.931627 -0.013292 4.92167e-06 0.510543 -1.96878e-20 7.28983e-24 -1.96805e-20 0.00139611 0.997816 8.59987e-05 0.152686 2.85251 0.00139611 0.997816 0.766697 0.00106246 0.00188094 0.000859987 0.455454 0.00188094 0.442783 0.000130485 1.02 0.888434 0.534469 0.287097 1.71864e-07 3.0773e-09 2375.81 3124.27 -0.0566758 0.482185 0.27736 0.253831 -0.593257 -0.169554 0.492495 -0.26643 -0.226074 2.356 1 0 296.717 0 2.19254 2.354 0.000299446 0.859105 0.687055 0.329984 0.427353 2.19273 136.897 83.8171 18.7149 60.8165 0.00402957 0 -40 10
1.455 4.21109e-08 2.5395e-06 0.136018 0.136017 0.0120305 1.91413e-05 0.00115432 0.170023 0.00065862 0.170677 0.925024 101.611 0.238164 0.815284 4.38866 0.0618356 0.0414025 0.958598 0.019591 0.00447195 0.0188517 0.00427765 0.00540901 0.00614834 0.21636 0.245934 58.0304 -87.898 126.218 15.9462 145.03 0.000141622 0.267258 192.776 0.31032 0.0673407 0.00409758 0.000562179 0.00138445 0.986968 0.991721 -2.98565e-06 -85.6598 0.0930593 31175.7 306.758 0.983504 0.319146 0.734665 0.734661 9.99958 2.98498e-06 1.19398e-05 0.132981 0.983263 0.931626 -0.013292 4.9217e-06 0.51056 -1.96891e-20 7.29037e-24 -1.96818e-20 0.00139611 0.997816 8.59988e-05 0.152686 2.85251 0.00139611 0.997816 0.766778 0.00106248 0.00188095 0.000859988 0.455454 0.00188094 0.442789 0.000130487 1.02 0.888435 0.534469 0.287099 1.71864e-07 3.07732e-09 2375.8 3124.31 -0.0566802 0.482185 0.27736 0.253834 -0.593257 -0.169555 0.492481 -0.266428 -0.226062 2.357 1 0 296.714 0 2.19268 2.355 0.000299445 0.859128 0.687099 0.329929 0.427376 2.19287 136.905 83.8166 18.7149 60.8162 0.00402959 0 -40 10
1.456 4.21397e-08 2.5395e-06 0.13606 0.136059 0.0120305 1.91544e-05 0.00115432 0.170075 0.000658621 0.170729 0.925109 101.611 0.238154 0.815411 4.38915 0.0618458 0.0414071 0.958593 0.0195905 0.00447234 0.0188512 0.00427798 0.00540948 0.00614882 0.216379 0.245953 58.0305 -87.898 126.217 15.9462 145.03 0.000141624 0.267258 192.776 0.310319 0.0673406 0.00409758 0.00056218 0.00138445 0.986968 0.991721 -2.98567e-06 -85.6598 0.0930593 31175.7 306.768 0.983504 0.319146 0.734675 0.734671 9.99958 2.98499e-06 1.19398e-05 0.132985 0.983264 0.931625 -0.013292 4.92173e-06 0.510576 -1.96904e-20 7.29092e-24 -1.96832e-20 0.00139612 0.997816 8.59988e-05 0.152686 2.85251 0.00139612 0.997816 0.766859 0.00106249 0.00188095 0.000859988 0.455454 0.00188095 0.442795 0.00013049 1.02 0.888436 0.534469 0.2871 1.71865e-07 3.07734e-09 2375.78 3124.35 -0.0566845 0.482185 0.277359 0.253837 -0.593256 -0.169555 0.492467 -0.266425 -0.226051 2.358 1 0 296.71 0 2.19282 2.356 0.000299444 0.859151 0.687144 0.329874 0.427399 2.19301 136.912 83.8161 18.7148 60.816 0.00402961 0 -40 10
1.457 4.21686e-08 2.5395e-06 0.136102 0.136101 0.0120305 1.91675e-05 0.00115432 0.170128 0.000658621 0.170782 0.925194 101.61 0.238144 0.815538 4.38964 0.061856 0.0414117 0.958588 0.01959 0.00447272 0.0188507 0.00427831 0.00540996 0.0061493 0.216398 0.245972 58.0306 -87.898 126.217 15.9461 145.03 0.000141626 0.267259 192.776 0.310319 0.0673406 0.00409758 0.00056218 0.00138445 0.986968 0.991721 -2.98568e-06 -85.6598 0.0930594 31175.7 306.779 0.983504 0.319146 0.734685 0.73468 9.99958 2.98499e-06 1.19399e-05 0.132988 0.983265 0.931624 -0.013292 4.92176e-06 0.510593 -1.96918e-20 7.29146e-24 -1.96845e-20 0.00139612 0.997816 8.59989e-05 0.152686 2.85251 0.00139612 0.997816 0.76694 0.00106251 0.00188095 0.000859989 0.455454 0.00188095 0.442801 0.000130492 1.02 0.888437 0.534468 0.287102 1.71865e-07 3.07737e-09 2375.76 3124.39 -0.0566889 0.482185 0.277359 0.253839 -0.593256 -0.169555 0.492453 -0.266423 -0.226039 2.359 1 0 296.706 0 2.19296 2.357 0.000299443 0.859174 0.687188 0.32982 0.427422 2.19315 136.92 83.8156 18.7148 60.8158 0.00402963 0 -40 10
1.458 4.21975e-08 2.5395e-06 0.136144 0.136143 0.0120305 1.91807e-05 0.00115432 0.17018 0.000658622 0.170834 0.925279 101.61 0.238134 0.815664 4.39013 0.0618662 0.0414163 0.958584 0.0195896 0.00447311 0.0188502 0.00427864 0.00541043 0.00614979 0.216417 0.245991 58.0306 -87.898 126.217 15.9461 145.03 0.000141628 0.267259 192.776 0.310318 0.0673405 0.00409759 0.000562181 0.00138445 0.986968 0.991721 -2.9857e-06 -85.6598 0.0930595 31175.7 306.789 0.983504 0.319146 0.734695 0.73469 9.99958 2.985e-06 1.19399e-05 0.132992 0.983266 0.931624 -0.013292 4.92179e-06 0.510609 -1.96931e-20 7.29201e-24 -1.96859e-20 0.00139612 0.997816 8.5999e-05 0.152686 2.85252 0.00139612 0.997816 0.767021 0.00106253 0.00188095 0.00085999 0.455454 0.00188095 0.442807 0.000130495 1.02 0.888438 0.534468 0.287103 1.71865e-07 3.07739e-09 2375.75 3124.43 -0.0566933 0.482185 0.277359 0.253842 -0.593255 -0.169555 0.492439 -0.266421 -0.226027 2.36 1 0 296.702 0 2.19311 2.358 0.000299442 0.859198 0.687232 0.329765 0.427445 2.19329 136.927 83.8151 18.7148 60.8155 0.00402965 0 -40 10
1.459 4.22264e-08 2.5395e-06 0.136186 0.136185 0.0120305 1.91938e-05 0.00115432 0.170233 0.000658623 0.170887 0.925364 101.609 0.238124 0.815791 4.39062 0.0618764 0.0414209 0.958579 0.0195891 0.00447349 0.0188497 0.00427897 0.00541091 0.00615027 0.216436 0.246011 58.0307 -87.898 126.217 15.9461 145.03 0.00014163 0.267259 192.775 0.310318 0.0673405 0.00409759 0.000562182 0.00138446 0.986968 0.991721 -2.98571e-06 -85.6598 0.0930596 31175.6 306.8 0.983503 0.319146 0.734704 0.7347 9.99958 2.985e-06 1.19399e-05 0.132996 0.983266 0.931623 -0.013292 4.92182e-06 0.510626 -1.96945e-20 7.29255e-24 -1.96872e-20 0.00139612 0.997816 8.59991e-05 0.152687 2.85252 0.00139612 0.997816 0.767102 0.00106255 0.00188095 0.000859991 0.455453 0.00188095 0.442813 0.000130498 1.02 0.888439 0.534468 0.287105 1.71865e-07 3.07741e-09 2375.73 3124.47 -0.0566976 0.482185 0.277358 0.253845 -0.593255 -0.169555 0.492425 -0.266419 -0.226015 2.361 1 0 296.698 0 2.19325 2.359 0.000299441 0.859221 0.687276 0.32971 0.427468 2.19343 136.935 83.8147 18.7148 60.8153 0.00402967 0 -40 10
1.46 4.22552e-08 2.5395e-06 0.136228 0.136227 0.0120305 1.92069e-05 0.00115432 0.170285 0.000658624 0.170939 0.925449 101.609 0.238113 0.815918 4.39111 0.0618866 0.0414255 0.958574 0.0195886 0.00447388 0.0188492 0.0042793 0.00541138 0.00615076 0.216455 0.24603 58.0308 -87.898 126.217 15.946 145.03 0.000141632 0.267259 192.775 0.310318 0.0673404 0.00409759 0.000562182 0.00138446 0.986968 0.991721 -2.98573e-06 -85.6598 0.0930597 31175.6 306.81 0.983503 0.319146 0.734714 0.73471 9.99958 2.98501e-06 1.19399e-05 0.133 0.983267 0.931622 -0.013292 4.92185e-06 0.510642 -1.96958e-20 7.29309e-24 -1.96886e-20 0.00139612 0.997816 8.59992e-05 0.152687 2.85252 0.00139612 0.997816 0.767183 0.00106256 0.00188095 0.000859992 0.455453 0.00188095 0.442819 0.0001305 1.02 0.88844 0.534467 0.287106 1.71866e-07 3.07744e-09 2375.71 3124.51 -0.056702 0.482186 0.277358 0.253847 -0.593254 -0.169555 0.492411 -0.266417 -0.226003 2.362 1 0 296.694 0 2.19339 2.36 0.00029944 0.859244 0.68732 0.329655 0.427491 2.19358 136.943 83.8142 18.7147 60.8151 0.00402969 0 -40 10
1.461 4.22841e-08 2.5395e-06 0.13627 0.136269 0.0120305 1.922e-05 0.00115432 0.170337 0.000658624 0.170991 0.925533 101.608 0.238103 0.816044 4.3916 0.0618968 0.0414302 0.95857 0.0195881 0.00447426 0.0188488 0.00427963 0.00541185 0.00615124 0.216474 0.24605 58.0308 -87.898 126.217 15.946 145.03 0.000141634 0.267259 192.775 0.310317 0.0673404 0.0040976 0.000562183 0.00138446 0.986968 0.991721 -2.98574e-06 -85.6598 0.0930598 31175.6 306.821 0.983503 0.319146 0.734724 0.73472 9.99958 2.98501e-06 1.19399e-05 0.133004 0.983268 0.931622 -0.013292 4.92188e-06 0.510659 -1.96972e-20 7.29364e-24 -1.96899e-20 0.00139612 0.997816 8.59992e-05 0.152687 2.85252 0.00139612 0.997816 0.767264 0.00106258 0.00188096 0.000859992 0.455453 0.00188095 0.442825 0.000130503 1.02 0.888442 0.534467 0.287108 1.71866e-07 3.07746e-09 2375.7 3124.55 -0.0567064 0.482186 0.277358 0.25385 -0.593254 -0.169555 0.492396 -0.266415 -0.225991 2.363 1 0 296.69 0 2.19353 2.361 0.00029944 0.859267 0.687364 0.329601 0.427514 2.19372 136.95 83.8137 18.7147 60.8148 0.00402971 0 -40 10
1.462 4.2313e-08 2.53951e-06 0.136312 0.136311 0.0120304 1.92332e-05 0.00115432 0.170389 0.000658625 0.171043 0.925618 101.608 0.238093 0.816171 4.39209 0.061907 0.0414348 0.958565 0.0195877 0.00447465 0.0188483 0.00427996 0.00541233 0.00615172 0.216493 0.246069 58.0309 -87.8981 126.216 15.9459 145.03 0.000141635 0.26726 192.775 0.310317 0.0673403 0.0040976 0.000562184 0.00138446 0.986968 0.991721 -2.98576e-06 -85.6598 0.0930599 31175.6 306.831 0.983503 0.319146 0.734734 0.73473 9.99958 2.98502e-06 1.194e-05 0.133008 0.983269 0.931621 -0.013292 4.92191e-06 0.510675 -1.96985e-20 7.29418e-24 -1.96913e-20 0.00139612 0.997816 8.59993e-05 0.152687 2.85252 0.00139612 0.997816 0.767344 0.0010626 0.00188096 0.000859993 0.455453 0.00188096 0.442831 0.000130506 1.02 0.888443 0.534467 0.287109 1.71866e-07 3.07748e-09 2375.68 3124.6 -0.0567108 0.482186 0.277358 0.253853 -0.593253 -0.169555 0.492382 -0.266413 -0.225979 2.364 1 0 296.686 0 2.19367 2.362 0.000299439 0.859291 0.687408 0.329546 0.427537 2.19386 136.958 83.8132 18.7147 60.8146 0.00402973 0 -40 10
1.463 4.23418e-08 2.53951e-06 0.136353 0.136353 0.0120304 1.92463e-05 0.00115432 0.170442 0.000658626 0.171096 0.925703 101.607 0.238083 0.816298 4.39258 0.0619172 0.0414394 0.958561 0.0195872 0.00447504 0.0188478 0.00428029 0.00541281 0.00615221 0.216512 0.246088 58.031 -87.8981 126.216 15.9459 145.03 0.000141637 0.26726 192.775 0.310316 0.0673403 0.0040976 0.000562184 0.00138446 0.986968 0.991721 -2.98577e-06 -85.6598 0.09306 31175.5 306.842 0.983503 0.319146 0.734744 0.73474 9.99958 2.98502e-06 1.194e-05 0.133012 0.983269 0.93162 -0.013292 4.92194e-06 0.510692 -1.96999e-20 7.29473e-24 -1.96926e-20 0.00139612 0.997816 8.59994e-05 0.152687 2.85252 0.00139612 0.997816 0.767425 0.00106261 0.00188096 0.000859994 0.455452 0.00188096 0.442837 0.000130508 1.02 0.888444 0.534467 0.287111 1.71866e-07 3.0775e-09 2375.66 3124.64 -0.0567151 0.482186 0.277357 0.253855 -0.593253 -0.169555 0.492368 -0.266411 -0.225967 2.365 1 0 296.682 0 2.19381 2.363 0.000299438 0.859314 0.687453 0.329492 0.42756 2.194 136.965 83.8127 18.7146 60.8144 0.00402975 0 -40 10
1.464 4.23707e-08 2.53951e-06 0.136395 0.136394 0.0120304 1.92594e-05 0.00115432 0.170494 0.000658627 0.171148 0.925788 101.607 0.238073 0.816425 4.39307 0.0619274 0.0414441 0.958556 0.0195867 0.00447542 0.0188473 0.00428062 0.00541328 0.00615269 0.216531 0.246108 58.031 -87.8981 126.216 15.9459 145.03 0.000141639 0.26726 192.775 0.310316 0.0673402 0.00409761 0.000562185 0.00138447 0.986968 0.991721 -2.98579e-06 -85.6597 0.09306 31175.5 306.852 0.983503 0.319146 0.734754 0.734749 9.99958 2.98503e-06 1.194e-05 0.133016 0.98327 0.931619 -0.013292 4.92197e-06 0.510709 -1.97013e-20 7.29528e-24 -1.9694e-20 0.00139613 0.997816 8.59995e-05 0.152687 2.85252 0.00139613 0.997816 0.767506 0.00106263 0.00188096 0.000859995 0.455452 0.00188096 0.442843 0.000130511 1.02 0.888445 0.534466 0.287112 1.71867e-07 3.07753e-09 2375.65 3124.68 -0.0567195 0.482186 0.277357 0.253858 -0.593252 -0.169555 0.492354 -0.266409 -0.225955 2.366 1 0 296.678 0 2.19395 2.364 0.000299437 0.859337 0.687497 0.329437 0.427583 2.19414 136.973 83.8122 18.7146 60.8141 0.00402977 0 -40 10
1.465 4.23996e-08 2.53951e-06 0.136437 0.136436 0.0120304 1.92725e-05 0.00115432 0.170546 0.000658628 0.1712 0.925873 101.606 0.238062 0.816552 4.39356 0.0619376 0.0414487 0.958551 0.0195862 0.00447581 0.0188468 0.00428095 0.00541376 0.00615318 0.21655 0.246127 58.0311 -87.8981 126.216 15.9458 145.03 0.000141641 0.26726 192.774 0.310315 0.0673402 0.00409761 0.000562186 0.00138447 0.986968 0.991721 -2.9858e-06 -85.6597 0.0930601 31175.5 306.863 0.983503 0.319146 0.734764 0.734759 9.99958 2.98503e-06 1.194e-05 0.13302 0.983271 0.931619 -0.013292 4.922e-06 0.510725 -1.97026e-20 7.29582e-24 -1.96953e-20 0.00139613 0.997816 8.59996e-05 0.152688 2.85252 0.00139613 0.997816 0.767587 0.00106265 0.00188096 0.000859996 0.455452 0.00188096 0.442849 0.000130514 1.02 0.888446 0.534466 0.287114 1.71867e-07 3.07755e-09 2375.63 3124.72 -0.0567239 0.482186 0.277357 0.253861 -0.593252 -0.169555 0.49234 -0.266406 -0.225943 2.367 1 0 296.674 0 2.19409 2.365 0.000299436 0.859361 0.687541 0.329383 0.427606 2.19428 136.98 83.8117 18.7146 60.8139 0.00402979 0 -40 10
1.466 4.24285e-08 2.53951e-06 0.136478 0.136478 0.0120304 1.92857e-05 0.00115432 0.170598 0.000658628 0.171252 0.925958 101.606 0.238052 0.816678 4.39406 0.0619478 0.0414534 0.958547 0.0195858 0.0044762 0.0188463 0.00428128 0.00541423 0.00615367 0.216569 0.246147 58.0311 -87.8981 126.216 15.9458 145.03 0.000141643 0.26726 192.774 0.310315 0.0673401 0.00409761 0.000562186 0.00138447 0.986967 0.991721 -2.98582e-06 -85.6597 0.0930602 31175.5 306.873 0.983503 0.319146 0.734774 0.734769 9.99958 2.98504e-06 1.194e-05 0.133024 0.983272 0.931618 -0.013292 4.92203e-06 0.510742 -1.9704e-20 7.29637e-24 -1.96967e-20 0.00139613 0.997816 8.59996e-05 0.152688 2.85252 0.00139613 0.997816 0.767667 0.00106267 0.00188096 0.000859996 0.455452 0.00188096 0.442855 0.000130516 1.02 0.888447 0.534466 0.287115 1.71867e-07 3.07757e-09 2375.61 3124.76 -0.0567283 0.482186 0.277356 0.253863 -0.593251 -0.169555 0.492326 -0.266404 -0.225931 2.368 1 0 296.671 0 2.19423 2.366 0.000299435 0.859384 0.687585 0.329329 0.427629 2.19442 136.988 83.8112 18.7146 60.8137 0.00402981 0 -40 10
1.467 4.24573e-08 2.53951e-06 0.13652 0.136519 0.0120304 1.92988e-05 0.00115432 0.17065 0.000658629 0.171304 0.926043 101.605 0.238042 0.816805 4.39455 0.0619581 0.041458 0.958542 0.0195853 0.00447658 0.0188458 0.00428162 0.00541471 0.00615415 0.216588 0.246166 58.0312 -87.8981 126.215 15.9458 145.03 0.000141645 0.26726 192.774 0.310315 0.0673401 0.00409762 0.000562187 0.00138447 0.986967 0.991721 -2.98583e-06 -85.6597 0.0930603 31175.4 306.884 0.983503 0.319146 0.734784 0.734779 9.99958 2.98504e-06 1.19401e-05 0.133028 0.983272 0.931617 -0.013292 4.92206e-06 0.510759 -1.97053e-20 7.29692e-24 -1.9698e-20 0.00139613 0.997816 8.59997e-05 0.152688 2.85252 0.00139613 0.997816 0.767748 0.00106268 0.00188096 0.000859997 0.455451 0.00188096 0.442861 0.000130519 1.02 0.888448 0.534465 0.287117 1.71867e-07 3.0776e-09 2375.6 3124.8 -0.0567327 0.482186 0.277356 0.253866 -0.59325 -0.169555 0.492312 -0.266402 -0.225919 2.369 1 0 296.667 0 2.19437 2.367 0.000299434 0.859408 0.687629 0.329274 0.427652 2.19456 136.995 83.8108 18.7145 60.8134 0.00402983 0 -40 10
1.468 4.24862e-08 2.53951e-06 0.136562 0.136561 0.0120304 1.93119e-05 0.00115432 0.170702 0.00065863 0.171356 0.926129 101.605 0.238032 0.816932 4.39504 0.0619683 0.0414627 0.958537 0.0195848 0.00447697 0.0188454 0.00428195 0.00541519 0.00615464 0.216608 0.246186 58.0313 -87.8981 126.215 15.9457 145.03 0.000141647 0.267261 192.774 0.310314 0.06734 0.00409762 0.000562188 0.00138448 0.986967 0.991721 -2.98585e-06 -85.6597 0.0930604 31175.4 306.894 0.983503 0.319146 0.734793 0.734789 9.99958 2.98505e-06 1.19401e-05 0.133032 0.983273 0.931616 -0.013292 4.92209e-06 0.510775 -1.97067e-20 7.29746e-24 -1.96994e-20 0.00139613 0.997816 8.59998e-05 0.152688 2.85253 0.00139613 0.997816 0.767829 0.0010627 0.00188097 0.000859998 0.455451 0.00188096 0.442867 0.000130522 1.02 0.888449 0.534465 0.287118 1.71868e-07 3.07762e-09 2375.58 3124.84 -0.0567371 0.482186 0.277356 0.253869 -0.59325 -0.169555 0.492298 -0.2664 -0.225907 2.37 1 0 296.663 0 2.19451 2.368 0.000299433 0.859431 0.687673 0.32922 0.427675 2.1947 137.003 83.8103 18.7145 60.8132 0.00402985 0 -40 10
1.469 4.25151e-08 2.53951e-06 0.136603 0.136602 0.0120304 1.9325e-05 0.00115432 0.170754 0.000658631 0.171408 0.926214 101.604 0.238021 0.817059 4.39554 0.0619785 0.0414673 0.958533 0.0195843 0.00447736 0.0188449 0.00428228 0.00541567 0.00615513 0.216627 0.246205 58.0313 -87.8981 126.215 15.9457 145.03 0.000141649 0.267261 192.774 0.310314 0.06734 0.00409762 0.000562188 0.00138448 0.986967 0.991721 -2.98586e-06 -85.6597 0.0930605 31175.4 306.905 0.983503 0.319146 0.734803 0.734799 9.99958 2.98505e-06 1.19401e-05 0.133036 0.983274 0.931616 -0.013292 4.92212e-06 0.510792 -1.9708e-20 7.29801e-24 -1.97007e-20 0.00139613 0.997816 8.59999e-05 0.152688 2.85253 0.00139613 0.997816 0.767909 0.00106272 0.00188097 0.000859999 0.455451 0.00188097 0.442873 0.000130524 1.02 0.88845 0.534465 0.28712 1.71868e-07 3.07764e-09 2375.56 3124.89 -0.0567415 0.482186 0.277356 0.253871 -0.593249 -0.169555 0.492284 -0.266398 -0.225895 2.371 1 0 296.659 0 2.19465 2.369 0.000299432 0.859455 0.687717 0.329166 0.427698 2.19484 137.011 83.8098 18.7145 60.8129 0.00402987 0 -40 10
1.47 4.25439e-08 2.53952e-06 0.136645 0.136644 0.0120303 1.93382e-05 0.00115433 0.170806 0.000658631 0.17146 0.926299 101.604 0.238011 0.817186 4.39603 0.0619887 0.041472 0.958528 0.0195839 0.00447775 0.0188444 0.00428261 0.00541614 0.00615562 0.216646 0.246225 58.0314 -87.8981 126.215 15.9456 145.03 0.000141651 0.267261 192.774 0.310313 0.0673399 0.00409762 0.000562189 0.00138448 0.986967 0.991721 -2.98588e-06 -85.6597 0.0930606 31175.4 306.915 0.983503 0.319146 0.734813 0.734809 9.99958 2.98506e-06 1.19401e-05 0.13304 0.983274 0.931615 -0.013292 4.92215e-06 0.510809 -1.97094e-20 7.29856e-24 -1.97021e-20 0.00139613 0.997816 8.6e-05 0.152688 2.85253 0.00139613 0.997816 0.76799 0.00106273 0.00188097 0.00086 0.455451 0.00188097 0.442879 0.000130527 1.02 0.888451 0.534464 0.287121 1.71868e-07 3.07766e-09 2375.55 3124.93 -0.0567459 0.482186 0.277355 0.253874 -0.593249 -0.169555 0.49227 -0.266396 -0.225883 2.372 1 0 296.655 0 2.1948 2.37 0.000299431 0.859478 0.687761 0.329112 0.427721 2.19498 137.018 83.8093 18.7145 60.8127 0.00402989 0 -40 10
1.471 4.25728e-08 2.53952e-06 0.136686 0.136685 0.0120303 1.93513e-05 0.00115433 0.170858 0.000658632 0.171512 0.926384 101.603 0.238001 0.817313 4.39653 0.061999 0.0414767 0.958523 0.0195834 0.00447814 0.0188439 0.00428295 0.00541662 0.0061561 0.216665 0.246244 58.0315 -87.8981 126.215 15.9456 145.03 0.000141653 0.267261 192.773 0.310313 0.0673399 0.00409763 0.00056219 0.00138448 0.986967 0.991721 -2.98589e-06 -85.6597 0.0930607 31175.4 306.926 0.983503 0.319146 0.734823 0.734819 9.99958 2.98506e-06 1.19401e-05 0.133044 0.983275 0.931614 -0.013292 4.92218e-06 0.510825 -1.97108e-20 7.29911e-24 -1.97035e-20 0.00139613 0.997816 8.6e-05 0.152688 2.85253 0.00139613 0.997816 0.76807 0.00106275 0.00188097 0.00086 0.455451 0.00188097 0.442885 0.000130529 1.02 0.888453 0.534464 0.287123 1.71869e-07 3.07769e-09 2375.53 3124.97 -0.0567503 0.482186 0.277355 0.253877 -0.593248 -0.169556 0.492256 -0.266394 -0.225871 2.373 1 0 296.651 0 2.19494 2.371 0.00029943 0.859502 0.687806 0.329058 0.427744 2.19512 137.026 83.8088 18.7144 60.8125 0.00402991 0 -40 10
1.472 4.26017e-08 2.53952e-06 0.136728 0.136727 0.0120303 1.93644e-05 0.00115433 0.17091 0.000658633 0.171564 0.926469 101.603 0.237991 0.81744 4.39702 0.0620092 0.0414813 0.958519 0.0195829 0.00447852 0.0188434 0.00428328 0.0054171 0.00615659 0.216684 0.246264 58.0315 -87.8981 126.215 15.9456 145.03 0.000141655 0.267261 192.773 0.310312 0.0673398 0.00409763 0.00056219 0.00138448 0.986967 0.991721 -2.98591e-06 -85.6597 0.0930607 31175.3 306.936 0.983503 0.319146 0.734833 0.734829 9.99958 2.98507e-06 1.19402e-05 0.133048 0.983276 0.931614 -0.013292 4.92221e-06 0.510842 -1.97121e-20 7.29966e-24 -1.97048e-20 0.00139613 0.997816 8.60001e-05 0.152689 2.85253 0.00139613 0.997816 0.768151 0.00106277 0.00188097 0.000860001 0.45545 0.00188097 0.442891 0.000130532 1.02 0.888454 0.534464 0.287124 1.71869e-07 3.07771e-09 2375.51 3125.01 -0.0567548 0.482186 0.277355 0.253879 -0.593248 -0.169556 0.492241 -0.266392 -0.225859 2.374 1 0 296.647 0 2.19508 2.372 0.000299429 0.859525 0.68785 0.329004 0.427767 2.19526 137.033 83.8083 18.7144 60.8122 0.00402993 0 -40 10
1.473 4.26306e-08 2.53952e-06 0.136769 0.136768 0.0120303 1.93775e-05 0.00115433 0.170961 0.000658634 0.171615 0.926554 101.602 0.237981 0.817567 4.39752 0.0620194 0.041486 0.958514 0.0195824 0.00447891 0.0188429 0.00428361 0.00541758 0.00615708 0.216703 0.246283 58.0316 -87.8981 126.214 15.9455 145.03 0.000141657 0.267262 192.773 0.310312 0.0673397 0.00409763 0.000562191 0.00138449 0.986967 0.991721 -2.98592e-06 -85.6597 0.0930608 31175.3 306.947 0.983503 0.319146 0.734843 0.734839 9.99958 2.98507e-06 1.19402e-05 0.133052 0.983277 0.931613 -0.013292 4.92224e-06 0.510859 -1.97135e-20 7.3002e-24 -1.97062e-20 0.00139614 0.997816 8.60002e-05 0.152689 2.85253 0.00139614 0.997816 0.768231 0.00106279 0.00188097 0.000860002 0.45545 0.00188097 0.442897 0.000130535 1.02 0.888455 0.534463 0.287126 1.71869e-07 3.07773e-09 2375.5 3125.05 -0.0567592 0.482186 0.277354 0.253882 -0.593247 -0.169556 0.492227 -0.26639 -0.225847 2.375 1 0 296.643 0 2.19522 2.373 0.000299428 0.859549 0.687894 0.32895 0.42779 2.19541 137.041 83.8078 18.7144 60.812 0.00402995 0 -40 10
1.474 4.26594e-08 2.53952e-06 0.136811 0.13681 0.0120303 1.93906e-05 0.00115433 0.171013 0.000658634 0.171667 0.926639 101.602 0.23797 0.817694 4.39802 0.0620297 0.0414907 0.958509 0.0195819 0.0044793 0.0188424 0.00428394 0.00541806 0.00615757 0.216722 0.246303 58.0316 -87.8981 126.214 15.9455 145.03 0.000141658 0.267262 192.773 0.310312 0.0673397 0.00409764 0.000562192 0.00138449 0.986967 0.991721 -2.98594e-06 -85.6597 0.0930609 31175.3 306.957 0.983503 0.319146 0.734853 0.734849 9.99958 2.98508e-06 1.19402e-05 0.133056 0.983277 0.931612 -0.013292 4.92227e-06 0.510876 -1.97148e-20 7.30075e-24 -1.97075e-20 0.00139614 0.997816 8.60003e-05 0.152689 2.85253 0.00139614 0.997816 0.768312 0.0010628 0.00188097 0.000860003 0.45545 0.00188097 0.442903 0.000130537 1.02 0.888456 0.534463 0.287127 1.71869e-07 3.07776e-09 2375.48 3125.09 -0.0567636 0.482187 0.277354 0.253885 -0.593247 -0.169556 0.492213 -0.266388 -0.225835 2.376 1 0 296.639 0 2.19536 2.374 0.000299427 0.859572 0.687938 0.328897 0.427813 2.19555 137.048 83.8073 18.7143 60.8118 0.00402997 0 -40 10
1.475 4.26883e-08 2.53952e-06 0.136852 0.136851 0.0120303 1.94038e-05 0.00115433 0.171065 0.000658635 0.171719 0.926725 101.601 0.23796 0.817821 4.39851 0.0620399 0.0414954 0.958505 0.0195815 0.00447969 0.0188419 0.00428428 0.00541854 0.00615806 0.216742 0.246322 58.0317 -87.8981 126.214 15.9455 145.03 0.00014166 0.267262 192.773 0.310311 0.0673396 0.00409764 0.000562192 0.00138449 0.986967 0.991721 -2.98595e-06 -85.6596 0.093061 31175.3 306.968 0.983503 0.319146 0.734863 0.734859 9.99958 2.98508e-06 1.19402e-05 0.13306 0.983278 0.931611 -0.013292 4.9223e-06 0.510892 -1.97162e-20 7.3013e-24 -1.97089e-20 0.00139614 0.997816 8.60004e-05 0.152689 2.85253 0.00139614 0.997816 0.768392 0.00106282 0.00188098 0.000860004 0.45545 0.00188097 0.442909 0.00013054 1.02 0.888457 0.534463 0.287129 1.7187e-07 3.07778e-09 2375.46 3125.14 -0.056768 0.482187 0.277354 0.253887 -0.593246 -0.169556 0.492199 -0.266385 -0.225823 2.377 1 0 296.635 0 2.1955 2.375 0.000299426 0.859596 0.687982 0.328843 0.427836 2.19569 137.056 83.8068 18.7143 60.8115 0.00402999 0 -40 10
1.476 4.27172e-08 2.53952e-06 0.136893 0.136892 0.0120303 1.94169e-05 0.00115433 0.171117 0.000658636 0.171771 0.92681 101.601 0.23795 0.817949 4.39901 0.0620502 0.0415001 0.9585 0.019581 0.00448008 0.0188415 0.00428461 0.00541902 0.00615855 0.216761 0.246342 58.0318 -87.8981 126.214 15.9454 145.03 0.000141662 0.267262 192.773 0.310311 0.0673396 0.00409764 0.000562193 0.00138449 0.986967 0.991721 -2.98597e-06 -85.6596 0.0930611 31175.2 306.979 0.983503 0.319146 0.734873 0.734869 9.99958 2.98509e-06 1.19402e-05 0.133063 0.983279 0.931611 -0.013292 4.92232e-06 0.510909 -1.97176e-20 7.30185e-24 -1.97103e-20 0.00139614 0.997816 8.60004e-05 0.152689 2.85253 0.00139614 0.997816 0.768473 0.00106284 0.00188098 0.000860004 0.455449 0.00188098 0.442915 0.000130543 1.02 0.888458 0.534463 0.287131 1.7187e-07 3.0778e-09 2375.45 3125.18 -0.0567724 0.482187 0.277354 0.25389 -0.593246 -0.169556 0.492185 -0.266383 -0.225811 2.378 1 0 296.631 0 2.19564 2.376 0.000299425 0.85962 0.688026 0.328789 0.427859 2.19583 137.063 83.8063 18.7143 60.8113 0.00403001 0 -40 10
1.477 4.2746e-08 2.53952e-06 0.136935 0.136934 0.0120302 1.943e-05 0.00115433 0.171168 0.000658637 0.171822 0.926895 101.6 0.23794 0.818076 4.39951 0.0620604 0.0415048 0.958495 0.0195805 0.00448047 0.018841 0.00428495 0.0054195 0.00615904 0.21678 0.246361 58.0318 -87.8981 126.214 15.9454 145.03 0.000141664 0.267262 192.772 0.31031 0.0673395 0.00409765 0.000562194 0.00138449 0.986967 0.991721 -2.98598e-06 -85.6596 0.0930612 31175.2 306.989 0.983503 0.319146 0.734883 0.734879 9.99958 2.98509e-06 1.19403e-05 0.133067 0.983279 0.93161 -0.013292 4.92235e-06 0.510926 -1.97189e-20 7.3024e-24 -1.97116e-20 0.00139614 0.997816 8.60005e-05 0.152689 2.85253 0.00139614 0.997816 0.768553 0.00106285 0.00188098 0.000860005 0.455449 0.00188098 0.442921 0.000130545 1.02 0.888459 0.534462 0.287132 1.7187e-07 3.07783e-09 2375.43 3125.22 -0.0567769 0.482187 0.277353 0.253893 -0.593245 -0.169556 0.49217 -0.266381 -0.225799 2.379 1 0 296.627 0 2.19578 2.377 0.000299424 0.859643 0.68807 0.328736 0.427882 2.19597 137.071 83.8058 18.7143 60.811 0.00403003 0 -40 10
1.478 4.27749e-08 2.53953e-06 0.136976 0.136975 0.0120302 1.94431e-05 0.00115433 0.17122 0.000658637 0.171874 0.92698 101.6 0.237929 0.818203 4.40001 0.0620707 0.0415095 0.958491 0.01958 0.00448086 0.0188405 0.00428528 0.00541998 0.00615953 0.216799 0.246381 58.0319 -87.8981 126.213 15.9453 145.03 0.000141666 0.267263 192.772 0.31031 0.0673395 0.00409765 0.000562194 0.0013845 0.986967 0.991721 -2.986e-06 -85.6596 0.0930613 31175.2 307 0.983503 0.319146 0.734893 0.734889 9.99958 2.9851e-06 1.19403e-05 0.133071 0.98328 0.931609 -0.013292 4.92238e-06 0.510943 -1.97203e-20 7.30295e-24 -1.9713e-20 0.00139614 0.997816 8.60006e-05 0.15269 2.85253 0.00139614 0.997816 0.768634 0.00106287 0.00188098 0.000860006 0.455449 0.00188098 0.442927 0.000130548 1.02 0.88846 0.534462 0.287134 1.7187e-07 3.07785e-09 2375.42 3125.26 -0.0567813 0.482187 0.277353 0.253895 -0.593245 -0.169556 0.492156 -0.266379 -0.225787 2.38 1 0 296.623 0 2.19592 2.378 0.000299423 0.859667 0.688114 0.328682 0.427905 2.19611 137.079 83.8053 18.7142 60.8108 0.00403005 0 -40 10
1.479 4.28038e-08 2.53953e-06 0.137017 0.137016 0.0120302 1.94563e-05 0.00115433 0.171271 0.000658638 0.171925 0.927066 101.599 0.237919 0.81833 4.4005 0.0620809 0.0415142 0.958486 0.0195795 0.00448125 0.01884 0.00428561 0.00542046 0.00616002 0.216818 0.246401 58.032 -87.8981 126.213 15.9453 145.03 0.000141668 0.267263 192.772 0.310309 0.0673394 0.00409765 0.000562195 0.0013845 0.986967 0.991721 -2.98601e-06 -85.6596 0.0930614 31175.2 307.01 0.983503 0.319146 0.734903 0.734899 9.99958 2.9851e-06 1.19403e-05 0.133075 0.983281 0.931608 -0.013292 4.92241e-06 0.51096 -1.97217e-20 7.3035e-24 -1.97144e-20 0.00139614 0.997816 8.60007e-05 0.15269 2.85254 0.00139614 0.997816 0.768714 0.00106289 0.00188098 0.000860007 0.455449 0.00188098 0.442933 0.00013055 1.02 0.888461 0.534462 0.287135 1.71871e-07 3.07787e-09 2375.4 3125.3 -0.0567858 0.482187 0.277353 0.253898 -0.593244 -0.169556 0.492142 -0.266377 -0.225774 2.381 1 0 296.619 0 2.19606 2.379 0.000299422 0.859691 0.688158 0.328629 0.427928 2.19625 137.086 83.8048 18.7142 60.8106 0.00403007 0 -40 10
1.48 4.28326e-08 2.53953e-06 0.137058 0.137058 0.0120302 1.94694e-05 0.00115433 0.171323 0.000658639 0.171977 0.927151 101.599 0.237909 0.818457 4.401 0.0620912 0.0415189 0.958481 0.0195791 0.00448164 0.0188395 0.00428595 0.00542094 0.00616051 0.216838 0.24642 58.032 -87.8981 126.213 15.9453 145.03 0.00014167 0.267263 192.772 0.310309 0.0673394 0.00409765 0.000562196 0.0013845 0.986967 0.991721 -2.98603e-06 -85.6596 0.0930614 31175.2 307.021 0.983503 0.319146 0.734913 0.734909 9.99958 2.98511e-06 1.19403e-05 0.133079 0.983281 0.931608 -0.013292 4.92244e-06 0.510976 -1.9723e-20 7.30405e-24 -1.97157e-20 0.00139614 0.997816 8.60008e-05 0.15269 2.85254 0.00139614 0.997816 0.768794 0.00106291 0.00188098 0.000860008 0.455449 0.00188098 0.442939 0.000130553 1.02 0.888462 0.534461 0.287137 1.71871e-07 3.07789e-09 2375.38 3125.35 -0.0567902 0.482187 0.277352 0.253901 -0.593244 -0.169556 0.492128 -0.266375 -0.225762 2.382 1 0 296.615 0 2.1962 2.38 0.000299421 0.859715 0.688202 0.328575 0.427951 2.19639 137.094 83.8043 18.7142 60.8103 0.00403009 0 -40 10
1.481 4.28615e-08 2.53953e-06 0.137099 0.137099 0.0120302 1.94825e-05 0.00115433 0.171374 0.00065864 0.172028 0.927236 101.598 0.237899 0.818585 4.4015 0.0621014 0.0415236 0.958476 0.0195786 0.00448203 0.018839 0.00428628 0.00542142 0.006161 0.216857 0.24644 58.0321 -87.8981 126.213 15.9452 145.03 0.000141672 0.267263 192.772 0.310309 0.0673393 0.00409766 0.000562196 0.0013845 0.986967 0.991721 -2.98604e-06 -85.6596 0.0930615 31175.1 307.032 0.983503 0.319146 0.734924 0.734919 9.99958 2.98511e-06 1.19403e-05 0.133083 0.983282 0.931607 -0.013292 4.92247e-06 0.510993 -1.97244e-20 7.30461e-24 -1.97171e-20 0.00139614 0.997816 8.60008e-05 0.15269 2.85254 0.00139614 0.997816 0.768874 0.00106292 0.00188099 0.000860008 0.455448 0.00188098 0.442944 0.000130556 1.02 0.888464 0.534461 0.287138 1.71871e-07 3.07792e-09 2375.37 3125.39 -0.0567946 0.482187 0.277352 0.253904 -0.593243 -0.169556 0.492114 -0.266373 -0.22575 2.383 1 0 296.611 0 2.19634 2.381 0.00029942 0.859738 0.688246 0.328522 0.427974 2.19653 137.101 83.8038 18.7141 60.8101 0.00403011 0 -40 10
1.482 4.28904e-08 2.53953e-06 0.137141 0.13714 0.0120302 1.94956e-05 0.00115433 0.171426 0.00065864 0.17208 0.927322 101.598 0.237888 0.818712 4.402 0.0621117 0.0415283 0.958472 0.0195781 0.00448242 0.0188385 0.00428662 0.0054219 0.00616149 0.216876 0.24646 58.0322 -87.8981 126.213 15.9452 145.03 0.000141674 0.267263 192.772 0.310308 0.0673393 0.00409766 0.000562197 0.00138451 0.986967 0.991721 -2.98606e-06 -85.6596 0.0930616 31175.1 307.042 0.983503 0.319146 0.734934 0.734929 9.99958 2.98512e-06 1.19404e-05 0.133087 0.983283 0.931606 -0.013292 4.9225e-06 0.51101 -1.97258e-20 7.30516e-24 -1.97185e-20 0.00139615 0.997816 8.60009e-05 0.15269 2.85254 0.00139615 0.997816 0.768955 0.00106294 0.00188099 0.000860009 0.455448 0.00188099 0.44295 0.000130558 1.02 0.888465 0.534461 0.28714 1.71872e-07 3.07794e-09 2375.35 3125.43 -0.0567991 0.482187 0.277352 0.253906 -0.593242 -0.169556 0.492099 -0.266371 -0.225738 2.384 1 0 296.607 0 2.19648 2.382 0.000299419 0.859762 0.68829 0.328469 0.427997 2.19667 137.109 83.8033 18.7141 60.8098 0.00403014 0 -40 10
1.483 4.29193e-08 2.53953e-06 0.137182 0.137181 0.0120302 1.95088e-05 0.00115433 0.171477 0.000658641 0.172131 0.927407 101.597 0.237878 0.818839 4.4025 0.0621219 0.041533 0.958467 0.0195776 0.00448282 0.018838 0.00428695 0.00542239 0.00616198 0.216895 0.246479 58.0322 -87.8981 126.213 15.9452 145.03 0.000141676 0.267264 192.771 0.310308 0.0673392 0.00409766 0.000562198 0.00138451 0.986967 0.991721 -2.98607e-06 -85.6596 0.0930617 31175.1 307.053 0.983503 0.319146 0.734944 0.734939 9.99958 2.98512e-06 1.19404e-05 0.133091 0.983284 0.931605 -0.013292 4.92253e-06 0.511027 -1.97271e-20 7.30571e-24 -1.97198e-20 0.00139615 0.997816 8.6001e-05 0.15269 2.85254 0.00139615 0.997816 0.769035 0.00106296 0.00188099 0.00086001 0.455448 0.00188099 0.442956 0.000130561 1.02 0.888466 0.53446 0.287141 1.71872e-07 3.07796e-09 2375.33 3125.47 -0.0568035 0.482187 0.277352 0.253909 -0.593242 -0.169556 0.492085 -0.266369 -0.225726 2.385 1 0 296.603 0 2.19662 2.383 0.000299418 0.859786 0.688334 0.328416 0.42802 2.19681 137.116 83.8028 18.7141 60.8096 0.00403016 0 -40 10
1.484 4.29481e-08 2.53953e-06 0.137223 0.137222 0.0120301 1.95219e-05 0.00115433 0.171528 0.000658642 0.172182 0.927493 101.597 0.237868 0.818966 4.403 0.0621322 0.0415378 0.958462 0.0195771 0.00448321 0.0188375 0.00428729 0.00542287 0.00616248 0.216915 0.246499 58.0323 -87.8981 126.212 15.9451 145.03 0.000141678 0.267264 192.771 0.310307 0.0673392 0.00409767 0.000562198 0.00138451 0.986967 0.991721 -2.98609e-06 -85.6596 0.0930618 31175.1 307.063 0.983503 0.319146 0.734954 0.734949 9.99958 2.98513e-06 1.19404e-05 0.133095 0.983284 0.931605 -0.013292 4.92256e-06 0.511044 -1.97285e-20 7.30626e-24 -1.97212e-20 0.00139615 0.997816 8.60011e-05 0.15269 2.85254 0.00139615 0.997816 0.769115 0.00106297 0.00188099 0.000860011 0.455448 0.00188099 0.442962 0.000130564 1.02 0.888467 0.53446 0.287143 1.71872e-07 3.07799e-09 2375.32 3125.51 -0.056808 0.482187 0.277351 0.253912 -0.593241 -0.169556 0.492071 -0.266366 -0.225714 2.386 1 0 296.599 0 2.19676 2.384 0.000299417 0.85981 0.688378 0.328362 0.428043 2.19695 137.124 83.8023 18.714 60.8094 0.00403018 0 -40 10
1.485 4.2977e-08 2.53953e-06 0.137264 0.137263 0.0120301 1.9535e-05 0.00115433 0.17158 0.000658643 0.172234 0.927578 101.596 0.237858 0.819094 4.40351 0.0621425 0.0415425 0.958457 0.0195767 0.0044836 0.018837 0.00428763 0.00542335 0.00616297 0.216934 0.246519 58.0323 -87.8981 126.212 15.9451 145.03 0.00014168 0.267264 192.771 0.310307 0.0673391 0.00409767 0.000562199 0.00138451 0.986967 0.991721 -2.9861e-06 -85.6596 0.0930619 31175 307.074 0.983503 0.319146 0.734964 0.73496 9.99958 2.98513e-06 1.19404e-05 0.133099 0.983285 0.931604 -0.013292 4.92259e-06 0.511061 -1.97299e-20 7.30681e-24 -1.97226e-20 0.00139615 0.997816 8.60012e-05 0.152691 2.85254 0.00139615 0.997816 0.769195 0.00106299 0.00188099 0.000860012 0.455447 0.00188099 0.442968 0.000130566 1.02 0.888468 0.53446 0.287144 1.71872e-07 3.07801e-09 2375.3 3125.56 -0.0568125 0.482187 0.277351 0.253914 -0.593241 -0.169556 0.492056 -0.266364 -0.225701 2.387 1 0 296.595 0 2.19691 2.385 0.000299416 0.859834 0.688422 0.328309 0.428066 2.19709 137.131 83.8018 18.714 60.8091 0.0040302 0 -40 10
1.486 4.30059e-08 2.53954e-06 0.137305 0.137304 0.0120301 1.95481e-05 0.00115433 0.171631 0.000658643 0.172285 0.927663 101.596 0.237847 0.819221 4.40401 0.0621527 0.0415472 0.958453 0.0195762 0.00448399 0.0188365 0.00428796 0.00542383 0.00616346 0.216953 0.246538 58.0324 -87.8981 126.212 15.945 145.03 0.000141682 0.267264 192.771 0.310306 0.0673391 0.00409767 0.0005622 0.00138451 0.986967 0.991721 -2.98612e-06 -85.6595 0.093062 31175 307.085 0.983503 0.319146 0.734974 0.73497 9.99958 2.98514e-06 1.19404e-05 0.133103 0.983286 0.931603 -0.013292 4.92262e-06 0.511077 -1.97312e-20 7.30737e-24 -1.97239e-20 0.00139615 0.997816 8.60013e-05 0.152691 2.85254 0.00139615 0.997816 0.769275 0.00106301 0.00188099 0.000860013 0.455447 0.00188099 0.442974 0.000130569 1.02 0.888469 0.534459 0.287146 1.71873e-07 3.07803e-09 2375.28 3125.6 -0.0568169 0.482187 0.277351 0.253917 -0.59324 -0.169556 0.492042 -0.266362 -0.225689 2.388 1 0 296.591 0 2.19705 2.386 0.000299415 0.859858 0.688466 0.328256 0.428089 2.19723 137.139 83.8013 18.714 60.8089 0.00403022 0 -40 10
1.487 4.30347e-08 2.53954e-06 0.137346 0.137345 0.0120301 1.95612e-05 0.00115433 0.171682 0.000658644 0.172336 0.927749 101.595 0.237837 0.819349 4.40451 0.062163 0.041552 0.958448 0.0195757 0.00448438 0.018836 0.0042883 0.00542432 0.00616395 0.216973 0.246558 58.0325 -87.8981 126.212 15.945 145.03 0.000141684 0.267264 192.771 0.310306 0.067339 0.00409768 0.0005622 0.00138452 0.986967 0.991721 -2.98613e-06 -85.6595 0.0930621 31175 307.095 0.983503 0.319146 0.734984 0.73498 9.99958 2.98514e-06 1.19405e-05 0.133107 0.983286 0.931602 -0.013292 4.92265e-06 0.511094 -1.97326e-20 7.30792e-24 -1.97253e-20 0.00139615 0.997816 8.60013e-05 0.152691 2.85254 0.00139615 0.997816 0.769355 0.00106303 0.00188099 0.000860013 0.455447 0.00188099 0.44298 0.000130571 1.02 0.88847 0.534459 0.287147 1.71873e-07 3.07805e-09 2375.27 3125.64 -0.0568214 0.482188 0.27735 0.25392 -0.59324 -0.169557 0.492028 -0.26636 -0.225677 2.389 1 0 296.587 0 2.19719 2.387 0.000299414 0.859882 0.68851 0.328203 0.428112 2.19737 137.146 83.8008 18.714 60.8086 0.00403024 0 -40 10
1.488 4.30636e-08 2.53954e-06 0.137387 0.137386 0.0120301 1.95744e-05 0.00115434 0.171733 0.000658645 0.172387 0.927834 101.595 0.237827 0.819476 4.40501 0.0621733 0.0415567 0.958443 0.0195752 0.00448478 0.0188356 0.00428863 0.0054248 0.00616445 0.216992 0.246578 58.0325 -87.8981 126.212 15.945 145.03 0.000141686 0.267264 192.771 0.310306 0.067339 0.00409768 0.000562201 0.00138452 0.986967 0.991721 -2.98615e-06 -85.6595 0.0930621 31175 307.106 0.983503 0.319146 0.734994 0.73499 9.99958 2.98515e-06 1.19405e-05 0.133111 0.983287 0.931602 -0.013292 4.92268e-06 0.511111 -1.9734e-20 7.30847e-24 -1.97267e-20 0.00139615 0.997816 8.60014e-05 0.152691 2.85254 0.00139615 0.997816 0.769436 0.00106304 0.001881 0.000860014 0.455447 0.00188099 0.442986 0.000130574 1.02 0.888471 0.534459 0.287149 1.71873e-07 3.07808e-09 2375.25 3125.68 -0.0568258 0.482188 0.27735 0.253923 -0.593239 -0.169557 0.492014 -0.266358 -0.225665 2.39 1 0 296.583 0 2.19733 2.388 0.000299414 0.859906 0.688554 0.328151 0.428135 2.19751 137.154 83.8003 18.7139 60.8084 0.00403026 0 -40 10
1.489 4.30925e-08 2.53954e-06 0.137428 0.137427 0.0120301 1.95875e-05 0.00115434 0.171784 0.000658646 0.172439 0.92792 101.594 0.237816 0.819603 4.40552 0.0621835 0.0415615 0.958439 0.0195747 0.00448517 0.0188351 0.00428897 0.00542528 0.00616494 0.217011 0.246598 58.0326 -87.8982 126.211 15.9449 145.03 0.000141688 0.267265 192.77 0.310305 0.0673389 0.00409768 0.000562202 0.00138452 0.986967 0.991721 -2.98616e-06 -85.6595 0.0930622 31175 307.117 0.983503 0.319146 0.735004 0.735 9.99958 2.98515e-06 1.19405e-05 0.133115 0.983288 0.931601 -0.013292 4.92271e-06 0.511128 -1.97354e-20 7.30903e-24 -1.9728e-20 0.00139615 0.997816 8.60015e-05 0.152691 2.85254 0.00139615 0.997816 0.769516 0.00106306 0.001881 0.000860015 0.455446 0.001881 0.442992 0.000130577 1.02 0.888472 0.534459 0.28715 1.71873e-07 3.0781e-09 2375.23 3125.73 -0.0568303 0.482188 0.27735 0.253925 -0.593239 -0.169557 0.491999 -0.266356 -0.225653 2.391 1 0 296.579 0 2.19747 2.389 0.000299413 0.85993 0.688598 0.328098 0.428158 2.19765 137.161 83.7998 18.7139 60.8082 0.00403028 0 -40 10
1.49 4.31213e-08 2.53954e-06 0.137468 0.137468 0.0120301 1.96006e-05 0.00115434 0.171836 0.000658646 0.17249 0.928005 101.594 0.237806 0.819731 4.40602 0.0621938 0.0415662 0.958434 0.0195742 0.00448556 0.0188346 0.00428931 0.00542577 0.00616544 0.217031 0.246617 58.0327 -87.8982 126.211 15.9449 145.031 0.00014169 0.267265 192.77 0.310305 0.0673388 0.00409769 0.000562202 0.00138452 0.986967 0.991721 -2.98618e-06 -85.6595 0.0930623 31174.9 307.127 0.983503 0.319146 0.735015 0.73501 9.99958 2.98516e-06 1.19405e-05 0.133119 0.983288 0.9316 -0.013292 4.92274e-06 0.511145 -1.97367e-20 7.30958e-24 -1.97294e-20 0.00139616 0.997816 8.60016e-05 0.152691 2.85255 0.00139615 0.997816 0.769596 0.00106308 0.001881 0.000860016 0.455446 0.001881 0.442998 0.000130579 1.02 0.888473 0.534458 0.287152 1.71874e-07 3.07812e-09 2375.22 3125.77 -0.0568348 0.482188 0.27735 0.253928 -0.593238 -0.169557 0.491985 -0.266354 -0.22564 2.392 1 0 296.575 0 2.19761 2.39 0.000299412 0.859954 0.688642 0.328045 0.428181 2.19779 137.169 83.7993 18.7139 60.8079 0.0040303 0 -40 10
1.491 4.31502e-08 2.53954e-06 0.137509 0.137509 0.01203 1.96137e-05 0.00115434 0.171887 0.000658647 0.172541 0.928091 101.593 0.237796 0.819858 4.40652 0.0622041 0.041571 0.958429 0.0195737 0.00448596 0.0188341 0.00428965 0.00542625 0.00616593 0.21705 0.246637 58.0327 -87.8982 126.211 15.9449 145.031 0.000141692 0.267265 192.77 0.310304 0.0673388 0.00409769 0.000562203 0.00138453 0.986967 0.99172 -2.98619e-06 -85.6595 0.0930624 31174.9 307.138 0.983503 0.319146 0.735025 0.73502 9.99958 2.98516e-06 1.19405e-05 0.133123 0.983289 0.931599 -0.013292 4.92277e-06 0.511162 -1.97381e-20 7.31013e-24 -1.97308e-20 0.00139616 0.997816 8.60017e-05 0.152692 2.85255 0.00139616 0.997816 0.769676 0.00106309 0.001881 0.000860017 0.455446 0.001881 0.443004 0.000130582 1.02 0.888475 0.534458 0.287153 1.71874e-07 3.07815e-09 2375.2 3125.81 -0.0568393 0.482188 0.277349 0.253931 -0.593238 -0.169557 0.49197 -0.266352 -0.225628 2.393 1 0 296.571 0 2.19775 2.391 0.000299411 0.859978 0.688686 0.327992 0.428204 2.19794 137.177 83.7988 18.7138 60.8077 0.00403032 0 -40 10
1.492 4.31791e-08 2.53954e-06 0.13755 0.137549 0.01203 1.96269e-05 0.00115434 0.171938 0.000658648 0.172592 0.928176 101.593 0.237786 0.819986 4.40703 0.0622144 0.0415757 0.958424 0.0195733 0.00448635 0.0188336 0.00428998 0.00542674 0.00616643 0.217069 0.246657 58.0328 -87.8982 126.211 15.9448 145.031 0.000141693 0.267265 192.77 0.310304 0.0673387 0.00409769 0.000562204 0.00138453 0.986967 0.99172 -2.98621e-06 -85.6595 0.0930625 31174.9 307.149 0.983503 0.319146 0.735035 0.735031 9.99958 2.98517e-06 1.19406e-05 0.133127 0.98329 0.931598 -0.013292 4.9228e-06 0.511179 -1.97395e-20 7.31069e-24 -1.97322e-20 0.00139616 0.997816 8.60017e-05 0.152692 2.85255 0.00139616 0.997816 0.769756 0.00106311 0.001881 0.000860017 0.455446 0.001881 0.44301 0.000130585 1.02 0.888476 0.534458 0.287155 1.71874e-07 3.07817e-09 2375.18 3125.85 -0.0568438 0.482188 0.277349 0.253934 -0.593237 -0.169557 0.491956 -0.26635 -0.225616 2.394 1 0 296.567 0 2.19789 2.392 0.00029941 0.860002 0.68873 0.32794 0.428227 2.19808 137.184 83.7983 18.7138 60.8074 0.00403034 0 -40 10
1.493 4.32079e-08 2.53954e-06 0.137591 0.13759 0.01203 1.964e-05 0.00115434 0.171989 0.000658649 0.172643 0.928262 101.592 0.237775 0.820114 4.40753 0.0622246 0.0415805 0.95842 0.0195728 0.00448674 0.0188331 0.00429032 0.00542722 0.00616692 0.217089 0.246677 58.0328 -87.8982 126.211 15.9448 145.031 0.000141695 0.267265 192.77 0.310303 0.0673387 0.00409769 0.000562204 0.00138453 0.986967 0.99172 -2.98622e-06 -85.6595 0.0930626 31174.9 307.159 0.983503 0.319146 0.735045 0.735041 9.99958 2.98517e-06 1.19406e-05 0.133131 0.98329 0.931598 -0.013292 4.92283e-06 0.511196 -1.97409e-20 7.31124e-24 -1.97335e-20 0.00139616 0.997815 8.60018e-05 0.152692 2.85255 0.00139616 0.997816 0.769836 0.00106313 0.001881 0.000860018 0.455446 0.001881 0.443016 0.000130587 1.02 0.888477 0.534457 0.287156 1.71875e-07 3.07819e-09 2375.17 3125.9 -0.0568482 0.482188 0.277349 0.253936 -0.593236 -0.169557 0.491942 -0.266348 -0.225604 2.395 1 0 296.563 0 2.19803 2.393 0.000299409 0.860026 0.688774 0.327887 0.42825 2.19822 137.192 83.7978 18.7138 60.8072 0.00403036 0 -40 10
1.494 4.32368e-08 2.53955e-06 0.137632 0.137631 0.01203 1.96531e-05 0.00115434 0.17204 0.000658649 0.172694 0.928348 101.592 0.237765 0.820241 4.40804 0.0622349 0.0415853 0.958415 0.0195723 0.00448714 0.0188326 0.00429066 0.00542771 0.00616742 0.217108 0.246697 58.0329 -87.8982 126.211 15.9447 145.031 0.000141697 0.267266 192.77 0.310303 0.0673386 0.0040977 0.000562205 0.00138453 0.986967 0.99172 -2.98624e-06 -85.6595 0.0930627 31174.8 307.17 0.983503 0.319146 0.735055 0.735051 9.99958 2.98518e-06 1.19406e-05 0.133135 0.983291 0.931597 -0.013292 4.92286e-06 0.511213 -1.97422e-20 7.3118e-24 -1.97349e-20 0.00139616 0.997815 8.60019e-05 0.152692 2.85255 0.00139616 0.997816 0.769915 0.00106315 0.001881 0.000860019 0.455445 0.001881 0.443022 0.00013059 1.02 0.888478 0.534457 0.287158 1.71875e-07 3.07821e-09 2375.15 3125.94 -0.0568527 0.482188 0.277349 0.253939 -0.593236 -0.169557 0.491927 -0.266345 -0.225591 2.396 1 0 296.559 0 2.19817 2.394 0.000299408 0.86005 0.688818 0.327834 0.428273 2.19836 137.199 83.7973 18.7138 60.807 0.00403038 0 -40 10
1.495 4.32657e-08 2.53955e-06 0.137672 0.137672 0.01203 1.96662e-05 0.00115434 0.17209 0.00065865 0.172744 0.928433 101.591 0.237755 0.820369 4.40854 0.0622452 0.04159 0.95841 0.0195718 0.00448753 0.0188321 0.004291 0.00542819 0.00616791 0.217128 0.246716 58.033 -87.8982 126.21 15.9447 145.031 0.000141699 0.267266 192.769 0.310303 0.0673386 0.0040977 0.000562206 0.00138453 0.986967 0.99172 -2.98625e-06 -85.6595 0.0930628 31174.8 307.181 0.983503 0.319146 0.735066 0.735061 9.99958 2.98518e-06 1.19406e-05 0.133139 0.983292 0.931596 -0.013292 4.92289e-06 0.51123 -1.97436e-20 7.31235e-24 -1.97363e-20 0.00139616 0.997815 8.6002e-05 0.152692 2.85255 0.00139616 0.997816 0.769995 0.00106316 0.00188101 0.00086002 0.455445 0.001881 0.443028 0.000130592 1.02 0.888479 0.534457 0.287159 1.71875e-07 3.07824e-09 2375.13 3125.98 -0.0568572 0.482188 0.277348 0.253942 -0.593235 -0.169557 0.491913 -0.266343 -0.225579 2.397 1 0 296.555 0 2.19831 2.395 0.000299407 0.860074 0.688862 0.327782 0.428295 2.1985 137.207 83.7968 18.7137 60.8067 0.0040304 0 -40 10
1.496 4.32945e-08 2.53955e-06 0.137713 0.137712 0.01203 1.96793e-05 0.00115434 0.172141 0.000658651 0.172795 0.928519 101.591 0.237745 0.820496 4.40905 0.0622555 0.0415948 0.958405 0.0195713 0.00448793 0.0188316 0.00429133 0.00542868 0.00616841 0.217147 0.246736 58.033 -87.8982 126.21 15.9447 145.031 0.000141701 0.267266 192.769 0.310302 0.0673385 0.0040977 0.000562207 0.00138454 0.986967 0.99172 -2.98627e-06 -85.6594 0.0930628 31174.8 307.192 0.983503 0.319146 0.735076 0.735071 9.99958 2.98519e-06 1.19406e-05 0.133144 0.983292 0.931595 -0.013292 4.92292e-06 0.511247 -1.9745e-20 7.31291e-24 -1.97377e-20 0.00139616 0.997815 8.60021e-05 0.152692 2.85255 0.00139616 0.997816 0.770075 0.00106318 0.00188101 0.000860021 0.455445 0.00188101 0.443033 0.000130595 1.02 0.88848 0.534456 0.287161 1.71875e-07 3.07826e-09 2375.12 3126.03 -0.0568617 0.482188 0.277348 0.253945 -0.593235 -0.169557 0.491899 -0.266341 -0.225567 2.398 1 0 296.551 0 2.19845 2.396 0.000299406 0.860098 0.688906 0.32773 0.428318 2.19864 137.214 83.7963 18.7137 60.8065 0.00403042 0 -40 10
1.497 4.33234e-08 2.53955e-06 0.137754 0.137753 0.01203 1.96925e-05 0.00115434 0.172192 0.000658652 0.172846 0.928605 101.59 0.237734 0.820624 4.40956 0.0622658 0.0415996 0.9584 0.0195708 0.00448832 0.0188311 0.00429167 0.00542916 0.00616891 0.217167 0.246756 58.0331 -87.8982 126.21 15.9446 145.031 0.000141703 0.267266 192.769 0.310302 0.0673385 0.00409771 0.000562207 0.00138454 0.986967 0.99172 -2.98628e-06 -85.6594 0.0930629 31174.8 307.202 0.983503 0.319146 0.735086 0.735082 9.99958 2.98519e-06 1.19407e-05 0.133148 0.983293 0.931595 -0.013292 4.92295e-06 0.511264 -1.97464e-20 7.31347e-24 -1.97391e-20 0.00139616 0.997815 8.60021e-05 0.152693 2.85255 0.00139616 0.997816 0.770155 0.0010632 0.00188101 0.000860021 0.455445 0.00188101 0.443039 0.000130598 1.02 0.888481 0.534456 0.287162 1.71876e-07 3.07828e-09 2375.1 3126.07 -0.0568662 0.482188 0.277348 0.253947 -0.593234 -0.169557 0.491884 -0.266339 -0.225555 2.399 1 0 296.547 0 2.19859 2.397 0.000299405 0.860122 0.68895 0.327677 0.428341 2.19878 137.222 83.7958 18.7137 60.8062 0.00403045 0 -40 10
1.498 4.33523e-08 2.53955e-06 0.137794 0.137794 0.01203 1.97056e-05 0.00115434 0.172243 0.000658652 0.172897 0.92869 101.59 0.237724 0.820752 4.41006 0.0622761 0.0416044 0.958396 0.0195703 0.00448872 0.0188306 0.00429201 0.00542965 0.0061694 0.217186 0.246776 58.0332 -87.8982 126.21 15.9446 145.031 0.000141705 0.267266 192.769 0.310301 0.0673384 0.00409771 0.000562208 0.00138454 0.986967 0.99172 -2.9863e-06 -85.6594 0.093063 31174.7 307.213 0.983503 0.319146 0.735096 0.735092 9.99958 2.9852e-06 1.19407e-05 0.133152 0.983294 0.931594 -0.013292 4.92298e-06 0.511281 -1.97478e-20 7.31402e-24 -1.97404e-20 0.00139616 0.997815 8.60022e-05 0.152693 2.85255 0.00139616 0.997816 0.770235 0.00106321 0.00188101 0.000860022 0.455444 0.00188101 0.443045 0.0001306 1.02 0.888482 0.534456 0.287164 1.71876e-07 3.07831e-09 2375.08 3126.11 -0.0568707 0.482188 0.277347 0.25395 -0.593234 -0.169557 0.49187 -0.266337 -0.225542 2.4 1 0 296.543 0 2.19873 2.398 0.000299404 0.860147 0.688994 0.327625 0.428364 2.19892 137.229 83.7953 18.7136 60.806 0.00403047 0 -40 10
1.499 4.33812e-08 2.53955e-06 0.137835 0.137834 0.0120299 1.97187e-05 0.00115434 0.172294 0.000658653 0.172948 0.928776 101.589 0.237714 0.820879 4.41057 0.0622864 0.0416092 0.958391 0.0195699 0.00448911 0.0188301 0.00429235 0.00543014 0.0061699 0.217206 0.246796 58.0332 -87.8982 126.21 15.9446 145.031 0.000141707 0.267267 192.769 0.310301 0.0673384 0.00409771 0.000562209 0.00138454 0.986967 0.99172 -2.98631e-06 -85.6594 0.0930631 31174.7 307.224 0.983503 0.319146 0.735107 0.735102 9.99958 2.9852e-06 1.19407e-05 0.133156 0.983294 0.931593 -0.013292 4.92301e-06 0.511298 -1.97491e-20 7.31458e-24 -1.97418e-20 0.00139617 0.997815 8.60023e-05 0.152693 2.85255 0.00139617 0.997816 0.770315 0.00106323 0.00188101 0.000860023 0.455444 0.00188101 0.443051 0.000130603 1.02 0.888483 0.534455 0.287166 1.71876e-07 3.07833e-09 2375.07 3126.15 -0.0568752 0.482188 0.277347 0.253953 -0.593233 -0.169557 0.491855 -0.266335 -0.22553 2.401 1 0 296.539 0 2.19887 2.399 0.000299403 0.860171 0.689038 0.327573 0.428387 2.19906 137.237 83.7948 18.7136 60.8057 0.00403049 0 -40 10
1.5 4.341e-08 2.53955e-06 0.137875 0.137875 0.0120299 1.97318e-05 0.00115434 0.172344 0.000658654 0.172998 0.928862 101.589 0.237703 0.821007 4.41108 0.0622967 0.041614 0.958386 0.0195694 0.00448951 0.0188296 0.00429269 0.00543063 0.0061704 0.217225 0.246816 58.0333 -87.8982 126.209 15.9445 145.031 0.000141709 0.267267 192.769 0.3103 0.0673383 0.00409772 0.000562209 0.00138454 0.986967 0.99172 -2.98633e-06 -85.6594 0.0930632 31174.7 307.235 0.983503 0.319146 0.735117 0.735112 9.99958 2.98521e-06 1.19407e-05 0.13316 0.983295 0.931592 -0.013292 4.92304e-06 0.511315 -1.97505e-20 7.31514e-24 -1.97432e-20 0.00139617 0.997815 8.60024e-05 0.152693 2.85255 0.00139617 0.997816 0.770394 0.00106325 0.00188101 0.000860024 0.455444 0.00188101 0.443057 0.000130605 1.02 0.888484 0.534455 0.287167 1.71876e-07 3.07835e-09 2375.05 3126.2 -0.0568797 0.482189 0.277347 0.253956 -0.593233 -0.169557 0.491841 -0.266333 -0.225518 2.402 1 0 296.535 0 2.19901 2.4 0.000299402 0.860195 0.689082 0.327521 0.42841 2.1992 137.244 83.7943 18.7136 60.8055 0.00403051 0 -40 10
1.501 4.34389e-08 2.53955e-06 0.137916 0.137915 0.0120299 1.97449e-05 0.00115434 0.172395 0.000658655 0.173049 0.928947 101.588 0.237693 0.821135 4.41159 0.062307 0.0416188 0.958381 0.0195689 0.0044899 0.0188291 0.00429303 0.00543111 0.00617089 0.217245 0.246836 58.0333 -87.8982 126.209 15.9445 145.031 0.000141711 0.267267 192.768 0.3103 0.0673383 0.00409772 0.00056221 0.00138455 0.986967 0.99172 -2.98634e-06 -85.6594 0.0930633 31174.7 307.245 0.983503 0.319146 0.735127 0.735123 9.99958 2.98521e-06 1.19407e-05 0.133164 0.983296 0.931592 -0.013292 4.92307e-06 0.511332 -1.97519e-20 7.31569e-24 -1.97446e-20 0.00139617 0.997815 8.60025e-05 0.152693 2.85256 0.00139617 0.997816 0.770474 0.00106326 0.00188101 0.000860025 0.455444 0.00188101 0.443063 0.000130608 1.02 0.888486 0.534455 0.287169 1.71877e-07 3.07838e-09 2375.04 3126.24 -0.0568842 0.482189 0.277347 0.253958 -0.593232 -0.169557 0.491827 -0.266331 -0.225505 2.403 1 0 296.531 0 2.19915 2.401 0.000299401 0.860219 0.689126 0.327468 0.428433 2.19934 137.252 83.7938 18.7136 60.8052 0.00403053 0 -40 10
1.502 4.34678e-08 2.53956e-06 0.137956 0.137956 0.0120299 1.97581e-05 0.00115434 0.172445 0.000658655 0.1731 0.929033 101.588 0.237683 0.821263 4.4121 0.0623173 0.0416236 0.958376 0.0195684 0.0044903 0.0188286 0.00429337 0.0054316 0.00617139 0.217264 0.246856 58.0334 -87.8982 126.209 15.9444 145.031 0.000141713 0.267267 192.768 0.3103 0.0673382 0.00409772 0.000562211 0.00138455 0.986967 0.99172 -2.98636e-06 -85.6594 0.0930634 31174.7 307.256 0.983503 0.319146 0.735137 0.735133 9.99958 2.98522e-06 1.19408e-05 0.133168 0.983296 0.931591 -0.013292 4.9231e-06 0.511349 -1.97533e-20 7.31625e-24 -1.9746e-20 0.00139617 0.997815 8.60025e-05 0.152693 2.85256 0.00139617 0.997816 0.770554 0.00106328 0.00188102 0.000860025 0.455444 0.00188102 0.443069 0.000130611 1.02 0.888487 0.534455 0.28717 1.71877e-07 3.0784e-09 2375.02 3126.28 -0.0568887 0.482189 0.277346 0.253961 -0.593232 -0.169558 0.491812 -0.266329 -0.225493 2.404 1 0 296.527 0 2.19929 2.402 0.0002994 0.860244 0.68917 0.327416 0.428456 2.19948 137.259 83.7933 18.7135 60.805 0.00403055 0 -40 10
1.503 4.34966e-08 2.53956e-06 0.137997 0.137996 0.0120299 1.97712e-05 0.00115434 0.172496 0.000658656 0.17315 0.929119 101.587 0.237672 0.821391 4.41261 0.0623276 0.0416284 0.958372 0.0195679 0.0044907 0.0188281 0.00429371 0.00543209 0.00617189 0.217284 0.246876 58.0335 -87.8982 126.209 15.9444 145.031 0.000141715 0.267267 192.768 0.310299 0.0673382 0.00409772 0.000562211 0.00138455 0.986966 0.99172 -2.98637e-06 -85.6594 0.0930635 31174.6 307.267 0.983503 0.319146 0.735148 0.735143 9.99958 2.98522e-06 1.19408e-05 0.133172 0.983297 0.93159 -0.013292 4.92313e-06 0.511366 -1.97547e-20 7.31681e-24 -1.97474e-20 0.00139617 0.997815 8.60026e-05 0.152693 2.85256 0.00139617 0.997816 0.770633 0.0010633 0.00188102 0.000860026 0.455443 0.00188102 0.443075 0.000130613 1.02 0.888488 0.534454 0.287172 1.71877e-07 3.07842e-09 2375 3126.33 -0.0568933 0.482189 0.277346 0.253964 -0.593231 -0.169558 0.491798 -0.266326 -0.225481 2.405 1 0 296.523 0 2.19943 2.403 0.000299399 0.860268 0.689214 0.327364 0.428479 2.19962 137.267 83.7928 18.7135 60.8048 0.00403057 0 -40 10
1.504 4.35255e-08 2.53956e-06 0.138037 0.138037 0.0120299 1.97843e-05 0.00115434 0.172547 0.000658657 0.173201 0.929205 101.587 0.237662 0.821518 4.41312 0.0623379 0.0416332 0.958367 0.0195674 0.00449109 0.0188276 0.00429405 0.00543258 0.00617239 0.217303 0.246896 58.0335 -87.8982 126.209 15.9444 145.031 0.000141717 0.267268 192.768 0.310299 0.0673381 0.00409773 0.000562212 0.00138455 0.986966 0.99172 -2.98639e-06 -85.6594 0.0930635 31174.6 307.278 0.983503 0.319146 0.735158 0.735154 9.99958 2.98523e-06 1.19408e-05 0.133176 0.983298 0.931589 -0.013292 4.92316e-06 0.511383 -1.97561e-20 7.31737e-24 -1.97487e-20 0.00139617 0.997815 8.60027e-05 0.152694 2.85256 0.00139617 0.997816 0.770713 0.00106332 0.00188102 0.000860027 0.455443 0.00188102 0.443081 0.000130616 1.02 0.888489 0.534454 0.287173 1.71877e-07 3.07844e-09 2374.99 3126.37 -0.0568978 0.482189 0.277346 0.253967 -0.59323 -0.169558 0.491783 -0.266324 -0.225468 2.406 1 0 296.519 0 2.19957 2.404 0.000299398 0.860292 0.689258 0.327313 0.428502 2.19976 137.274 83.7923 18.7135 60.8045 0.00403059 0 -40 10
1.505 4.35544e-08 2.53956e-06 0.138078 0.138077 0.0120299 1.97974e-05 0.00115435 0.172597 0.000658658 0.173251 0.929291 101.586 0.237652 0.821646 4.41363 0.0623482 0.041638 0.958362 0.0195669 0.00449149 0.0188271 0.00429439 0.00543307 0.00617289 0.217323 0.246916 58.0336 -87.8982 126.208 15.9443 145.031 0.000141719 0.267268 192.768 0.310298 0.0673381 0.00409773 0.000562213 0.00138456 0.986966 0.99172 -2.9864e-06 -85.6594 0.0930636 31174.6 307.288 0.983503 0.319146 0.735168 0.735164 9.99958 2.98523e-06 1.19408e-05 0.13318 0.983298 0.931588 -0.013292 4.92319e-06 0.5114 -1.97574e-20 7.31792e-24 -1.97501e-20 0.00139617 0.997815 8.60028e-05 0.152694 2.85256 0.00139617 0.997816 0.770793 0.00106333 0.00188102 0.000860028 0.455443 0.00188102 0.443087 0.000130619 1.02 0.88849 0.534454 0.287175 1.71878e-07 3.07847e-09 2374.97 3126.41 -0.0569023 0.482189 0.277345 0.253969 -0.59323 -0.169558 0.491769 -0.266322 -0.225456 2.407 1 0 296.515 0 2.19971 2.405 0.000299397 0.860317 0.689302 0.327261 0.428525 2.1999 137.282 83.7918 18.7134 60.8043 0.00403061 0 -40 10
1.506 4.35832e-08 2.53956e-06 0.138118 0.138117 0.0120298 1.98106e-05 0.00115435 0.172647 0.000658658 0.173302 0.929376 101.586 0.237642 0.821774 4.41414 0.0623585 0.0416428 0.958357 0.0195664 0.00449189 0.0188266 0.00429473 0.00543356 0.00617339 0.217342 0.246936 58.0337 -87.8982 126.208 15.9443 145.031 0.000141721 0.267268 192.768 0.310298 0.067338 0.00409773 0.000562213 0.00138456 0.986966 0.99172 -2.98642e-06 -85.6594 0.0930637 31174.6 307.299 0.983503 0.319146 0.735179 0.735174 9.99958 2.98524e-06 1.19408e-05 0.133184 0.983299 0.931588 -0.013292 4.92322e-06 0.511417 -1.97588e-20 7.31848e-24 -1.97515e-20 0.00139617 0.997815 8.60029e-05 0.152694 2.85256 0.00139617 0.997816 0.770872 0.00106335 0.00188102 0.000860029 0.455443 0.00188102 0.443092 0.000130621 1.02 0.888491 0.534453 0.287176 1.71878e-07 3.07849e-09 2374.95 3126.46 -0.0569068 0.482189 0.277345 0.253972 -0.593229 -0.169558 0.491754 -0.26632 -0.225443 2.408 1 0 296.511 0 2.19985 2.406 0.000299396 0.860341 0.689346 0.327209 0.428548 2.20004 137.289 83.7912 18.7134 60.804 0.00403063 0 -40 10
1.507 4.36121e-08 2.53956e-06 0.138158 0.138158 0.0120298 1.98237e-05 0.00115435 0.172698 0.000658659 0.173352 0.929462 101.585 0.237631 0.821902 4.41465 0.0623688 0.0416477 0.958352 0.019566 0.00449228 0.0188261 0.00429507 0.00543404 0.00617389 0.217362 0.246956 58.0337 -87.8982 126.208 15.9443 145.031 0.000141723 0.267268 192.767 0.310297 0.067338 0.00409774 0.000562214 0.00138456 0.986966 0.99172 -2.98643e-06 -85.6593 0.0930638 31174.5 307.31 0.983503 0.319146 0.735189 0.735185 9.99958 2.98524e-06 1.19409e-05 0.133188 0.983299 0.931587 -0.013292 4.92325e-06 0.511435 -1.97602e-20 7.31904e-24 -1.97529e-20 0.00139617 0.997815 8.60029e-05 0.152694 2.85256 0.00139617 0.997816 0.770952 0.00106337 0.00188102 0.000860029 0.455442 0.00188102 0.443098 0.000130624 1.02 0.888492 0.534453 0.287178 1.71878e-07 3.07851e-09 2374.94 3126.5 -0.0569113 0.482189 0.277345 0.253975 -0.593229 -0.169558 0.49174 -0.266318 -0.225431 2.409 1 0 296.507 0 2.19999 2.407 0.000299395 0.860365 0.68939 0.327157 0.42857 2.20018 137.297 83.7907 18.7134 60.8038 0.00403066 0 -40 10
1.508 4.3641e-08 2.53956e-06 0.138199 0.138198 0.0120298 1.98368e-05 0.00115435 0.172748 0.00065866 0.173402 0.929548 101.585 0.237621 0.82203 4.41516 0.0623791 0.0416525 0.958348 0.0195655 0.00449268 0.0188256 0.00429541 0.00543453 0.00617439 0.217381 0.246976 58.0338 -87.8982 126.208 15.9442 145.031 0.000141725 0.267268 192.767 0.310297 0.0673379 0.00409774 0.000562215 0.00138456 0.986966 0.99172 -2.98645e-06 -85.6593 0.0930639 31174.5 307.321 0.983503 0.319146 0.735199 0.735195 9.99958 2.98525e-06 1.19409e-05 0.133192 0.9833 0.931586 -0.013292 4.92327e-06 0.511452 -1.97616e-20 7.3196e-24 -1.97543e-20 0.00139618 0.997815 8.6003e-05 0.152694 2.85256 0.00139618 0.997816 0.771031 0.00106338 0.00188103 0.00086003 0.455442 0.00188102 0.443104 0.000130626 1.02 0.888493 0.534453 0.287179 1.71879e-07 3.07854e-09 2374.92 3126.54 -0.0569159 0.482189 0.277345 0.253978 -0.593228 -0.169558 0.491725 -0.266316 -0.225419 2.41 1 0 296.502 0 2.20013 2.408 0.000299394 0.86039 0.689434 0.327105 0.428593 2.20032 137.305 83.7902 18.7133 60.8035 0.00403068 0 -40 10
1.509 4.36698e-08 2.53956e-06 0.138239 0.138238 0.0120298 1.98499e-05 0.00115435 0.172799 0.00065866 0.173453 0.929634 101.584 0.237611 0.822158 4.41568 0.0623894 0.0416573 0.958343 0.019565 0.00449308 0.0188251 0.00429575 0.00543502 0.00617489 0.217401 0.246996 58.0339 -87.8982 126.208 15.9442 145.031 0.000141727 0.267269 192.767 0.310297 0.0673378 0.00409774 0.000562215 0.00138456 0.986966 0.99172 -2.98646e-06 -85.6593 0.093064 31174.5 307.332 0.983502 0.319146 0.73521 0.735205 9.99958 2.98525e-06 1.19409e-05 0.133196 0.983301 0.931585 -0.013292 4.9233e-06 0.511469 -1.9763e-20 7.32016e-24 -1.97557e-20 0.00139618 0.997815 8.60031e-05 0.152694 2.85256 0.00139618 0.997816 0.771111 0.0010634 0.00188103 0.000860031 0.455442 0.00188103 0.44311 0.000130629 1.02 0.888494 0.534452 0.287181 1.71879e-07 3.07856e-09 2374.9 3126.58 -0.0569204 0.482189 0.277344 0.253981 -0.593228 -0.169558 0.491711 -0.266314 -0.225406 2.411 1 0 296.498 0 2.20027 2.409 0.000299393 0.860414 0.689478 0.327054 0.428616 2.20046 137.312 83.7897 18.7133 60.8033 0.0040307 0 -40 10
1.51 4.36987e-08 2.53957e-06 0.138279 0.138278 0.0120298 1.9863e-05 0.00115435 0.172849 0.000658661 0.173503 0.92972 101.584 0.2376 0.822286 4.41619 0.0623997 0.0416622 0.958338 0.0195645 0.00449348 0.0188246 0.00429609 0.00543551 0.00617539 0.217421 0.247016 58.0339 -87.8982 126.208 15.9441 145.031 0.000141729 0.267269 192.767 0.310296 0.0673378 0.00409775 0.000562216 0.00138457 0.986966 0.99172 -2.98648e-06 -85.6593 0.0930641 31174.5 307.342 0.983502 0.319146 0.73522 0.735216 9.99958 2.98526e-06 1.19409e-05 0.1332 0.983301 0.931584 -0.013292 4.92333e-06 0.511486 -1.97644e-20 7.32072e-24 -1.97571e-20 0.00139618 0.997815 8.60032e-05 0.152695 2.85256 0.00139618 0.997816 0.77119 0.00106342 0.00188103 0.000860032 0.455442 0.00188103 0.443116 0.000130632 1.02 0.888495 0.534452 0.287182 1.71879e-07 3.07858e-09 2374.89 3126.63 -0.0569249 0.482189 0.277344 0.253983 -0.593227 -0.169558 0.491696 -0.266312 -0.225394 2.412 1 0 296.494 0 2.20041 2.41 0.000299392 0.860439 0.689522 0.327002 0.428639 2.2006 137.32 83.7892 18.7133 60.803 0.00403072 0 -40 10
1.511 4.37276e-08 2.53957e-06 0.138319 0.138319 0.0120298 1.98762e-05 0.00115435 0.172899 0.000658662 0.173553 0.929806 101.583 0.23759 0.822414 4.4167 0.06241 0.041667 0.958333 0.019564 0.00449388 0.0188241 0.00429644 0.00543601 0.00617589 0.21744 0.247036 58.034 -87.8982 126.207 15.9441 145.031 0.000141731 0.267269 192.767 0.310296 0.0673377 0.00409775 0.000562217 0.00138457 0.986966 0.99172 -2.98649e-06 -85.6593 0.0930642 31174.5 307.353 0.983502 0.319146 0.73523 0.735226 9.99958 2.98526e-06 1.19409e-05 0.133204 0.983302 0.931584 -0.013292 4.92336e-06 0.511503 -1.97658e-20 7.32128e-24 -1.97585e-20 0.00139618 0.997815 8.60033e-05 0.152695 2.85256 0.00139618 0.997816 0.77127 0.00106343 0.00188103 0.000860033 0.455442 0.00188103 0.443122 0.000130634 1.02 0.888497 0.534452 0.287184 1.71879e-07 3.0786e-09 2374.87 3126.67 -0.0569295 0.482189 0.277344 0.253986 -0.593227 -0.169558 0.491682 -0.26631 -0.225381 2.413 1 0 296.49 0 2.20055 2.411 0.000299391 0.860463 0.689565 0.326951 0.428662 2.20074 137.327 83.7887 18.7133 60.8028 0.00403074 0 -40 10
1.512 4.37564e-08 2.53957e-06 0.138359 0.138359 0.0120298 1.98893e-05 0.00115435 0.172949 0.000658663 0.173603 0.929892 101.583 0.23758 0.822542 4.41721 0.0624204 0.0416718 0.958328 0.0195635 0.00449427 0.0188236 0.00429678 0.0054365 0.00617639 0.21746 0.247056 58.034 -87.8982 126.207 15.9441 145.031 0.000141733 0.267269 192.767 0.310295 0.0673377 0.00409775 0.000562217 0.00138457 0.986966 0.99172 -2.98651e-06 -85.6593 0.0930642 31174.4 307.364 0.983502 0.319146 0.735241 0.735236 9.99958 2.98527e-06 1.1941e-05 0.133208 0.983303 0.931583 -0.0132919 4.92339e-06 0.51152 -1.97672e-20 7.32184e-24 -1.97598e-20 0.00139618 0.997815 8.60034e-05 0.152695 2.85257 0.00139618 0.997816 0.771349 0.00106345 0.00188103 0.000860034 0.455441 0.00188103 0.443128 0.000130637 1.02 0.888498 0.534451 0.287185 1.7188e-07 3.07863e-09 2374.85 3126.71 -0.056934 0.482189 0.277343 0.253989 -0.593226 -0.169558 0.491667 -0.266307 -0.225369 2.414 1 0 296.486 0 2.20069 2.412 0.00029939 0.860488 0.689609 0.326899 0.428685 2.20088 137.335 83.7882 18.7132 60.8025 0.00403076 0 -40 10
1.513 4.37853e-08 2.53957e-06 0.1384 0.138399 0.0120297 1.99024e-05 0.00115435 0.172999 0.000658663 0.173653 0.929978 101.582 0.237569 0.82267 4.41773 0.0624307 0.0416767 0.958323 0.019563 0.00449467 0.0188231 0.00429712 0.00543699 0.0061769 0.21748 0.247076 58.0341 -87.8982 126.207 15.944 145.031 0.000141735 0.267269 192.766 0.310295 0.0673376 0.00409776 0.000562218 0.00138457 0.986966 0.99172 -2.98652e-06 -85.6593 0.0930643 31174.4 307.375 0.983502 0.319146 0.735251 0.735247 9.99958 2.98527e-06 1.1941e-05 0.133212 0.983303 0.931582 -0.0132919 4.92342e-06 0.511538 -1.97686e-20 7.3224e-24 -1.97612e-20 0.00139618 0.997815 8.60034e-05 0.152695 2.85257 0.00139618 0.997816 0.771428 0.00106347 0.00188103 0.000860034 0.455441 0.00188103 0.443134 0.000130639 1.02 0.888499 0.534451 0.287187 1.7188e-07 3.07865e-09 2374.84 3126.76 -0.0569386 0.482189 0.277343 0.253992 -0.593225 -0.169558 0.491653 -0.266305 -0.225357 2.415 1 0 296.482 0 2.20083 2.413 0.000299389 0.860512 0.689653 0.326848 0.428708 2.20102 137.342 83.7877 18.7132 60.8023 0.00403078 0 -40 10
1.514 4.38142e-08 2.53957e-06 0.13844 0.138439 0.0120297 1.99155e-05 0.00115435 0.17305 0.000658664 0.173704 0.930064 101.582 0.237559 0.822798 4.41824 0.062441 0.0416815 0.958318 0.0195625 0.00449507 0.0188226 0.00429746 0.00543748 0.0061774 0.217499 0.247096 58.0342 -87.8982 126.207 15.944 145.031 0.000141737 0.267269 192.766 0.310294 0.0673376 0.00409776 0.000562219 0.00138458 0.986966 0.99172 -2.98654e-06 -85.6593 0.0930644 31174.4 307.386 0.983502 0.319146 0.735261 0.735257 9.99958 2.98528e-06 1.1941e-05 0.133216 0.983304 0.931581 -0.0132919 4.92345e-06 0.511555 -1.977e-20 7.32296e-24 -1.97626e-20 0.00139618 0.997815 8.60035e-05 0.152695 2.85257 0.00139618 0.997816 0.771508 0.00106349 0.00188103 0.000860035 0.455441 0.00188103 0.443139 0.000130642 1.02 0.8885 0.534451 0.287188 1.7188e-07 3.07867e-09 2374.82 3126.8 -0.0569431 0.48219 0.277343 0.253995 -0.593225 -0.169558 0.491638 -0.266303 -0.225344 2.416 1 0 296.478 0 2.20097 2.414 0.000299388 0.860537 0.689697 0.326797 0.428731 2.20116 137.35 83.7872 18.7132 60.8021 0.0040308 0 -40 10
1.515 4.3843e-08 2.53957e-06 0.13848 0.138479 0.0120297 1.99287e-05 0.00115435 0.1731 0.000658665 0.173754 0.93015 101.581 0.237549 0.822926 4.41876 0.0624513 0.0416864 0.958314 0.019562 0.00449547 0.0188221 0.0042978 0.00543797 0.0061779 0.217519 0.247116 58.0342 -87.8982 126.207 15.944 145.031 0.000141739 0.26727 192.766 0.310294 0.0673375 0.00409776 0.000562219 0.00138458 0.986966 0.99172 -2.98655e-06 -85.6593 0.0930645 31174.4 307.396 0.983502 0.319146 0.735272 0.735267 9.99958 2.98528e-06 1.1941e-05 0.13322 0.983304 0.931581 -0.0132919 4.92348e-06 0.511572 -1.97714e-20 7.32353e-24 -1.9764e-20 0.00139618 0.997815 8.60036e-05 0.152695 2.85257 0.00139618 0.997816 0.771587 0.0010635 0.00188104 0.000860036 0.455441 0.00188103 0.443145 0.000130645 1.02 0.888501 0.534451 0.28719 1.7188e-07 3.0787e-09 2374.8 3126.85 -0.0569477 0.48219 0.277343 0.253997 -0.593224 -0.169558 0.491623 -0.266301 -0.225332 2.417 1 0 296.474 0 2.20111 2.415 0.000299387 0.860561 0.689741 0.326745 0.428753 2.2013 137.357 83.7866 18.7131 60.8018 0.00403082 0 -40 10
1.516 4.38719e-08 2.53957e-06 0.13852 0.138519 0.0120297 1.99418e-05 0.00115435 0.17315 0.000658666 0.173804 0.930236 101.581 0.237538 0.823054 4.41927 0.0624617 0.0416913 0.958309 0.0195615 0.00449587 0.0188216 0.00429815 0.00543846 0.0061784 0.217539 0.247136 58.0343 -87.8983 126.206 15.9439 145.031 0.000141741 0.26727 192.766 0.310294 0.0673375 0.00409776 0.00056222 0.00138458 0.986966 0.99172 -2.98657e-06 -85.6593 0.0930646 31174.3 307.407 0.983502 0.319146 0.735282 0.735278 9.99958 2.98529e-06 1.1941e-05 0.133225 0.983305 0.93158 -0.0132919 4.92351e-06 0.511589 -1.97727e-20 7.32409e-24 -1.97654e-20 0.00139618 0.997815 8.60037e-05 0.152695 2.85257 0.00139618 0.997816 0.771666 0.00106352 0.00188104 0.000860037 0.45544 0.00188104 0.443151 0.000130647 1.02 0.888502 0.53445 0.287191 1.71881e-07 3.07872e-09 2374.79 3126.89 -0.0569522 0.48219 0.277342 0.254 -0.593224 -0.169558 0.491609 -0.266299 -0.225319 2.418 1 0 296.47 0 2.20125 2.416 0.000299386 0.860586 0.689785 0.326694 0.428776 2.20144 137.365 83.7861 18.7131 60.8016 0.00403085 0 -40 10
1.517 4.39008e-08 2.53958e-06 0.13856 0.138559 0.0120297 1.99549e-05 0.00115435 0.1732 0.000658666 0.173854 0.930322 101.58 0.237528 0.823182 4.41979 0.062472 0.0416961 0.958304 0.019561 0.00449627 0.0188211 0.00429849 0.00543896 0.00617891 0.217558 0.247156 58.0344 -87.8983 126.206 15.9439 145.031 0.000141743 0.26727 192.766 0.310293 0.0673374 0.00409777 0.000562221 0.00138458 0.986966 0.99172 -2.98658e-06 -85.6593 0.0930647 31174.3 307.418 0.983502 0.319146 0.735293 0.735288 9.99958 2.98529e-06 1.19411e-05 0.133229 0.983306 0.931579 -0.0132919 4.92354e-06 0.511606 -1.97741e-20 7.32465e-24 -1.97668e-20 0.00139619 0.997815 8.60038e-05 0.152696 2.85257 0.00139619 0.997816 0.771746 0.00106354 0.00188104 0.000860038 0.45544 0.00188104 0.443157 0.00013065 1.02 0.888503 0.53445 0.287193 1.71881e-07 3.07874e-09 2374.77 3126.93 -0.0569568 0.48219 0.277342 0.254003 -0.593223 -0.169558 0.491594 -0.266297 -0.225307 2.419 1 0 296.466 0 2.2014 2.417 0.000299385 0.860611 0.689829 0.326643 0.428799 2.20158 137.372 83.7856 18.7131 60.8013 0.00403087 0 -40 10
1.518 4.39296e-08 2.53958e-06 0.1386 0.138599 0.0120297 1.9968e-05 0.00115435 0.17325 0.000658667 0.173904 0.930408 101.58 0.237518 0.82331 4.42031 0.0624823 0.041701 0.958299 0.0195606 0.00449667 0.0188206 0.00429883 0.00543945 0.00617941 0.217578 0.247176 58.0344 -87.8983 126.206 15.9438 145.031 0.000141745 0.26727 192.766 0.310293 0.0673374 0.00409777 0.000562221 0.00138458 0.986966 0.99172 -2.9866e-06 -85.6592 0.0930648 31174.3 307.429 0.983502 0.319146 0.735303 0.735299 9.99958 2.9853e-06 1.19411e-05 0.133233 0.983306 0.931578 -0.0132919 4.92357e-06 0.511624 -1.97755e-20 7.32521e-24 -1.97682e-20 0.00139619 0.997815 8.60038e-05 0.152696 2.85257 0.00139619 0.997816 0.771825 0.00106355 0.00188104 0.000860038 0.45544 0.00188104 0.443163 0.000130652 1.02 0.888504 0.53445 0.287194 1.71881e-07 3.07876e-09 2374.75 3126.98 -0.0569614 0.48219 0.277342 0.254006 -0.593223 -0.169559 0.49158 -0.266295 -0.225294 2.42 1 0 296.462 0 2.20154 2.418 0.000299384 0.860635 0.689873 0.326592 0.428822 2.20172 137.38 83.7851 18.713 60.8011 0.00403089 0 -40 10
1.519 4.39585e-08 2.53958e-06 0.13864 0.138639 0.0120297 1.99811e-05 0.00115435 0.173299 0.000658668 0.173954 0.930494 101.579 0.237507 0.823439 4.42082 0.0624927 0.0417059 0.958294 0.0195601 0.00449707 0.0188201 0.00429918 0.00543994 0.00617991 0.217598 0.247197 58.0345 -87.8983 126.206 15.9438 145.031 0.000141747 0.26727 192.765 0.310292 0.0673373 0.00409777 0.000562222 0.00138459 0.986966 0.99172 -2.98661e-06 -85.6592 0.0930649 31174.3 307.44 0.983502 0.319146 0.735314 0.735309 9.99958 2.9853e-06 1.19411e-05 0.133237 0.983307 0.931577 -0.0132919 4.9236e-06 0.511641 -1.97769e-20 7.32577e-24 -1.97696e-20 0.00139619 0.997815 8.60039e-05 0.152696 2.85257 0.00139619 0.997816 0.771904 0.00106357 0.00188104 0.000860039 0.45544 0.00188104 0.443169 0.000130655 1.02 0.888505 0.534449 0.287196 1.71882e-07 3.07879e-09 2374.74 3127.02 -0.0569659 0.48219 0.277341 0.254009 -0.593222 -0.169559 0.491565 -0.266293 -0.225282 2.421 1 0 296.458 0 2.20168 2.419 0.000299383 0.86066 0.689917 0.326541 0.428845 2.20186 137.387 83.7846 18.713 60.8008 0.00403091 0 -40 10
1.52 4.39874e-08 2.53958e-06 0.138679 0.138679 0.0120297 1.99943e-05 0.00115435 0.173349 0.000658668 0.174003 0.93058 101.579 0.237497 0.823567 4.42134 0.062503 0.0417108 0.958289 0.0195596 0.00449747 0.0188196 0.00429952 0.00544043 0.00618042 0.217617 0.247217 58.0345 -87.8983 126.206 15.9438 145.031 0.000141749 0.267271 192.765 0.310292 0.0673373 0.00409778 0.000562223 0.00138459 0.986966 0.99172 -2.98663e-06 -85.6592 0.0930649 31174.3 307.451 0.983502 0.319146 0.735324 0.73532 9.99958 2.98531e-06 1.19411e-05 0.133241 0.983308 0.931577 -0.0132919 4.92363e-06 0.511658 -1.97783e-20 7.32634e-24 -1.9771e-20 0.00139619 0.997815 8.6004e-05 0.152696 2.85257 0.00139619 0.997816 0.771983 0.00106359 0.00188104 0.00086004 0.455439 0.00188104 0.443174 0.000130657 1.02 0.888506 0.534449 0.287197 1.71882e-07 3.07881e-09 2374.72 3127.06 -0.0569705 0.48219 0.277341 0.254011 -0.593222 -0.169559 0.49155 -0.266291 -0.225269 2.422 1 0 296.453 0 2.20182 2.42 0.000299382 0.860685 0.68996 0.32649 0.428868 2.202 137.395 83.7841 18.713 60.8006 0.00403093 0 -40 10
1.521 4.40162e-08 2.53958e-06 0.138719 0.138719 0.0120296 2.00074e-05 0.00115435 0.173399 0.000658669 0.174053 0.930666 101.578 0.237487 0.823695 4.42186 0.0625134 0.0417156 0.958284 0.0195591 0.00449787 0.0188191 0.00429986 0.00544093 0.00618092 0.217637 0.247237 58.0346 -87.8983 126.205 15.9437 145.031 0.000141751 0.267271 192.765 0.310291 0.0673372 0.00409778 0.000562223 0.00138459 0.986966 0.99172 -2.98664e-06 -85.6592 0.093065 31174.2 307.462 0.983502 0.319146 0.735335 0.73533 9.99958 2.98531e-06 1.19411e-05 0.133245 0.983308 0.931576 -0.0132919 4.92366e-06 0.511675 -1.97797e-20 7.3269e-24 -1.97724e-20 0.00139619 0.997815 8.60041e-05 0.152696 2.85257 0.00139619 0.997816 0.772062 0.00106361 0.00188104 0.000860041 0.455439 0.00188104 0.44318 0.00013066 1.02 0.888508 0.534449 0.287199 1.71882e-07 3.07883e-09 2374.71 3127.11 -0.0569751 0.48219 0.277341 0.254014 -0.593221 -0.169559 0.491536 -0.266289 -0.225257 2.423 1 0 296.449 0 2.20196 2.421 0.000299381 0.860709 0.690004 0.326439 0.428891 2.20214 137.402 83.7836 18.713 60.8003 0.00403095 0 -40 10
1.522 4.40451e-08 2.53958e-06 0.138759 0.138758 0.0120296 2.00205e-05 0.00115436 0.173449 0.00065867 0.174103 0.930753 101.578 0.237476 0.823823 4.42238 0.0625237 0.0417205 0.958279 0.0195586 0.00449827 0.0188186 0.00430021 0.00544142 0.00618143 0.217657 0.247257 58.0347 -87.8983 126.205 15.9437 145.031 0.000141753 0.267271 192.765 0.310291 0.0673372 0.00409778 0.000562224 0.00138459 0.986966 0.99172 -2.98666e-06 -85.6592 0.0930651 31174.2 307.473 0.983502 0.319146 0.735345 0.735341 9.99958 2.98532e-06 1.19412e-05 0.133249 0.983309 0.931575 -0.0132919 4.92369e-06 0.511693 -1.97811e-20 7.32746e-24 -1.97738e-20 0.00139619 0.997815 8.60042e-05 0.152696 2.85257 0.00139619 0.997816 0.772141 0.00106362 0.00188105 0.000860042 0.455439 0.00188105 0.443186 0.000130663 1.02 0.888509 0.534448 0.287201 1.71882e-07 3.07886e-09 2374.69 3127.15 -0.0569796 0.48219 0.277341 0.254017 -0.59322 -0.169559 0.491521 -0.266286 -0.225244 2.424 1 0 296.445 0 2.2021 2.422 0.00029938 0.860734 0.690048 0.326388 0.428913 2.20228 137.41 83.783 18.7129 60.8001 0.00403097 0 -40 10
1.523 4.4074e-08 2.53958e-06 0.138799 0.138798 0.0120296 2.00336e-05 0.00115436 0.173499 0.000658671 0.174153 0.930839 101.577 0.237466 0.823952 4.4229 0.062534 0.0417254 0.958275 0.0195581 0.00449868 0.0188181 0.00430055 0.00544192 0.00618193 0.217677 0.247277 58.0347 -87.8983 126.205 15.9437 145.031 0.000141755 0.267271 192.765 0.310291 0.0673371 0.00409779 0.000562225 0.00138459 0.986966 0.99172 -2.98667e-06 -85.6592 0.0930652 31174.2 307.483 0.983502 0.319146 0.735355 0.735351 9.99958 2.98532e-06 1.19412e-05 0.133253 0.983309 0.931574 -0.0132919 4.92372e-06 0.51171 -1.97825e-20 7.32803e-24 -1.97752e-20 0.00139619 0.997815 8.60042e-05 0.152697 2.85258 0.00139619 0.997816 0.772221 0.00106364 0.00188105 0.000860042 0.455439 0.00188105 0.443192 0.000130665 1.02 0.88851 0.534448 0.287202 1.71883e-07 3.07888e-09 2374.67 3127.2 -0.0569842 0.48219 0.27734 0.25402 -0.59322 -0.169559 0.491507 -0.266284 -0.225232 2.425 1 0 296.441 0 2.20224 2.423 0.000299379 0.860759 0.690092 0.326337 0.428936 2.20242 137.417 83.7825 18.7129 60.7998 0.00403099 0 -40 10
1.524 4.41028e-08 2.53958e-06 0.138839 0.138838 0.0120296 2.00467e-05 0.00115436 0.173548 0.000658671 0.174203 0.930925 101.577 0.237456 0.82408 4.42341 0.0625444 0.0417303 0.95827 0.0195576 0.00449908 0.0188176 0.0043009 0.00544241 0.00618244 0.217696 0.247297 58.0348 -87.8983 126.205 15.9436 145.031 0.000141757 0.267271 192.765 0.31029 0.0673371 0.00409779 0.000562225 0.0013846 0.986966 0.99172 -2.98669e-06 -85.6592 0.0930653 31174.2 307.494 0.983502 0.319146 0.735366 0.735362 9.99958 2.98533e-06 1.19412e-05 0.133257 0.98331 0.931573 -0.0132919 4.92375e-06 0.511727 -1.97839e-20 7.32859e-24 -1.97766e-20 0.00139619 0.997815 8.60043e-05 0.152697 2.85258 0.00139619 0.997816 0.7723 0.00106366 0.00188105 0.000860043 0.455439 0.00188105 0.443198 0.000130668 1.02 0.888511 0.534448 0.287204 1.71883e-07 3.0789e-09 2374.66 3127.24 -0.0569888 0.48219 0.27734 0.254023 -0.593219 -0.169559 0.491492 -0.266282 -0.225219 2.426 1 0 296.437 0 2.20238 2.424 0.000299378 0.860784 0.690136 0.326286 0.428959 2.20256 137.425 83.782 18.7129 60.7996 0.00403102 0 -40 10
1.525 4.41317e-08 2.53959e-06 0.138878 0.138878 0.0120296 2.00599e-05 0.00115436 0.173598 0.000658672 0.174252 0.931011 101.576 0.237445 0.824208 4.42393 0.0625547 0.0417352 0.958265 0.0195571 0.00449948 0.0188171 0.00430124 0.00544291 0.00618294 0.217716 0.247318 58.0349 -87.8983 126.205 15.9436 145.031 0.000141759 0.267272 192.764 0.31029 0.067337 0.00409779 0.000562226 0.0013846 0.986966 0.99172 -2.9867e-06 -85.6592 0.0930654 31174.1 307.505 0.983502 0.319146 0.735376 0.735372 9.99958 2.98533e-06 1.19412e-05 0.133261 0.983311 0.931572 -0.0132919 4.92378e-06 0.511745 -1.97853e-20 7.32916e-24 -1.9778e-20 0.0013962 0.997815 8.60044e-05 0.152697 2.85258 0.0013962 0.997816 0.772379 0.00106367 0.00188105 0.000860044 0.455438 0.00188105 0.443204 0.00013067 1.02 0.888512 0.534447 0.287205 1.71883e-07 3.07893e-09 2374.64 3127.28 -0.0569934 0.48219 0.27734 0.254025 -0.593219 -0.169559 0.491477 -0.26628 -0.225207 2.427 1 0 296.433 0 2.20252 2.425 0.000299377 0.860808 0.69018 0.326236 0.428982 2.2027 137.432 83.7815 18.7128 60.7993 0.00403104 0 -40 10
1.526 4.41606e-08 2.53959e-06 0.138918 0.138917 0.0120296 2.0073e-05 0.00115436 0.173648 0.000658673 0.174302 0.931097 101.576 0.237435 0.824337 4.42445 0.0625651 0.0417401 0.95826 0.0195566 0.00449988 0.0188166 0.00430159 0.0054434 0.00618345 0.217736 0.247338 58.0349 -87.8983 126.204 15.9435 145.031 0.000141761 0.267272 192.764 0.310289 0.067337 0.00409779 0.000562227 0.0013846 0.986966 0.99172 -2.98672e-06 -85.6592 0.0930655 31174.1 307.516 0.983502 0.319146 0.735387 0.735383 9.99958 2.98534e-06 1.19412e-05 0.133265 0.983311 0.931572 -0.0132919 4.92381e-06 0.511762 -1.97867e-20 7.32972e-24 -1.97794e-20 0.0013962 0.997815 8.60045e-05 0.152697 2.85258 0.0013962 0.997816 0.772458 0.00106369 0.00188105 0.000860045 0.455438 0.00188105 0.443209 0.000130673 1.02 0.888513 0.534447 0.287207 1.71883e-07 3.07895e-09 2374.62 3127.33 -0.0569979 0.48219 0.277339 0.254028 -0.593218 -0.169559 0.491463 -0.266278 -0.225194 2.428 1 0 296.429 0 2.20266 2.426 0.000299376 0.860833 0.690224 0.326185 0.429005 2.20284 137.44 83.781 18.7128 60.7991 0.00403106 0 -40 10
1.527 4.41894e-08 2.53959e-06 0.138958 0.138957 0.0120296 2.00861e-05 0.00115436 0.173697 0.000658673 0.174351 0.931184 101.575 0.237425 0.824465 4.42498 0.0625754 0.041745 0.958255 0.0195561 0.00450028 0.018816 0.00430193 0.0054439 0.00618396 0.217756 0.247358 58.035 -87.8983 126.204 15.9435 145.031 0.000141763 0.267272 192.764 0.310289 0.0673369 0.0040978 0.000562227 0.0013846 0.986966 0.99172 -2.98673e-06 -85.6592 0.0930656 31174.1 307.527 0.983502 0.319146 0.735397 0.735393 9.99958 2.98534e-06 1.19413e-05 0.13327 0.983312 0.931571 -0.0132919 4.92384e-06 0.511779 -1.97881e-20 7.33029e-24 -1.97808e-20 0.0013962 0.997815 8.60046e-05 0.152697 2.85258 0.0013962 0.997816 0.772537 0.00106371 0.00188105 0.000860046 0.455438 0.00188105 0.443215 0.000130676 1.02 0.888514 0.534447 0.287208 1.71884e-07 3.07897e-09 2374.61 3127.37 -0.0570025 0.482191 0.277339 0.254031 -0.593218 -0.169559 0.491448 -0.266276 -0.225181 2.429 1 0 296.425 0 2.20279 2.427 0.000299375 0.860858 0.690267 0.326134 0.429028 2.20298 137.447 83.7804 18.7128 60.7988 0.00403108 0 -40 10
1.528 4.42183e-08 2.53959e-06 0.138998 0.138997 0.0120295 2.00992e-05 0.00115436 0.173747 0.000658674 0.174401 0.93127 101.575 0.237414 0.824593 4.4255 0.0625858 0.04175 0.95825 0.0195556 0.00450069 0.0188155 0.00430228 0.00544439 0.00618446 0.217776 0.247378 58.035 -87.8983 126.204 15.9435 145.031 0.000141765 0.267272 192.764 0.310288 0.0673368 0.0040978 0.000562228 0.00138461 0.986966 0.99172 -2.98675e-06 -85.6591 0.0930656 31174.1 307.538 0.983502 0.319146 0.735408 0.735404 9.99958 2.98535e-06 1.19413e-05 0.133274 0.983312 0.93157 -0.0132919 4.92387e-06 0.511797 -1.97896e-20 7.33085e-24 -1.97822e-20 0.0013962 0.997815 8.60046e-05 0.152697 2.85258 0.0013962 0.997816 0.772616 0.00106372 0.00188106 0.000860046 0.455438 0.00188105 0.443221 0.000130678 1.02 0.888515 0.534447 0.28721 1.71884e-07 3.07899e-09 2374.59 3127.41 -0.0570071 0.482191 0.277339 0.254034 -0.593217 -0.169559 0.491433 -0.266274 -0.225169 2.43 1 0 296.421 0 2.20293 2.428 0.000299374 0.860883 0.690311 0.326084 0.42905 2.20312 137.455 83.7799 18.7127 60.7986 0.0040311 0 -40 10
1.529 4.42472e-08 2.53959e-06 0.139037 0.139036 0.0120295 2.01123e-05 0.00115436 0.173796 0.000658675 0.17445 0.931356 101.574 0.237404 0.824722 4.42602 0.0625962 0.0417549 0.958245 0.0195551 0.00450109 0.018815 0.00430262 0.00544489 0.00618497 0.217796 0.247399 58.0351 -87.8983 126.204 15.9434 145.031 0.000141767 0.267272 192.764 0.310288 0.0673368 0.0040978 0.000562229 0.00138461 0.986966 0.99172 -2.98676e-06 -85.6591 0.0930657 31174 307.549 0.983502 0.319146 0.735419 0.735414 9.99958 2.98535e-06 1.19413e-05 0.133278 0.983313 0.931569 -0.0132919 4.9239e-06 0.511814 -1.9791e-20 7.33142e-24 -1.97836e-20 0.0013962 0.997815 8.60047e-05 0.152697 2.85258 0.0013962 0.997816 0.772695 0.00106374 0.00188106 0.000860047 0.455437 0.00188106 0.443227 0.000130681 1.02 0.888516 0.534446 0.287211 1.71884e-07 3.07902e-09 2374.57 3127.46 -0.0570117 0.482191 0.277339 0.254037 -0.593217 -0.169559 0.491419 -0.266272 -0.225156 2.431 1 0 296.416 0 2.20307 2.429 0.000299373 0.860908 0.690355 0.326033 0.429073 2.20326 137.462 83.7794 18.7127 60.7983 0.00403112 0 -40 10
1.53 4.4276e-08 2.53959e-06 0.139077 0.139076 0.0120295 2.01255e-05 0.00115436 0.173846 0.000658675 0.1745 0.931442 101.573 0.237393 0.82485 4.42654 0.0626065 0.0417598 0.95824 0.0195546 0.00450149 0.0188145 0.00430297 0.00544538 0.00618548 0.217815 0.247419 58.0352 -87.8983 126.204 15.9434 145.031 0.000141769 0.267273 192.764 0.310288 0.0673367 0.00409781 0.000562229 0.00138461 0.986966 0.99172 -2.98678e-06 -85.6591 0.0930658 31174 307.56 0.983502 0.319146 0.735429 0.735425 9.99958 2.98536e-06 1.19413e-05 0.133282 0.983314 0.931568 -0.0132919 4.92393e-06 0.511831 -1.97924e-20 7.33198e-24 -1.9785e-20 0.0013962 0.997815 8.60048e-05 0.152698 2.85258 0.0013962 0.997816 0.772774 0.00106376 0.00188106 0.000860048 0.455437 0.00188106 0.443233 0.000130683 1.02 0.888517 0.534446 0.287213 1.71885e-07 3.07904e-09 2374.56 3127.5 -0.0570163 0.482191 0.277338 0.25404 -0.593216 -0.169559 0.491404 -0.26627 -0.225144 2.432 1 0 296.412 0 2.20321 2.43 0.000299372 0.860933 0.690399 0.325983 0.429096 2.2034 137.47 83.7789 18.7127 60.7981 0.00403114 0 -40 10
1.531 4.43049e-08 2.53959e-06 0.139116 0.139116 0.0120295 2.01386e-05 0.00115436 0.173895 0.000658676 0.174549 0.931529 101.573 0.237383 0.824979 4.42706 0.0626169 0.0417647 0.958235 0.0195541 0.00450189 0.018814 0.00430331 0.00544588 0.00618598 0.217835 0.247439 58.0352 -87.8983 126.204 15.9434 145.031 0.000141771 0.267273 192.763 0.310287 0.0673367 0.00409781 0.00056223 0.00138461 0.986966 0.99172 -2.98679e-06 -85.6591 0.0930659 31174 307.571 0.983502 0.319146 0.73544 0.735435 9.99958 2.98536e-06 1.19413e-05 0.133286 0.983314 0.931568 -0.0132919 4.92396e-06 0.511849 -1.97938e-20 7.33255e-24 -1.97864e-20 0.0013962 0.997815 8.60049e-05 0.152698 2.85258 0.0013962 0.997816 0.772852 0.00106377 0.00188106 0.000860049 0.455437 0.00188106 0.443239 0.000130686 1.02 0.888519 0.534446 0.287214 1.71885e-07 3.07906e-09 2374.54 3127.55 -0.0570209 0.482191 0.277338 0.254042 -0.593215 -0.169559 0.491389 -0.266267 -0.225131 2.433 1 0 296.408 0 2.20335 2.431 0.000299371 0.860958 0.690443 0.325933 0.429119 2.20354 137.477 83.7784 18.7127 60.7978 0.00403117 0 -40 10
1.532 4.43337e-08 2.53959e-06 0.139156 0.139155 0.0120295 2.01517e-05 0.00115436 0.173945 0.000658677 0.174599 0.931615 101.572 0.237373 0.825107 4.42758 0.0626272 0.0417697 0.95823 0.0195536 0.0045023 0.0188135 0.00430366 0.00544638 0.00618649 0.217855 0.24746 58.0353 -87.8983 126.203 15.9433 145.031 0.000141774 0.267273 192.763 0.310287 0.0673366 0.00409781 0.000562231 0.00138461 0.986966 0.99172 -2.98681e-06 -85.6591 0.093066 31174 307.582 0.983502 0.319146 0.73545 0.735446 9.99958 2.98536e-06 1.19414e-05 0.13329 0.983315 0.931567 -0.0132919 4.92399e-06 0.511866 -1.97952e-20 7.33312e-24 -1.97878e-20 0.0013962 0.997815 8.6005e-05 0.152698 2.85258 0.0013962 0.997816 0.772931 0.00106379 0.00188106 0.00086005 0.455437 0.00188106 0.443244 0.000130689 1.02 0.88852 0.534445 0.287216 1.71885e-07 3.07909e-09 2374.52 3127.59 -0.0570255 0.482191 0.277338 0.254045 -0.593215 -0.169559 0.491375 -0.266265 -0.225119 2.434 1 0 296.404 0 2.20349 2.432 0.00029937 0.860983 0.690486 0.325882 0.429142 2.20368 137.485 83.7778 18.7126 60.7976 0.00403119 0 -40 10
1.533 4.43626e-08 2.5396e-06 0.139195 0.139195 0.0120295 2.01648e-05 0.00115436 0.173994 0.000658678 0.174648 0.931701 101.572 0.237362 0.825236 4.42811 0.0626376 0.0417746 0.958225 0.0195531 0.0045027 0.018813 0.00430401 0.00544688 0.006187 0.217875 0.24748 58.0354 -87.8983 126.203 15.9433 145.031 0.000141776 0.267273 192.763 0.310286 0.0673366 0.00409782 0.000562231 0.00138462 0.986966 0.99172 -2.98682e-06 -85.6591 0.0930661 31174 307.593 0.983502 0.319146 0.735461 0.735456 9.99958 2.98537e-06 1.19414e-05 0.133294 0.983315 0.931566 -0.0132919 4.92402e-06 0.511884 -1.97966e-20 7.33368e-24 -1.97893e-20 0.0013962 0.997815 8.6005e-05 0.152698 2.85259 0.0013962 0.997816 0.77301 0.00106381 0.00188106 0.00086005 0.455437 0.00188106 0.44325 0.000130691 1.02 0.888521 0.534445 0.287217 1.71885e-07 3.07911e-09 2374.51 3127.64 -0.0570301 0.482191 0.277338 0.254048 -0.593214 -0.169559 0.49136 -0.266263 -0.225106 2.435 1 0 296.4 0 2.20363 2.433 0.000299369 0.861008 0.69053 0.325832 0.429165 2.20382 137.492 83.7773 18.7126 60.7973 0.00403121 0 -40 10
1.534 4.43915e-08 2.5396e-06 0.139235 0.139234 0.0120295 2.01779e-05 0.00115436 0.174043 0.000658678 0.174697 0.931788 101.571 0.237352 0.825364 4.42863 0.062648 0.0417795 0.95822 0.0195526 0.00450311 0.0188125 0.00430435 0.00544737 0.00618751 0.217895 0.2475 58.0354 -87.8983 126.203 15.9432 145.031 0.000141778 0.267273 192.763 0.310286 0.0673365 0.00409782 0.000562232 0.00138462 0.986966 0.99172 -2.98684e-06 -85.6591 0.0930662 31173.9 307.604 0.983502 0.319146 0.735471 0.735467 9.99958 2.98537e-06 1.19414e-05 0.133298 0.983316 0.931565 -0.0132919 4.92405e-06 0.511901 -1.9798e-20 7.33425e-24 -1.97907e-20 0.00139621 0.997815 8.60051e-05 0.152698 2.85259 0.00139621 0.997816 0.773089 0.00106383 0.00188106 0.000860051 0.455436 0.00188106 0.443256 0.000130694 1.02 0.888522 0.534445 0.287219 1.71886e-07 3.07913e-09 2374.49 3127.68 -0.0570347 0.482191 0.277337 0.254051 -0.593214 -0.16956 0.491345 -0.266261 -0.225093 2.436 1 0 296.396 0 2.20377 2.434 0.000299368 0.861033 0.690574 0.325782 0.429187 2.20396 137.5 83.7768 18.7126 60.7971 0.00403123 0 -40 10
1.535 4.44203e-08 2.5396e-06 0.139274 0.139273 0.0120294 2.01911e-05 0.00115436 0.174093 0.000658679 0.174747 0.931874 101.571 0.237342 0.825493 4.42916 0.0626583 0.0417845 0.958216 0.0195521 0.00450351 0.018812 0.0043047 0.00544787 0.00618802 0.217915 0.247521 58.0355 -87.8983 126.203 15.9432 145.031 0.00014178 0.267273 192.763 0.310285 0.0673365 0.00409782 0.000562233 0.00138462 0.986966 0.99172 -2.98685e-06 -85.6591 0.0930663 31173.9 307.615 0.983502 0.319146 0.735482 0.735477 9.99958 2.98538e-06 1.19414e-05 0.133302 0.983316 0.931564 -0.0132919 4.92408e-06 0.511918 -1.97994e-20 7.33482e-24 -1.97921e-20 0.00139621 0.997815 8.60052e-05 0.152698 2.85259 0.00139621 0.997816 0.773168 0.00106384 0.00188107 0.000860052 0.455436 0.00188106 0.443262 0.000130696 1.02 0.888523 0.534444 0.28722 1.71886e-07 3.07915e-09 2374.47 3127.72 -0.0570393 0.482191 0.277337 0.254054 -0.593213 -0.16956 0.49133 -0.266259 -0.225081 2.437 1 0 296.392 0 2.20391 2.435 0.000299367 0.861058 0.690618 0.325732 0.42921 2.2041 137.507 83.7763 18.7125 60.7968 0.00403125 0 -40 10
1.536 4.44492e-08 2.5396e-06 0.139314 0.139313 0.0120294 2.02042e-05 0.00115436 0.174142 0.00065868 0.174796 0.931961 101.57 0.237331 0.825621 4.42968 0.0626687 0.0417894 0.958211 0.0195516 0.00450391 0.0188115 0.00430505 0.00544837 0.00618853 0.217935 0.247541 58.0356 -87.8983 126.203 15.9432 145.031 0.000141782 0.267274 192.763 0.310285 0.0673364 0.00409783 0.000562233 0.00138462 0.986966 0.99172 -2.98687e-06 -85.6591 0.0930663 31173.9 307.626 0.983502 0.319146 0.735492 0.735488 9.99958 2.98538e-06 1.19414e-05 0.133307 0.983317 0.931564 -0.0132919 4.92411e-06 0.511936 -1.98008e-20 7.33539e-24 -1.97935e-20 0.00139621 0.997815 8.60053e-05 0.152699 2.85259 0.00139621 0.997816 0.773246 0.00106386 0.00188107 0.000860053 0.455436 0.00188107 0.443268 0.000130699 1.02 0.888524 0.534444 0.287222 1.71886e-07 3.07918e-09 2374.46 3127.77 -0.0570439 0.482191 0.277337 0.254057 -0.593213 -0.16956 0.491316 -0.266257 -0.225068 2.438 1 0 296.388 0 2.20405 2.436 0.000299366 0.861083 0.690662 0.325681 0.429233 2.20424 137.515 83.7758 18.7125 60.7966 0.00403127 0 -40 10
1.537 4.44781e-08 2.5396e-06 0.139353 0.139352 0.0120294 2.02173e-05 0.00115436 0.174191 0.00065868 0.174845 0.932047 101.57 0.237321 0.82575 4.43021 0.0626791 0.0417944 0.958206 0.0195511 0.00450432 0.018811 0.0043054 0.00544887 0.00618904 0.217955 0.247562 58.0356 -87.8983 126.202 15.9431 145.031 0.000141784 0.267274 192.762 0.310285 0.0673364 0.00409783 0.000562234 0.00138463 0.986966 0.99172 -2.98688e-06 -85.6591 0.0930664 31173.9 307.637 0.983502 0.319146 0.735503 0.735499 9.99958 2.98539e-06 1.19415e-05 0.133311 0.983318 0.931563 -0.0132919 4.92414e-06 0.511953 -1.98022e-20 7.33595e-24 -1.97949e-20 0.00139621 0.997815 8.60054e-05 0.152699 2.85259 0.00139621 0.997816 0.773325 0.00106388 0.00188107 0.000860054 0.455436 0.00188107 0.443273 0.000130701 1.02 0.888525 0.534444 0.287223 1.71886e-07 3.0792e-09 2374.44 3127.81 -0.0570485 0.482191 0.277336 0.25406 -0.593212 -0.16956 0.491301 -0.266255 -0.225055 2.439 1 0 296.383 0 2.20419 2.437 0.000299365 0.861108 0.690705 0.325631 0.429256 2.20438 137.522 83.7752 18.7125 60.7963 0.00403129 0 -40 10
1.538 4.45069e-08 2.5396e-06 0.139392 0.139391 0.0120294 2.02304e-05 0.00115436 0.17424 0.000658681 0.174894 0.932134 101.569 0.237311 0.825879 4.43073 0.0626895 0.0417993 0.958201 0.0195506 0.00450472 0.0188105 0.00430574 0.00544937 0.00618955 0.217975 0.247582 58.0357 -87.8983 126.202 15.9431 145.031 0.000141786 0.267274 192.762 0.310284 0.0673363 0.00409783 0.000562235 0.00138463 0.986966 0.99172 -2.9869e-06 -85.6591 0.0930665 31173.8 307.648 0.983502 0.319146 0.735514 0.735509 9.99958 2.98539e-06 1.19415e-05 0.133315 0.983318 0.931562 -0.0132919 4.92417e-06 0.511971 -1.98036e-20 7.33652e-24 -1.97963e-20 0.00139621 0.997815 8.60055e-05 0.152699 2.85259 0.00139621 0.997816 0.773404 0.00106389 0.00188107 0.000860055 0.455435 0.00188107 0.443279 0.000130704 1.02 0.888526 0.534443 0.287225 1.71887e-07 3.07922e-09 2374.42 3127.86 -0.0570532 0.482191 0.277336 0.254062 -0.593211 -0.16956 0.491286 -0.266253 -0.225043 2.44 1 0 296.379 0 2.20433 2.438 0.000299364 0.861133 0.690749 0.325581 0.429279 2.20452 137.53 83.7747 18.7124 60.7961 0.00403132 0 -40 10
1.539 4.45358e-08 2.5396e-06 0.139431 0.139431 0.0120294 2.02435e-05 0.00115437 0.174289 0.000658682 0.174943 0.93222 101.569 0.2373 0.826007 4.43126 0.0626998 0.0418043 0.958196 0.0195501 0.00450513 0.0188099 0.00430609 0.00544987 0.00619006 0.217995 0.247602 58.0357 -87.8983 126.202 15.9431 145.032 0.000141788 0.267274 192.762 0.310284 0.0673363 0.00409783 0.000562235 0.00138463 0.986965 0.99172 -2.98691e-06 -85.659 0.0930666 31173.8 307.659 0.983502 0.319146 0.735524 0.73552 9.99958 2.9854e-06 1.19415e-05 0.133319 0.983319 0.931561 -0.0132919 4.92419e-06 0.511988 -1.98051e-20 7.33709e-24 -1.97977e-20 0.00139621 0.997815 8.60055e-05 0.152699 2.85259 0.00139621 0.997816 0.773482 0.00106391 0.00188107 0.000860055 0.455435 0.00188107 0.443285 0.000130707 1.02 0.888527 0.534443 0.287226 1.71887e-07 3.07925e-09 2374.41 3127.9 -0.0570578 0.482191 0.277336 0.254065 -0.593211 -0.16956 0.491271 -0.266251 -0.22503 2.441 1 0 296.375 0 2.20447 2.439 0.000299363 0.861158 0.690793 0.325531 0.429301 2.20466 137.537 83.7742 18.7124 60.7958 0.00403134 0 -40 10
1.54 4.45647e-08 2.53961e-06 0.139471 0.13947 0.0120294 2.02567e-05 0.00115437 0.174338 0.000658682 0.174993 0.932307 101.568 0.23729 0.826136 4.43178 0.0627102 0.0418093 0.958191 0.0195496 0.00450553 0.0188094 0.00430644 0.00545037 0.00619057 0.218015 0.247623 58.0358 -87.8983 126.202 15.943 145.032 0.00014179 0.267274 192.762 0.310283 0.0673362 0.00409784 0.000562236 0.00138463 0.986965 0.99172 -2.98693e-06 -85.659 0.0930667 31173.8 307.67 0.983502 0.319146 0.735535 0.735531 9.99958 2.9854e-06 1.19415e-05 0.133323 0.983319 0.93156 -0.0132919 4.92422e-06 0.512006 -1.98065e-20 7.33766e-24 -1.97991e-20 0.00139621 0.997815 8.60056e-05 0.152699 2.85259 0.00139621 0.997816 0.773561 0.00106393 0.00188107 0.000860056 0.455435 0.00188107 0.443291 0.000130709 1.02 0.888528 0.534443 0.287228 1.71887e-07 3.07927e-09 2374.39 3127.95 -0.0570624 0.482192 0.277336 0.254068 -0.59321 -0.16956 0.491257 -0.266249 -0.225017 2.442 1 0 296.371 0 2.20461 2.44 0.000299362 0.861183 0.690837 0.325482 0.429324 2.2048 137.545 83.7737 18.7124 60.7955 0.00403136 0 -40 10
1.541 4.45935e-08 2.53961e-06 0.13951 0.139509 0.0120294 2.02698e-05 0.00115437 0.174387 0.000658683 0.175042 0.932393 101.568 0.237279 0.826265 4.43231 0.0627206 0.0418142 0.958186 0.0195491 0.00450594 0.0188089 0.00430679 0.00545086 0.00619108 0.218035 0.247643 58.0359 -87.8983 126.202 15.943 145.032 0.000141792 0.267275 192.762 0.310283 0.0673362 0.00409784 0.000562237 0.00138463 0.986965 0.99172 -2.98694e-06 -85.659 0.0930668 31173.8 307.681 0.983502 0.319146 0.735546 0.735541 9.99958 2.98541e-06 1.19415e-05 0.133327 0.98332 0.931559 -0.0132919 4.92425e-06 0.512023 -1.98079e-20 7.33823e-24 -1.98006e-20 0.00139621 0.997815 8.60057e-05 0.152699 2.85259 0.00139621 0.997816 0.77364 0.00106394 0.00188107 0.000860057 0.455435 0.00188107 0.443296 0.000130712 1.02 0.88853 0.534443 0.287229 1.71887e-07 3.07929e-09 2374.38 3127.99 -0.057067 0.482192 0.277335 0.254071 -0.59321 -0.16956 0.491242 -0.266246 -0.225005 2.443 1 0 296.367 0 2.20475 2.441 0.000299361 0.861208 0.690881 0.325432 0.429347 2.20494 137.552 83.7731 18.7124 60.7953 0.00403138 0 -40 10
1.542 4.46224e-08 2.53961e-06 0.139549 0.139548 0.0120293 2.02829e-05 0.00115437 0.174436 0.000658684 0.175091 0.93248 101.567 0.237269 0.826393 4.43284 0.062731 0.0418192 0.958181 0.0195486 0.00450635 0.0188084 0.00430714 0.00545136 0.00619159 0.218055 0.247664 58.0359 -87.8984 126.201 15.9429 145.032 0.000141794 0.267275 192.762 0.310282 0.0673361 0.00409784 0.000562237 0.00138464 0.986965 0.99172 -2.98696e-06 -85.659 0.0930669 31173.8 307.692 0.983502 0.319146 0.735556 0.735552 9.99958 2.98541e-06 1.19416e-05 0.133331 0.98332 0.931559 -0.0132919 4.92428e-06 0.512041 -1.98093e-20 7.3388e-24 -1.9802e-20 0.00139621 0.997815 8.60058e-05 0.152699 2.85259 0.00139621 0.997816 0.773718 0.00106396 0.00188108 0.000860058 0.455434 0.00188107 0.443302 0.000130714 1.02 0.888531 0.534442 0.287231 1.71888e-07 3.07931e-09 2374.36 3128.04 -0.0570717 0.482192 0.277335 0.254074 -0.593209 -0.16956 0.491227 -0.266244 -0.224992 2.444 1 0 296.363 0 2.20489 2.442 0.00029936 0.861233 0.690924 0.325382 0.42937 2.20508 137.56 83.7726 18.7123 60.795 0.0040314 0 -40 10
1.543 4.46513e-08 2.53961e-06 0.139588 0.139588 0.0120293 2.0296e-05 0.00115437 0.174485 0.000658685 0.17514 0.932566 101.567 0.237259 0.826522 4.43337 0.0627414 0.0418242 0.958176 0.0195481 0.00450675 0.0188079 0.00430749 0.00545187 0.0061921 0.218075 0.247684 58.036 -87.8984 126.201 15.9429 145.032 0.000141796 0.267275 192.762 0.310282 0.0673361 0.00409785 0.000562238 0.00138464 0.986965 0.99172 -2.98697e-06 -85.659 0.093067 31173.7 307.703 0.983502 0.319146 0.735567 0.735562 9.99958 2.98542e-06 1.19416e-05 0.133335 0.983321 0.931558 -0.0132919 4.92431e-06 0.512058 -1.98107e-20 7.33937e-24 -1.98034e-20 0.00139622 0.997815 8.60059e-05 0.1527 2.85259 0.00139622 0.997816 0.773797 0.00106398 0.00188108 0.000860059 0.455434 0.00188108 0.443308 0.000130717 1.02 0.888532 0.534442 0.287232 1.71888e-07 3.07934e-09 2374.34 3128.08 -0.0570763 0.482192 0.277335 0.254077 -0.593209 -0.16956 0.491212 -0.266242 -0.224979 2.445 1 0 296.358 0 2.20503 2.443 0.000299359 0.861258 0.690968 0.325332 0.429392 2.20522 137.567 83.7721 18.7123 60.7948 0.00403142 0 -40 10
1.544 4.46801e-08 2.53961e-06 0.139627 0.139627 0.0120293 2.03091e-05 0.00115437 0.174534 0.000658685 0.175188 0.932653 101.566 0.237248 0.826651 4.43389 0.0627518 0.0418292 0.958171 0.0195476 0.00450716 0.0188074 0.00430783 0.00545237 0.00619261 0.218095 0.247705 58.0361 -87.8984 126.201 15.9429 145.032 0.000141798 0.267275 192.761 0.310282 0.067336 0.00409785 0.000562239 0.00138464 0.986965 0.99172 -2.98699e-06 -85.659 0.093067 31173.7 307.714 0.983502 0.319146 0.735578 0.735573 9.99958 2.98542e-06 1.19416e-05 0.13334 0.983322 0.931557 -0.0132919 4.92434e-06 0.512076 -1.98121e-20 7.33994e-24 -1.98048e-20 0.00139622 0.997815 8.60059e-05 0.1527 2.8526 0.00139622 0.997816 0.773875 0.00106399 0.00188108 0.000860059 0.455434 0.00188108 0.443314 0.000130719 1.02 0.888533 0.534442 0.287234 1.71888e-07 3.07936e-09 2374.33 3128.12 -0.0570809 0.482192 0.277334 0.25408 -0.593208 -0.16956 0.491197 -0.26624 -0.224967 2.446 1 0 296.354 0 2.20517 2.444 0.000299358 0.861284 0.691012 0.325283 0.429415 2.20536 137.575 83.7716 18.7123 60.7945 0.00403145 0 -40 10
1.545 4.4709e-08 2.53961e-06 0.139667 0.139666 0.0120293 2.03223e-05 0.00115437 0.174583 0.000658686 0.175237 0.932739 101.566 0.237238 0.82678 4.43442 0.0627622 0.0418342 0.958166 0.0195471 0.00450757 0.0188069 0.00430818 0.00545287 0.00619313 0.218115 0.247725 58.0361 -87.8984 126.201 15.9428 145.032 0.0001418 0.267275 192.761 0.310281 0.0673359 0.00409785 0.000562239 0.00138464 0.986965 0.99172 -2.987e-06 -85.659 0.0930671 31173.7 307.725 0.983502 0.319146 0.735588 0.735584 9.99958 2.98543e-06 1.19416e-05 0.133344 0.983322 0.931556 -0.0132919 4.92437e-06 0.512093 -1.98136e-20 7.34051e-24 -1.98062e-20 0.00139622 0.997815 8.6006e-05 0.1527 2.8526 0.00139622 0.997816 0.773954 0.00106401 0.00188108 0.00086006 0.455434 0.00188108 0.44332 0.000130722 1.02 0.888534 0.534441 0.287236 1.71889e-07 3.07938e-09 2374.31 3128.17 -0.0570856 0.482192 0.277334 0.254082 -0.593207 -0.16956 0.491183 -0.266238 -0.224954 2.447 1 0 296.35 0 2.20531 2.445 0.000299357 0.861309 0.691056 0.325233 0.429438 2.2055 137.582 83.771 18.7122 60.7943 0.00403147 0 -40 10
1.546 4.47378e-08 2.53961e-06 0.139706 0.139705 0.0120293 2.03354e-05 0.00115437 0.174632 0.000658687 0.175286 0.932826 101.565 0.237227 0.826909 4.43495 0.0627725 0.0418392 0.958161 0.0195466 0.00450797 0.0188064 0.00430853 0.00545337 0.00619364 0.218135 0.247746 58.0362 -87.8984 126.201 15.9428 145.032 0.000141802 0.267276 192.761 0.310281 0.0673359 0.00409786 0.00056224 0.00138464 0.986965 0.99172 -2.98702e-06 -85.659 0.0930672 31173.7 307.736 0.983502 0.319146 0.735599 0.735594 9.99958 2.98543e-06 1.19416e-05 0.133348 0.983323 0.931555 -0.0132919 4.9244e-06 0.512111 -1.9815e-20 7.34108e-24 -1.98076e-20 0.00139622 0.997815 8.60061e-05 0.1527 2.8526 0.00139622 0.997816 0.774032 0.00106403 0.00188108 0.000860061 0.455434 0.00188108 0.443325 0.000130725 1.02 0.888535 0.534441 0.287237 1.71889e-07 3.07941e-09 2374.29 3128.21 -0.0570902 0.482192 0.277334 0.254085 -0.593207 -0.16956 0.491168 -0.266236 -0.224941 2.448 1 0 296.346 0 2.20545 2.446 0.000299356 0.861334 0.691099 0.325183 0.429461 2.20564 137.59 83.7705 18.7122 60.794 0.00403149 0 -40 10
1.547 4.47667e-08 2.53961e-06 0.139745 0.139744 0.0120293 2.03485e-05 0.00115437 0.174681 0.000658687 0.175335 0.932913 101.565 0.237217 0.827037 4.43548 0.0627829 0.0418442 0.958156 0.0195461 0.00450838 0.0188058 0.00430888 0.00545387 0.00619415 0.218155 0.247766 58.0362 -87.8984 126.2 15.9428 145.032 0.000141804 0.267276 192.761 0.31028 0.0673358 0.00409786 0.000562241 0.00138465 0.986965 0.99172 -2.98703e-06 -85.659 0.0930673 31173.6 307.747 0.983502 0.319146 0.73561 0.735605 9.99958 2.98544e-06 1.19417e-05 0.133352 0.983323 0.931555 -0.0132919 4.92443e-06 0.512129 -1.98164e-20 7.34165e-24 -1.98091e-20 0.00139622 0.997815 8.60062e-05 0.1527 2.8526 0.00139622 0.997816 0.774111 0.00106405 0.00188108 0.000860062 0.455433 0.00188108 0.443331 0.000130727 1.02 0.888536 0.534441 0.287239 1.71889e-07 3.07943e-09 2374.28 3128.26 -0.0570948 0.482192 0.277334 0.254088 -0.593206 -0.16956 0.491153 -0.266234 -0.224928 2.449 1 0 296.342 0 2.20559 2.447 0.000299355 0.861359 0.691143 0.325134 0.429484 2.20578 137.597 83.77 18.7122 60.7938 0.00403151 0 -40 10
1.548 4.47956e-08 2.53962e-06 0.139784 0.139783 0.0120293 2.03616e-05 0.00115437 0.17473 0.000658688 0.175384 0.932999 101.564 0.237207 0.827166 4.43601 0.0627933 0.0418492 0.958151 0.0195456 0.00450879 0.0188053 0.00430923 0.00545437 0.00619467 0.218175 0.247787 58.0363 -87.8984 126.2 15.9427 145.032 0.000141806 0.267276 192.761 0.31028 0.0673358 0.00409786 0.000562241 0.00138465 0.986965 0.99172 -2.98705e-06 -85.659 0.0930674 31173.6 307.758 0.983502 0.319146 0.73562 0.735616 9.99958 2.98544e-06 1.19417e-05 0.133356 0.983324 0.931554 -0.0132919 4.92446e-06 0.512146 -1.98178e-20 7.34222e-24 -1.98105e-20 0.00139622 0.997815 8.60063e-05 0.1527 2.8526 0.00139622 0.997816 0.774189 0.00106406 0.00188109 0.000860063 0.455433 0.00188108 0.443337 0.00013073 1.02 0.888537 0.53444 0.28724 1.71889e-07 3.07945e-09 2374.26 3128.3 -0.0570995 0.482192 0.277333 0.254091 -0.593206 -0.16956 0.491138 -0.266232 -0.224916 2.45 1 0 296.338 0 2.20573 2.448 0.000299353 0.861385 0.691187 0.325084 0.429506 2.20592 137.605 83.7695 18.7121 60.7935 0.00403153 0 -40 10
1.549 4.48244e-08 2.53962e-06 0.139823 0.139822 0.0120293 2.03747e-05 0.00115437 0.174778 0.000658689 0.175432 0.933086 101.563 0.237196 0.827295 4.43654 0.0628037 0.0418542 0.958146 0.0195451 0.00450919 0.0188048 0.00430958 0.00545487 0.00619518 0.218195 0.247807 58.0364 -87.8984 126.2 15.9427 145.032 0.000141808 0.267276 192.761 0.310279 0.0673357 0.00409786 0.000562242 0.00138465 0.986965 0.99172 -2.98706e-06 -85.6589 0.0930675 31173.6 307.769 0.983502 0.319146 0.735631 0.735627 9.99958 2.98545e-06 1.19417e-05 0.13336 0.983324 0.931553 -0.0132919 4.92449e-06 0.512164 -1.98192e-20 7.3428e-24 -1.98119e-20 0.00139622 0.997815 8.60063e-05 0.152701 2.8526 0.00139622 0.997816 0.774267 0.00106408 0.00188109 0.000860063 0.455433 0.00188109 0.443343 0.000130732 1.02 0.888538 0.53444 0.287242 1.7189e-07 3.07948e-09 2374.24 3128.35 -0.0571041 0.482192 0.277333 0.254094 -0.593205 -0.16956 0.491123 -0.26623 -0.224903 2.451 1 0 296.333 0 2.20587 2.449 0.000299352 0.86141 0.691231 0.325035 0.429529 2.20606 137.612 83.7689 18.7121 60.7933 0.00403156 0 -40 10
1.55 4.48533e-08 2.53962e-06 0.139862 0.139861 0.0120292 2.03879e-05 0.00115437 0.174827 0.000658689 0.175481 0.933173 101.563 0.237186 0.827424 4.43707 0.0628141 0.0418592 0.958141 0.0195446 0.0045096 0.0188043 0.00430993 0.00545538 0.00619569 0.218215 0.247828 58.0364 -87.8984 126.2 15.9426 145.032 0.00014181 0.267276 192.76 0.310279 0.0673357 0.00409787 0.000562243 0.00138465 0.986965 0.99172 -2.98708e-06 -85.6589 0.0930676 31173.6 307.78 0.983502 0.319146 0.735642 0.735637 9.99958 2.98545e-06 1.19417e-05 0.133365 0.983325 0.931552 -0.0132919 4.92452e-06 0.512181 -1.98207e-20 7.34337e-24 -1.98133e-20 0.00139622 0.997815 8.60064e-05 0.152701 2.8526 0.00139622 0.997816 0.774346 0.0010641 0.00188109 0.000860064 0.455433 0.00188109 0.443348 0.000130735 1.02 0.888539 0.53444 0.287243 1.7189e-07 3.0795e-09 2374.23 3128.39 -0.0571088 0.482192 0.277333 0.254097 -0.593205 -0.169561 0.491108 -0.266228 -0.22489 2.452 1 0 296.329 0 2.20601 2.45 0.000299351 0.861435 0.691274 0.324986 0.429552 2.20619 137.62 83.7684 18.7121 60.793 0.00403158 0 -40 10
1.551 4.48822e-08 2.53962e-06 0.139901 0.1399 0.0120292 2.0401e-05 0.00115437 0.174876 0.00065869 0.17553 0.933259 101.562 0.237175 0.827553 4.4376 0.0628245 0.0418642 0.958136 0.0195441 0.00451001 0.0188038 0.00431028 0.00545588 0.00619621 0.218235 0.247848 58.0365 -87.8984 126.2 15.9426 145.032 0.000141813 0.267277 192.76 0.310279 0.0673356 0.00409787 0.000562243 0.00138466 0.986965 0.99172 -2.98709e-06 -85.6589 0.0930677 31173.6 307.791 0.983502 0.319146 0.735652 0.735648 9.99958 2.98546e-06 1.19417e-05 0.133369 0.983326 0.931551 -0.0132919 4.92455e-06 0.512199 -1.98221e-20 7.34394e-24 -1.98147e-20 0.00139623 0.997815 8.60065e-05 0.152701 2.8526 0.00139622 0.997816 0.774424 0.00106411 0.00188109 0.000860065 0.455432 0.00188109 0.443354 0.000130737 1.02 0.888541 0.534439 0.287245 1.7189e-07 3.07952e-09 2374.21 3128.44 -0.0571134 0.482192 0.277332 0.2541 -0.593204 -0.169561 0.491093 -0.266225 -0.224877 2.453 1 0 296.325 0 2.20615 2.451 0.00029935 0.861461 0.691318 0.324936 0.429575 2.20633 137.627 83.7679 18.7121 60.7928 0.0040316 0 -40 10
1.552 4.4911e-08 2.53962e-06 0.139939 0.139939 0.0120292 2.04141e-05 0.00115437 0.174924 0.000658691 0.175578 0.933346 101.562 0.237165 0.827682 4.43814 0.0628349 0.0418692 0.958131 0.0195436 0.00451042 0.0188033 0.00431063 0.00545638 0.00619672 0.218255 0.247869 58.0366 -87.8984 126.199 15.9426 145.032 0.000141815 0.267277 192.76 0.310278 0.0673356 0.00409787 0.000562244 0.00138466 0.986965 0.99172 -2.98711e-06 -85.6589 0.0930677 31173.5 307.802 0.983502 0.319146 0.735663 0.735659 9.99958 2.98546e-06 1.19417e-05 0.133373 0.983326 0.93155 -0.0132919 4.92458e-06 0.512217 -1.98235e-20 7.34451e-24 -1.98162e-20 0.00139623 0.997815 8.60066e-05 0.152701 2.8526 0.00139623 0.997816 0.774502 0.00106413 0.00188109 0.000860066 0.455432 0.00188109 0.44336 0.00013074 1.02 0.888542 0.534439 0.287246 1.7189e-07 3.07954e-09 2374.19 3128.48 -0.0571181 0.482192 0.277332 0.254103 -0.593203 -0.169561 0.491079 -0.266223 -0.224865 2.454 1 0 296.321 0 2.20629 2.452 0.000299349 0.861486 0.691362 0.324887 0.429597 2.20647 137.635 83.7673 18.712 60.7925 0.00403162 0 -40 10
1.553 4.49399e-08 2.53962e-06 0.139978 0.139978 0.0120292 2.04272e-05 0.00115437 0.174973 0.000658691 0.175627 0.933433 101.561 0.237155 0.827811 4.43867 0.0628453 0.0418742 0.958126 0.0195431 0.00451083 0.0188028 0.00431098 0.00545688 0.00619724 0.218275 0.247889 58.0366 -87.8984 126.199 15.9425 145.032 0.000141817 0.267277 192.76 0.310278 0.0673355 0.00409788 0.000562245 0.00138466 0.986965 0.991719 -2.98712e-06 -85.6589 0.0930678 31173.5 307.813 0.983502 0.319146 0.735674 0.735669 9.99958 2.98547e-06 1.19418e-05 0.133377 0.983327 0.93155 -0.0132919 4.92461e-06 0.512234 -1.98249e-20 7.34508e-24 -1.98176e-20 0.00139623 0.997815 8.60067e-05 0.152701 2.8526 0.00139623 0.997816 0.774581 0.00106415 0.00188109 0.000860067 0.455432 0.00188109 0.443366 0.000130743 1.02 0.888543 0.534439 0.287248 1.71891e-07 3.07957e-09 2374.18 3128.53 -0.0571227 0.482193 0.277332 0.254106 -0.593203 -0.169561 0.491064 -0.266221 -0.224852 2.455 1 0 296.317 0 2.20643 2.453 0.000299348 0.861511 0.691406 0.324838 0.42962 2.20661 137.642 83.7668 18.712 60.7922 0.00403164 0 -40 10
1.554 4.49688e-08 2.53962e-06 0.140017 0.140016 0.0120292 2.04403e-05 0.00115437 0.175021 0.000658692 0.175675 0.933519 101.561 0.237144 0.82794 4.4392 0.0628558 0.0418793 0.958121 0.0195426 0.00451124 0.0188022 0.00431134 0.00545739 0.00619775 0.218296 0.24791 58.0367 -87.8984 126.199 15.9425 145.032 0.000141819 0.267277 192.76 0.310277 0.0673355 0.00409788 0.000562245 0.00138466 0.986965 0.991719 -2.98714e-06 -85.6589 0.0930679 31173.5 307.825 0.983502 0.319146 0.735685 0.73568 9.99958 2.98547e-06 1.19418e-05 0.133381 0.983327 0.931549 -0.0132919 4.92464e-06 0.512252 -1.98264e-20 7.34566e-24 -1.9819e-20 0.00139623 0.997815 8.60067e-05 0.152701 2.8526 0.00139623 0.997816 0.774659 0.00106416 0.00188109 0.000860067 0.455432 0.00188109 0.443371 0.000130745 1.02 0.888544 0.534439 0.287249 1.71891e-07 3.07959e-09 2374.16 3128.57 -0.0571274 0.482193 0.277332 0.254108 -0.593202 -0.169561 0.491049 -0.266219 -0.224839 2.456 1 0 296.313 0 2.20657 2.454 0.000299347 0.861537 0.691449 0.324789 0.429643 2.20675 137.65 83.7663 18.712 60.792 0.00403166 0 -40 10
1.555 4.49976e-08 2.53963e-06 0.140056 0.140055 0.0120292 2.04535e-05 0.00115438 0.17507 0.000658693 0.175724 0.933606 101.56 0.237134 0.828069 4.43974 0.0628662 0.0418843 0.958116 0.0195421 0.00451165 0.0188017 0.00431169 0.00545789 0.00619827 0.218316 0.247931 58.0367 -87.8984 126.199 15.9425 145.032 0.000141821 0.267277 192.76 0.310277 0.0673354 0.00409788 0.000562246 0.00138466 0.986965 0.991719 -2.98715e-06 -85.6589 0.093068 31173.5 307.836 0.983502 0.319146 0.735695 0.735691 9.99958 2.98548e-06 1.19418e-05 0.133385 0.983328 0.931548 -0.0132919 4.92467e-06 0.512269 -1.98278e-20 7.34623e-24 -1.98204e-20 0.00139623 0.997815 8.60068e-05 0.152701 2.85261 0.00139623 0.997816 0.774737 0.00106418 0.0018811 0.000860068 0.455432 0.00188109 0.443377 0.000130748 1.02 0.888545 0.534438 0.287251 1.71891e-07 3.07961e-09 2374.14 3128.62 -0.057132 0.482193 0.277331 0.254111 -0.593202 -0.169561 0.491034 -0.266217 -0.224826 2.457 1 0 296.308 0 2.20671 2.455 0.000299346 0.861562 0.691493 0.32474 0.429666 2.20689 137.657 83.7657 18.7119 60.7917 0.00403169 0 -40 10
1.556 4.50265e-08 2.53963e-06 0.140095 0.140094 0.0120292 2.04666e-05 0.00115438 0.175118 0.000658693 0.175772 0.933693 101.56 0.237123 0.828198 4.44027 0.0628766 0.0418893 0.958111 0.0195416 0.00451205 0.0188012 0.00431204 0.0054584 0.00619878 0.218336 0.247951 58.0368 -87.8984 126.199 15.9424 145.032 0.000141823 0.267278 192.759 0.310276 0.0673354 0.00409789 0.000562247 0.00138467 0.986965 0.991719 -2.98717e-06 -85.6589 0.0930681 31173.4 307.847 0.983502 0.319146 0.735706 0.735702 9.99958 2.98548e-06 1.19418e-05 0.13339 0.983328 0.931547 -0.0132919 4.9247e-06 0.512287 -1.98292e-20 7.34681e-24 -1.98219e-20 0.00139623 0.997815 8.60069e-05 0.152702 2.85261 0.00139623 0.997816 0.774815 0.0010642 0.0018811 0.000860069 0.455431 0.0018811 0.443383 0.00013075 1.02 0.888546 0.534438 0.287252 1.71892e-07 3.07964e-09 2374.13 3128.66 -0.0571367 0.482193 0.277331 0.254114 -0.593201 -0.169561 0.491019 -0.266215 -0.224814 2.458 1 0 296.304 0 2.20685 2.456 0.000299345 0.861588 0.691537 0.324691 0.429688 2.20703 137.665 83.7652 18.7119 60.7915 0.00403171 0 -40 10
1.557 4.50553e-08 2.53963e-06 0.140133 0.140133 0.0120291 2.04797e-05 0.00115438 0.175167 0.000658694 0.175821 0.93378 101.559 0.237113 0.828327 4.4408 0.062887 0.0418944 0.958106 0.0195411 0.00451246 0.0188007 0.00431239 0.0054589 0.0061993 0.218356 0.247972 58.0369 -87.8984 126.198 15.9424 145.032 0.000141825 0.267278 192.759 0.310276 0.0673353 0.00409789 0.000562247 0.00138467 0.986965 0.991719 -2.98718e-06 -85.6589 0.0930682 31173.4 307.858 0.983502 0.319146 0.735717 0.735712 9.99958 2.98549e-06 1.19418e-05 0.133394 0.983329 0.931546 -0.0132919 4.92473e-06 0.512305 -1.98306e-20 7.34738e-24 -1.98233e-20 0.00139623 0.997815 8.6007e-05 0.152702 2.85261 0.00139623 0.997816 0.774893 0.00106421 0.0018811 0.00086007 0.455431 0.0018811 0.443389 0.000130753 1.02 0.888547 0.534438 0.287254 1.71892e-07 3.07966e-09 2374.11 3128.71 -0.0571414 0.482193 0.277331 0.254117 -0.593201 -0.169561 0.491004 -0.266213 -0.224801 2.459 1 0 296.3 0 2.20699 2.457 0.000299344 0.861613 0.69158 0.324642 0.429711 2.20717 137.672 83.7647 18.7119 60.7912 0.00403173 0 -40 10
1.558 4.50842e-08 2.53963e-06 0.140172 0.140171 0.0120291 2.04928e-05 0.00115438 0.175215 0.000658695 0.175869 0.933867 101.559 0.237103 0.828456 4.44134 0.0628974 0.0418994 0.958101 0.0195406 0.00451287 0.0188002 0.00431274 0.00545941 0.00619982 0.218376 0.247993 58.0369 -87.8984 126.198 15.9423 145.032 0.000141827 0.267278 192.759 0.310276 0.0673353 0.00409789 0.000562248 0.00138467 0.986965 0.991719 -2.9872e-06 -85.6589 0.0930683 31173.4 307.869 0.983501 0.319146 0.735728 0.735723 9.99958 2.98549e-06 1.19419e-05 0.133398 0.983329 0.931545 -0.0132919 4.92476e-06 0.512322 -1.98321e-20 7.34795e-24 -1.98247e-20 0.00139623 0.997815 8.60071e-05 0.152702 2.85261 0.00139623 0.997816 0.774972 0.00106423 0.0018811 0.000860071 0.455431 0.0018811 0.443394 0.000130755 1.02 0.888548 0.534437 0.287255 1.71892e-07 3.07968e-09 2374.1 3128.75 -0.057146 0.482193 0.27733 0.25412 -0.5932 -0.169561 0.490989 -0.266211 -0.224788 2.46 1 0 296.296 0 2.20713 2.458 0.000299343 0.861638 0.691624 0.324593 0.429734 2.20731 137.68 83.7642 18.7118 60.791 0.00403175 0 -40 10
1.559 4.51131e-08 2.53963e-06 0.140211 0.14021 0.0120291 2.05059e-05 0.00115438 0.175263 0.000658696 0.175918 0.933954 101.558 0.237092 0.828585 4.44187 0.0629078 0.0419045 0.958096 0.0195401 0.00451328 0.0187997 0.00431309 0.00545991 0.00620033 0.218396 0.248013 58.037 -87.8984 126.198 15.9423 145.032 0.000141829 0.267278 192.759 0.310275 0.0673352 0.0040979 0.000562249 0.00138467 0.986965 0.991719 -2.98721e-06 -85.6589 0.0930684 31173.4 307.88 0.983501 0.319146 0.735738 0.735734 9.99958 2.9855e-06 1.19419e-05 0.133402 0.98333 0.931544 -0.0132919 4.92479e-06 0.51234 -1.98335e-20 7.34853e-24 -1.98261e-20 0.00139623 0.997815 8.60071e-05 0.152702 2.85261 0.00139623 0.997816 0.77505 0.00106425 0.0018811 0.000860071 0.455431 0.0018811 0.4434 0.000130758 1.02 0.888549 0.534437 0.287257 1.71892e-07 3.0797e-09 2374.08 3128.8 -0.0571507 0.482193 0.27733 0.254123 -0.593199 -0.169561 0.490974 -0.266209 -0.224775 2.461 1 0 296.292 0 2.20727 2.459 0.000299342 0.861664 0.691668 0.324544 0.429757 2.20745 137.687 83.7636 18.7118 60.7907 0.00403177 0 -40 10
1.56 4.51419e-08 2.53963e-06 0.140249 0.140249 0.0120291 2.05191e-05 0.00115438 0.175312 0.000658696 0.175966 0.93404 101.558 0.237082 0.828714 4.44241 0.0629182 0.0419095 0.95809 0.0195396 0.00451369 0.0187992 0.00431345 0.00546042 0.00620085 0.218417 0.248034 58.0371 -87.8984 126.198 15.9423 145.032 0.000141831 0.267278 192.759 0.310275 0.0673352 0.0040979 0.000562249 0.00138468 0.986965 0.991719 -2.98723e-06 -85.6588 0.0930684 31173.4 307.891 0.983501 0.319146 0.735749 0.735745 9.99958 2.9855e-06 1.19419e-05 0.133406 0.98333 0.931544 -0.0132919 4.92482e-06 0.512358 -1.98349e-20 7.3491e-24 -1.98276e-20 0.00139624 0.997815 8.60072e-05 0.152702 2.85261 0.00139624 0.997816 0.775128 0.00106427 0.0018811 0.000860072 0.45543 0.0018811 0.443406 0.000130761 1.02 0.88855 0.534437 0.287258 1.71893e-07 3.07973e-09 2374.06 3128.84 -0.0571554 0.482193 0.27733 0.254126 -0.593199 -0.169561 0.490959 -0.266206 -0.224762 2.462 1 0 296.287 0 2.2074 2.46 0.000299341 0.861689 0.691711 0.324495 0.429779 2.20759 137.695 83.7631 18.7118 60.7905 0.0040318 0 -40 10
1.561 4.51708e-08 2.53963e-06 0.140288 0.140287 0.0120291 2.05322e-05 0.00115438 0.17536 0.000658697 0.176014 0.934127 101.557 0.237071 0.828843 4.44294 0.0629287 0.0419146 0.958085 0.0195391 0.00451411 0.0187986 0.0043138 0.00546092 0.00620137 0.218437 0.248055 58.0371 -87.8984 126.198 15.9422 145.032 0.000141833 0.267278 192.759 0.310274 0.0673351 0.0040979 0.00056225 0.00138468 0.986965 0.991719 -2.98724e-06 -85.6588 0.0930685 31173.3 307.902 0.983501 0.319146 0.73576 0.735756 9.99958 2.98551e-06 1.19419e-05 0.13341 0.983331 0.931543 -0.0132919 4.92485e-06 0.512376 -1.98364e-20 7.34968e-24 -1.9829e-20 0.00139624 0.997815 8.60073e-05 0.152702 2.85261 0.00139624 0.997816 0.775206 0.00106428 0.0018811 0.000860073 0.45543 0.0018811 0.443412 0.000130763 1.02 0.888551 0.534436 0.28726 1.71893e-07 3.07975e-09 2374.05 3128.89 -0.0571601 0.482193 0.27733 0.254129 -0.593198 -0.169561 0.490944 -0.266204 -0.224749 2.463 1 0 296.283 0 2.20754 2.461 0.00029934 0.861715 0.691755 0.324446 0.429802 2.20773 137.702 83.7626 18.7117 60.7902 0.00403182 0 -40 10
1.562 4.51997e-08 2.53964e-06 0.140327 0.140326 0.0120291 2.05453e-05 0.00115438 0.175408 0.000658698 0.176062 0.934214 101.557 0.237061 0.828973 4.44348 0.0629391 0.0419196 0.95808 0.0195386 0.00451452 0.0187981 0.00431415 0.00546143 0.00620188 0.218457 0.248075 58.0372 -87.8984 126.198 15.9422 145.032 0.000141835 0.267279 192.758 0.310274 0.0673351 0.0040979 0.000562251 0.00138468 0.986965 0.991719 -2.98726e-06 -85.6588 0.0930686 31173.3 307.914 0.983501 0.319146 0.735771 0.735766 9.99958 2.98551e-06 1.19419e-05 0.133415 0.983331 0.931542 -0.0132919 4.92488e-06 0.512393 -1.98378e-20 7.35025e-24 -1.98304e-20 0.00139624 0.997815 8.60074e-05 0.152703 2.85261 0.00139624 0.997816 0.775284 0.0010643 0.00188111 0.000860074 0.45543 0.0018811 0.443417 0.000130766 1.02 0.888553 0.534436 0.287261 1.71893e-07 3.07977e-09 2374.03 3128.93 -0.0571647 0.482193 0.277329 0.254132 -0.593198 -0.169561 0.49093 -0.266202 -0.224737 2.464 1 0 296.279 0 2.20768 2.462 0.000299339 0.861741 0.691799 0.324398 0.429825 2.20787 137.71 83.762 18.7117 60.7899 0.00403184 0 -40 10
1.563 4.52285e-08 2.53964e-06 0.140365 0.140364 0.0120291 2.05584e-05 0.00115438 0.175456 0.000658698 0.17611 0.934301 101.556 0.23705 0.829102 4.44402 0.0629495 0.0419247 0.958075 0.0195381 0.00451493 0.0187976 0.0043145 0.00546193 0.0062024 0.218477 0.248096 58.0372 -87.8984 126.197 15.9422 145.032 0.000141837 0.267279 192.758 0.310273 0.067335 0.00409791 0.000562251 0.00138468 0.986965 0.991719 -2.98727e-06 -85.6588 0.0930687 31173.3 307.925 0.983501 0.319146 0.735782 0.735777 9.99958 2.98552e-06 1.1942e-05 0.133419 0.983332 0.931541 -0.0132919 4.92491e-06 0.512411 -1.98392e-20 7.35083e-24 -1.98319e-20 0.00139624 0.997815 8.60075e-05 0.152703 2.85261 0.00139624 0.997816 0.775362 0.00106432 0.00188111 0.000860075 0.45543 0.00188111 0.443423 0.000130768 1.02 0.888554 0.534436 0.287263 1.71893e-07 3.0798e-09 2374.01 3128.98 -0.0571694 0.482193 0.277329 0.254135 -0.593197 -0.169561 0.490915 -0.2662 -0.224724 2.465 1 0 296.275 0 2.20782 2.463 0.000299338 0.861766 0.691842 0.324349 0.429847 2.20801 137.717 83.7615 18.7117 60.7897 0.00403186 0 -40 10
1.564 4.52574e-08 2.53964e-06 0.140404 0.140403 0.012029 2.05715e-05 0.00115438 0.175505 0.000658699 0.176159 0.934388 101.555 0.23704 0.829231 4.44456 0.0629599 0.0419298 0.95807 0.0195376 0.00451534 0.0187971 0.00431486 0.00546244 0.00620292 0.218498 0.248117 58.0373 -87.8984 126.197 15.9421 145.032 0.00014184 0.267279 192.758 0.310273 0.0673349 0.00409791 0.000562252 0.00138468 0.986965 0.991719 -2.98729e-06 -85.6588 0.0930688 31173.3 307.936 0.983501 0.319146 0.735792 0.735788 9.99958 2.98552e-06 1.1942e-05 0.133423 0.983333 0.93154 -0.0132919 4.92494e-06 0.512429 -1.98407e-20 7.35141e-24 -1.98333e-20 0.00139624 0.997815 8.60076e-05 0.152703 2.85261 0.00139624 0.997816 0.77544 0.00106433 0.00188111 0.000860076 0.45543 0.00188111 0.443429 0.000130771 1.02 0.888555 0.534435 0.287264 1.71894e-07 3.07982e-09 2374 3129.02 -0.0571741 0.482193 0.277329 0.254137 -0.593197 -0.169561 0.4909 -0.266198 -0.224711 2.466 1 0 296.271 0 2.20796 2.464 0.000299337 0.861792 0.691886 0.3243 0.42987 2.20815 137.725 83.761 18.7116 60.7894 0.00403188 0 -40 10
1.565 4.52862e-08 2.53964e-06 0.140442 0.140441 0.012029 2.05847e-05 0.00115438 0.175553 0.0006587 0.176207 0.934475 101.555 0.23703 0.82936 4.44509 0.0629704 0.0419348 0.958065 0.0195371 0.00451575 0.0187966 0.00431521 0.00546295 0.00620344 0.218518 0.248138 58.0374 -87.8984 126.197 15.9421 145.032 0.000141842 0.267279 192.758 0.310273 0.0673349 0.00409791 0.000562253 0.00138469 0.986965 0.991719 -2.9873e-06 -85.6588 0.0930689 31173.2 307.947 0.983501 0.319146 0.735803 0.735799 9.99958 2.98553e-06 1.1942e-05 0.133427 0.983333 0.931539 -0.0132919 4.92497e-06 0.512447 -1.98421e-20 7.35198e-24 -1.98347e-20 0.00139624 0.997815 8.60076e-05 0.152703 2.85261 0.00139624 0.997816 0.775518 0.00106435 0.00188111 0.000860076 0.455429 0.00188111 0.443434 0.000130773 1.02 0.888556 0.534435 0.287266 1.71894e-07 3.07984e-09 2373.98 3129.07 -0.0571788 0.482193 0.277329 0.25414 -0.593196 -0.169561 0.490885 -0.266196 -0.224698 2.467 1 0 296.266 0 2.2081 2.465 0.000299336 0.861817 0.69193 0.324252 0.429893 2.20829 137.732 83.7604 18.7116 60.7892 0.00403191 0 -40 10
1.566 4.53151e-08 2.53964e-06 0.140481 0.14048 0.012029 2.05978e-05 0.00115438 0.175601 0.0006587 0.176255 0.934562 101.554 0.237019 0.829489 4.44563 0.0629808 0.0419399 0.95806 0.0195365 0.00451616 0.018796 0.00431557 0.00546345 0.00620396 0.218538 0.248158 58.0374 -87.8984 126.197 15.942 145.032 0.000141844 0.267279 192.758 0.310272 0.0673348 0.00409792 0.000562254 0.00138469 0.986965 0.991719 -2.98732e-06 -85.6588 0.093069 31173.2 307.958 0.983501 0.319146 0.735814 0.73581 9.99958 2.98553e-06 1.1942e-05 0.133431 0.983334 0.931539 -0.0132919 4.925e-06 0.512464 -1.98435e-20 7.35256e-24 -1.98362e-20 0.00139624 0.997815 8.60077e-05 0.152703 2.85262 0.00139624 0.997816 0.775596 0.00106437 0.00188111 0.000860077 0.455429 0.00188111 0.44344 0.000130776 1.02 0.888557 0.534435 0.287267 1.71894e-07 3.07987e-09 2373.96 3129.11 -0.0571835 0.482193 0.277328 0.254143 -0.593195 -0.169562 0.49087 -0.266194 -0.224685 2.468 1 0 296.262 0 2.20824 2.466 0.000299335 0.861843 0.691973 0.324203 0.429916 2.20843 137.739 83.7599 18.7116 60.7889 0.00403193 0 -40 10
1.567 4.5344e-08 2.53964e-06 0.140519 0.140518 0.012029 2.06109e-05 0.00115438 0.175649 0.000658701 0.176303 0.934649 101.554 0.237009 0.829619 4.44617 0.0629912 0.041945 0.958055 0.019536 0.00451657 0.0187955 0.00431592 0.00546396 0.00620448 0.218558 0.248179 58.0375 -87.8984 126.197 15.942 145.032 0.000141846 0.26728 192.758 0.310272 0.0673348 0.00409792 0.000562254 0.00138469 0.986965 0.991719 -2.98733e-06 -85.6588 0.0930691 31173.2 307.97 0.983501 0.319146 0.735825 0.735821 9.99958 2.98554e-06 1.1942e-05 0.133436 0.983334 0.931538 -0.0132919 4.92503e-06 0.512482 -1.9845e-20 7.35314e-24 -1.98376e-20 0.00139624 0.997815 8.60078e-05 0.152703 2.85262 0.00139624 0.997816 0.775674 0.00106438 0.00188111 0.000860078 0.455429 0.00188111 0.443446 0.000130778 1.02 0.888558 0.534435 0.287269 1.71895e-07 3.07989e-09 2373.95 3129.16 -0.0571882 0.482194 0.277328 0.254146 -0.593195 -0.169562 0.490855 -0.266192 -0.224672 2.469 1 0 296.258 0 2.20838 2.467 0.000299334 0.861869 0.692017 0.324155 0.429938 2.20857 137.747 83.7594 18.7116 60.7887 0.00403195 0 -40 10
1.568 4.53728e-08 2.53964e-06 0.140557 0.140557 0.012029 2.0624e-05 0.00115438 0.175697 0.000658702 0.176351 0.934736 101.553 0.236998 0.829748 4.44671 0.0630017 0.0419501 0.95805 0.0195355 0.00451699 0.018795 0.00431627 0.00546447 0.006205 0.218579 0.2482 58.0376 -87.8984 126.196 15.942 145.032 0.000141848 0.26728 192.757 0.310271 0.0673347 0.00409792 0.000562255 0.00138469 0.986965 0.991719 -2.98735e-06 -85.6588 0.0930691 31173.2 307.981 0.983501 0.319146 0.735836 0.735831 9.99958 2.98554e-06 1.19421e-05 0.13344 0.983335 0.931537 -0.0132919 4.92506e-06 0.5125 -1.98464e-20 7.35371e-24 -1.9839e-20 0.00139624 0.997815 8.60079e-05 0.152703 2.85262 0.00139624 0.997816 0.775751 0.0010644 0.00188112 0.000860079 0.455429 0.00188111 0.443451 0.000130781 1.02 0.888559 0.534434 0.28727 1.71895e-07 3.07991e-09 2373.93 3129.21 -0.0571929 0.482194 0.277328 0.254149 -0.593194 -0.169562 0.49084 -0.26619 -0.224659 2.47 1 0 296.254 0 2.20852 2.468 0.000299333 0.861894 0.692061 0.324106 0.429961 2.2087 137.754 83.7588 18.7115 60.7884 0.00403197 0 -40 10
1.569 4.54017e-08 2.53964e-06 0.140596 0.140595 0.012029 2.06371e-05 0.00115438 0.175745 0.000658702 0.176399 0.934823 101.553 0.236988 0.829877 4.44725 0.0630121 0.0419552 0.958045 0.019535 0.0045174 0.0187945 0.00431663 0.00546498 0.00620552 0.218599 0.248221 58.0376 -87.8985 126.196 15.9419 145.032 0.00014185 0.26728 192.757 0.310271 0.0673347 0.00409793 0.000562256 0.00138469 0.986965 0.991719 -2.98736e-06 -85.6588 0.0930692 31173.1 307.992 0.983501 0.319146 0.735847 0.735842 9.99958 2.98555e-06 1.19421e-05 0.133444 0.983335 0.931536 -0.0132919 4.92509e-06 0.512518 -1.98478e-20 7.35429e-24 -1.98405e-20 0.00139625 0.997815 8.6008e-05 0.152704 2.85262 0.00139625 0.997816 0.775829 0.00106442 0.00188112 0.00086008 0.455428 0.00188112 0.443457 0.000130784 1.02 0.88856 0.534434 0.287272 1.71895e-07 3.07993e-09 2373.91 3129.25 -0.0571976 0.482194 0.277327 0.254152 -0.593194 -0.169562 0.490825 -0.266188 -0.224647 2.471 1 0 296.249 0 2.20866 2.469 0.000299332 0.86192 0.692104 0.324058 0.429984 2.20884 137.762 83.7583 18.7115 60.7881 0.00403199 0 -40 10
1.57 4.54305e-08 2.53965e-06 0.140634 0.140633 0.012029 2.06502e-05 0.00115438 0.175793 0.000658703 0.176447 0.93491 101.552 0.236977 0.830007 4.44779 0.0630226 0.0419603 0.95804 0.0195345 0.00451781 0.018794 0.00431698 0.00546549 0.00620604 0.218619 0.248242 58.0377 -87.8985 126.196 15.9419 145.032 0.000141852 0.26728 192.757 0.31027 0.0673346 0.00409793 0.000562256 0.0013847 0.986965 0.991719 -2.98738e-06 -85.6588 0.0930693 31173.1 308.003 0.983501 0.319146 0.735858 0.735853 9.99958 2.98555e-06 1.19421e-05 0.133448 0.983336 0.931535 -0.0132919 4.92511e-06 0.512536 -1.98493e-20 7.35487e-24 -1.98419e-20 0.00139625 0.997815 8.6008e-05 0.152704 2.85262 0.00139625 0.997816 0.775907 0.00106443 0.00188112 0.00086008 0.455428 0.00188112 0.443463 0.000130786 1.02 0.888561 0.534434 0.287274 1.71895e-07 3.07996e-09 2373.9 3129.3 -0.0572023 0.482194 0.277327 0.254155 -0.593193 -0.169562 0.49081 -0.266185 -0.224634 2.472 1 0 296.245 0 2.2088 2.47 0.000299331 0.861946 0.692148 0.32401 0.430006 2.20898 137.769 83.7577 18.7115 60.7879 0.00403202 0 -40 10
1.571 4.54594e-08 2.53965e-06 0.140672 0.140672 0.012029 2.06634e-05 0.00115439 0.17584 0.000658704 0.176494 0.934997 101.552 0.236967 0.830136 4.44833 0.063033 0.0419654 0.958035 0.019534 0.00451822 0.0187934 0.00431734 0.00546599 0.00620656 0.21864 0.248262 58.0378 -87.8985 126.196 15.9419 145.032 0.000141854 0.26728 192.757 0.31027 0.0673346 0.00409793 0.000562257 0.0013847 0.986965 0.991719 -2.98739e-06 -85.6587 0.0930694 31173.1 308.014 0.983501 0.319146 0.735868 0.735864 9.99958 2.98556e-06 1.19421e-05 0.133452 0.983336 0.931534 -0.0132919 4.92514e-06 0.512553 -1.98507e-20 7.35545e-24 -1.98434e-20 0.00139625 0.997815 8.60081e-05 0.152704 2.85262 0.00139625 0.997816 0.775985 0.00106445 0.00188112 0.000860081 0.455428 0.00188112 0.443469 0.000130789 1.02 0.888562 0.534433 0.287275 1.71896e-07 3.07998e-09 2373.88 3129.34 -0.057207 0.482194 0.277327 0.254158 -0.593193 -0.169562 0.490795 -0.266183 -0.224621 2.473 1 0 296.241 0 2.20894 2.471 0.00029933 0.861971 0.692192 0.323961 0.430029 2.20912 137.777 83.7572 18.7114 60.7876 0.00403204 0 -40 10
1.572 4.54883e-08 2.53965e-06 0.140711 0.14071 0.0120289 2.06765e-05 0.00115439 0.175888 0.000658704 0.176542 0.935084 101.551 0.236957 0.830265 4.44887 0.0630434 0.0419705 0.95803 0.0195335 0.00451864 0.0187929 0.00431769 0.0054665 0.00620708 0.21866 0.248283 58.0378 -87.8985 126.196 15.9418 145.032 0.000141856 0.267281 192.757 0.31027 0.0673345 0.00409793 0.000562258 0.0013847 0.986965 0.991719 -2.98741e-06 -85.6587 0.0930695 31173.1 308.026 0.983501 0.319146 0.735879 0.735875 9.99958 2.98556e-06 1.19421e-05 0.133457 0.983337 0.931533 -0.0132919 4.92517e-06 0.512571 -1.98521e-20 7.35603e-24 -1.98448e-20 0.00139625 0.997815 8.60082e-05 0.152704 2.85262 0.00139625 0.997816 0.776063 0.00106447 0.00188112 0.000860082 0.455428 0.00188112 0.443474 0.000130791 1.02 0.888564 0.534433 0.287277 1.71896e-07 3.08e-09 2373.86 3129.39 -0.0572117 0.482194 0.277327 0.254161 -0.593192 -0.169562 0.49078 -0.266181 -0.224608 2.474 1 0 296.237 0 2.20908 2.472 0.000299329 0.861997 0.692235 0.323913 0.430052 2.20926 137.784 83.7567 18.7114 60.7874 0.00403206 0 -40 10
1.573 4.55171e-08 2.53965e-06 0.140749 0.140748 0.0120289 2.06896e-05 0.00115439 0.175936 0.000658705 0.17659 0.935171 101.551 0.236946 0.830395 4.44941 0.0630539 0.0419756 0.958024 0.019533 0.00451905 0.0187924 0.00431805 0.00546701 0.0062076 0.21868 0.248304 58.0379 -87.8985 126.195 15.9418 145.032 0.000141858 0.267281 192.757 0.310269 0.0673345 0.00409794 0.000562258 0.0013847 0.986965 0.991719 -2.98742e-06 -85.6587 0.0930696 31173.1 308.037 0.983501 0.319146 0.73589 0.735886 9.99958 2.98557e-06 1.19422e-05 0.133461 0.983337 0.931533 -0.0132919 4.9252e-06 0.512589 -1.98536e-20 7.3566e-24 -1.98462e-20 0.00139625 0.997815 8.60083e-05 0.152704 2.85262 0.00139625 0.997816 0.77614 0.00106448 0.00188112 0.000860083 0.455427 0.00188112 0.44348 0.000130794 1.02 0.888565 0.534433 0.287278 1.71896e-07 3.08003e-09 2373.85 3129.43 -0.0572164 0.482194 0.277326 0.254164 -0.593191 -0.169562 0.490765 -0.266179 -0.224595 2.475 1 0 296.233 0 2.20922 2.473 0.000299328 0.862023 0.692279 0.323865 0.430075 2.2094 137.792 83.7561 18.7114 60.7871 0.00403208 0 -40 10
1.574 4.5546e-08 2.53965e-06 0.140787 0.140786 0.0120289 2.07027e-05 0.00115439 0.175984 0.000658706 0.176638 0.935259 101.55 0.236936 0.830524 4.44995 0.0630643 0.0419807 0.958019 0.0195325 0.00451946 0.0187919 0.0043184 0.00546752 0.00620812 0.218701 0.248325 58.0379 -87.8985 126.195 15.9417 145.032 0.00014186 0.267281 192.756 0.310269 0.0673344 0.00409794 0.000562259 0.00138471 0.986965 0.991719 -2.98744e-06 -85.6587 0.0930697 31173 308.048 0.983501 0.319146 0.735901 0.735897 9.99958 2.98557e-06 1.19422e-05 0.133465 0.983338 0.931532 -0.0132919 4.92523e-06 0.512607 -1.9855e-20 7.35718e-24 -1.98477e-20 0.00139625 0.997815 8.60084e-05 0.152704 2.85262 0.00139625 0.997816 0.776218 0.0010645 0.00188112 0.000860084 0.455427 0.00188112 0.443486 0.000130796 1.02 0.888566 0.534432 0.28728 1.71896e-07 3.08005e-09 2373.83 3129.48 -0.0572211 0.482194 0.277326 0.254167 -0.593191 -0.169562 0.49075 -0.266177 -0.224582 2.476 1 0 296.228 0 2.20936 2.474 0.000299326 0.862049 0.692323 0.323817 0.430097 2.20954 137.799 83.7556 18.7113 60.7868 0.00403211 0 -40 10
1.575 4.55748e-08 2.53965e-06 0.140825 0.140825 0.0120289 2.07158e-05 0.00115439 0.176031 0.000658706 0.176686 0.935346 101.55 0.236925 0.830654 4.4505 0.0630748 0.0419858 0.958014 0.019532 0.00451988 0.0187914 0.00431876 0.00546803 0.00620864 0.218721 0.248346 58.038 -87.8985 126.195 15.9417 145.032 0.000141863 0.267281 192.756 0.310268 0.0673344 0.00409794 0.00056226 0.00138471 0.986965 0.991719 -2.98745e-06 -85.6587 0.0930698 31173 308.059 0.983501 0.319146 0.735912 0.735908 9.99958 2.98558e-06 1.19422e-05 0.133469 0.983338 0.931531 -0.0132919 4.92526e-06 0.512625 -1.98565e-20 7.35776e-24 -1.98491e-20 0.00139625 0.997815 8.60084e-05 0.152705 2.85262 0.00139625 0.997816 0.776296 0.00106452 0.00188113 0.000860084 0.455427 0.00188112 0.443491 0.000130799 1.02 0.888567 0.534432 0.287281 1.71897e-07 3.08007e-09 2373.82 3129.52 -0.0572258 0.482194 0.277326 0.25417 -0.59319 -0.169562 0.490735 -0.266175 -0.224569 2.477 1 0 296.224 0 2.2095 2.475 0.000299325 0.862075 0.692366 0.323769 0.43012 2.20968 137.807 83.7551 18.7113 60.7866 0.00403213 0 -40 10
1.576 4.56037e-08 2.53965e-06 0.140863 0.140863 0.0120289 2.0729e-05 0.00115439 0.176079 0.000658707 0.176733 0.935433 101.549 0.236915 0.830783 4.45104 0.0630852 0.0419909 0.958009 0.0195315 0.00452029 0.0187908 0.00431911 0.00546854 0.00620917 0.218742 0.248367 58.0381 -87.8985 126.195 15.9417 145.032 0.000141865 0.267281 192.756 0.310268 0.0673343 0.00409795 0.00056226 0.00138471 0.986964 0.991719 -2.98747e-06 -85.6587 0.0930698 31173 308.07 0.983501 0.319146 0.735923 0.735918 9.99958 2.98558e-06 1.19422e-05 0.133474 0.983339 0.93153 -0.0132919 4.92529e-06 0.512643 -1.98579e-20 7.35834e-24 -1.98506e-20 0.00139625 0.997815 8.60085e-05 0.152705 2.85262 0.00139625 0.997816 0.776373 0.00106453 0.00188113 0.000860085 0.455427 0.00188113 0.443497 0.000130801 1.02 0.888568 0.534432 0.287283 1.71897e-07 3.08009e-09 2373.8 3129.57 -0.0572305 0.482194 0.277325 0.254173 -0.59319 -0.169562 0.49072 -0.266173 -0.224556 2.478 1 0 296.22 0 2.20963 2.476 0.000299324 0.8621 0.69241 0.323721 0.430143 2.20982 137.814 83.7545 18.7113 60.7863 0.00403215 0 -40 10
1.577 4.56326e-08 2.53966e-06 0.140901 0.140901 0.0120289 2.07421e-05 0.00115439 0.176127 0.000658708 0.176781 0.93552 101.548 0.236904 0.830913 4.45158 0.0630957 0.0419961 0.958004 0.0195309 0.00452071 0.0187903 0.00431947 0.00546905 0.00620969 0.218762 0.248388 58.0381 -87.8985 126.195 15.9416 145.032 0.000141867 0.267282 192.756 0.310267 0.0673343 0.00409795 0.000562261 0.00138471 0.986964 0.991719 -2.98748e-06 -85.6587 0.0930699 31173 308.082 0.983501 0.319146 0.735934 0.735929 9.99958 2.98559e-06 1.19422e-05 0.133478 0.983339 0.931529 -0.0132919 4.92532e-06 0.512661 -1.98594e-20 7.35892e-24 -1.9852e-20 0.00139625 0.997815 8.60086e-05 0.152705 2.85263 0.00139625 0.997816 0.776451 0.00106455 0.00188113 0.000860086 0.455427 0.00188113 0.443503 0.000130804 1.02 0.888569 0.534431 0.287284 1.71897e-07 3.08012e-09 2373.78 3129.62 -0.0572352 0.482194 0.277325 0.254175 -0.593189 -0.169562 0.490704 -0.266171 -0.224543 2.479 1 0 296.216 0 2.20977 2.477 0.000299323 0.862126 0.692454 0.323673 0.430165 2.20996 137.822 83.754 18.7112 60.7861 0.00403217 0 -40 10
1.578 4.56614e-08 2.53966e-06 0.14094 0.140939 0.0120289 2.07552e-05 0.00115439 0.176174 0.000658708 0.176829 0.935607 101.548 0.236894 0.831042 4.45213 0.0631061 0.0420012 0.957999 0.0195304 0.00452112 0.0187898 0.00431983 0.00546956 0.00621021 0.218783 0.248408 58.0382 -87.8985 126.194 15.9416 145.032 0.000141869 0.267282 192.756 0.310267 0.0673342 0.00409795 0.000562262 0.00138471 0.986964 0.991719 -2.9875e-06 -85.6587 0.09307 31172.9 308.093 0.983501 0.319146 0.735945 0.73594 9.99958 2.98559e-06 1.19423e-05 0.133482 0.98334 0.931528 -0.0132919 4.92535e-06 0.512678 -1.98608e-20 7.3595e-24 -1.98534e-20 0.00139626 0.997815 8.60087e-05 0.152705 2.85263 0.00139626 0.997816 0.776529 0.00106457 0.00188113 0.000860087 0.455426 0.00188113 0.443508 0.000130807 1.02 0.88857 0.534431 0.287286 1.71897e-07 3.08014e-09 2373.77 3129.66 -0.0572399 0.482194 0.277325 0.254178 -0.593188 -0.169562 0.490689 -0.266169 -0.22453 2.48 1 0 296.211 0 2.20991 2.478 0.000299322 0.862152 0.692497 0.323625 0.430188 2.2101 137.829 83.7534 18.7112 60.7858 0.00403219 0 -40 10
1.579 4.56903e-08 2.53966e-06 0.140978 0.140977 0.0120288 2.07683e-05 0.00115439 0.176222 0.000658709 0.176876 0.935694 101.547 0.236883 0.831172 4.45267 0.0631166 0.0420063 0.957994 0.0195299 0.00452153 0.0187893 0.00432018 0.00547007 0.00621073 0.218803 0.248429 58.0383 -87.8985 126.194 15.9416 145.032 0.000141871 0.267282 192.756 0.310267 0.0673342 0.00409796 0.000562262 0.00138472 0.986964 0.991719 -2.98751e-06 -85.6587 0.0930701 31172.9 308.104 0.983501 0.319146 0.735956 0.735951 9.99958 2.9856e-06 1.19423e-05 0.133486 0.98334 0.931527 -0.0132919 4.92538e-06 0.512696 -1.98622e-20 7.36008e-24 -1.98549e-20 0.00139626 0.997815 8.60088e-05 0.152705 2.85263 0.00139626 0.997816 0.776606 0.00106458 0.00188113 0.000860088 0.455426 0.00188113 0.443514 0.000130809 1.02 0.888571 0.534431 0.287287 1.71898e-07 3.08016e-09 2373.75 3129.71 -0.0572447 0.482194 0.277325 0.254181 -0.593188 -0.169562 0.490674 -0.266167 -0.224517 2.481 1 0 296.207 0 2.21005 2.479 0.000299321 0.862178 0.692541 0.323577 0.430211 2.21024 137.837 83.7529 18.7112 60.7855 0.00403222 0 -40 10
1.58 4.57192e-08 2.53966e-06 0.141016 0.141015 0.0120288 2.07814e-05 0.00115439 0.176269 0.00065871 0.176924 0.935782 101.547 0.236873 0.831301 4.45322 0.0631271 0.0420115 0.957989 0.0195294 0.00452195 0.0187887 0.00432054 0.00547058 0.00621126 0.218823 0.24845 58.0383 -87.8985 126.194 15.9415 145.032 0.000141873 0.267282 192.755 0.310266 0.0673341 0.00409796 0.000562263 0.00138472 0.986964 0.991719 -2.98753e-06 -85.6587 0.0930702 31172.9 308.116 0.983501 0.319146 0.735967 0.735962 9.99958 2.9856e-06 1.19423e-05 0.13349 0.983341 0.931527 -0.0132919 4.92541e-06 0.512714 -1.98637e-20 7.36066e-24 -1.98563e-20 0.00139626 0.997815 8.60088e-05 0.152705 2.85263 0.00139626 0.997816 0.776684 0.0010646 0.00188113 0.000860088 0.455426 0.00188113 0.44352 0.000130812 1.02 0.888572 0.534431 0.287289 1.71898e-07 3.08019e-09 2373.73 3129.75 -0.0572494 0.482195 0.277324 0.254184 -0.593187 -0.169562 0.490659 -0.266164 -0.224504 2.482 1 0 296.203 0 2.21019 2.48 0.00029932 0.862204 0.692584 0.323529 0.430233 2.21038 137.844 83.7524 18.7112 60.7853 0.00403224 0 -40 10
1.581 4.5748e-08 2.53966e-06 0.141054 0.141053 0.0120288 2.07946e-05 0.00115439 0.176317 0.00065871 0.176971 0.935869 101.546 0.236862 0.831431 4.45376 0.0631375 0.0420166 0.957983 0.0195289 0.00452237 0.0187882 0.0043209 0.0054711 0.00621178 0.218844 0.248471 58.0384 -87.8985 126.194 15.9415 145.032 0.000141875 0.267282 192.755 0.310266 0.0673341 0.00409796 0.000562264 0.00138472 0.986964 0.991719 -2.98755e-06 -85.6586 0.0930703 31172.9 308.127 0.983501 0.319146 0.735978 0.735973 9.99958 2.98561e-06 1.19423e-05 0.133495 0.983341 0.931526 -0.0132919 4.92544e-06 0.512732 -1.98651e-20 7.36125e-24 -1.98578e-20 0.00139626 0.997815 8.60089e-05 0.152705 2.85263 0.00139626 0.997816 0.776761 0.00106462 0.00188113 0.000860089 0.455426 0.00188113 0.443525 0.000130814 1.02 0.888573 0.53443 0.28729 1.71898e-07 3.08021e-09 2373.72 3129.8 -0.0572541 0.482195 0.277324 0.254187 -0.593187 -0.169562 0.490644 -0.266162 -0.224491 2.483 1 0 296.199 0 2.21033 2.481 0.000299319 0.86223 0.692628 0.323481 0.430256 2.21051 137.852 83.7518 18.7111 60.785 0.00403226 0 -40 10
1.582 4.57769e-08 2.53966e-06 0.141092 0.141091 0.0120288 2.08077e-05 0.00115439 0.176364 0.000658711 0.177019 0.935956 101.546 0.236852 0.83156 4.45431 0.063148 0.0420218 0.957978 0.0195284 0.00452278 0.0187877 0.00432125 0.00547161 0.00621231 0.218864 0.248492 58.0384 -87.8985 126.194 15.9414 145.032 0.000141877 0.267282 192.755 0.310265 0.067334 0.00409797 0.000562264 0.00138472 0.986964 0.991719 -2.98756e-06 -85.6586 0.0930704 31172.9 308.138 0.983501 0.319146 0.735989 0.735984 9.99958 2.98561e-06 1.19423e-05 0.133499 0.983342 0.931525 -0.0132918 4.92547e-06 0.51275 -1.98666e-20 7.36183e-24 -1.98592e-20 0.00139626 0.997815 8.6009e-05 0.152706 2.85263 0.00139626 0.997816 0.776839 0.00106464 0.00188114 0.00086009 0.455425 0.00188113 0.443531 0.000130817 1.02 0.888575 0.53443 0.287292 1.71899e-07 3.08023e-09 2373.7 3129.85 -0.0572588 0.482195 0.277324 0.25419 -0.593186 -0.169563 0.490629 -0.26616 -0.224478 2.484 1 0 296.194 0 2.21047 2.482 0.000299318 0.862256 0.692672 0.323434 0.430279 2.21065 137.859 83.7513 18.7111 60.7848 0.00403228 0 -40 10
1.583 4.58057e-08 2.53966e-06 0.141129 0.141129 0.0120288 2.08208e-05 0.00115439 0.176412 0.000658712 0.177066 0.936043 101.545 0.236842 0.83169 4.45485 0.0631584 0.0420269 0.957973 0.0195279 0.0045232 0.0187872 0.00432161 0.00547212 0.00621283 0.218885 0.248513 58.0385 -87.8985 126.193 15.9414 145.032 0.000141879 0.267283 192.755 0.310265 0.0673339 0.00409797 0.000562265 0.00138473 0.986964 0.991719 -2.98758e-06 -85.6586 0.0930705 31172.8 308.149 0.983501 0.319146 0.735999 0.735995 9.99958 2.98562e-06 1.19424e-05 0.133503 0.983342 0.931524 -0.0132918 4.9255e-06 0.512768 -1.9868e-20 7.36241e-24 -1.98607e-20 0.00139626 0.997815 8.60091e-05 0.152706 2.85263 0.00139626 0.997816 0.776916 0.00106465 0.00188114 0.000860091 0.455425 0.00188114 0.443537 0.000130819 1.02 0.888576 0.53443 0.287293 1.71899e-07 3.08025e-09 2373.68 3129.89 -0.0572636 0.482195 0.277323 0.254193 -0.593186 -0.169563 0.490614 -0.266158 -0.224465 2.485 1 0 296.19 0 2.21061 2.483 0.000299317 0.862282 0.692715 0.323386 0.430301 2.21079 137.867 83.7507 18.7111 60.7845 0.00403231 0 -40 10
1.584 4.58346e-08 2.53967e-06 0.141167 0.141167 0.0120288 2.08339e-05 0.00115439 0.176459 0.000658712 0.177113 0.936131 101.545 0.236831 0.83182 4.4554 0.0631689 0.0420321 0.957968 0.0195274 0.00452361 0.0187866 0.00432197 0.00547263 0.00621335 0.218905 0.248534 58.0386 -87.8985 126.193 15.9414 145.032 0.000141882 0.267283 192.755 0.310264 0.0673339 0.00409797 0.000562266 0.00138473 0.986964 0.991719 -2.98759e-06 -85.6586 0.0930705 31172.8 308.161 0.983501 0.319146 0.73601 0.736006 9.99958 2.98562e-06 1.19424e-05 0.133507 0.983343 0.931523 -0.0132918 4.92553e-06 0.512786 -1.98695e-20 7.36299e-24 -1.98621e-20 0.00139626 0.997815 8.60092e-05 0.152706 2.85263 0.00139626 0.997816 0.776993 0.00106467 0.00188114 0.000860092 0.455425 0.00188114 0.443542 0.000130822 1.02 0.888577 0.534429 0.287295 1.71899e-07 3.08028e-09 2373.67 3129.94 -0.0572683 0.482195 0.277323 0.254196 -0.593185 -0.169563 0.490599 -0.266156 -0.224452 2.486 1 0 296.186 0 2.21075 2.484 0.000299316 0.862308 0.692759 0.323338 0.430324 2.21093 137.874 83.7502 18.711 60.7842 0.00403233 0 -40 10
1.585 4.58635e-08 2.53967e-06 0.141205 0.141205 0.0120288 2.0847e-05 0.00115439 0.176507 0.000658713 0.177161 0.936218 101.544 0.236821 0.831949 4.45595 0.0631794 0.0420372 0.957963 0.0195269 0.00452403 0.0187861 0.00432233 0.00547315 0.00621388 0.218926 0.248555 58.0386 -87.8985 126.193 15.9413 145.032 0.000141884 0.267283 192.755 0.310264 0.0673338 0.00409797 0.000562266 0.00138473 0.986964 0.991719 -2.98761e-06 -85.6586 0.0930706 31172.8 308.172 0.983501 0.319146 0.736021 0.736017 9.99958 2.98563e-06 1.19424e-05 0.133512 0.983343 0.931522 -0.0132918 4.92556e-06 0.512804 -1.98709e-20 7.36357e-24 -1.98636e-20 0.00139626 0.997815 8.60092e-05 0.152706 2.85263 0.00139626 0.997816 0.777071 0.00106469 0.00188114 0.000860092 0.455425 0.00188114 0.443548 0.000130824 1.02 0.888578 0.534429 0.287296 1.71899e-07 3.0803e-09 2373.65 3129.98 -0.057273 0.482195 0.277323 0.254199 -0.593184 -0.169563 0.490584 -0.266154 -0.224439 2.487 1 0 296.182 0 2.21089 2.485 0.000299315 0.862334 0.692802 0.323291 0.430347 2.21107 137.881 83.7497 18.711 60.784 0.00403235 0 -40 10
1.586 4.58923e-08 2.53967e-06 0.141243 0.141242 0.0120287 2.08601e-05 0.00115439 0.176554 0.000658714 0.177208 0.936305 101.544 0.23681 0.832079 4.45649 0.0631898 0.0420424 0.957958 0.0195263 0.00452444 0.0187856 0.00432268 0.00547366 0.00621441 0.218946 0.248576 58.0387 -87.8985 126.193 15.9413 145.032 0.000141886 0.267283 192.754 0.310264 0.0673338 0.00409798 0.000562267 0.00138473 0.986964 0.991719 -2.98762e-06 -85.6586 0.0930707 31172.8 308.183 0.983501 0.319146 0.736032 0.736028 9.99958 2.98563e-06 1.19424e-05 0.133516 0.983344 0.931521 -0.0132918 4.92559e-06 0.512822 -1.98724e-20 7.36416e-24 -1.9865e-20 0.00139627 0.997815 8.60093e-05 0.152706 2.85263 0.00139627 0.997816 0.777148 0.0010647 0.00188114 0.000860093 0.455425 0.00188114 0.443554 0.000130827 1.02 0.888579 0.534429 0.287298 1.719e-07 3.08032e-09 2373.63 3130.03 -0.0572778 0.482195 0.277323 0.254202 -0.593184 -0.169563 0.490569 -0.266152 -0.224426 2.488 1 0 296.177 0 2.21103 2.486 0.000299314 0.86236 0.692846 0.323243 0.430369 2.21121 137.889 83.7491 18.711 60.7837 0.00403237 0 -40 10
1.587 4.59212e-08 2.53967e-06 0.141281 0.14128 0.0120287 2.08733e-05 0.0011544 0.176601 0.000658714 0.177255 0.936393 101.543 0.2368 0.832209 4.45704 0.0632003 0.0420476 0.957952 0.0195258 0.00452486 0.0187851 0.00432304 0.00547417 0.00621493 0.218967 0.248597 58.0388 -87.8985 126.193 15.9413 145.032 0.000141888 0.267283 192.754 0.310263 0.0673337 0.00409798 0.000562268 0.00138473 0.986964 0.991719 -2.98764e-06 -85.6586 0.0930708 31172.7 308.195 0.983501 0.319146 0.736043 0.736039 9.99958 2.98564e-06 1.19424e-05 0.13352 0.983344 0.931521 -0.0132918 4.92562e-06 0.51284 -1.98738e-20 7.36474e-24 -1.98665e-20 0.00139627 0.997815 8.60094e-05 0.152706 2.85263 0.00139627 0.997816 0.777226 0.00106472 0.00188114 0.000860094 0.455424 0.00188114 0.443559 0.000130829 1.02 0.88858 0.534428 0.287299 1.719e-07 3.08035e-09 2373.62 3130.07 -0.0572825 0.482195 0.277322 0.254205 -0.593183 -0.169563 0.490554 -0.26615 -0.224413 2.489 1 0 296.173 0 2.21117 2.487 0.000299313 0.862386 0.69289 0.323196 0.430392 2.21135 137.896 83.7486 18.7109 60.7835 0.0040324 0 -40 10
1.588 4.595e-08 2.53967e-06 0.141319 0.141318 0.0120287 2.08864e-05 0.0011544 0.176648 0.000658715 0.177302 0.93648 101.542 0.236789 0.832338 4.45759 0.0632108 0.0420527 0.957947 0.0195253 0.00452528 0.0187845 0.0043234 0.00547469 0.00621546 0.218987 0.248618 58.0388 -87.8985 126.192 15.9412 145.032 0.00014189 0.267284 192.754 0.310263 0.0673337 0.00409798 0.000562268 0.00138474 0.986964 0.991719 -2.98765e-06 -85.6586 0.0930709 31172.7 308.206 0.983501 0.319146 0.736054 0.73605 9.99958 2.98564e-06 1.19425e-05 0.133524 0.983345 0.93152 -0.0132918 4.92565e-06 0.512858 -1.98753e-20 7.36532e-24 -1.98679e-20 0.00139627 0.997815 8.60095e-05 0.152707 2.85264 0.00139627 0.997816 0.777303 0.00106474 0.00188114 0.000860095 0.455424 0.00188114 0.443565 0.000130832 1.02 0.888581 0.534428 0.287301 1.719e-07 3.08037e-09 2373.6 3130.12 -0.0572872 0.482195 0.277322 0.254208 -0.593183 -0.169563 0.490538 -0.266148 -0.2244 2.49 1 0 296.169 0 2.2113 2.488 0.000299312 0.862412 0.692933 0.323148 0.430415 2.21149 137.904 83.748 18.7109 60.7832 0.00403242 0 -40 10
1.589 4.59789e-08 2.53967e-06 0.141356 0.141356 0.0120287 2.08995e-05 0.0011544 0.176695 0.000658715 0.17735 0.936568 101.542 0.236779 0.832468 4.45814 0.0632213 0.0420579 0.957942 0.0195248 0.0045257 0.018784 0.00432376 0.0054752 0.00621598 0.219008 0.248639 58.0389 -87.8985 126.192 15.9412 145.033 0.000141892 0.267284 192.754 0.310262 0.0673336 0.00409799 0.000562269 0.00138474 0.986964 0.991719 -2.98767e-06 -85.6586 0.093071 31172.7 308.217 0.983501 0.319146 0.736065 0.736061 9.99958 2.98565e-06 1.19425e-05 0.133529 0.983345 0.931519 -0.0132918 4.92568e-06 0.512876 -1.98767e-20 7.36591e-24 -1.98694e-20 0.00139627 0.997815 8.60096e-05 0.152707 2.85264 0.00139627 0.997816 0.77738 0.00106475 0.00188115 0.000860096 0.455424 0.00188115 0.443571 0.000130834 1.02 0.888582 0.534428 0.287302 1.719e-07 3.08039e-09 2373.58 3130.17 -0.057292 0.482195 0.277322 0.254211 -0.593182 -0.169563 0.490523 -0.266145 -0.224387 2.491 1 0 296.165 0 2.21144 2.489 0.000299311 0.862438 0.692977 0.323101 0.430437 2.21163 137.911 83.7475 18.7109 60.7829 0.00403244 0 -40 10
1.59 4.60077e-08 2.53967e-06 0.141394 0.141393 0.0120287 2.09126e-05 0.0011544 0.176743 0.000658716 0.177397 0.936655 101.541 0.236768 0.832598 4.45869 0.0632317 0.0420631 0.957937 0.0195243 0.00452611 0.0187835 0.00432412 0.00547571 0.00621651 0.219029 0.24866 58.0389 -87.8985 126.192 15.9411 145.033 0.000141894 0.267284 192.754 0.310262 0.0673336 0.00409799 0.00056227 0.00138474 0.986964 0.991719 -2.98768e-06 -85.6586 0.0930711 31172.7 308.229 0.983501 0.319146 0.736076 0.736072 9.99958 2.98565e-06 1.19425e-05 0.133533 0.983346 0.931518 -0.0132918 4.92571e-06 0.512894 -1.98782e-20 7.36649e-24 -1.98708e-20 0.00139627 0.997815 8.60096e-05 0.152707 2.85264 0.00139627 0.997816 0.777457 0.00106477 0.00188115 0.000860096 0.455424 0.00188115 0.443576 0.000130837 1.02 0.888583 0.534427 0.287304 1.71901e-07 3.08042e-09 2373.57 3130.21 -0.0572967 0.482195 0.277321 0.254214 -0.593181 -0.169563 0.490508 -0.266143 -0.224374 2.492 1 0 296.16 0 2.21158 2.49 0.00029931 0.862464 0.69302 0.323054 0.43046 2.21177 137.919 83.747 18.7108 60.7827 0.00403246 0 -40 10
1.591 4.60366e-08 2.53968e-06 0.141432 0.141431 0.0120287 2.09257e-05 0.0011544 0.17679 0.000658717 0.177444 0.936742 101.541 0.236758 0.832728 4.45924 0.0632422 0.0420683 0.957932 0.0195238 0.00452653 0.018783 0.00432448 0.00547623 0.00621704 0.219049 0.248681 58.039 -87.8985 126.192 15.9411 145.033 0.000141896 0.267284 192.754 0.310261 0.0673335 0.00409799 0.00056227 0.00138474 0.986964 0.991719 -2.9877e-06 -85.6586 0.0930712 31172.7 308.24 0.983501 0.319146 0.736087 0.736083 9.99958 2.98566e-06 1.19425e-05 0.133537 0.983346 0.931517 -0.0132918 4.92574e-06 0.512912 -1.98796e-20 7.36707e-24 -1.98723e-20 0.00139627 0.997815 8.60097e-05 0.152707 2.85264 0.00139627 0.997816 0.777535 0.00106479 0.00188115 0.000860097 0.455423 0.00188115 0.443582 0.00013084 1.02 0.888584 0.534427 0.287305 1.71901e-07 3.08044e-09 2373.55 3130.26 -0.0573015 0.482195 0.277321 0.254217 -0.593181 -0.169563 0.490493 -0.266141 -0.224361 2.493 1 0 296.156 0 2.21172 2.491 0.000299309 0.86249 0.693064 0.323006 0.430482 2.21191 137.926 83.7464 18.7108 60.7824 0.00403249 0 -40 10
1.592 4.60655e-08 2.53968e-06 0.141469 0.141469 0.0120287 2.09388e-05 0.0011544 0.176837 0.000658717 0.177491 0.93683 101.54 0.236747 0.832857 4.45979 0.0632527 0.0420735 0.957927 0.0195233 0.00452695 0.0187824 0.00432484 0.00547674 0.00621756 0.21907 0.248703 58.0391 -87.8985 126.192 15.9411 145.033 0.000141899 0.267284 192.753 0.310261 0.0673335 0.004098 0.000562271 0.00138474 0.986964 0.991719 -2.98771e-06 -85.6585 0.0930712 31172.6 308.251 0.983501 0.319146 0.736098 0.736094 9.99958 2.98566e-06 1.19425e-05 0.133541 0.983347 0.931516 -0.0132918 4.92577e-06 0.51293 -1.98811e-20 7.36766e-24 -1.98737e-20 0.00139627 0.997815 8.60098e-05 0.152707 2.85264 0.00139627 0.997816 0.777612 0.0010648 0.00188115 0.000860098 0.455423 0.00188115 0.443588 0.000130842 1.02 0.888586 0.534427 0.287307 1.71901e-07 3.08046e-09 2373.54 3130.31 -0.0573062 0.482195 0.277321 0.25422 -0.59318 -0.169563 0.490478 -0.266139 -0.224348 2.494 1 0 296.152 0 2.21186 2.492 0.000299307 0.862516 0.693107 0.322959 0.430505 2.21204 137.934 83.7459 18.7108 60.7822 0.00403251 0 -40 10
1.593 4.60943e-08 2.53968e-06 0.141507 0.141506 0.0120286 2.0952e-05 0.0011544 0.176884 0.000658718 0.177538 0.936917 101.54 0.236737 0.832987 4.46034 0.0632632 0.0420787 0.957921 0.0195227 0.00452737 0.0187819 0.0043252 0.00547726 0.00621809 0.21909 0.248724 58.0391 -87.8985 126.191 15.941 145.033 0.000141901 0.267285 192.753 0.310261 0.0673334 0.004098 0.000562272 0.00138475 0.986964 0.991719 -2.98773e-06 -85.6585 0.0930713 31172.6 308.263 0.983501 0.319146 0.73611 0.736105 9.99958 2.98567e-06 1.19426e-05 0.133546 0.983347 0.931515 -0.0132918 4.9258e-06 0.512948 -1.98826e-20 7.36824e-24 -1.98752e-20 0.00139627 0.997815 8.60099e-05 0.152707 2.85264 0.00139627 0.997816 0.777689 0.00106482 0.00188115 0.000860099 0.455423 0.00188115 0.443593 0.000130845 1.02 0.888587 0.534427 0.287309 1.71902e-07 3.08048e-09 2373.52 3130.35 -0.057311 0.482196 0.277321 0.254223 -0.59318 -0.169563 0.490463 -0.266137 -0.224335 2.495 1 0 296.147 0 2.212 2.493 0.000299306 0.862542 0.693151 0.322912 0.430528 2.21218 137.941 83.7453 18.7107 60.7819 0.00403253 0 -40 10
1.594 4.61232e-08 2.53968e-06 0.141545 0.141544 0.0120286 2.09651e-05 0.0011544 0.176931 0.000658719 0.177585 0.937005 101.539 0.236726 0.833117 4.46089 0.0632737 0.0420839 0.957916 0.0195222 0.00452778 0.0187814 0.00432556 0.00547777 0.00621862 0.219111 0.248745 58.0392 -87.8985 126.191 15.941 145.033 0.000141903 0.267285 192.753 0.31026 0.0673334 0.004098 0.000562272 0.00138475 0.986964 0.991719 -2.98774e-06 -85.6585 0.0930714 31172.6 308.274 0.983501 0.319146 0.736121 0.736116 9.99958 2.98567e-06 1.19426e-05 0.13355 0.983348 0.931514 -0.0132918 4.92583e-06 0.512966 -1.9884e-20 7.36883e-24 -1.98766e-20 0.00139627 0.997815 8.601e-05 0.152707 2.85264 0.00139627 0.997816 0.777766 0.00106484 0.00188115 0.0008601 0.455423 0.00188115 0.443599 0.000130847 1.02 0.888588 0.534426 0.28731 1.71902e-07 3.08051e-09 2373.5 3130.4 -0.0573157 0.482196 0.27732 0.254226 -0.593179 -0.169563 0.490448 -0.266135 -0.224322 2.496 1 0 296.143 0 2.21214 2.494 0.000299305 0.862568 0.693194 0.322865 0.43055 2.21232 137.949 83.7448 18.7107 60.7816 0.00403255 0 -40 10
1.595 4.6152e-08 2.53968e-06 0.141582 0.141582 0.0120286 2.09782e-05 0.0011544 0.176978 0.000658719 0.177632 0.937092 101.539 0.236716 0.833247 4.46144 0.0632842 0.0420891 0.957911 0.0195217 0.0045282 0.0187809 0.00432592 0.00547829 0.00621915 0.219132 0.248766 58.0393 -87.8985 126.191 15.941 145.033 0.000141905 0.267285 192.753 0.31026 0.0673333 0.004098 0.000562273 0.00138475 0.986964 0.991719 -2.98776e-06 -85.6585 0.0930715 31172.6 308.285 0.983501 0.319146 0.736132 0.736127 9.99958 2.98568e-06 1.19426e-05 0.133554 0.983348 0.931514 -0.0132918 4.92586e-06 0.512984 -1.98855e-20 7.36941e-24 -1.98781e-20 0.00139628 0.997815 8.60101e-05 0.152708 2.85264 0.00139628 0.997816 0.777843 0.00106485 0.00188116 0.000860101 0.455422 0.00188115 0.443604 0.00013085 1.02 0.888589 0.534426 0.287312 1.71902e-07 3.08053e-09 2373.49 3130.44 -0.0573205 0.482196 0.27732 0.254229 -0.593179 -0.169563 0.490432 -0.266133 -0.224309 2.497 1 0 296.139 0 2.21228 2.495 0.000299304 0.862594 0.693238 0.322818 0.430573 2.21246 137.956 83.7442 18.7107 60.7814 0.00403258 0 -40 10
1.596 4.61809e-08 2.53968e-06 0.14162 0.141619 0.0120286 2.09913e-05 0.0011544 0.177025 0.00065872 0.177679 0.93718 101.538 0.236705 0.833377 4.46199 0.0632947 0.0420943 0.957906 0.0195212 0.00452862 0.0187803 0.00432628 0.0054788 0.00621968 0.219152 0.248787 58.0393 -87.8986 126.191 15.9409 145.033 0.000141907 0.267285 192.753 0.310259 0.0673333 0.00409801 0.000562274 0.00138475 0.986964 0.991719 -2.98777e-06 -85.6585 0.0930716 31172.5 308.297 0.983501 0.319146 0.736143 0.736138 9.99958 2.98568e-06 1.19426e-05 0.133558 0.983349 0.931513 -0.0132918 4.92589e-06 0.513003 -1.98869e-20 7.37e-24 -1.98796e-20 0.00139628 0.997815 8.60101e-05 0.152708 2.85264 0.00139628 0.997816 0.77792 0.00106487 0.00188116 0.000860101 0.455422 0.00188116 0.44361 0.000130852 1.02 0.88859 0.534426 0.287313 1.71902e-07 3.08055e-09 2373.47 3130.49 -0.0573252 0.482196 0.27732 0.254232 -0.593178 -0.169563 0.490417 -0.266131 -0.224296 2.498 1 0 296.135 0 2.21242 2.496 0.000299303 0.862621 0.693282 0.322771 0.430596 2.2126 137.964 83.7437 18.7106 60.7811 0.0040326 0 -40 10
1.597 4.62098e-08 2.53968e-06 0.141657 0.141657 0.0120286 2.10044e-05 0.0011544 0.177072 0.000658721 0.177726 0.937267 101.537 0.236695 0.833507 4.46255 0.0633051 0.0420995 0.957901 0.0195207 0.00452904 0.0187798 0.00432664 0.00547932 0.0062202 0.219173 0.248808 58.0394 -87.8986 126.191 15.9409 145.033 0.000141909 0.267285 192.753 0.310259 0.0673332 0.00409801 0.000562274 0.00138476 0.986964 0.991719 -2.98779e-06 -85.6585 0.0930717 31172.5 308.308 0.983501 0.319146 0.736154 0.736149 9.99958 2.98569e-06 1.19426e-05 0.133563 0.983349 0.931512 -0.0132918 4.92592e-06 0.513021 -1.98884e-20 7.37058e-24 -1.9881e-20 0.00139628 0.997815 8.60102e-05 0.152708 2.85264 0.00139628 0.997816 0.777998 0.00106489 0.00188116 0.000860102 0.455422 0.00188116 0.443616 0.000130855 1.02 0.888591 0.534425 0.287315 1.71903e-07 3.08058e-09 2373.45 3130.54 -0.05733 0.482196 0.277319 0.254235 -0.593177 -0.169564 0.490402 -0.266129 -0.224283 2.499 1 0 296.13 0 2.21256 2.497 0.000299302 0.862647 0.693325 0.322724 0.430618 2.21274 137.971 83.7431 18.7106 60.7808 0.00403262 0 -40 10
1.598 4.62386e-08 2.53969e-06 0.141695 0.141694 0.0120286 2.10176e-05 0.0011544 0.177118 0.000658721 0.177773 0.937355 101.537 0.236684 0.833637 4.4631 0.0633156 0.0421047 0.957895 0.0195202 0.00452946 0.0187793 0.004327 0.00547984 0.00622073 0.219193 0.248829 58.0394 -87.8986 126.19 15.9408 145.033 0.000141911 0.267286 192.752 0.310258 0.0673332 0.00409801 0.000562275 0.00138476 0.986964 0.991719 -2.9878e-06 -85.6585 0.0930718 31172.5 308.32 0.983501 0.319146 0.736165 0.73616 9.99958 2.98569e-06 1.19427e-05 0.133567 0.98335 0.931511 -0.0132918 4.92595e-06 0.513039 -1.98898e-20 7.37117e-24 -1.98825e-20 0.00139628 0.997815 8.60103e-05 0.152708 2.85264 0.00139628 0.997816 0.778075 0.0010649 0.00188116 0.000860103 0.455422 0.00188116 0.443621 0.000130857 1.02 0.888592 0.534425 0.287316 1.71903e-07 3.0806e-09 2373.44 3130.58 -0.0573347 0.482196 0.277319 0.254238 -0.593177 -0.169564 0.490387 -0.266127 -0.22427 2.5 1 0 296.126 0 2.21269 2.498 0.000299301 0.862673 0.693369 0.322677 0.430641 2.21288 137.978 83.7426 18.7106 60.7806 0.00403264 0 -40 10
1.599 4.62675e-08 2.53969e-06 0.141732 0.141732 0.0120286 2.10307e-05 0.0011544 0.177165 0.000658722 0.177819 0.937443 101.536 0.236674 0.833767 4.46365 0.0633261 0.0421099 0.95789 0.0195196 0.00452988 0.0187787 0.00432736 0.00548035 0.00622126 0.219214 0.248851 58.0395 -87.8986 126.19 15.9408 145.033 0.000141913 0.267286 192.752 0.310258 0.0673331 0.00409802 0.000562276 0.00138476 0.986964 0.991719 -2.98782e-06 -85.6585 0.0930719 31172.5 308.331 0.983501 0.319146 0.736176 0.736171 9.99958 2.9857e-06 1.19427e-05 0.133571 0.98335 0.93151 -0.0132918 4.92598e-06 0.513057 -1.98913e-20 7.37176e-24 -1.98839e-20 0.00139628 0.997815 8.60104e-05 0.152708 2.85265 0.00139628 0.997816 0.778152 0.00106492 0.00188116 0.000860104 0.455422 0.00188116 0.443627 0.00013086 1.02 0.888593 0.534425 0.287318 1.71903e-07 3.08062e-09 2373.42 3130.63 -0.0573395 0.482196 0.277319 0.254241 -0.593176 -0.169564 0.490372 -0.266124 -0.224257 2.501 1 0 296.122 0 2.21283 2.499 0.0002993 0.862699 0.693412 0.32263 0.430663 2.21302 137.986 83.742 18.7106 60.7803 0.00403267 0 -40 10
1.6 4.62963e-08 2.53969e-06 0.14177 0.141769 0.0120286 2.10438e-05 0.0011544 0.177212 0.000658723 0.177866 0.93753 101.536 0.236663 0.833897 4.46421 0.0633366 0.0421152 0.957885 0.0195191 0.0045303 0.0187782 0.00432772 0.00548087 0.00622179 0.219235 0.248872 58.0396 -87.8986 126.19 15.9408 145.033 0.000141916 0.267286 192.752 0.310258 0.067333 0.00409802 0.000562276 0.00138476 0.986964 0.991719 -2.98783e-06 -85.6585 0.0930719 31172.4 308.342 0.983501 0.319146 0.736187 0.736183 9.99958 2.9857e-06 1.19427e-05 0.133576 0.983351 0.931509 -0.0132918 4.926e-06 0.513075 -1.98928e-20 7.37234e-24 -1.98854e-20 0.00139628 0.997815 8.60105e-05 0.152708 2.85265 0.00139628 0.997816 0.778229 0.00106494 0.00188116 0.000860105 0.455421 0.00188116 0.443633 0.000130862 1.02 0.888594 0.534424 0.287319 1.71903e-07 3.08064e-09 2373.4 3130.68 -0.0573443 0.482196 0.277319 0.254244 -0.593176 -0.169564 0.490356 -0.266122 -0.224243 2.502 1 0 296.117 0 2.21297 2.5 0.000299299 0.862726 0.693456 0.322583 0.430686 2.21316 137.993 83.7415 18.7105 60.78 0.00403269 0 -40 10
1.601 4.63252e-08 2.53969e-06 0.141807 0.141806 0.0120285 2.10569e-05 0.0011544 0.177259 0.000658723 0.177913 0.937618 101.535 0.236653 0.834027 4.46476 0.0633471 0.0421204 0.95788 0.0195186 0.00453072 0.0187777 0.00432808 0.00548139 0.00622232 0.219256 0.248893 58.0396 -87.8986 126.19 15.9407 145.033 0.000141918 0.267286 192.752 0.310257 0.067333 0.00409802 0.000562277 0.00138476 0.986964 0.991719 -2.98785e-06 -85.6585 0.093072 31172.4 308.354 0.983501 0.319146 0.736198 0.736194 9.99958 2.98571e-06 1.19427e-05 0.13358 0.983351 0.931508 -0.0132918 4.92603e-06 0.513093 -1.98942e-20 7.37293e-24 -1.98869e-20 0.00139628 0.997815 8.60105e-05 0.152709 2.85265 0.00139628 0.997816 0.778306 0.00106495 0.00188116 0.000860105 0.455421 0.00188116 0.443638 0.000130865 1.02 0.888595 0.534424 0.287321 1.71904e-07 3.08067e-09 2373.39 3130.72 -0.057349 0.482196 0.277318 0.254247 -0.593175 -0.169564 0.490341 -0.26612 -0.22423 2.503 1 0 296.113 0 2.21311 2.501 0.000299298 0.862752 0.693499 0.322536 0.430709 2.2133 138.001 83.741 18.7105 60.7798 0.00403271 0 -40 10
1.602 4.63541e-08 2.53969e-06 0.141844 0.141844 0.0120285 2.107e-05 0.00115441 0.177305 0.000658724 0.177959 0.937705 101.535 0.236642 0.834157 4.46532 0.0633576 0.0421256 0.957874 0.0195181 0.00453114 0.0187771 0.00432844 0.00548191 0.00622285 0.219276 0.248914 58.0397 -87.8986 126.19 15.9407 145.033 0.00014192 0.267286 192.752 0.310257 0.0673329 0.00409803 0.000562278 0.00138477 0.986964 0.991719 -2.98786e-06 -85.6585 0.0930721 31172.4 308.365 0.983501 0.319146 0.736209 0.736205 9.99958 2.98571e-06 1.19427e-05 0.133584 0.983351 0.931507 -0.0132918 4.92606e-06 0.513111 -1.98957e-20 7.37352e-24 -1.98883e-20 0.00139628 0.997815 8.60106e-05 0.152709 2.85265 0.00139628 0.997816 0.778382 0.00106497 0.00188117 0.000860106 0.455421 0.00188116 0.443644 0.000130867 1.02 0.888597 0.534424 0.287322 1.71904e-07 3.08069e-09 2373.37 3130.77 -0.0573538 0.482196 0.277318 0.25425 -0.593174 -0.169564 0.490326 -0.266118 -0.224217 2.504 1 0 296.109 0 2.21325 2.502 0.000299297 0.862778 0.693543 0.322489 0.430731 2.21343 138.008 83.7404 18.7105 60.7795 0.00403273 0 -40 10
1.603 4.63829e-08 2.53969e-06 0.141882 0.141881 0.0120285 2.10831e-05 0.00115441 0.177352 0.000658724 0.178006 0.937793 101.534 0.236632 0.834287 4.46587 0.0633681 0.0421309 0.957869 0.0195176 0.00453156 0.0187766 0.0043288 0.00548242 0.00622338 0.219297 0.248935 58.0398 -87.8986 126.189 15.9407 145.033 0.000141922 0.267287 192.752 0.310256 0.0673329 0.00409803 0.000562278 0.00138477 0.986964 0.991719 -2.98788e-06 -85.6584 0.0930722 31172.4 308.377 0.983501 0.319146 0.73622 0.736216 9.99958 2.98572e-06 1.19428e-05 0.133588 0.983352 0.931506 -0.0132918 4.92609e-06 0.51313 -1.98972e-20 7.37411e-24 -1.98898e-20 0.00139628 0.997815 8.60107e-05 0.152709 2.85265 0.00139628 0.997816 0.778459 0.00106499 0.00188117 0.000860107 0.455421 0.00188117 0.443649 0.00013087 1.02 0.888598 0.534423 0.287324 1.71904e-07 3.08071e-09 2373.35 3130.82 -0.0573586 0.482196 0.277318 0.254253 -0.593174 -0.169564 0.490311 -0.266116 -0.224204 2.505 1 0 296.105 0 2.21339 2.503 0.000299296 0.862804 0.693586 0.322443 0.430754 2.21357 138.016 83.7399 18.7104 60.7793 0.00403276 0 -40 10
1.604 4.64118e-08 2.53969e-06 0.141919 0.141918 0.0120285 2.10963e-05 0.00115441 0.177399 0.000658725 0.178053 0.937881 101.534 0.236621 0.834417 4.46643 0.0633786 0.0421361 0.957864 0.0195171 0.00453198 0.0187761 0.00432916 0.00548294 0.00622391 0.219318 0.248957 58.0398 -87.8986 126.189 15.9406 145.033 0.000141924 0.267287 192.751 0.310256 0.0673328 0.00409803 0.000562279 0.00138477 0.986964 0.991719 -2.98789e-06 -85.6584 0.0930723 31172.4 308.388 0.983501 0.319146 0.736231 0.736227 9.99958 2.98572e-06 1.19428e-05 0.133593 0.983352 0.931506 -0.0132918 4.92612e-06 0.513148 -1.98986e-20 7.37469e-24 -1.98912e-20 0.00139629 0.997815 8.60108e-05 0.152709 2.85265 0.00139629 0.997816 0.778536 0.001065 0.00188117 0.000860108 0.45542 0.00188117 0.443655 0.000130872 1.02 0.888599 0.534423 0.287325 1.71905e-07 3.08074e-09 2373.34 3130.86 -0.0573634 0.482196 0.277318 0.254255 -0.593173 -0.169564 0.490296 -0.266114 -0.224191 2.506 1 0 296.1 0 2.21353 2.504 0.000299295 0.862831 0.69363 0.322396 0.430777 2.21371 138.023 83.7393 18.7104 60.779 0.00403278 0 -40 10
1.605 4.64406e-08 2.5397e-06 0.141956 0.141956 0.0120285 2.11094e-05 0.00115441 0.177445 0.000658726 0.178099 0.937968 101.533 0.236611 0.834547 4.46698 0.0633891 0.0421413 0.957859 0.0195165 0.0045324 0.0187756 0.00432953 0.00548346 0.00622445 0.219338 0.248978 58.0399 -87.8986 126.189 15.9406 145.033 0.000141926 0.267287 192.751 0.310255 0.0673328 0.00409804 0.00056228 0.00138477 0.986964 0.991719 -2.98791e-06 -85.6584 0.0930724 31172.3 308.399 0.983501 0.319146 0.736242 0.736238 9.99958 2.98573e-06 1.19428e-05 0.133597 0.983353 0.931505 -0.0132918 4.92615e-06 0.513166 -1.99001e-20 7.37528e-24 -1.98927e-20 0.00139629 0.997815 8.60109e-05 0.152709 2.85265 0.00139629 0.997816 0.778613 0.00106502 0.00188117 0.000860109 0.45542 0.00188117 0.443661 0.000130875 1.02 0.8886 0.534423 0.287327 1.71905e-07 3.08076e-09 2373.32 3130.91 -0.0573681 0.482196 0.277317 0.254258 -0.593173 -0.169564 0.49028 -0.266112 -0.224178 2.507 1 0 296.096 0 2.21367 2.505 0.000299294 0.862857 0.693673 0.322349 0.430799 2.21385 138.031 83.7388 18.7104 60.7787 0.0040328 0 -40 10
1.606 4.64695e-08 2.5397e-06 0.141993 0.141993 0.0120285 2.11225e-05 0.00115441 0.177492 0.000658726 0.178146 0.938056 101.532 0.2366 0.834677 4.46754 0.0633996 0.0421466 0.957853 0.019516 0.00453282 0.018775 0.00432989 0.00548398 0.00622498 0.219359 0.248999 58.04 -87.8986 126.189 15.9405 145.033 0.000141928 0.267287 192.751 0.310255 0.0673327 0.00409804 0.00056228 0.00138478 0.986964 0.991719 -2.98792e-06 -85.6584 0.0930725 31172.3 308.411 0.983501 0.319146 0.736254 0.736249 9.99958 2.98573e-06 1.19428e-05 0.133601 0.983353 0.931504 -0.0132918 4.92618e-06 0.513184 -1.99016e-20 7.37587e-24 -1.98942e-20 0.00139629 0.997815 8.60109e-05 0.152709 2.85265 0.00139629 0.997816 0.77869 0.00106504 0.00188117 0.000860109 0.45542 0.00188117 0.443666 0.000130877 1.02 0.888601 0.534423 0.287328 1.71905e-07 3.08078e-09 2373.31 3130.96 -0.0573729 0.482196 0.277317 0.254261 -0.593172 -0.169564 0.490265 -0.26611 -0.224165 2.508 1 0 296.092 0 2.21381 2.506 0.000299292 0.862883 0.693717 0.322303 0.430822 2.21399 138.038 83.7382 18.7103 60.7785 0.00403282 0 -40 10
1.607 4.64983e-08 2.5397e-06 0.142031 0.14203 0.0120285 2.11356e-05 0.00115441 0.177538 0.000658727 0.178192 0.938144 101.532 0.23659 0.834807 4.4681 0.0634101 0.0421518 0.957848 0.0195155 0.00453324 0.0187745 0.00433025 0.0054845 0.00622551 0.21938 0.24902 58.04 -87.8986 126.189 15.9405 145.033 0.000141931 0.267287 192.751 0.310255 0.0673327 0.00409804 0.000562281 0.00138478 0.986964 0.991719 -2.98794e-06 -85.6584 0.0930726 31172.3 308.422 0.9835 0.319146 0.736265 0.73626 9.99958 2.98574e-06 1.19428e-05 0.133606 0.983354 0.931503 -0.0132918 4.92621e-06 0.513202 -1.9903e-20 7.37646e-24 -1.98956e-20 0.00139629 0.997815 8.6011e-05 0.152709 2.85265 0.00139629 0.997816 0.778767 0.00106505 0.00188117 0.00086011 0.45542 0.00188117 0.443672 0.00013088 1.02 0.888602 0.534422 0.28733 1.71905e-07 3.0808e-09 2373.29 3131 -0.0573777 0.482197 0.277317 0.254264 -0.593171 -0.169564 0.49025 -0.266108 -0.224152 2.509 1 0 296.087 0 2.21394 2.507 0.000299291 0.86291 0.69376 0.322256 0.430844 2.21413 138.046 83.7377 18.7103 60.7782 0.00403285 0 -40 10
1.608 4.65272e-08 2.5397e-06 0.142068 0.142067 0.0120284 2.11487e-05 0.00115441 0.177585 0.000658728 0.178239 0.938231 101.531 0.236579 0.834937 4.46865 0.0634207 0.0421571 0.957843 0.019515 0.00453367 0.018774 0.00433061 0.00548502 0.00622604 0.219401 0.249042 58.0401 -87.8986 126.188 15.9405 145.033 0.000141933 0.267287 192.751 0.310254 0.0673326 0.00409804 0.000562282 0.00138478 0.986964 0.991719 -2.98795e-06 -85.6584 0.0930726 31172.3 308.434 0.9835 0.319146 0.736276 0.736271 9.99958 2.98574e-06 1.19429e-05 0.13361 0.983354 0.931502 -0.0132918 4.92624e-06 0.513221 -1.99045e-20 7.37705e-24 -1.98971e-20 0.00139629 0.997815 8.60111e-05 0.15271 2.85265 0.00139629 0.997816 0.778844 0.00106507 0.00188117 0.000860111 0.45542 0.00188117 0.443677 0.000130883 1.02 0.888603 0.534422 0.287331 1.71906e-07 3.08083e-09 2373.27 3131.05 -0.0573825 0.482197 0.277316 0.254267 -0.593171 -0.169564 0.490235 -0.266106 -0.224138 2.51 1 0 296.083 0 2.21408 2.508 0.00029929 0.862936 0.693804 0.32221 0.430867 2.21427 138.053 83.7371 18.7103 60.7779 0.00403287 0 -40 10
1.609 4.65561e-08 2.5397e-06 0.142105 0.142104 0.0120284 2.11618e-05 0.00115441 0.177631 0.000658728 0.178285 0.938319 101.531 0.236569 0.835067 4.46921 0.0634312 0.0421624 0.957838 0.0195145 0.00453409 0.0187734 0.00433098 0.00548554 0.00622657 0.219421 0.249063 58.0401 -87.8986 126.188 15.9404 145.033 0.000141935 0.267288 192.751 0.310254 0.0673326 0.00409805 0.000562282 0.00138478 0.986964 0.991719 -2.98797e-06 -85.6584 0.0930727 31172.2 308.445 0.9835 0.319146 0.736287 0.736283 9.99958 2.98575e-06 1.19429e-05 0.133614 0.983355 0.931501 -0.0132918 4.92627e-06 0.513239 -1.9906e-20 7.37764e-24 -1.98986e-20 0.00139629 0.997815 8.60112e-05 0.15271 2.85266 0.00139629 0.997816 0.77892 0.00106509 0.00188118 0.000860112 0.455419 0.00188117 0.443683 0.000130885 1.02 0.888604 0.534422 0.287333 1.71906e-07 3.08085e-09 2373.26 3131.09 -0.0573873 0.482197 0.277316 0.25427 -0.59317 -0.169564 0.490219 -0.266103 -0.224125 2.511 1 0 296.079 0 2.21422 2.509 0.000299289 0.862963 0.693847 0.322163 0.43089 2.21441 138.06 83.7366 18.7102 60.7777 0.00403289 0 -40 10
1.61 4.65849e-08 2.5397e-06 0.142142 0.142141 0.0120284 2.1175e-05 0.00115441 0.177678 0.000658729 0.178332 0.938407 101.53 0.236558 0.835197 4.46977 0.0634417 0.0421676 0.957832 0.0195139 0.00453451 0.0187729 0.00433134 0.00548606 0.00622711 0.219442 0.249084 58.0402 -87.8986 126.188 15.9404 145.033 0.000141937 0.267288 192.75 0.310253 0.0673325 0.00409805 0.000562283 0.00138478 0.986964 0.991719 -2.98798e-06 -85.6584 0.0930728 31172.2 308.457 0.9835 0.319146 0.736298 0.736294 9.99958 2.98575e-06 1.19429e-05 0.133618 0.983355 0.9315 -0.0132918 4.9263e-06 0.513257 -1.99074e-20 7.37823e-24 -1.99e-20 0.00139629 0.997815 8.60113e-05 0.15271 2.85266 0.00139629 0.997816 0.778997 0.0010651 0.00188118 0.000860113 0.455419 0.00188118 0.443689 0.000130888 1.02 0.888605 0.534421 0.287334 1.71906e-07 3.08087e-09 2373.24 3131.14 -0.0573921 0.482197 0.277316 0.254273 -0.59317 -0.169564 0.490204 -0.266101 -0.224112 2.512 1 0 296.074 0 2.21436 2.51 0.000299288 0.862989 0.693891 0.322117 0.430912 2.21454 138.068 83.736 18.7102 60.7774 0.00403291 0 -40 10
1.611 4.66138e-08 2.5397e-06 0.142179 0.142178 0.0120284 2.11881e-05 0.00115441 0.177724 0.00065873 0.178378 0.938495 101.53 0.236548 0.835327 4.47033 0.0634522 0.0421729 0.957827 0.0195134 0.00453493 0.0187724 0.0043317 0.00548658 0.00622764 0.219463 0.249106 58.0403 -87.8986 126.188 15.9404 145.033 0.000141939 0.267288 192.75 0.310253 0.0673325 0.00409805 0.000562284 0.00138479 0.986964 0.991719 -2.988e-06 -85.6584 0.0930729 31172.2 308.468 0.9835 0.319146 0.736309 0.736305 9.99958 2.98576e-06 1.19429e-05 0.133623 0.983356 0.931499 -0.0132918 4.92633e-06 0.513275 -1.99089e-20 7.37882e-24 -1.99015e-20 0.00139629 0.997815 8.60113e-05 0.15271 2.85266 0.00139629 0.997816 0.779074 0.00106512 0.00188118 0.000860113 0.455419 0.00188118 0.443694 0.00013089 1.02 0.888606 0.534421 0.287336 1.71906e-07 3.0809e-09 2373.22 3131.19 -0.0573968 0.482197 0.277316 0.254276 -0.593169 -0.169564 0.490189 -0.266099 -0.224099 2.513 1 0 296.07 0 2.2145 2.511 0.000299287 0.863016 0.693934 0.322071 0.430935 2.21468 138.075 83.7355 18.7102 60.7771 0.00403294 0 -40 10
1.612 4.66426e-08 2.53971e-06 0.142216 0.142216 0.0120284 2.12012e-05 0.00115441 0.17777 0.00065873 0.178424 0.938583 101.529 0.236537 0.835458 4.47089 0.0634627 0.0421782 0.957822 0.0195129 0.00453535 0.0187718 0.00433207 0.0054871 0.00622817 0.219484 0.249127 58.0403 -87.8986 126.188 15.9403 145.033 0.000141941 0.267288 192.75 0.310252 0.0673324 0.00409806 0.000562284 0.00138479 0.986964 0.991719 -2.98801e-06 -85.6584 0.093073 31172.2 308.48 0.9835 0.319146 0.73632 0.736316 9.99958 2.98576e-06 1.19429e-05 0.133627 0.983356 0.931498 -0.0132918 4.92636e-06 0.513294 -1.99104e-20 7.37941e-24 -1.9903e-20 0.0013963 0.997815 8.60114e-05 0.15271 2.85266 0.00139629 0.997816 0.77915 0.00106514 0.00188118 0.000860114 0.455419 0.00188118 0.4437 0.000130893 1.02 0.888608 0.534421 0.287337 1.71907e-07 3.08092e-09 2373.21 3131.24 -0.0574016 0.482197 0.277315 0.254279 -0.593168 -0.169564 0.490173 -0.266097 -0.224086 2.514 1 0 296.066 0 2.21464 2.512 0.000299286 0.863042 0.693978 0.322024 0.430957 2.21482 138.083 83.7349 18.7101 60.7769 0.00403296 0 -40 10
1.613 4.66715e-08 2.53971e-06 0.142253 0.142253 0.0120284 2.12143e-05 0.00115441 0.177816 0.000658731 0.178471 0.93867 101.529 0.236527 0.835588 4.47145 0.0634732 0.0421835 0.957817 0.0195124 0.00453578 0.0187713 0.00433243 0.00548762 0.00622871 0.219505 0.249148 58.0404 -87.8986 126.187 15.9403 145.033 0.000141943 0.267288 192.75 0.310252 0.0673324 0.00409806 0.000562285 0.00138479 0.986963 0.991719 -2.98803e-06 -85.6583 0.0930731 31172.2 308.491 0.9835 0.319146 0.736332 0.736327 9.99958 2.98577e-06 1.1943e-05 0.133631 0.983356 0.931498 -0.0132918 4.92639e-06 0.513312 -1.99118e-20 7.38e-24 -1.99045e-20 0.0013963 0.997815 8.60115e-05 0.15271 2.85266 0.0013963 0.997816 0.779227 0.00106515 0.00188118 0.000860115 0.455418 0.00188118 0.443705 0.000130895 1.02 0.888609 0.53442 0.287339 1.71907e-07 3.08094e-09 2373.19 3131.28 -0.0574064 0.482197 0.277315 0.254282 -0.593168 -0.169565 0.490158 -0.266095 -0.224073 2.515 1 0 296.062 0 2.21478 2.513 0.000299285 0.863068 0.694021 0.321978 0.43098 2.21496 138.09 83.7344 18.7101 60.7766 0.00403298 0 -40 10
1.614 4.67003e-08 2.53971e-06 0.14229 0.14229 0.0120284 2.12274e-05 0.00115441 0.177863 0.000658731 0.178517 0.938758 101.528 0.236516 0.835718 4.47201 0.0634838 0.0421888 0.957811 0.0195119 0.0045362 0.0187708 0.00433279 0.00548814 0.00622924 0.219526 0.24917 58.0405 -87.8986 126.187 15.9402 145.033 0.000141946 0.267289 192.75 0.310252 0.0673323 0.00409806 0.000562286 0.00138479 0.986963 0.991718 -2.98804e-06 -85.6583 0.0930732 31172.1 308.503 0.9835 0.319146 0.736343 0.736338 9.99958 2.98577e-06 1.1943e-05 0.133636 0.983357 0.931497 -0.0132918 4.92642e-06 0.51333 -1.99133e-20 7.38059e-24 -1.99059e-20 0.0013963 0.997815 8.60116e-05 0.152711 2.85266 0.0013963 0.997816 0.779304 0.00106517 0.00188118 0.000860116 0.455418 0.00188118 0.443711 0.000130898 1.02 0.88861 0.53442 0.28734 1.71907e-07 3.08097e-09 2373.17 3131.33 -0.0574112 0.482197 0.277315 0.254285 -0.593167 -0.169565 0.490143 -0.266093 -0.224059 2.516 1 0 296.057 0 2.21492 2.514 0.000299284 0.863095 0.694065 0.321932 0.431002 2.2151 138.098 83.7338 18.7101 60.7763 0.00403301 0 -40 10
1.615 4.67292e-08 2.53971e-06 0.142327 0.142327 0.0120283 2.12405e-05 0.00115441 0.177909 0.000658732 0.178563 0.938846 101.527 0.236506 0.835848 4.47257 0.0634943 0.042194 0.957806 0.0195113 0.00453662 0.0187702 0.00433316 0.00548866 0.00622978 0.219546 0.249191 58.0405 -87.8986 126.187 15.9402 145.033 0.000141948 0.267289 192.75 0.310251 0.0673323 0.00409807 0.000562286 0.00138479 0.986963 0.991718 -2.98806e-06 -85.6583 0.0930733 31172.1 308.514 0.9835 0.319146 0.736354 0.73635 9.99958 2.98578e-06 1.1943e-05 0.13364 0.983357 0.931496 -0.0132918 4.92645e-06 0.513348 -1.99148e-20 7.38118e-24 -1.99074e-20 0.0013963 0.997815 8.60117e-05 0.152711 2.85266 0.0013963 0.997816 0.77938 0.00106519 0.00188119 0.000860117 0.455418 0.00188118 0.443716 0.0001309 1.02 0.888611 0.53442 0.287342 1.71907e-07 3.08099e-09 2373.16 3131.38 -0.057416 0.482197 0.277314 0.254288 -0.593167 -0.169565 0.490128 -0.266091 -0.224046 2.517 1 0 296.053 0 2.21506 2.515 0.000299283 0.863121 0.694108 0.321886 0.431025 2.21524 138.105 83.7333 18.71 60.7761 0.00403303 0 -40 10
1.616 4.67581e-08 2.53971e-06 0.142364 0.142363 0.0120283 2.12537e-05 0.00115441 0.177955 0.000658733 0.178609 0.938934 101.527 0.236495 0.835979 4.47313 0.0635048 0.0421993 0.957801 0.0195108 0.00453705 0.0187697 0.00433352 0.00548918 0.00623031 0.219567 0.249212 58.0406 -87.8986 126.187 15.9402 145.033 0.00014195 0.267289 192.749 0.310251 0.0673322 0.00409807 0.000562287 0.0013848 0.986963 0.991718 -2.98807e-06 -85.6583 0.0930733 31172.1 308.526 0.9835 0.319146 0.736365 0.736361 9.99958 2.98578e-06 1.1943e-05 0.133644 0.983358 0.931495 -0.0132918 4.92648e-06 0.513367 -1.99163e-20 7.38177e-24 -1.99089e-20 0.0013963 0.997815 8.60117e-05 0.152711 2.85266 0.0013963 0.997816 0.779457 0.0010652 0.00188119 0.000860117 0.455418 0.00188119 0.443722 0.000130903 1.02 0.888612 0.534419 0.287343 1.71908e-07 3.08101e-09 2373.14 3131.42 -0.0574208 0.482197 0.277314 0.254291 -0.593166 -0.169565 0.490112 -0.266089 -0.224033 2.518 1 0 296.049 0 2.21519 2.516 0.000299282 0.863148 0.694152 0.321839 0.431048 2.21538 138.113 83.7327 18.71 60.7758 0.00403305 0 -40 10
1.617 4.67869e-08 2.53971e-06 0.142401 0.1424 0.0120283 2.12668e-05 0.00115441 0.178001 0.000658733 0.178655 0.939022 101.526 0.236485 0.836109 4.47369 0.0635153 0.0422046 0.957795 0.0195103 0.00453747 0.0187692 0.00433389 0.0054897 0.00623084 0.219588 0.249234 58.0406 -87.8986 126.187 15.9401 145.033 0.000141952 0.267289 192.749 0.31025 0.0673322 0.00409807 0.000562288 0.0013848 0.986963 0.991718 -2.98809e-06 -85.6583 0.0930734 31172.1 308.537 0.9835 0.319146 0.736376 0.736372 9.99958 2.98579e-06 1.1943e-05 0.133649 0.983358 0.931494 -0.0132918 4.92651e-06 0.513385 -1.99177e-20 7.38236e-24 -1.99103e-20 0.0013963 0.997815 8.60118e-05 0.152711 2.85266 0.0013963 0.997816 0.779533 0.00106522 0.00188119 0.000860118 0.455418 0.00188119 0.443728 0.000130905 1.02 0.888613 0.534419 0.287345 1.71908e-07 3.08103e-09 2373.12 3131.47 -0.0574256 0.482197 0.277314 0.254294 -0.593166 -0.169565 0.490097 -0.266087 -0.22402 2.519 1 0 296.044 0 2.21533 2.517 0.000299281 0.863175 0.694195 0.321793 0.43107 2.21552 138.12 83.7322 18.71 60.7755 0.00403307 0 -40 10
1.618 4.68158e-08 2.53971e-06 0.142438 0.142437 0.0120283 2.12799e-05 0.00115442 0.178047 0.000658734 0.178701 0.93911 101.526 0.236474 0.836239 4.47425 0.0635259 0.0422099 0.95779 0.0195098 0.00453789 0.0187686 0.00433425 0.00549023 0.00623138 0.219609 0.249255 58.0407 -87.8986 126.186 15.9401 145.033 0.000141954 0.267289 192.749 0.31025 0.0673321 0.00409807 0.000562288 0.0013848 0.986963 0.991718 -2.9881e-06 -85.6583 0.0930735 31172 308.549 0.9835 0.319146 0.736388 0.736383 9.99958 2.98579e-06 1.19431e-05 0.133653 0.983359 0.931493 -0.0132918 4.92654e-06 0.513403 -1.99192e-20 7.38295e-24 -1.99118e-20 0.0013963 0.997815 8.60119e-05 0.152711 2.85266 0.0013963 0.997816 0.77961 0.00106524 0.00188119 0.000860119 0.455417 0.00188119 0.443733 0.000130908 1.02 0.888614 0.534419 0.287347 1.71908e-07 3.08106e-09 2373.11 3131.52 -0.0574304 0.482197 0.277314 0.254298 -0.593165 -0.169565 0.490082 -0.266084 -0.224007 2.52 1 0 296.04 0 2.21547 2.518 0.000299279 0.863201 0.694238 0.321747 0.431093 2.21565 138.127 83.7316 18.7099 60.7753 0.0040331 0 -40 10
1.619 4.68446e-08 2.53972e-06 0.142475 0.142474 0.0120283 2.1293e-05 0.00115442 0.178093 0.000658735 0.178747 0.939198 101.525 0.236464 0.83637 4.47482 0.0635364 0.0422152 0.957785 0.0195093 0.00453832 0.0187681 0.00433462 0.00549075 0.00623192 0.21963 0.249277 58.0408 -87.8986 126.186 15.9401 145.033 0.000141956 0.26729 192.749 0.310249 0.067332 0.00409808 0.000562289 0.0013848 0.986963 0.991718 -2.98812e-06 -85.6583 0.0930736 31172 308.56 0.9835 0.319146 0.736399 0.736394 9.99958 2.9858e-06 1.19431e-05 0.133657 0.983359 0.931492 -0.0132918 4.92657e-06 0.513422 -1.99207e-20 7.38355e-24 -1.99133e-20 0.0013963 0.997815 8.6012e-05 0.152711 2.85266 0.0013963 0.997816 0.779686 0.00106525 0.00188119 0.00086012 0.455417 0.00188119 0.443739 0.00013091 1.02 0.888615 0.534419 0.287348 1.71909e-07 3.08108e-09 2373.09 3131.56 -0.0574352 0.482197 0.277313 0.254301 -0.593164 -0.169565 0.490066 -0.266082 -0.223993 2.521 1 0 296.036 0 2.21561 2.519 0.000299278 0.863228 0.694282 0.321701 0.431115 2.21579 138.135 83.7311 18.7099 60.775 0.00403312 0 -40 10
1.62 4.68735e-08 2.53972e-06 0.142511 0.142511 0.0120283 2.13061e-05 0.00115442 0.178139 0.000658735 0.178794 0.939286 101.525 0.236453 0.8365 4.47538 0.0635469 0.0422206 0.957779 0.0195087 0.00453874 0.0187675 0.00433498 0.00549127 0.00623245 0.219651 0.249298 58.0408 -87.8986 126.186 15.94 145.033 0.000141959 0.26729 192.749 0.310249 0.067332 0.00409808 0.00056229 0.00138481 0.986963 0.991718 -2.98813e-06 -85.6583 0.0930737 31172 308.572 0.9835 0.319146 0.73641 0.736406 9.99958 2.9858e-06 1.19431e-05 0.133662 0.98336 0.931491 -0.0132918 4.9266e-06 0.51344 -1.99222e-20 7.38414e-24 -1.99148e-20 0.0013963 0.997815 8.60121e-05 0.152711 2.85267 0.0013963 0.997816 0.779763 0.00106527 0.00188119 0.000860121 0.455417 0.00188119 0.443744 0.000130913 1.02 0.888616 0.534418 0.28735 1.71909e-07 3.0811e-09 2373.08 3131.61 -0.05744 0.482198 0.277313 0.254304 -0.593164 -0.169565 0.490051 -0.26608 -0.22398 2.522 1 0 296.031 0 2.21575 2.52 0.000299277 0.863254 0.694325 0.321655 0.431138 2.21593 138.142 83.7305 18.7099 60.7747 0.00403314 0 -40 10
1.621 4.69023e-08 2.53972e-06 0.142548 0.142548 0.0120283 2.13192e-05 0.00115442 0.178185 0.000658736 0.178839 0.939374 101.524 0.236443 0.83663 4.47594 0.0635575 0.0422259 0.957774 0.0195082 0.00453917 0.018767 0.00433535 0.00549179 0.00623299 0.219672 0.24932 58.0409 -87.8986 126.186 15.94 145.033 0.000141961 0.26729 192.749 0.310249 0.0673319 0.00409808 0.00056229 0.00138481 0.986963 0.991718 -2.98815e-06 -85.6583 0.0930738 31172 308.583 0.9835 0.319146 0.736421 0.736417 9.99958 2.98581e-06 1.19431e-05 0.133666 0.98336 0.93149 -0.0132918 4.92663e-06 0.513458 -1.99236e-20 7.38473e-24 -1.99162e-20 0.00139631 0.997815 8.60122e-05 0.152712 2.85267 0.00139631 0.997816 0.779839 0.00106529 0.00188119 0.000860122 0.455417 0.00188119 0.44375 0.000130915 1.02 0.888617 0.534418 0.287351 1.71909e-07 3.08113e-09 2373.06 3131.66 -0.0574448 0.482198 0.277313 0.254307 -0.593163 -0.169565 0.490036 -0.266078 -0.223967 2.523 1 0 296.027 0 2.21589 2.521 0.000299276 0.863281 0.694369 0.32161 0.43116 2.21607 138.15 83.73 18.7099 60.7745 0.00403316 0 -40 10
1.622 4.69312e-08 2.53972e-06 0.142585 0.142584 0.0120282 2.13324e-05 0.00115442 0.178231 0.000658736 0.178885 0.939462 101.523 0.236432 0.836761 4.47651 0.063568 0.0422312 0.957769 0.0195077 0.00453959 0.0187665 0.00433571 0.00549232 0.00623352 0.219693 0.249341 58.041 -87.8987 126.186 15.9399 145.033 0.000141963 0.26729 192.748 0.310248 0.0673319 0.00409809 0.000562291 0.00138481 0.986963 0.991718 -2.98816e-06 -85.6583 0.0930739 31172 308.595 0.9835 0.319146 0.736432 0.736428 9.99958 2.98581e-06 1.19431e-05 0.13367 0.98336 0.93149 -0.0132918 4.92666e-06 0.513477 -1.99251e-20 7.38533e-24 -1.99177e-20 0.00139631 0.997815 8.60122e-05 0.152712 2.85267 0.00139631 0.997816 0.779916 0.0010653 0.0018812 0.000860122 0.455416 0.00188119 0.443755 0.000130918 1.02 0.888619 0.534418 0.287353 1.71909e-07 3.08115e-09 2373.04 3131.7 -0.0574497 0.482198 0.277312 0.25431 -0.593163 -0.169565 0.49002 -0.266076 -0.223954 2.524 1 0 296.023 0 2.21603 2.522 0.000299275 0.863307 0.694412 0.321564 0.431183 2.21621 138.157 83.7294 18.7098 60.7742 0.00403319 0 -40 10
1.623 4.69601e-08 2.53972e-06 0.142622 0.142621 0.0120282 2.13455e-05 0.00115442 0.178277 0.000658737 0.178931 0.93955 101.523 0.236421 0.836891 4.47707 0.0635785 0.0422365 0.957763 0.0195072 0.00454002 0.0187659 0.00433608 0.00549284 0.00623406 0.219714 0.249362 58.041 -87.8987 126.185 15.9399 145.033 0.000141965 0.26729 192.748 0.310248 0.0673318 0.00409809 0.000562292 0.00138481 0.986963 0.991718 -2.98818e-06 -85.6583 0.093074 31171.9 308.606 0.9835 0.319146 0.736444 0.736439 9.99958 2.98582e-06 1.19432e-05 0.133675 0.983361 0.931489 -0.0132918 4.92669e-06 0.513495 -1.99266e-20 7.38592e-24 -1.99192e-20 0.00139631 0.997815 8.60123e-05 0.152712 2.85267 0.00139631 0.997816 0.779992 0.00106532 0.0018812 0.000860123 0.455416 0.0018812 0.443761 0.00013092 1.02 0.88862 0.534417 0.287354 1.7191e-07 3.08117e-09 2373.03 3131.75 -0.0574545 0.482198 0.277312 0.254313 -0.593162 -0.169565 0.490005 -0.266074 -0.22394 2.525 1 0 296.018 0 2.21616 2.523 0.000299274 0.863334 0.694456 0.321518 0.431205 2.21635 138.165 83.7288 18.7098 60.7739 0.00403321 0 -40 10
1.624 4.69889e-08 2.53972e-06 0.142658 0.142658 0.0120282 2.13586e-05 0.00115442 0.178323 0.000658738 0.178977 0.939638 101.522 0.236411 0.837022 4.47764 0.0635891 0.0422418 0.957758 0.0195066 0.00454044 0.0187654 0.00433644 0.00549336 0.0062346 0.219735 0.249384 58.0411 -87.8987 126.185 15.9399 145.033 0.000141967 0.267291 192.748 0.310247 0.0673318 0.00409809 0.000562292 0.00138481 0.986963 0.991718 -2.98819e-06 -85.6582 0.093074 31171.9 308.618 0.9835 0.319146 0.736455 0.73645 9.99958 2.98582e-06 1.19432e-05 0.133679 0.983361 0.931488 -0.0132918 4.92672e-06 0.513514 -1.99281e-20 7.38651e-24 -1.99207e-20 0.00139631 0.997815 8.60124e-05 0.152712 2.85267 0.00139631 0.997816 0.780068 0.00106534 0.0018812 0.000860124 0.455416 0.0018812 0.443766 0.000130923 1.02 0.888621 0.534417 0.287356 1.7191e-07 3.08119e-09 2373.01 3131.8 -0.0574593 0.482198 0.277312 0.254316 -0.593161 -0.169565 0.48999 -0.266072 -0.223927 2.526 1 0 296.014 0 2.2163 2.524 0.000299273 0.863361 0.694499 0.321472 0.431228 2.21649 138.172 83.7283 18.7098 60.7737 0.00403323 0 -40 10
1.625 4.70178e-08 2.53972e-06 0.142695 0.142695 0.0120282 2.13717e-05 0.00115442 0.178369 0.000658738 0.179023 0.939726 101.522 0.2364 0.837152 4.4782 0.0635996 0.0422472 0.957753 0.0195061 0.00454087 0.0187649 0.00433681 0.00549389 0.00623514 0.219756 0.249405 58.0411 -87.8987 126.185 15.9398 145.033 0.000141969 0.267291 192.748 0.310247 0.0673317 0.0040981 0.000562293 0.00138482 0.986963 0.991718 -2.98821e-06 -85.6582 0.0930741 31171.9 308.629 0.9835 0.319146 0.736466 0.736462 9.99958 2.98583e-06 1.19432e-05 0.133683 0.983362 0.931487 -0.0132918 4.92675e-06 0.513532 -1.99296e-20 7.38711e-24 -1.99222e-20 0.00139631 0.997815 8.60125e-05 0.152712 2.85267 0.00139631 0.997816 0.780145 0.00106535 0.0018812 0.000860125 0.455416 0.0018812 0.443772 0.000130925 1.02 0.888622 0.534417 0.287357 1.7191e-07 3.08122e-09 2372.99 3131.85 -0.0574641 0.482198 0.277312 0.254319 -0.593161 -0.169565 0.489974 -0.26607 -0.223914 2.527 1 0 296.01 0 2.21644 2.525 0.000299272 0.863387 0.694543 0.321426 0.431251 2.21663 138.18 83.7277 18.7097 60.7734 0.00403326 0 -40 10
1.626 4.70466e-08 2.53973e-06 0.142732 0.142731 0.0120282 2.13848e-05 0.00115442 0.178415 0.000658739 0.179069 0.939814 101.521 0.23639 0.837283 4.47877 0.0636102 0.0422525 0.957747 0.0195056 0.00454129 0.0187643 0.00433718 0.00549441 0.00623567 0.219777 0.249427 58.0412 -87.8987 126.185 15.9398 145.033 0.000141972 0.267291 192.748 0.310246 0.0673317 0.0040981 0.000562294 0.00138482 0.986963 0.991718 -2.98822e-06 -85.6582 0.0930742 31171.9 308.641 0.9835 0.319146 0.736477 0.736473 9.99958 2.98583e-06 1.19432e-05 0.133688 0.983362 0.931486 -0.0132918 4.92678e-06 0.51355 -1.9931e-20 7.3877e-24 -1.99236e-20 0.00139631 0.997815 8.60126e-05 0.152712 2.85267 0.00139631 0.997816 0.780221 0.00106537 0.0018812 0.000860126 0.455415 0.0018812 0.443778 0.000130928 1.02 0.888623 0.534416 0.287359 1.7191e-07 3.08124e-09 2372.98 3131.89 -0.0574689 0.482198 0.277311 0.254322 -0.59316 -0.169565 0.489959 -0.266068 -0.223901 2.528 1 0 296.005 0 2.21658 2.526 0.000299271 0.863414 0.694586 0.321381 0.431273 2.21676 138.187 83.7272 18.7097 60.7731 0.00403328 0 -40 10
1.627 4.70755e-08 2.53973e-06 0.142768 0.142768 0.0120282 2.13979e-05 0.00115442 0.17846 0.00065874 0.179115 0.939902 101.521 0.236379 0.837413 4.47933 0.0636207 0.0422579 0.957742 0.0195051 0.00454172 0.0187638 0.00433754 0.00549494 0.00623621 0.219798 0.249448 58.0413 -87.8987 126.184 15.9398 145.033 0.000141974 0.267291 192.748 0.310246 0.0673316 0.0040981 0.000562294 0.00138482 0.986963 0.991718 -2.98824e-06 -85.6582 0.0930743 31171.8 308.652 0.9835 0.319146 0.736489 0.736484 9.99958 2.98584e-06 1.19432e-05 0.133692 0.983363 0.931485 -0.0132918 4.92681e-06 0.513569 -1.99325e-20 7.3883e-24 -1.99251e-20 0.00139631 0.997815 8.60126e-05 0.152713 2.85267 0.00139631 0.997816 0.780297 0.00106539 0.0018812 0.000860126 0.455415 0.0018812 0.443783 0.00013093 1.02 0.888624 0.534416 0.28736 1.71911e-07 3.08126e-09 2372.96 3131.94 -0.0574737 0.482198 0.277311 0.254325 -0.59316 -0.169565 0.489944 -0.266066 -0.223887 2.529 1 0 296.001 0 2.21672 2.527 0.00029927 0.863441 0.694629 0.321335 0.431296 2.2169 138.194 83.7266 18.7097 60.7729 0.0040333 0 -40 10
1.628 4.71043e-08 2.53973e-06 0.142805 0.142804 0.0120282 2.14111e-05 0.00115442 0.178506 0.00065874 0.17916 0.93999 101.52 0.236369 0.837544 4.4799 0.0636312 0.0422632 0.957737 0.0195045 0.00454214 0.0187633 0.00433791 0.00549546 0.00623675 0.219819 0.24947 58.0413 -87.8987 126.184 15.9397 145.033 0.000141976 0.267291 192.748 0.310246 0.0673316 0.00409811 0.000562295 0.00138482 0.986963 0.991718 -2.98825e-06 -85.6582 0.0930744 31171.8 308.664 0.9835 0.319146 0.7365 0.736495 9.99958 2.98584e-06 1.19433e-05 0.133696 0.983363 0.931484 -0.0132918 4.92684e-06 0.513587 -1.9934e-20 7.38889e-24 -1.99266e-20 0.00139631 0.997815 8.60127e-05 0.152713 2.85267 0.00139631 0.997816 0.780373 0.0010654 0.0018812 0.000860127 0.455415 0.0018812 0.443789 0.000130933 1.02 0.888625 0.534416 0.287362 1.71911e-07 3.08129e-09 2372.94 3131.99 -0.0574786 0.482198 0.277311 0.254328 -0.593159 -0.169565 0.489928 -0.266063 -0.223874 2.53 1 0 295.997 0 2.21686 2.528 0.000299268 0.863468 0.694673 0.321289 0.431318 2.21704 138.202 83.7261 18.7096 60.7726 0.00403333 0 -40 10
1.629 4.71332e-08 2.53973e-06 0.142841 0.142841 0.0120282 2.14242e-05 0.00115442 0.178552 0.000658741 0.179206 0.940078 101.52 0.236358 0.837674 4.48047 0.0636418 0.0422685 0.957731 0.019504 0.00454257 0.0187627 0.00433828 0.00549599 0.00623729 0.21984 0.249492 58.0414 -87.8987 126.184 15.9397 145.033 0.000141978 0.267291 192.747 0.310245 0.0673315 0.00409811 0.000562296 0.00138482 0.986963 0.991718 -2.98827e-06 -85.6582 0.0930745 31171.8 308.676 0.9835 0.319146 0.736511 0.736507 9.99958 2.98585e-06 1.19433e-05 0.133701 0.983364 0.931483 -0.0132918 4.92687e-06 0.513606 -1.99355e-20 7.38949e-24 -1.99281e-20 0.00139631 0.997815 8.60128e-05 0.152713 2.85267 0.00139631 0.997816 0.78045 0.00106542 0.00188121 0.000860128 0.455415 0.0018812 0.443794 0.000130935 1.02 0.888626 0.534415 0.287363 1.71911e-07 3.08131e-09 2372.93 3132.03 -0.0574834 0.482198 0.27731 0.254331 -0.593158 -0.169566 0.489913 -0.266061 -0.223861 2.531 1 0 295.992 0 2.217 2.529 0.000299267 0.863494 0.694716 0.321244 0.431341 2.21718 138.209 83.7255 18.7096 60.7723 0.00403335 0 -40 10
1.63 4.7162e-08 2.53973e-06 0.142878 0.142877 0.0120281 2.14373e-05 0.00115442 0.178598 0.000658741 0.179252 0.940166 101.519 0.236348 0.837805 4.48103 0.0636523 0.0422739 0.957726 0.0195035 0.004543 0.0187622 0.00433864 0.00549651 0.00623783 0.219861 0.249513 58.0415 -87.8987 126.184 15.9396 145.033 0.00014198 0.267292 192.747 0.310245 0.0673315 0.00409811 0.000562296 0.00138483 0.986963 0.991718 -2.98828e-06 -85.6582 0.0930746 31171.8 308.687 0.9835 0.319146 0.736522 0.736518 9.99958 2.98585e-06 1.19433e-05 0.133705 0.983364 0.931482 -0.0132918 4.92689e-06 0.513624 -1.9937e-20 7.39008e-24 -1.99296e-20 0.00139632 0.997815 8.60129e-05 0.152713 2.85267 0.00139632 0.997816 0.780526 0.00106544 0.00188121 0.000860129 0.455415 0.00188121 0.4438 0.000130938 1.02 0.888627 0.534415 0.287365 1.71912e-07 3.08133e-09 2372.91 3132.08 -0.0574882 0.482198 0.27731 0.254334 -0.593158 -0.169566 0.489897 -0.266059 -0.223848 2.532 1 0 295.988 0 2.21713 2.53 0.000299266 0.863521 0.69476 0.321198 0.431363 2.21732 138.217 83.725 18.7096 60.7721 0.00403337 0 -40 10
1.631 4.71909e-08 2.53973e-06 0.142915 0.142914 0.0120281 2.14504e-05 0.00115442 0.178643 0.000658742 0.179297 0.940254 101.518 0.236337 0.837935 4.4816 0.0636629 0.0422793 0.957721 0.019503 0.00454342 0.0187616 0.00433901 0.00549704 0.00623837 0.219882 0.249535 58.0415 -87.8987 126.184 15.9396 145.033 0.000141982 0.267292 192.747 0.310244 0.0673314 0.00409811 0.000562297 0.00138483 0.986963 0.991718 -2.9883e-06 -85.6582 0.0930747 31171.8 308.699 0.9835 0.319146 0.736534 0.736529 9.99958 2.98586e-06 1.19433e-05 0.133709 0.983364 0.931481 -0.0132918 4.92692e-06 0.513643 -1.99385e-20 7.39068e-24 -1.99311e-20 0.00139632 0.997815 8.6013e-05 0.152713 2.85268 0.00139632 0.997816 0.780602 0.00106545 0.00188121 0.00086013 0.455414 0.00188121 0.443805 0.00013094 1.02 0.888628 0.534415 0.287366 1.71912e-07 3.08135e-09 2372.89 3132.13 -0.057493 0.482198 0.27731 0.254337 -0.593157 -0.169566 0.489882 -0.266057 -0.223834 2.533 1 0 295.984 0 2.21727 2.531 0.000299265 0.863548 0.694803 0.321153 0.431386 2.21746 138.224 83.7244 18.7095 60.7718 0.00403339 0 -40 10
1.632 4.72198e-08 2.53973e-06 0.142951 0.14295 0.0120281 2.14635e-05 0.00115442 0.178689 0.000658743 0.179343 0.940342 101.518 0.236327 0.838066 4.48217 0.0636735 0.0422846 0.957715 0.0195024 0.00454385 0.0187611 0.00433938 0.00549757 0.00623891 0.219903 0.249556 58.0416 -87.8987 126.183 15.9396 145.033 0.000141985 0.267292 192.747 0.310244 0.0673314 0.00409812 0.000562298 0.00138483 0.986963 0.991718 -2.98831e-06 -85.6582 0.0930747 31171.7 308.71 0.9835 0.319146 0.736545 0.736541 9.99958 2.98586e-06 1.19433e-05 0.133714 0.983365 0.931481 -0.0132918 4.92695e-06 0.513661 -1.99399e-20 7.39127e-24 -1.99325e-20 0.00139632 0.997815 8.6013e-05 0.152713 2.85268 0.00139632 0.997816 0.780678 0.00106547 0.00188121 0.00086013 0.455414 0.00188121 0.443811 0.000130943 1.02 0.888629 0.534415 0.287368 1.71912e-07 3.08138e-09 2372.88 3132.18 -0.0574979 0.482198 0.27731 0.25434 -0.593157 -0.169566 0.489867 -0.266055 -0.223821 2.534 1 0 295.979 0 2.21741 2.532 0.000299264 0.863575 0.694846 0.321107 0.431408 2.21759 138.232 83.7238 18.7095 60.7715 0.00403342 0 -40 10
1.633 4.72486e-08 2.53974e-06 0.142987 0.142987 0.0120281 2.14766e-05 0.00115443 0.178734 0.000658743 0.179388 0.94043 101.517 0.236316 0.838196 4.48274 0.063684 0.04229 0.95771 0.0195019 0.00454428 0.0187606 0.00433975 0.00549809 0.00623945 0.219924 0.249578 58.0416 -87.8987 126.183 15.9395 145.033 0.000141987 0.267292 192.747 0.310243 0.0673313 0.00409812 0.000562298 0.00138483 0.986963 0.991718 -2.98833e-06 -85.6582 0.0930748 31171.7 308.722 0.9835 0.319146 0.736556 0.736552 9.99958 2.98587e-06 1.19434e-05 0.133718 0.983365 0.93148 -0.0132918 4.92698e-06 0.51368 -1.99414e-20 7.39187e-24 -1.9934e-20 0.00139632 0.997815 8.60131e-05 0.152713 2.85268 0.00139632 0.997816 0.780754 0.00106549 0.00188121 0.000860131 0.455414 0.00188121 0.443816 0.000130945 1.02 0.888631 0.534414 0.287369 1.71912e-07 3.0814e-09 2372.86 3132.22 -0.0575027 0.482199 0.277309 0.254343 -0.593156 -0.169566 0.489851 -0.266053 -0.223808 2.535 1 0 295.975 0 2.21755 2.533 0.000299263 0.863601 0.69489 0.321062 0.431431 2.21773 138.239 83.7233 18.7095 60.7713 0.00403344 0 -40 10
1.634 4.72775e-08 2.53974e-06 0.143024 0.143023 0.0120281 2.14898e-05 0.00115443 0.17878 0.000658744 0.179434 0.940519 101.517 0.236305 0.838327 4.48331 0.0636946 0.0422954 0.957705 0.0195014 0.00454471 0.01876 0.00434012 0.00549862 0.00623999 0.219945 0.249599 58.0417 -87.8987 126.183 15.9395 145.033 0.000141989 0.267292 192.747 0.310243 0.0673313 0.00409812 0.000562299 0.00138484 0.986963 0.991718 -2.98834e-06 -85.6582 0.0930749 31171.7 308.734 0.9835 0.319146 0.736568 0.736563 9.99958 2.98587e-06 1.19434e-05 0.133722 0.983366 0.931479 -0.0132918 4.92701e-06 0.513698 -1.99429e-20 7.39247e-24 -1.99355e-20 0.00139632 0.997815 8.60132e-05 0.152714 2.85268 0.00139632 0.997816 0.78083 0.0010655 0.00188121 0.000860132 0.455414 0.00188121 0.443822 0.000130948 1.02 0.888632 0.534414 0.287371 1.71913e-07 3.08142e-09 2372.85 3132.27 -0.0575075 0.482199 0.277309 0.254346 -0.593155 -0.169566 0.489836 -0.266051 -0.223794 2.536 1 0 295.97 0 2.21769 2.534 0.000299262 0.863628 0.694933 0.321017 0.431453 2.21787 138.246 83.7227 18.7094 60.771 0.00403346 0 -40 10
1.635 4.73063e-08 2.53974e-06 0.14306 0.14306 0.0120281 2.15029e-05 0.00115443 0.178825 0.000658745 0.179479 0.940607 101.516 0.236295 0.838458 4.48388 0.0637051 0.0423007 0.957699 0.0195009 0.00454513 0.0187595 0.00434048 0.00549915 0.00624053 0.219966 0.249621 58.0418 -87.8987 126.183 15.9395 145.033 0.000141991 0.267293 192.746 0.310243 0.0673312 0.00409813 0.0005623 0.00138484 0.986963 0.991718 -2.98836e-06 -85.6581 0.093075 31171.7 308.745 0.9835 0.319146 0.736579 0.736574 9.99958 2.98588e-06 1.19434e-05 0.133727 0.983366 0.931478 -0.0132918 4.92704e-06 0.513717 -1.99444e-20 7.39306e-24 -1.9937e-20 0.00139632 0.997815 8.60133e-05 0.152714 2.85268 0.00139632 0.997816 0.780906 0.00106552 0.00188122 0.000860133 0.455413 0.00188121 0.443827 0.00013095 1.02 0.888633 0.534414 0.287372 1.71913e-07 3.08145e-09 2372.83 3132.32 -0.0575124 0.482199 0.277309 0.254349 -0.593155 -0.169566 0.48982 -0.266049 -0.223781 2.537 1 0 295.966 0 2.21783 2.535 0.000299261 0.863655 0.694977 0.320971 0.431476 2.21801 138.254 83.7222 18.7094 60.7707 0.00403349 0 -40 10
1.636 4.73352e-08 2.53974e-06 0.143097 0.143096 0.0120281 2.1516e-05 0.00115443 0.178871 0.000658745 0.179525 0.940695 101.516 0.236284 0.838588 4.48445 0.0637157 0.0423061 0.957694 0.0195003 0.00454556 0.0187589 0.00434085 0.00549967 0.00624107 0.219987 0.249643 58.0418 -87.8987 126.183 15.9394 145.033 0.000141993 0.267293 192.746 0.310242 0.0673312 0.00409813 0.000562301 0.00138484 0.986963 0.991718 -2.98837e-06 -85.6581 0.0930751 31171.6 308.757 0.9835 0.319146 0.73659 0.736586 9.99958 2.98588e-06 1.19434e-05 0.133731 0.983366 0.931477 -0.0132918 4.92707e-06 0.513735 -1.99459e-20 7.39366e-24 -1.99385e-20 0.00139632 0.997815 8.60134e-05 0.152714 2.85268 0.00139632 0.997816 0.780982 0.00106554 0.00188122 0.000860134 0.455413 0.00188122 0.443833 0.000130953 1.02 0.888634 0.534413 0.287374 1.71913e-07 3.08147e-09 2372.81 3132.37 -0.0575172 0.482199 0.277309 0.254352 -0.593154 -0.169566 0.489805 -0.266047 -0.223768 2.538 1 0 295.962 0 2.21797 2.536 0.00029926 0.863682 0.69502 0.320926 0.431498 2.21815 138.261 83.7216 18.7094 60.7705 0.00403351 0 -40 10
1.637 4.7364e-08 2.53974e-06 0.143133 0.143132 0.012028 2.15291e-05 0.00115443 0.178916 0.000658746 0.17957 0.940783 101.515 0.236274 0.838719 4.48502 0.0637262 0.0423115 0.957689 0.0194998 0.00454599 0.0187584 0.00434122 0.0055002 0.00624161 0.220008 0.249664 58.0419 -87.8987 126.182 15.9394 145.033 0.000141995 0.267293 192.746 0.310242 0.0673311 0.00409813 0.000562301 0.00138484 0.986963 0.991718 -2.98839e-06 -85.6581 0.0930752 31171.6 308.769 0.9835 0.319146 0.736601 0.736597 9.99958 2.98589e-06 1.19434e-05 0.133735 0.983367 0.931476 -0.0132918 4.9271e-06 0.513754 -1.99474e-20 7.39426e-24 -1.994e-20 0.00139632 0.997815 8.60134e-05 0.152714 2.85268 0.00139632 0.997816 0.781058 0.00106555 0.00188122 0.000860134 0.455413 0.00188122 0.443838 0.000130955 1.02 0.888635 0.534413 0.287375 1.71913e-07 3.08149e-09 2372.8 3132.41 -0.057522 0.482199 0.277308 0.254355 -0.593154 -0.169566 0.48979 -0.266045 -0.223754 2.539 1 0 295.957 0 2.2181 2.537 0.000299259 0.863709 0.695063 0.320881 0.431521 2.21829 138.269 83.7211 18.7093 60.7702 0.00403353 0 -40 10
1.638 4.73929e-08 2.53974e-06 0.143169 0.143169 0.012028 2.15422e-05 0.00115443 0.178961 0.000658746 0.179616 0.940871 101.514 0.236263 0.83885 4.48559 0.0637368 0.0423169 0.957683 0.0194993 0.00454642 0.0187579 0.00434159 0.00550073 0.00624215 0.220029 0.249686 58.042 -87.8987 126.182 15.9393 145.034 0.000141998 0.267293 192.746 0.310241 0.067331 0.00409814 0.000562302 0.00138484 0.986963 0.991718 -2.9884e-06 -85.6581 0.0930753 31171.6 308.78 0.9835 0.319146 0.736613 0.736608 9.99958 2.98589e-06 1.19435e-05 0.13374 0.983367 0.931475 -0.0132918 4.92713e-06 0.513772 -1.99489e-20 7.39486e-24 -1.99415e-20 0.00139632 0.997815 8.60135e-05 0.152714 2.85268 0.00139632 0.997816 0.781134 0.00106557 0.00188122 0.000860135 0.455413 0.00188122 0.443844 0.000130958 1.02 0.888636 0.534413 0.287377 1.71914e-07 3.08152e-09 2372.78 3132.46 -0.0575269 0.482199 0.277308 0.254358 -0.593153 -0.169566 0.489774 -0.266042 -0.223741 2.54 1 0 295.953 0 2.21824 2.538 0.000299257 0.863736 0.695107 0.320836 0.431543 2.21843 138.276 83.7205 18.7093 60.7699 0.00403356 0 -40 10
1.639 4.74217e-08 2.53974e-06 0.143205 0.143205 0.012028 2.15553e-05 0.00115443 0.179007 0.000658747 0.179661 0.94096 101.514 0.236253 0.83898 4.48616 0.0637474 0.0423223 0.957678 0.0194987 0.00454685 0.0187573 0.00434196 0.00550126 0.00624269 0.22005 0.249708 58.042 -87.8987 126.182 15.9393 145.034 0.000142 0.267293 192.746 0.310241 0.067331 0.00409814 0.000562303 0.00138485 0.986963 0.991718 -2.98842e-06 -85.6581 0.0930754 31171.6 308.792 0.9835 0.319146 0.736624 0.73662 9.99958 2.9859e-06 1.19435e-05 0.133744 0.983368 0.931474 -0.0132918 4.92716e-06 0.513791 -1.99504e-20 7.39545e-24 -1.9943e-20 0.00139633 0.997815 8.60136e-05 0.152714 2.85268 0.00139633 0.997816 0.78121 0.00106559 0.00188122 0.000860136 0.455413 0.00188122 0.443849 0.00013096 1.02 0.888637 0.534412 0.287378 1.71914e-07 3.08154e-09 2372.76 3132.51 -0.0575317 0.482199 0.277308 0.254361 -0.593152 -0.169566 0.489759 -0.26604 -0.223728 2.541 1 0 295.949 0 2.21838 2.539 0.000299256 0.863763 0.69515 0.320791 0.431566 2.21856 138.284 83.7199 18.7093 60.7697 0.00403358 0 -40 10
1.64 4.74506e-08 2.53975e-06 0.143242 0.143241 0.012028 2.15685e-05 0.00115443 0.179052 0.000658748 0.179706 0.941048 101.513 0.236242 0.839111 4.48673 0.0637579 0.0423277 0.957672 0.0194982 0.00454727 0.0187568 0.00434233 0.00550178 0.00624323 0.220071 0.249729 58.0421 -87.8987 126.182 15.9393 145.034 0.000142002 0.267294 192.746 0.31024 0.0673309 0.00409814 0.000562303 0.00138485 0.986963 0.991718 -2.98843e-06 -85.6581 0.0930754 31171.5 308.803 0.9835 0.319146 0.736635 0.736631 9.99958 2.9859e-06 1.19435e-05 0.133749 0.983368 0.931473 -0.0132918 4.92719e-06 0.513809 -1.99519e-20 7.39605e-24 -1.99445e-20 0.00139633 0.997815 8.60137e-05 0.152715 2.85268 0.00139633 0.997816 0.781286 0.0010656 0.00188122 0.000860137 0.455412 0.00188122 0.443855 0.000130963 1.02 0.888638 0.534412 0.28738 1.71914e-07 3.08156e-09 2372.75 3132.55 -0.0575366 0.482199 0.277307 0.254364 -0.593152 -0.169566 0.489743 -0.266038 -0.223714 2.542 1 0 295.944 0 2.21852 2.54 0.000299255 0.863789 0.695193 0.320746 0.431588 2.2187 138.291 83.7194 18.7092 60.7694 0.0040336 0 -40 10
1.641 4.74794e-08 2.53975e-06 0.143278 0.143277 0.012028 2.15816e-05 0.00115443 0.179097 0.000658748 0.179751 0.941136 101.513 0.236231 0.839242 4.48731 0.0637685 0.0423331 0.957667 0.0194977 0.0045477 0.0187562 0.0043427 0.00550231 0.00624378 0.220093 0.249751 58.0421 -87.8987 126.182 15.9392 145.034 0.000142004 0.267294 192.745 0.31024 0.0673309 0.00409814 0.000562304 0.00138485 0.986963 0.991718 -2.98845e-06 -85.6581 0.0930755 31171.5 308.815 0.9835 0.319146 0.736647 0.736642 9.99958 2.98591e-06 1.19435e-05 0.133753 0.983369 0.931472 -0.0132918 4.92722e-06 0.513828 -1.99533e-20 7.39665e-24 -1.99459e-20 0.00139633 0.997815 8.60138e-05 0.152715 2.85268 0.00139633 0.997816 0.781362 0.00106562 0.00188122 0.000860138 0.455412 0.00188122 0.44386 0.000130965 1.02 0.888639 0.534412 0.287382 1.71915e-07 3.08158e-09 2372.73 3132.6 -0.0575414 0.482199 0.277307 0.254367 -0.593151 -0.169566 0.489728 -0.266036 -0.223701 2.543 1 0 295.94 0 2.21866 2.541 0.000299254 0.863816 0.695237 0.320701 0.431611 2.21884 138.298 83.7188 18.7092 60.7691 0.00403362 0 -40 10
1.642 4.75083e-08 2.53975e-06 0.143314 0.143313 0.012028 2.15947e-05 0.00115443 0.179142 0.000658749 0.179797 0.941225 101.512 0.236221 0.839373 4.48788 0.0637791 0.0423385 0.957662 0.0194972 0.00454813 0.0187557 0.00434307 0.00550284 0.00624432 0.220114 0.249773 58.0422 -87.8987 126.181 15.9392 145.034 0.000142006 0.267294 192.745 0.31024 0.0673308 0.00409815 0.000562305 0.00138485 0.986963 0.991718 -2.98846e-06 -85.6581 0.0930756 31171.5 308.827 0.9835 0.319146 0.736658 0.736654 9.99958 2.98591e-06 1.19435e-05 0.133757 0.983369 0.931471 -0.0132918 4.92725e-06 0.513847 -1.99548e-20 7.39725e-24 -1.99474e-20 0.00139633 0.997815 8.60138e-05 0.152715 2.85269 0.00139633 0.997816 0.781438 0.00106564 0.00188123 0.000860138 0.455412 0.00188122 0.443866 0.000130968 1.02 0.88864 0.534411 0.287383 1.71915e-07 3.08161e-09 2372.71 3132.65 -0.0575463 0.482199 0.277307 0.25437 -0.593151 -0.169566 0.489712 -0.266034 -0.223688 2.544 1 0 295.936 0 2.2188 2.542 0.000299253 0.863843 0.69528 0.320656 0.431633 2.21898 138.306 83.7183 18.7092 60.7689 0.00403365 0 -40 10
1.643 4.75372e-08 2.53975e-06 0.14335 0.143349 0.012028 2.16078e-05 0.00115443 0.179188 0.000658749 0.179842 0.941313 101.512 0.23621 0.839504 4.48845 0.0637897 0.0423439 0.957656 0.0194966 0.00454856 0.0187551 0.00434344 0.00550337 0.00624486 0.220135 0.249794 58.0423 -87.8987 126.181 15.9392 145.034 0.000142009 0.267294 192.745 0.310239 0.0673308 0.00409815 0.000562305 0.00138486 0.986963 0.991718 -2.98848e-06 -85.6581 0.0930757 31171.5 308.838 0.9835 0.319146 0.736669 0.736665 9.99958 2.98592e-06 1.19436e-05 0.133762 0.983369 0.93147 -0.0132918 4.92728e-06 0.513865 -1.99563e-20 7.39785e-24 -1.99489e-20 0.00139633 0.997815 8.60139e-05 0.152715 2.85269 0.00139633 0.997816 0.781514 0.00106565 0.00188123 0.000860139 0.455412 0.00188123 0.443871 0.00013097 1.02 0.888642 0.534411 0.287385 1.71915e-07 3.08163e-09 2372.7 3132.7 -0.0575511 0.482199 0.277307 0.254373 -0.59315 -0.169566 0.489697 -0.266032 -0.223674 2.545 1 0 295.931 0 2.21893 2.543 0.000299252 0.86387 0.695324 0.320611 0.431656 2.21912 138.313 83.7177 18.7091 60.7686 0.00403367 0 -40 10
1.644 4.7566e-08 2.53975e-06 0.143386 0.143386 0.0120279 2.16209e-05 0.00115443 0.179233 0.00065875 0.179887 0.941401 101.511 0.2362 0.839634 4.48903 0.0638002 0.0423493 0.957651 0.0194961 0.00454899 0.0187546 0.00434381 0.0055039 0.0062454 0.220156 0.249816 58.0423 -87.8987 126.181 15.9391 145.034 0.000142011 0.267294 192.745 0.310239 0.0673307 0.00409815 0.000562306 0.00138486 0.986963 0.991718 -2.98849e-06 -85.6581 0.0930758 31171.5 308.85 0.9835 0.319146 0.736681 0.736676 9.99958 2.98592e-06 1.19436e-05 0.133766 0.98337 0.93147 -0.0132918 4.92731e-06 0.513884 -1.99578e-20 7.39845e-24 -1.99504e-20 0.00139633 0.997815 8.6014e-05 0.152715 2.85269 0.00139633 0.997816 0.78159 0.00106567 0.00188123 0.00086014 0.455411 0.00188123 0.443877 0.000130973 1.02 0.888643 0.534411 0.287386 1.71915e-07 3.08165e-09 2372.68 3132.74 -0.057556 0.482199 0.277306 0.254376 -0.593149 -0.169566 0.489681 -0.26603 -0.223661 2.546 1 0 295.927 0 2.21907 2.544 0.000299251 0.863897 0.695367 0.320566 0.431678 2.21926 138.321 83.7171 18.7091 60.7683 0.00403369 0 -40 10
1.645 4.75949e-08 2.53975e-06 0.143422 0.143422 0.0120279 2.1634e-05 0.00115443 0.179278 0.000658751 0.179932 0.94149 101.51 0.236189 0.839765 4.4896 0.0638108 0.0423547 0.957645 0.0194956 0.00454942 0.0187541 0.00434418 0.00550443 0.00624595 0.220177 0.249838 58.0424 -87.8987 126.181 15.9391 145.034 0.000142013 0.267295 192.745 0.310238 0.0673307 0.00409816 0.000562307 0.00138486 0.986963 0.991718 -2.98851e-06 -85.658 0.0930759 31171.4 308.862 0.9835 0.319146 0.736692 0.736688 9.99958 2.98593e-06 1.19436e-05 0.13377 0.98337 0.931469 -0.0132918 4.92734e-06 0.513902 -1.99593e-20 7.39905e-24 -1.99519e-20 0.00139633 0.997815 8.60141e-05 0.152715 2.85269 0.00139633 0.997816 0.781665 0.00106569 0.00188123 0.000860141 0.455411 0.00188123 0.443882 0.000130975 1.02 0.888644 0.534411 0.287388 1.71916e-07 3.08168e-09 2372.66 3132.79 -0.0575608 0.482199 0.277306 0.254379 -0.593149 -0.169567 0.489666 -0.266028 -0.223648 2.547 1 0 295.922 0 2.21921 2.545 0.00029925 0.863924 0.69541 0.320521 0.431701 2.21939 138.328 83.7166 18.7091 60.768 0.00403372 0 -40 10
1.646 4.76237e-08 2.53975e-06 0.143458 0.143458 0.0120279 2.16471e-05 0.00115443 0.179323 0.000658751 0.179977 0.941578 101.51 0.236179 0.839896 4.49018 0.0638214 0.0423601 0.95764 0.019495 0.00454985 0.0187535 0.00434455 0.00550496 0.00624649 0.220198 0.24986 58.0425 -87.8987 126.181 15.939 145.034 0.000142015 0.267295 192.745 0.310238 0.0673306 0.00409816 0.000562307 0.00138486 0.986963 0.991718 -2.98852e-06 -85.658 0.093076 31171.4 308.873 0.9835 0.319146 0.736704 0.736699 9.99958 2.98593e-06 1.19436e-05 0.133775 0.983371 0.931468 -0.0132918 4.92737e-06 0.513921 -1.99608e-20 7.39965e-24 -1.99534e-20 0.00139633 0.997815 8.60142e-05 0.152715 2.85269 0.00139633 0.997816 0.781741 0.0010657 0.00188123 0.000860142 0.455411 0.00188123 0.443888 0.000130978 1.02 0.888645 0.53441 0.287389 1.71916e-07 3.0817e-09 2372.65 3132.84 -0.0575657 0.4822 0.277306 0.254383 -0.593148 -0.169567 0.489651 -0.266026 -0.223634 2.548 1 0 295.918 0 2.21935 2.546 0.000299249 0.863951 0.695454 0.320476 0.431723 2.21953 138.336 83.716 18.709 60.7678 0.00403374 0 -40 10
1.647 4.76526e-08 2.53976e-06 0.143494 0.143494 0.0120279 2.16603e-05 0.00115443 0.179368 0.000658752 0.180022 0.941666 101.509 0.236168 0.840027 4.49075 0.063832 0.0423656 0.957634 0.0194945 0.00455028 0.018753 0.00434492 0.00550549 0.00624704 0.22022 0.249881 58.0425 -87.8987 126.18 15.939 145.034 0.000142017 0.267295 192.744 0.310237 0.0673306 0.00409816 0.000562308 0.00138486 0.986963 0.991718 -2.98854e-06 -85.658 0.0930761 31171.4 308.885 0.9835 0.319146 0.736715 0.736711 9.99958 2.98594e-06 1.19436e-05 0.133779 0.983371 0.931467 -0.0132918 4.9274e-06 0.51394 -1.99623e-20 7.40025e-24 -1.99549e-20 0.00139634 0.997815 8.60143e-05 0.152716 2.85269 0.00139634 0.997816 0.781817 0.00106572 0.00188123 0.000860143 0.455411 0.00188123 0.443893 0.00013098 1.02 0.888646 0.53441 0.287391 1.71916e-07 3.08172e-09 2372.63 3132.89 -0.0575705 0.4822 0.277305 0.254386 -0.593148 -0.169567 0.489635 -0.266024 -0.223621 2.549 1 0 295.914 0 2.21949 2.547 0.000299247 0.863978 0.695497 0.320431 0.431746 2.21967 138.343 83.7155 18.709 60.7675 0.00403376 0 -40 10
1.648 4.76814e-08 2.53976e-06 0.14353 0.14353 0.0120279 2.16734e-05 0.00115444 0.179413 0.000658752 0.180067 0.941755 101.509 0.236157 0.840158 4.49133 0.0638425 0.042371 0.957629 0.019494 0.00455071 0.0187524 0.00434529 0.00550602 0.00624758 0.220241 0.249903 58.0426 -87.8987 126.18 15.939 145.034 0.00014202 0.267295 192.744 0.310237 0.0673305 0.00409817 0.000562309 0.00138487 0.986963 0.991718 -2.98855e-06 -85.658 0.0930761 31171.4 308.897 0.9835 0.319146 0.736726 0.736722 9.99958 2.98594e-06 1.19437e-05 0.133784 0.983371 0.931466 -0.0132918 4.92743e-06 0.513958 -1.99638e-20 7.40085e-24 -1.99564e-20 0.00139634 0.997815 8.60143e-05 0.152716 2.85269 0.00139634 0.997816 0.781893 0.00106574 0.00188123 0.000860143 0.45541 0.00188123 0.443899 0.000130983 1.02 0.888647 0.53441 0.287392 1.71916e-07 3.08174e-09 2372.62 3132.94 -0.0575754 0.4822 0.277305 0.254389 -0.593147 -0.169567 0.48962 -0.266021 -0.223608 2.55 1 0 295.909 0 2.21963 2.548 0.000299246 0.864005 0.69554 0.320386 0.431768 2.21981 138.35 83.7149 18.709 60.7672 0.00403379 0 -40 10
1.649 4.77103e-08 2.53976e-06 0.143566 0.143566 0.0120279 2.16865e-05 0.00115444 0.179458 0.000658753 0.180112 0.941843 101.508 0.236147 0.840289 4.4919 0.0638531 0.0423764 0.957624 0.0194934 0.00455114 0.0187519 0.00434566 0.00550655 0.00624812 0.220262 0.249925 58.0427 -87.8988 126.18 15.9389 145.034 0.000142022 0.267295 192.744 0.310237 0.0673305 0.00409817 0.000562309 0.00138487 0.986962 0.991718 -2.98857e-06 -85.658 0.0930762 31171.3 308.909 0.9835 0.319146 0.736738 0.736733 9.99958 2.98595e-06 1.19437e-05 0.133788 0.983372 0.931465 -0.0132918 4.92746e-06 0.513977 -1.99653e-20 7.40145e-24 -1.99579e-20 0.00139634 0.997815 8.60144e-05 0.152716 2.85269 0.00139634 0.997816 0.781968 0.00106575 0.00188124 0.000860144 0.45541 0.00188123 0.443904 0.000130985 1.02 0.888648 0.534409 0.287394 1.71917e-07 3.08177e-09 2372.6 3132.98 -0.0575802 0.4822 0.277305 0.254392 -0.593146 -0.169567 0.489604 -0.266019 -0.223594 2.551 1 0 295.905 0 2.21977 2.549 0.000299245 0.864032 0.695584 0.320342 0.431791 2.21995 138.358 83.7143 18.7089 60.767 0.00403381 0 -40 10
1.65 4.77391e-08 2.53976e-06 0.143602 0.143602 0.0120279 2.16996e-05 0.00115444 0.179503 0.000658754 0.180157 0.941932 101.508 0.236136 0.84042 4.49248 0.0638637 0.0423819 0.957618 0.0194929 0.00455158 0.0187513 0.00434603 0.00550708 0.00624867 0.220283 0.249947 58.0427 -87.8988 126.18 15.9389 145.034 0.000142024 0.267296 192.744 0.310236 0.0673304 0.00409817 0.00056231 0.00138487 0.986962 0.991718 -2.98858e-06 -85.658 0.0930763 31171.3 308.92 0.9835 0.319146 0.736749 0.736745 9.99958 2.98595e-06 1.19437e-05 0.133792 0.983372 0.931464 -0.0132918 4.92749e-06 0.513996 -1.99668e-20 7.40205e-24 -1.99594e-20 0.00139634 0.997815 8.60145e-05 0.152716 2.85269 0.00139634 0.997816 0.782044 0.00106577 0.00188124 0.000860145 0.45541 0.00188124 0.44391 0.000130988 1.02 0.888649 0.534409 0.287395 1.71917e-07 3.08179e-09 2372.58 3133.03 -0.0575851 0.4822 0.277305 0.254395 -0.593146 -0.169567 0.489589 -0.266017 -0.223581 2.552 1 0 295.901 0 2.2199 2.55 0.000299244 0.864059 0.695627 0.320297 0.431813 2.22009 138.365 83.7138 18.7089 60.7667 0.00403383 0 -40 10
1.651 4.7768e-08 2.53976e-06 0.143638 0.143638 0.0120278 2.17127e-05 0.00115444 0.179548 0.000658754 0.180202 0.94202 101.507 0.236126 0.840551 4.49306 0.0638743 0.0423873 0.957613 0.0194924 0.00455201 0.0187508 0.0043464 0.00550761 0.00624921 0.220305 0.249969 58.0428 -87.8988 126.18 15.9389 145.034 0.000142026 0.267296 192.744 0.310236 0.0673304 0.00409818 0.000562311 0.00138487 0.986962 0.991718 -2.9886e-06 -85.658 0.0930764 31171.3 308.932 0.9835 0.319146 0.73676 0.736756 9.99958 2.98596e-06 1.19437e-05 0.133797 0.983373 0.931463 -0.0132917 4.92752e-06 0.514014 -1.99683e-20 7.40265e-24 -1.99609e-20 0.00139634 0.997815 8.60146e-05 0.152716 2.85269 0.00139634 0.997816 0.782119 0.00106579 0.00188124 0.000860146 0.45541 0.00188124 0.443915 0.00013099 1.02 0.88865 0.534409 0.287397 1.71917e-07 3.08181e-09 2372.57 3133.08 -0.05759 0.4822 0.277304 0.254398 -0.593145 -0.169567 0.489573 -0.266015 -0.223567 2.553 1 0 295.896 0 2.22004 2.551 0.000299243 0.864087 0.69567 0.320252 0.431836 2.22022 138.373 83.7132 18.7089 60.7664 0.00403386 0 -40 10
1.652 4.77968e-08 2.53976e-06 0.143674 0.143673 0.0120278 2.17258e-05 0.00115444 0.179593 0.000658755 0.180247 0.942109 101.506 0.236115 0.840681 4.49363 0.0638849 0.0423928 0.957607 0.0194919 0.00455244 0.0187502 0.00434678 0.00550815 0.00624976 0.220326 0.24999 58.0428 -87.8988 126.179 15.9388 145.034 0.000142028 0.267296 192.744 0.310235 0.0673303 0.00409818 0.000562311 0.00138487 0.986962 0.991718 -2.98861e-06 -85.658 0.0930765 31171.3 308.944 0.9835 0.319146 0.736772 0.736767 9.99958 2.98596e-06 1.19437e-05 0.133801 0.983373 0.931462 -0.0132917 4.92755e-06 0.514033 -1.99698e-20 7.40326e-24 -1.99624e-20 0.00139634 0.997815 8.60147e-05 0.152716 2.85269 0.00139634 0.997816 0.782195 0.0010658 0.00188124 0.000860147 0.45541 0.00188124 0.443921 0.000130993 1.02 0.888651 0.534408 0.287398 1.71917e-07 3.08184e-09 2372.55 3133.13 -0.0575948 0.4822 0.277304 0.254401 -0.593145 -0.169567 0.489558 -0.266013 -0.223554 2.554 1 0 295.892 0 2.22018 2.552 0.000299242 0.864114 0.695714 0.320208 0.431858 2.22036 138.38 83.7127 18.7088 60.7661 0.00403388 0 -40 10
1.653 4.78257e-08 2.53977e-06 0.14371 0.143709 0.0120278 2.1739e-05 0.00115444 0.179637 0.000658755 0.180292 0.942197 101.506 0.236105 0.840812 4.49421 0.0638955 0.0423982 0.957602 0.0194913 0.00455287 0.0187497 0.00434715 0.00550868 0.00625031 0.220347 0.250012 58.0429 -87.8988 126.179 15.9388 145.034 0.000142031 0.267296 192.743 0.310235 0.0673303 0.00409818 0.000562312 0.00138488 0.986962 0.991718 -2.98863e-06 -85.658 0.0930766 31171.3 308.955 0.9835 0.319146 0.736783 0.736779 9.99958 2.98597e-06 1.19438e-05 0.133806 0.983373 0.931461 -0.0132917 4.92758e-06 0.514052 -1.99713e-20 7.40386e-24 -1.99639e-20 0.00139634 0.997815 8.60147e-05 0.152717 2.8527 0.00139634 0.997816 0.782271 0.00106582 0.00188124 0.000860147 0.455409 0.00188124 0.443926 0.000130995 1.02 0.888653 0.534408 0.2874 1.71918e-07 3.08186e-09 2372.53 3133.17 -0.0575997 0.4822 0.277304 0.254404 -0.593144 -0.169567 0.489542 -0.266011 -0.223541 2.555 1 0 295.887 0 2.22032 2.553 0.000299241 0.864141 0.695757 0.320163 0.431881 2.2205 138.388 83.7121 18.7088 60.7659 0.0040339 0 -40 10
1.654 4.78545e-08 2.53977e-06 0.143746 0.143745 0.0120278 2.17521e-05 0.00115444 0.179682 0.000658756 0.180336 0.942286 101.505 0.236094 0.840943 4.49479 0.0639061 0.0424037 0.957596 0.0194908 0.0045533 0.0187491 0.00434752 0.00550921 0.00625085 0.220368 0.250034 58.043 -87.8988 126.179 15.9387 145.034 0.000142033 0.267296 192.743 0.310234 0.0673302 0.00409818 0.000562313 0.00138488 0.986962 0.991718 -2.98864e-06 -85.658 0.0930767 31171.2 308.967 0.9835 0.319146 0.736795 0.73679 9.99958 2.98597e-06 1.19438e-05 0.13381 0.983374 0.93146 -0.0132917 4.92761e-06 0.51407 -1.99728e-20 7.40446e-24 -1.99654e-20 0.00139634 0.997815 8.60148e-05 0.152717 2.8527 0.00139634 0.997816 0.782346 0.00106584 0.00188124 0.000860148 0.455409 0.00188124 0.443932 0.000130998 1.02 0.888654 0.534408 0.287401 1.71918e-07 3.08188e-09 2372.52 3133.22 -0.0576046 0.4822 0.277303 0.254407 -0.593143 -0.169567 0.489527 -0.266009 -0.223527 2.556 1 0 295.883 0 2.22046 2.554 0.00029924 0.864168 0.6958 0.320119 0.431903 2.22064 138.395 83.7115 18.7088 60.7656 0.00403393 0 -40 10
1.655 4.78834e-08 2.53977e-06 0.143782 0.143781 0.0120278 2.17652e-05 0.00115444 0.179727 0.000658757 0.180381 0.942374 101.505 0.236083 0.841074 4.49537 0.0639167 0.0424091 0.957591 0.0194903 0.00455373 0.0187486 0.00434789 0.00550974 0.0062514 0.22039 0.250056 58.043 -87.8988 126.179 15.9387 145.034 0.000142035 0.267296 192.743 0.310234 0.0673301 0.00409819 0.000562313 0.00138488 0.986962 0.991718 -2.98866e-06 -85.658 0.0930768 31171.2 308.979 0.9835 0.319146 0.736806 0.736802 9.99958 2.98598e-06 1.19438e-05 0.133814 0.983374 0.931459 -0.0132917 4.92764e-06 0.514089 -1.99743e-20 7.40506e-24 -1.99669e-20 0.00139634 0.997815 8.60149e-05 0.152717 2.8527 0.00139634 0.997816 0.782422 0.00106585 0.00188124 0.000860149 0.455409 0.00188124 0.443937 0.000131 1.02 0.888655 0.534407 0.287403 1.71918e-07 3.08191e-09 2372.5 3133.27 -0.0576094 0.4822 0.277303 0.25441 -0.593143 -0.169567 0.489511 -0.266007 -0.223514 2.557 1 0 295.879 0 2.22059 2.555 0.000299239 0.864195 0.695844 0.320074 0.431926 2.22078 138.402 83.711 18.7088 60.7653 0.00403395 0 -40 10
1.656 4.79123e-08 2.53977e-06 0.143817 0.143817 0.0120278 2.17783e-05 0.00115444 0.179772 0.000658757 0.180426 0.942463 101.504 0.236073 0.841205 4.49595 0.0639272 0.0424146 0.957585 0.0194897 0.00455417 0.0187481 0.00434826 0.00551028 0.00625195 0.220411 0.250078 58.0431 -87.8988 126.179 15.9387 145.034 0.000142037 0.267297 192.743 0.310234 0.0673301 0.00409819 0.000562314 0.00138488 0.986962 0.991718 -2.98867e-06 -85.6579 0.0930768 31171.2 308.991 0.983499 0.319146 0.736818 0.736813 9.99958 2.98598e-06 1.19438e-05 0.133819 0.983375 0.931459 -0.0132917 4.92767e-06 0.514108 -1.99758e-20 7.40567e-24 -1.99684e-20 0.00139635 0.997815 8.6015e-05 0.152717 2.8527 0.00139635 0.997816 0.782497 0.00106587 0.00188125 0.00086015 0.455409 0.00188125 0.443943 0.000131003 1.02 0.888656 0.534407 0.287404 1.71919e-07 3.08193e-09 2372.48 3133.32 -0.0576143 0.4822 0.277303 0.254413 -0.593142 -0.169567 0.489496 -0.266005 -0.2235 2.558 1 0 295.874 0 2.22073 2.556 0.000299237 0.864222 0.695887 0.32003 0.431948 2.22092 138.41 83.7104 18.7087 60.7651 0.00403397 0 -40 10
1.657 4.79411e-08 2.53977e-06 0.143853 0.143852 0.0120278 2.17914e-05 0.00115444 0.179816 0.000658758 0.18047 0.942551 101.503 0.236062 0.841337 4.49653 0.0639378 0.0424201 0.95758 0.0194892 0.0045546 0.0187475 0.00434864 0.00551081 0.00625249 0.220432 0.2501 58.0432 -87.8988 126.178 15.9386 145.034 0.000142039 0.267297 192.743 0.310233 0.06733 0.00409819 0.000562315 0.00138489 0.986962 0.991718 -2.98869e-06 -85.6579 0.0930769 31171.2 309.002 0.983499 0.319146 0.736829 0.736825 9.99958 2.98599e-06 1.19438e-05 0.133823 0.983375 0.931458 -0.0132917 4.9277e-06 0.514126 -1.99773e-20 7.40627e-24 -1.99699e-20 0.00139635 0.997815 8.60151e-05 0.152717 2.8527 0.00139635 0.997816 0.782573 0.00106589 0.00188125 0.000860151 0.455408 0.00188125 0.443948 0.000131005 1.02 0.888657 0.534407 0.287406 1.71919e-07 3.08195e-09 2372.47 3133.37 -0.0576192 0.4822 0.277303 0.254416 -0.593141 -0.169567 0.48948 -0.266003 -0.223487 2.559 1 0 295.87 0 2.22087 2.557 0.000299236 0.864249 0.69593 0.319986 0.43197 2.22105 138.417 83.7098 18.7087 60.7648 0.004034 0 -40 10
1.658 4.797e-08 2.53977e-06 0.143889 0.143888 0.0120278 2.18045e-05 0.00115444 0.179861 0.000658758 0.180515 0.94264 101.503 0.236052 0.841468 4.49711 0.0639484 0.0424256 0.957574 0.0194887 0.00455503 0.018747 0.00434901 0.00551134 0.00625304 0.220454 0.250122 58.0432 -87.8988 126.178 15.9386 145.034 0.000142042 0.267297 192.743 0.310233 0.06733 0.0040982 0.000562315 0.00138489 0.986962 0.991718 -2.9887e-06 -85.6579 0.093077 31171.1 309.014 0.983499 0.319146 0.73684 0.736836 9.99958 2.98599e-06 1.19439e-05 0.133828 0.983375 0.931457 -0.0132917 4.92773e-06 0.514145 -1.99788e-20 7.40687e-24 -1.99714e-20 0.00139635 0.997815 8.60151e-05 0.152717 2.8527 0.00139635 0.997816 0.782648 0.0010659 0.00188125 0.000860151 0.455408 0.00188125 0.443954 0.000131008 1.02 0.888658 0.534407 0.287407 1.71919e-07 3.08197e-09 2372.45 3133.41 -0.0576241 0.4822 0.277302 0.254419 -0.593141 -0.169567 0.489464 -0.266 -0.223473 2.56 1 0 295.865 0 2.22101 2.558 0.000299235 0.864276 0.695973 0.319941 0.431993 2.22119 138.425 83.7093 18.7087 60.7645 0.00403402 0 -40 10
1.659 4.79988e-08 2.53977e-06 0.143924 0.143924 0.0120277 2.18176e-05 0.00115444 0.179905 0.000658759 0.18056 0.942728 101.502 0.236041 0.841599 4.49769 0.063959 0.042431 0.957569 0.0194881 0.00455546 0.0187464 0.00434938 0.00551188 0.00625359 0.220475 0.250144 58.0433 -87.8988 126.178 15.9386 145.034 0.000142044 0.267297 192.742 0.310232 0.0673299 0.0040982 0.000562316 0.00138489 0.986962 0.991718 -2.98872e-06 -85.6579 0.0930771 31171.1 309.026 0.983499 0.319146 0.736852 0.736847 9.99958 2.986e-06 1.19439e-05 0.133832 0.983376 0.931456 -0.0132917 4.92776e-06 0.514164 -1.99803e-20 7.40748e-24 -1.99729e-20 0.00139635 0.997815 8.60152e-05 0.152717 2.8527 0.00139635 0.997816 0.782723 0.00106592 0.00188125 0.000860152 0.455408 0.00188125 0.443959 0.00013101 1.02 0.888659 0.534406 0.287409 1.71919e-07 3.082e-09 2372.43 3133.46 -0.0576289 0.4822 0.277302 0.254422 -0.59314 -0.169567 0.489449 -0.265998 -0.22346 2.561 1 0 295.861 0 2.22115 2.559 0.000299234 0.864304 0.696017 0.319897 0.432015 2.22133 138.432 83.7087 18.7086 60.7642 0.00403404 0 -40 10
1.66 4.80277e-08 2.53978e-06 0.14396 0.143959 0.0120277 2.18308e-05 0.00115444 0.17995 0.00065876 0.180604 0.942817 101.502 0.23603 0.84173 4.49827 0.0639696 0.0424365 0.957563 0.0194876 0.0045559 0.0187459 0.00434976 0.00551241 0.00625414 0.220496 0.250165 58.0433 -87.8988 126.178 15.9385 145.034 0.000142046 0.267297 192.742 0.310232 0.0673299 0.0040982 0.000562317 0.00138489 0.986962 0.991718 -2.98873e-06 -85.6579 0.0930772 31171.1 309.038 0.983499 0.319146 0.736863 0.736859 9.99958 2.986e-06 1.19439e-05 0.133836 0.983376 0.931455 -0.0132917 4.92778e-06 0.514183 -1.99818e-20 7.40808e-24 -1.99744e-20 0.00139635 0.997815 8.60153e-05 0.152718 2.8527 0.00139635 0.997815 0.782799 0.00106593 0.00188125 0.000860153 0.455408 0.00188125 0.443964 0.000131013 1.02 0.88866 0.534406 0.28741 1.7192e-07 3.08202e-09 2372.42 3133.51 -0.0576338 0.482201 0.277302 0.254425 -0.59314 -0.169567 0.489433 -0.265996 -0.223447 2.562 1 0 295.857 0 2.22129 2.56 0.000299233 0.864331 0.69606 0.319853 0.432038 2.22147 138.44 83.7082 18.7086 60.764 0.00403407 0 -40 10
1.661 4.80565e-08 2.53978e-06 0.143996 0.143995 0.0120277 2.18439e-05 0.00115444 0.179995 0.00065876 0.180649 0.942906 101.501 0.23602 0.841861 4.49885 0.0639802 0.042442 0.957558 0.0194871 0.00455633 0.0187453 0.00435013 0.00551294 0.00625468 0.220518 0.250187 58.0434 -87.8988 126.177 15.9385 145.034 0.000142048 0.267298 192.742 0.310231 0.0673298 0.00409821 0.000562317 0.00138489 0.986962 0.991718 -2.98875e-06 -85.6579 0.0930773 31171.1 309.049 0.983499 0.319146 0.736875 0.73687 9.99958 2.98601e-06 1.19439e-05 0.133841 0.983377 0.931454 -0.0132917 4.92781e-06 0.514202 -1.99834e-20 7.40868e-24 -1.99759e-20 0.00139635 0.997815 8.60154e-05 0.152718 2.8527 0.00139635 0.997815 0.782874 0.00106595 0.00188125 0.000860154 0.455408 0.00188125 0.44397 0.000131015 1.02 0.888661 0.534406 0.287412 1.7192e-07 3.08204e-09 2372.4 3133.56 -0.0576387 0.482201 0.277301 0.254429 -0.593139 -0.169568 0.489418 -0.265994 -0.223433 2.563 1 0 295.852 0 2.22142 2.561 0.000299232 0.864358 0.696103 0.319809 0.43206 2.22161 138.447 83.7076 18.7086 60.7637 0.00403409 0 -40 10
1.662 4.80854e-08 2.53978e-06 0.144031 0.144031 0.0120277 2.1857e-05 0.00115444 0.180039 0.000658761 0.180693 0.942994 101.501 0.236009 0.841992 4.49943 0.0639908 0.0424475 0.957553 0.0194865 0.00455677 0.0187448 0.0043505 0.00551348 0.00625523 0.220539 0.250209 58.0435 -87.8988 126.177 15.9384 145.034 0.00014205 0.267298 192.742 0.310231 0.0673298 0.00409821 0.000562318 0.0013849 0.986962 0.991718 -2.98876e-06 -85.6579 0.0930774 31171.1 309.061 0.983499 0.319146 0.736886 0.736882 9.99958 2.98601e-06 1.19439e-05 0.133845 0.983377 0.931453 -0.0132917 4.92784e-06 0.51422 -1.99849e-20 7.40929e-24 -1.99775e-20 0.00139635 0.997815 8.60155e-05 0.152718 2.8527 0.00139635 0.997815 0.78295 0.00106597 0.00188126 0.000860155 0.455407 0.00188125 0.443975 0.000131018 1.02 0.888662 0.534405 0.287413 1.7192e-07 3.08207e-09 2372.39 3133.61 -0.0576436 0.482201 0.277301 0.254432 -0.593138 -0.169568 0.489402 -0.265992 -0.22342 2.564 1 0 295.848 0 2.22156 2.562 0.000299231 0.864385 0.696147 0.319764 0.432083 2.22174 138.454 83.707 18.7085 60.7634 0.00403411 0 -40 10
1.663 4.81142e-08 2.53978e-06 0.144067 0.144066 0.0120277 2.18701e-05 0.00115445 0.180084 0.000658761 0.180738 0.943083 101.5 0.235999 0.842123 4.50002 0.0640015 0.042453 0.957547 0.019486 0.0045572 0.0187442 0.00435088 0.00551401 0.00625578 0.220561 0.250231 58.0435 -87.8988 126.177 15.9384 145.034 0.000142053 0.267298 192.742 0.310231 0.0673297 0.00409821 0.000562319 0.0013849 0.986962 0.991718 -2.98878e-06 -85.6579 0.0930775 31171 309.073 0.983499 0.319146 0.736898 0.736893 9.99958 2.98602e-06 1.1944e-05 0.13385 0.983377 0.931452 -0.0132917 4.92787e-06 0.514239 -1.99864e-20 7.40989e-24 -1.9979e-20 0.00139635 0.997815 8.60155e-05 0.152718 2.8527 0.00139635 0.997815 0.783025 0.00106598 0.00188126 0.000860155 0.455407 0.00188126 0.443981 0.00013102 1.02 0.888664 0.534405 0.287415 1.7192e-07 3.08209e-09 2372.37 3133.65 -0.0576485 0.482201 0.277301 0.254435 -0.593138 -0.169568 0.489387 -0.26599 -0.223406 2.565 1 0 295.843 0 2.2217 2.563 0.00029923 0.864413 0.69619 0.31972 0.432105 2.22188 138.462 83.7065 18.7085 60.7632 0.00403414 0 -40 10
1.664 4.81431e-08 2.53978e-06 0.144102 0.144102 0.0120277 2.18832e-05 0.00115445 0.180128 0.000658762 0.180782 0.943172 101.499 0.235988 0.842254 4.5006 0.0640121 0.0424585 0.957542 0.0194855 0.00455763 0.0187437 0.00435125 0.00551455 0.00625633 0.220582 0.250253 58.0436 -87.8988 126.177 15.9384 145.034 0.000142055 0.267298 192.742 0.31023 0.0673297 0.00409821 0.000562319 0.0013849 0.986962 0.991718 -2.98879e-06 -85.6579 0.0930775 31171 309.085 0.983499 0.319146 0.736909 0.736905 9.99958 2.98602e-06 1.1944e-05 0.133854 0.983378 0.931451 -0.0132917 4.9279e-06 0.514258 -1.99879e-20 7.4105e-24 -1.99805e-20 0.00139635 0.997815 8.60156e-05 0.152718 2.85271 0.00139635 0.997815 0.7831 0.001066 0.00188126 0.000860156 0.455407 0.00188126 0.443986 0.000131022 1.02 0.888665 0.534405 0.287416 1.71921e-07 3.08211e-09 2372.35 3133.7 -0.0576534 0.482201 0.277301 0.254438 -0.593137 -0.169568 0.489371 -0.265988 -0.223393 2.566 1 0 295.839 0 2.22184 2.564 0.000299228 0.86444 0.696233 0.319676 0.432128 2.22202 138.469 83.7059 18.7085 60.7629 0.00403416 0 -40 10
1.665 4.81719e-08 2.53978e-06 0.144138 0.144137 0.0120277 2.18963e-05 0.00115445 0.180172 0.000658763 0.180826 0.94326 101.499 0.235977 0.842386 4.50118 0.0640227 0.042464 0.957536 0.0194849 0.00455807 0.0187431 0.00435163 0.00551508 0.00625688 0.220603 0.250275 58.0437 -87.8988 126.177 15.9383 145.034 0.000142057 0.267298 192.741 0.31023 0.0673296 0.00409822 0.00056232 0.0013849 0.986962 0.991718 -2.98881e-06 -85.6579 0.0930776 31171 309.097 0.983499 0.319146 0.736921 0.736916 9.99958 2.98603e-06 1.1944e-05 0.133858 0.983378 0.93145 -0.0132917 4.92793e-06 0.514277 -1.99894e-20 7.4111e-24 -1.9982e-20 0.00139636 0.997815 8.60157e-05 0.152718 2.85271 0.00139636 0.997815 0.783175 0.00106602 0.00188126 0.000860157 0.455407 0.00188126 0.443992 0.000131025 1.02 0.888666 0.534404 0.287418 1.71921e-07 3.08213e-09 2372.34 3133.75 -0.0576582 0.482201 0.2773 0.254441 -0.593137 -0.169568 0.489356 -0.265986 -0.223379 2.567 1 0 295.835 0 2.22198 2.565 0.000299227 0.864467 0.696276 0.319632 0.43215 2.22216 138.477 83.7053 18.7084 60.7626 0.00403418 0 -40 10
1.666 4.82008e-08 2.53978e-06 0.144173 0.144173 0.0120276 2.19094e-05 0.00115445 0.180217 0.000658763 0.180871 0.943349 101.498 0.235967 0.842517 4.50177 0.0640333 0.0424695 0.95753 0.0194844 0.0045585 0.0187426 0.004352 0.00551562 0.00625743 0.220625 0.250297 58.0437 -87.8988 126.176 15.9383 145.034 0.000142059 0.267299 192.741 0.310229 0.0673296 0.00409822 0.000562321 0.00138491 0.986962 0.991718 -2.98882e-06 -85.6578 0.0930777 31171 309.108 0.983499 0.319146 0.736932 0.736928 9.99958 2.98603e-06 1.1944e-05 0.133863 0.983378 0.931449 -0.0132917 4.92796e-06 0.514296 -1.99909e-20 7.41171e-24 -1.99835e-20 0.00139636 0.997815 8.60158e-05 0.152719 2.85271 0.00139636 0.997815 0.783251 0.00106603 0.00188126 0.000860158 0.455406 0.00188126 0.443997 0.000131027 1.02 0.888667 0.534404 0.28742 1.71921e-07 3.08216e-09 2372.32 3133.8 -0.0576631 0.482201 0.2773 0.254444 -0.593136 -0.169568 0.48934 -0.265984 -0.223366 2.568 1 0 295.83 0 2.22211 2.566 0.000299226 0.864494 0.69632 0.319588 0.432172 2.2223 138.484 83.7048 18.7084 60.7623 0.00403421 0 -40 10
1.667 4.82296e-08 2.53979e-06 0.144209 0.144208 0.0120276 2.19226e-05 0.00115445 0.180261 0.000658764 0.180915 0.943438 101.498 0.235956 0.842648 4.50235 0.0640439 0.042475 0.957525 0.0194838 0.00455894 0.018742 0.00435238 0.00551615 0.00625798 0.220646 0.250319 58.0438 -87.8988 126.176 15.9383 145.034 0.000142061 0.267299 192.741 0.310229 0.0673295 0.00409822 0.000562321 0.00138491 0.986962 0.991718 -2.98884e-06 -85.6578 0.0930778 31170.9 309.12 0.983499 0.319146 0.736944 0.736939 9.99958 2.98604e-06 1.1944e-05 0.133867 0.983379 0.931448 -0.0132917 4.92799e-06 0.514314 -1.99924e-20 7.41232e-24 -1.9985e-20 0.00139636 0.997815 8.60159e-05 0.152719 2.85271 0.00139636 0.997815 0.783326 0.00106605 0.00188126 0.000860159 0.455406 0.00188126 0.444003 0.00013103 1.02 0.888668 0.534404 0.287421 1.71922e-07 3.08218e-09 2372.3 3133.85 -0.057668 0.482201 0.2773 0.254447 -0.593135 -0.169568 0.489324 -0.265982 -0.223352 2.569 1 0 295.826 0 2.22225 2.567 0.000299225 0.864522 0.696363 0.319544 0.432195 2.22243 138.491 83.7042 18.7084 60.7621 0.00403423 0 -40 10
1.668 4.82585e-08 2.53979e-06 0.144244 0.144244 0.0120276 2.19357e-05 0.00115445 0.180305 0.000658764 0.180959 0.943526 101.497 0.235945 0.842779 4.50294 0.0640545 0.0424805 0.957519 0.0194833 0.00455937 0.0187415 0.00435275 0.00551669 0.00625853 0.220668 0.250341 58.0438 -87.8988 126.176 15.9382 145.034 0.000142064 0.267299 192.741 0.310228 0.0673295 0.00409823 0.000562322 0.00138491 0.986962 0.991718 -2.98885e-06 -85.6578 0.0930779 31170.9 309.132 0.983499 0.319146 0.736955 0.736951 9.99958 2.98604e-06 1.19441e-05 0.133872 0.983379 0.931447 -0.0132917 4.92802e-06 0.514333 -1.99939e-20 7.41292e-24 -1.99865e-20 0.00139636 0.997815 8.60159e-05 0.152719 2.85271 0.00139636 0.997815 0.783401 0.00106607 0.00188126 0.000860159 0.455406 0.00188126 0.444008 0.000131032 1.02 0.888669 0.534403 0.287423 1.71922e-07 3.0822e-09 2372.29 3133.89 -0.0576729 0.482201 0.2773 0.25445 -0.593135 -0.169568 0.489309 -0.265979 -0.223339 2.57 1 0 295.821 0 2.22239 2.568 0.000299224 0.864549 0.696406 0.3195 0.432217 2.22257 138.499 83.7036 18.7083 60.7618 0.00403425 0 -40 10
1.669 4.82873e-08 2.53979e-06 0.14428 0.144279 0.0120276 2.19488e-05 0.00115445 0.180349 0.000658765 0.181004 0.943615 101.496 0.235935 0.842911 4.50352 0.0640651 0.0424861 0.957514 0.0194828 0.00455981 0.0187409 0.00435313 0.00551723 0.00625908 0.220689 0.250363 58.0439 -87.8988 126.176 15.9382 145.034 0.000142066 0.267299 192.741 0.310228 0.0673294 0.00409823 0.000562323 0.00138491 0.986962 0.991718 -2.98887e-06 -85.6578 0.093078 31170.9 309.144 0.983499 0.319146 0.736966 0.736962 9.99958 2.98605e-06 1.19441e-05 0.133876 0.98338 0.931446 -0.0132917 4.92805e-06 0.514352 -1.99954e-20 7.41353e-24 -1.9988e-20 0.00139636 0.997815 8.6016e-05 0.152719 2.85271 0.00139636 0.997815 0.783476 0.00106608 0.00188127 0.00086016 0.455406 0.00188126 0.444013 0.000131035 1.02 0.88867 0.534403 0.287424 1.71922e-07 3.08223e-09 2372.27 3133.94 -0.0576778 0.482201 0.277299 0.254453 -0.593134 -0.169568 0.489293 -0.265977 -0.223325 2.571 1 0 295.817 0 2.22253 2.569 0.000299223 0.864576 0.696449 0.319456 0.43224 2.22271 138.506 83.7031 18.7083 60.7615 0.00403428 0 -40 10
1.67 4.83162e-08 2.53979e-06 0.144315 0.144314 0.0120276 2.19619e-05 0.00115445 0.180394 0.000658765 0.181048 0.943704 101.496 0.235924 0.843042 4.50411 0.0640757 0.0424916 0.957508 0.0194822 0.00456024 0.0187404 0.0043535 0.00551776 0.00625963 0.220711 0.250385 58.044 -87.8988 126.176 15.9381 145.034 0.000142068 0.267299 192.741 0.310228 0.0673294 0.00409823 0.000562323 0.00138491 0.986962 0.991718 -2.98888e-06 -85.6578 0.0930781 31170.9 309.156 0.983499 0.319146 0.736978 0.736974 9.99958 2.98605e-06 1.19441e-05 0.133881 0.98338 0.931446 -0.0132917 4.92808e-06 0.514371 -1.9997e-20 7.41414e-24 -1.99895e-20 0.00139636 0.997815 8.60161e-05 0.152719 2.85271 0.00139636 0.997815 0.783551 0.0010661 0.00188127 0.000860161 0.455406 0.00188127 0.444019 0.000131037 1.02 0.888671 0.534403 0.287426 1.71922e-07 3.08225e-09 2372.25 3133.99 -0.0576827 0.482201 0.277299 0.254456 -0.593134 -0.169568 0.489278 -0.265975 -0.223312 2.572 1 0 295.813 0 2.22267 2.57 0.000299222 0.864604 0.696493 0.319412 0.432262 2.22285 138.514 83.7025 18.7083 60.7613 0.0040343 0 -40 10
1.671 4.8345e-08 2.53979e-06 0.14435 0.14435 0.0120276 2.1975e-05 0.00115445 0.180438 0.000658766 0.181092 0.943793 101.495 0.235914 0.843173 4.50469 0.0640864 0.0424971 0.957503 0.0194817 0.00456068 0.0187398 0.00435388 0.0055183 0.00626018 0.220732 0.250407 58.044 -87.8988 126.175 15.9381 145.034 0.00014207 0.2673 192.74 0.310227 0.0673293 0.00409824 0.000562324 0.00138492 0.986962 0.991718 -2.9889e-06 -85.6578 0.0930782 31170.8 309.168 0.983499 0.319146 0.736989 0.736985 9.99958 2.98606e-06 1.19441e-05 0.133885 0.98338 0.931445 -0.0132917 4.92811e-06 0.51439 -1.99985e-20 7.41474e-24 -1.99911e-20 0.00139636 0.997815 8.60162e-05 0.152719 2.85271 0.00139636 0.997815 0.783626 0.00106612 0.00188127 0.000860162 0.455405 0.00188127 0.444024 0.00013104 1.02 0.888672 0.534403 0.287427 1.71923e-07 3.08227e-09 2372.24 3134.04 -0.0576876 0.482201 0.277299 0.254459 -0.593133 -0.169568 0.489262 -0.265973 -0.223298 2.573 1 0 295.808 0 2.22281 2.571 0.00029922 0.864631 0.696536 0.319369 0.432285 2.22299 138.521 83.7019 18.7082 60.761 0.00403432 0 -40 10
1.672 4.83739e-08 2.53979e-06 0.144386 0.144385 0.0120276 2.19881e-05 0.00115445 0.180482 0.000658767 0.181136 0.943882 101.495 0.235903 0.843304 4.50528 0.064097 0.0425026 0.957497 0.0194812 0.00456111 0.0187393 0.00435425 0.00551884 0.00626073 0.220753 0.250429 58.0441 -87.8988 126.175 15.9381 145.034 0.000142072 0.2673 192.74 0.310227 0.0673293 0.00409824 0.000562325 0.00138492 0.986962 0.991718 -2.98891e-06 -85.6578 0.0930782 31170.8 309.179 0.983499 0.319146 0.737001 0.736997 9.99958 2.98606e-06 1.19441e-05 0.13389 0.983381 0.931444 -0.0132917 4.92814e-06 0.514409 -2e-20 7.41535e-24 -1.99926e-20 0.00139636 0.997815 8.60163e-05 0.152719 2.85271 0.00139636 0.997815 0.783701 0.00106613 0.00188127 0.000860163 0.455405 0.00188127 0.44403 0.000131042 1.02 0.888673 0.534402 0.287429 1.71923e-07 3.08229e-09 2372.22 3134.09 -0.0576925 0.482201 0.277298 0.254462 -0.593132 -0.169568 0.489246 -0.265971 -0.223285 2.574 1 0 295.804 0 2.22294 2.572 0.000299219 0.864659 0.696579 0.319325 0.432307 2.22313 138.528 83.7014 18.7082 60.7607 0.00403435 0 -40 10
1.673 4.84027e-08 2.5398e-06 0.144421 0.14442 0.0120275 2.20012e-05 0.00115445 0.180526 0.000658767 0.18118 0.94397 101.494 0.235892 0.843436 4.50587 0.0641076 0.0425082 0.957492 0.0194806 0.00456155 0.0187387 0.00435463 0.00551937 0.00626129 0.220775 0.250451 58.0442 -87.8988 126.175 15.938 145.034 0.000142075 0.2673 192.74 0.310226 0.0673292 0.00409824 0.000562325 0.00138492 0.986962 0.991718 -2.98893e-06 -85.6578 0.0930783 31170.8 309.191 0.983499 0.319146 0.737012 0.737008 9.99958 2.98607e-06 1.19442e-05 0.133894 0.983381 0.931443 -0.0132917 4.92817e-06 0.514428 -2.00015e-20 7.41596e-24 -1.99941e-20 0.00139637 0.997815 8.60163e-05 0.15272 2.85271 0.00139636 0.997815 0.783776 0.00106615 0.00188127 0.000860163 0.455405 0.00188127 0.444035 0.000131045 1.02 0.888675 0.534402 0.28743 1.71923e-07 3.08232e-09 2372.2 3134.13 -0.0576974 0.482202 0.277298 0.254466 -0.593132 -0.169568 0.489231 -0.265969 -0.223271 2.575 1 0 295.799 0 2.22308 2.573 0.000299218 0.864686 0.696622 0.319281 0.432329 2.22326 138.536 83.7008 18.7082 60.7604 0.00403437 0 -40 10
1.674 4.84316e-08 2.5398e-06 0.144456 0.144456 0.0120275 2.20144e-05 0.00115445 0.18057 0.000658768 0.181224 0.944059 101.494 0.235882 0.843567 4.50645 0.0641182 0.0425137 0.957486 0.0194801 0.00456199 0.0187382 0.004355 0.00551991 0.00626184 0.220796 0.250474 58.0442 -87.8988 126.175 15.938 145.034 0.000142077 0.2673 192.74 0.310226 0.0673291 0.00409825 0.000562326 0.00138492 0.986962 0.991718 -2.98894e-06 -85.6578 0.0930784 31170.8 309.203 0.983499 0.319146 0.737024 0.73702 9.99958 2.98607e-06 1.19442e-05 0.133898 0.983381 0.931442 -0.0132917 4.9282e-06 0.514447 -2.0003e-20 7.41657e-24 -1.99956e-20 0.00139637 0.997815 8.60164e-05 0.15272 2.85271 0.00139637 0.997815 0.783852 0.00106617 0.00188127 0.000860164 0.455405 0.00188127 0.44404 0.000131047 1.02 0.888676 0.534402 0.287432 1.71923e-07 3.08234e-09 2372.19 3134.18 -0.0577023 0.482202 0.277298 0.254469 -0.593131 -0.169568 0.489215 -0.265967 -0.223258 2.576 1 0 295.795 0 2.22322 2.574 0.000299217 0.864713 0.696666 0.319237 0.432352 2.2234 138.543 83.7002 18.7081 60.7602 0.00403439 0 -40 10
1.675 4.84604e-08 2.5398e-06 0.144491 0.144491 0.0120275 2.20275e-05 0.00115445 0.180614 0.000658768 0.181268 0.944148 101.493 0.235871 0.843698 4.50704 0.0641288 0.0425193 0.957481 0.0194795 0.00456242 0.0187376 0.00435538 0.00552045 0.00626239 0.220818 0.250496 58.0443 -87.8988 126.175 15.938 145.034 0.000142079 0.2673 192.74 0.310225 0.0673291 0.00409825 0.000562327 0.00138492 0.986962 0.991718 -2.98896e-06 -85.6578 0.0930785 31170.8 309.215 0.983499 0.319146 0.737036 0.737031 9.99958 2.98607e-06 1.19442e-05 0.133903 0.983382 0.931441 -0.0132917 4.92823e-06 0.514465 -2.00045e-20 7.41718e-24 -1.99971e-20 0.00139637 0.997815 8.60165e-05 0.15272 2.85272 0.00139637 0.997815 0.783927 0.00106618 0.00188127 0.000860165 0.455404 0.00188127 0.444046 0.00013105 1.02 0.888677 0.534401 0.287433 1.71924e-07 3.08236e-09 2372.17 3134.23 -0.0577072 0.482202 0.277298 0.254472 -0.593131 -0.169568 0.4892 -0.265965 -0.223244 2.577 1 0 295.791 0 2.22336 2.575 0.000299216 0.864741 0.696709 0.319194 0.432374 2.22354 138.551 83.6997 18.7081 60.7599 0.00403442 0 -40 10
1.676 4.84893e-08 2.5398e-06 0.144527 0.144526 0.0120275 2.20406e-05 0.00115445 0.180658 0.000658769 0.181312 0.944237 101.492 0.235861 0.84383 4.50763 0.0641395 0.0425248 0.957475 0.019479 0.00456286 0.0187371 0.00435576 0.00552099 0.00626294 0.22084 0.250518 58.0443 -87.8989 126.174 15.9379 145.034 0.000142081 0.2673 192.74 0.310225 0.067329 0.00409825 0.000562327 0.00138493 0.986962 0.991717 -2.98897e-06 -85.6578 0.0930786 31170.7 309.227 0.983499 0.319146 0.737047 0.737043 9.99958 2.98608e-06 1.19442e-05 0.133907 0.983382 0.93144 -0.0132917 4.92826e-06 0.514484 -2.00061e-20 7.41778e-24 -1.99986e-20 0.00139637 0.997815 8.60166e-05 0.15272 2.85272 0.00139637 0.997815 0.784001 0.0010662 0.00188128 0.000860166 0.455404 0.00188127 0.444051 0.000131052 1.02 0.888678 0.534401 0.287435 1.71924e-07 3.08239e-09 2372.16 3134.28 -0.0577121 0.482202 0.277297 0.254475 -0.59313 -0.169568 0.489184 -0.265963 -0.223231 2.578 1 0 295.786 0 2.2235 2.576 0.000299215 0.864768 0.696752 0.31915 0.432397 2.22368 138.558 83.6991 18.7081 60.7596 0.00403444 0 -40 10
1.677 4.85181e-08 2.5398e-06 0.144562 0.144561 0.0120275 2.20537e-05 0.00115446 0.180702 0.00065877 0.181356 0.944326 101.492 0.23585 0.843961 4.50822 0.0641501 0.0425304 0.95747 0.0194785 0.0045633 0.0187365 0.00435613 0.00552153 0.0062635 0.220861 0.25054 58.0444 -87.8989 126.174 15.9379 145.034 0.000142084 0.267301 192.739 0.310225 0.067329 0.00409825 0.000562328 0.00138493 0.986962 0.991717 -2.98899e-06 -85.6577 0.0930787 31170.7 309.239 0.983499 0.319146 0.737059 0.737054 9.99958 2.98608e-06 1.19442e-05 0.133912 0.983383 0.931439 -0.0132917 4.92829e-06 0.514503 -2.00076e-20 7.41839e-24 -2.00002e-20 0.00139637 0.997815 8.60167e-05 0.15272 2.85272 0.00139637 0.997815 0.784076 0.00106622 0.00188128 0.000860167 0.455404 0.00188128 0.444057 0.000131055 1.02 0.888679 0.534401 0.287436 1.71924e-07 3.08241e-09 2372.14 3134.33 -0.057717 0.482202 0.277297 0.254478 -0.593129 -0.169569 0.489168 -0.265961 -0.223217 2.579 1 0 295.782 0 2.22363 2.577 0.000299214 0.864796 0.696795 0.319107 0.432419 2.22382 138.565 83.6985 18.708 60.7593 0.00403446 0 -40 10
1.678 4.8547e-08 2.5398e-06 0.144597 0.144596 0.0120275 2.20668e-05 0.00115446 0.180746 0.00065877 0.1814 0.944415 101.491 0.235839 0.844093 4.50881 0.0641607 0.0425359 0.957464 0.0194779 0.00456373 0.0187359 0.00435651 0.00552207 0.00626405 0.220883 0.250562 58.0445 -87.8989 126.174 15.9378 145.034 0.000142086 0.267301 192.739 0.310224 0.0673289 0.00409826 0.000562329 0.00138493 0.986962 0.991717 -2.989e-06 -85.6577 0.0930788 31170.7 309.251 0.983499 0.319146 0.73707 0.737066 9.99958 2.98609e-06 1.19443e-05 0.133916 0.983383 0.931438 -0.0132917 4.92832e-06 0.514522 -2.00091e-20 7.419e-24 -2.00017e-20 0.00139637 0.997815 8.60168e-05 0.15272 2.85272 0.00139637 0.997815 0.784151 0.00106623 0.00188128 0.000860168 0.455404 0.00188128 0.444062 0.000131057 1.02 0.88868 0.5344 0.287438 1.71925e-07 3.08243e-09 2372.12 3134.38 -0.0577219 0.482202 0.277297 0.254481 -0.593129 -0.169569 0.489153 -0.265958 -0.223204 2.58 1 0 295.777 0 2.22377 2.578 0.000299212 0.864823 0.696839 0.319063 0.432441 2.22395 138.573 83.698 18.708 60.7591 0.00403449 0 -40 10
1.679 4.85758e-08 2.5398e-06 0.144632 0.144631 0.0120275 2.20799e-05 0.00115446 0.18079 0.000658771 0.181444 0.944504 101.491 0.235829 0.844224 4.5094 0.0641714 0.0425415 0.957458 0.0194774 0.00456417 0.0187354 0.00435689 0.0055226 0.0062646 0.220904 0.250584 58.0445 -87.8989 126.174 15.9378 145.034 0.000142088 0.267301 192.739 0.310224 0.0673289 0.00409826 0.000562329 0.00138493 0.986962 0.991717 -2.98902e-06 -85.6577 0.0930789 31170.7 309.262 0.983499 0.319146 0.737082 0.737077 9.99958 2.98609e-06 1.19443e-05 0.133921 0.983383 0.931437 -0.0132917 4.92835e-06 0.514541 -2.00106e-20 7.41961e-24 -2.00032e-20 0.00139637 0.997815 8.60168e-05 0.152721 2.85272 0.00139637 0.997815 0.784226 0.00106625 0.00188128 0.000860168 0.455403 0.00188128 0.444067 0.00013106 1.02 0.888681 0.5344 0.287439 1.71925e-07 3.08246e-09 2372.11 3134.42 -0.0577268 0.482202 0.277296 0.254484 -0.593128 -0.169569 0.489137 -0.265956 -0.22319 2.581 1 0 295.773 0 2.22391 2.579 0.000299211 0.864851 0.696882 0.31902 0.432464 2.22409 138.58 83.6974 18.708 60.7588 0.00403451 0 -40 10
1.68 4.86047e-08 2.53981e-06 0.144667 0.144666 0.0120274 2.2093e-05 0.00115446 0.180834 0.000658771 0.181488 0.944593 101.49 0.235818 0.844356 4.50999 0.064182 0.0425471 0.957453 0.0194769 0.00456461 0.0187348 0.00435727 0.00552314 0.00626516 0.220926 0.250606 58.0446 -87.8989 126.174 15.9378 145.034 0.00014209 0.267301 192.739 0.310223 0.0673288 0.00409826 0.00056233 0.00138494 0.986962 0.991717 -2.98903e-06 -85.6577 0.0930789 31170.6 309.274 0.983499 0.319146 0.737093 0.737089 9.99958 2.9861e-06 1.19443e-05 0.133925 0.983384 0.931436 -0.0132917 4.92838e-06 0.51456 -2.00121e-20 7.42022e-24 -2.00047e-20 0.00139637 0.997815 8.60169e-05 0.152721 2.85272 0.00139637 0.997815 0.784301 0.00106626 0.00188128 0.000860169 0.455403 0.00188128 0.444073 0.000131062 1.02 0.888682 0.5344 0.287441 1.71925e-07 3.08248e-09 2372.09 3134.47 -0.0577317 0.482202 0.277296 0.254487 -0.593127 -0.169569 0.489122 -0.265954 -0.223177 2.582 1 0 295.768 0 2.22405 2.58 0.00029921 0.864878 0.696925 0.318976 0.432486 2.22423 138.588 83.6968 18.7079 60.7585 0.00403453 0 -40 10
1.681 4.86335e-08 2.53981e-06 0.144702 0.144701 0.0120274 2.21062e-05 0.00115446 0.180878 0.000658772 0.181532 0.944682 101.489 0.235807 0.844487 4.51058 0.0641926 0.0425526 0.957447 0.0194763 0.00456505 0.0187343 0.00435764 0.00552368 0.00626571 0.220947 0.250628 58.0447 -87.8989 126.173 15.9377 145.034 0.000142092 0.267301 192.739 0.310223 0.0673288 0.00409827 0.000562331 0.00138494 0.986962 0.991717 -2.98905e-06 -85.6577 0.093079 31170.6 309.286 0.983499 0.319146 0.737105 0.7371 9.99958 2.9861e-06 1.19443e-05 0.13393 0.983384 0.931435 -0.0132917 4.92841e-06 0.514579 -2.00137e-20 7.42083e-24 -2.00062e-20 0.00139637 0.997815 8.6017e-05 0.152721 2.85272 0.00139637 0.997815 0.784376 0.00106628 0.00188128 0.00086017 0.455403 0.00188128 0.444078 0.000131064 1.02 0.888683 0.534399 0.287442 1.71925e-07 3.0825e-09 2372.07 3134.52 -0.0577367 0.482202 0.277296 0.25449 -0.593127 -0.169569 0.489106 -0.265952 -0.223163 2.583 1 0 295.764 0 2.22419 2.581 0.000299209 0.864906 0.696968 0.318933 0.432509 2.22437 138.595 83.6963 18.7079 60.7582 0.00403456 0 -40 10
1.682 4.86624e-08 2.53981e-06 0.144737 0.144736 0.0120274 2.21193e-05 0.00115446 0.180921 0.000658772 0.181576 0.944771 101.489 0.235797 0.844618 4.51117 0.0642033 0.0425582 0.957442 0.0194758 0.00456549 0.0187337 0.00435802 0.00552422 0.00626627 0.220969 0.250651 58.0447 -87.8989 126.173 15.9377 145.034 0.000142095 0.267302 192.739 0.310222 0.0673287 0.00409827 0.000562331 0.00138494 0.986962 0.991717 -2.98906e-06 -85.6577 0.0930791 31170.6 309.298 0.983499 0.319146 0.737116 0.737112 9.99958 2.98611e-06 1.19443e-05 0.133934 0.983384 0.931434 -0.0132917 4.92844e-06 0.514598 -2.00152e-20 7.42144e-24 -2.00078e-20 0.00139638 0.997815 8.60171e-05 0.152721 2.85272 0.00139638 0.997815 0.784451 0.0010663 0.00188129 0.000860171 0.455403 0.00188128 0.444084 0.000131067 1.02 0.888684 0.534399 0.287444 1.71926e-07 3.08252e-09 2372.06 3134.57 -0.0577416 0.482202 0.277296 0.254493 -0.593126 -0.169569 0.48909 -0.26595 -0.22315 2.584 1 0 295.76 0 2.22432 2.582 0.000299208 0.864933 0.697012 0.318889 0.432531 2.2245 138.603 83.6957 18.7079 60.758 0.00403458 0 -40 10
1.683 4.86912e-08 2.53981e-06 0.144772 0.144771 0.0120274 2.21324e-05 0.00115446 0.180965 0.000658773 0.181619 0.944859 101.488 0.235786 0.84475 4.51176 0.0642139 0.0425638 0.957436 0.0194752 0.00456592 0.0187332 0.0043584 0.00552476 0.00626682 0.220991 0.250673 58.0448 -87.8989 126.173 15.9377 145.034 0.000142097 0.267302 192.738 0.310222 0.0673287 0.00409827 0.000562332 0.00138494 0.986962 0.991717 -2.98908e-06 -85.6577 0.0930792 31170.6 309.31 0.983499 0.319146 0.737128 0.737123 9.99958 2.98611e-06 1.19444e-05 0.133939 0.983385 0.931433 -0.0132917 4.92847e-06 0.514617 -2.00167e-20 7.42205e-24 -2.00093e-20 0.00139638 0.997815 8.60172e-05 0.152721 2.85272 0.00139638 0.997815 0.784525 0.00106631 0.00188129 0.000860172 0.455403 0.00188129 0.444089 0.000131069 1.02 0.888686 0.534399 0.287445 1.71926e-07 3.08255e-09 2372.04 3134.62 -0.0577465 0.482202 0.277295 0.254497 -0.593126 -0.169569 0.489075 -0.265948 -0.223136 2.585 1 0 295.755 0 2.22446 2.583 0.000299207 0.864961 0.697055 0.318846 0.432553 2.22464 138.61 83.6951 18.7078 60.7577 0.0040346 0 -40 10
1.684 4.87201e-08 2.53981e-06 0.144807 0.144806 0.0120274 2.21455e-05 0.00115446 0.181009 0.000658774 0.181663 0.944948 101.488 0.235775 0.844881 4.51236 0.0642245 0.0425694 0.957431 0.0194747 0.00456636 0.0187326 0.00435878 0.0055253 0.00626738 0.221012 0.250695 58.0448 -87.8989 126.173 15.9376 145.034 0.000142099 0.267302 192.738 0.310222 0.0673286 0.00409828 0.000562333 0.00138494 0.986962 0.991717 -2.98909e-06 -85.6577 0.0930793 31170.6 309.322 0.983499 0.319146 0.737139 0.737135 9.99958 2.98612e-06 1.19444e-05 0.133943 0.983385 0.931432 -0.0132917 4.9285e-06 0.514636 -2.00182e-20 7.42266e-24 -2.00108e-20 0.00139638 0.997815 8.60172e-05 0.152721 2.85272 0.00139638 0.997815 0.7846 0.00106633 0.00188129 0.000860172 0.455402 0.00188129 0.444094 0.000131072 1.02 0.888687 0.534399 0.287447 1.71926e-07 3.08257e-09 2372.02 3134.67 -0.0577514 0.482202 0.277295 0.2545 -0.593125 -0.169569 0.489059 -0.265946 -0.223123 2.586 1 0 295.751 0 2.2246 2.584 0.000299206 0.864988 0.697098 0.318803 0.432576 2.22478 138.617 83.6946 18.7078 60.7574 0.00403463 0 -40 10
1.685 4.87489e-08 2.53981e-06 0.144842 0.144841 0.0120274 2.21586e-05 0.00115446 0.181052 0.000658774 0.181707 0.945037 101.487 0.235765 0.845013 4.51295 0.0642352 0.042575 0.957425 0.0194742 0.0045668 0.0187321 0.00435916 0.00552584 0.00626793 0.221034 0.250717 58.0449 -87.8989 126.172 15.9376 145.034 0.000142101 0.267302 192.738 0.310221 0.0673286 0.00409828 0.000562333 0.00138495 0.986962 0.991717 -2.98911e-06 -85.6577 0.0930794 31170.5 309.334 0.983499 0.319146 0.737151 0.737147 9.99958 2.98612e-06 1.19444e-05 0.133947 0.983385 0.931431 -0.0132917 4.92853e-06 0.514655 -2.00198e-20 7.42328e-24 -2.00123e-20 0.00139638 0.997815 8.60173e-05 0.152721 2.85273 0.00139638 0.997815 0.784675 0.00106635 0.00188129 0.000860173 0.455402 0.00188129 0.4441 0.000131074 1.02 0.888688 0.534398 0.287448 1.71926e-07 3.08259e-09 2372.01 3134.71 -0.0577563 0.482202 0.277295 0.254503 -0.593124 -0.169569 0.489043 -0.265944 -0.223109 2.587 1 0 295.746 0 2.22474 2.585 0.000299204 0.865016 0.697141 0.318759 0.432598 2.22492 138.625 83.694 18.7078 60.7571 0.00403465 0 -40 10
1.686 4.87778e-08 2.53982e-06 0.144877 0.144876 0.0120274 2.21717e-05 0.00115446 0.181096 0.000658775 0.18175 0.945127 101.486 0.235754 0.845145 4.51354 0.0642458 0.0425806 0.957419 0.0194736 0.00456724 0.0187315 0.00435953 0.00552639 0.00626849 0.221055 0.250739 58.045 -87.8989 126.172 15.9375 145.034 0.000142104 0.267302 192.738 0.310221 0.0673285 0.00409828 0.000562334 0.00138495 0.986961 0.991717 -2.98912e-06 -85.6577 0.0930795 31170.5 309.346 0.983499 0.319146 0.737163 0.737158 9.99958 2.98613e-06 1.19444e-05 0.133952 0.983386 0.93143 -0.0132917 4.92856e-06 0.514674 -2.00213e-20 7.42389e-24 -2.00139e-20 0.00139638 0.997815 8.60174e-05 0.152722 2.85273 0.00139638 0.997815 0.78475 0.00106636 0.00188129 0.000860174 0.455402 0.00188129 0.444105 0.000131077 1.02 0.888689 0.534398 0.28745 1.71927e-07 3.08262e-09 2371.99 3134.76 -0.0577612 0.482203 0.277294 0.254506 -0.593124 -0.169569 0.489028 -0.265942 -0.223095 2.588 1 0 295.742 0 2.22487 2.586 0.000299203 0.865043 0.697184 0.318716 0.432621 2.22506 138.632 83.6934 18.7077 60.7569 0.00403468 0 -40 10
1.687 4.88066e-08 2.53982e-06 0.144912 0.144911 0.0120274 2.21848e-05 0.00115446 0.18114 0.000658775 0.181794 0.945216 101.486 0.235744 0.845276 4.51413 0.0642565 0.0425862 0.957414 0.0194731 0.00456768 0.018731 0.00435991 0.00552693 0.00626904 0.221077 0.250762 58.045 -87.8989 126.172 15.9375 145.035 0.000142106 0.267303 192.738 0.31022 0.0673285 0.00409828 0.000562335 0.00138495 0.986961 0.991717 -2.98914e-06 -85.6577 0.0930796 31170.5 309.358 0.983499 0.319146 0.737174 0.73717 9.99958 2.98613e-06 1.19444e-05 0.133956 0.983386 0.93143 -0.0132917 4.92859e-06 0.514693 -2.00228e-20 7.4245e-24 -2.00154e-20 0.00139638 0.997815 8.60175e-05 0.152722 2.85273 0.00139638 0.997815 0.784824 0.00106638 0.00188129 0.000860175 0.455402 0.00188129 0.444111 0.000131079 1.02 0.88869 0.534398 0.287451 1.71927e-07 3.08264e-09 2371.98 3134.81 -0.0577662 0.482203 0.277294 0.254509 -0.593123 -0.169569 0.489012 -0.26594 -0.223082 2.589 1 0 295.737 0 2.22501 2.587 0.000299202 0.865071 0.697228 0.318673 0.432643 2.22519 138.64 83.6928 18.7077 60.7566 0.0040347 0 -40 10
1.688 4.88355e-08 2.53982e-06 0.144947 0.144946 0.0120273 2.2198e-05 0.00115446 0.181183 0.000658776 0.181837 0.945305 101.485 0.235733 0.845408 4.51473 0.0642671 0.0425918 0.957408 0.0194725 0.00456812 0.0187304 0.00436029 0.00552747 0.0062696 0.221099 0.250784 58.0451 -87.8989 126.172 15.9375 145.035 0.000142108 0.267303 192.738 0.31022 0.0673284 0.00409829 0.000562335 0.00138495 0.986961 0.991717 -2.98915e-06 -85.6576 0.0930796 31170.5 309.37 0.983499 0.319146 0.737186 0.737181 9.99958 2.98614e-06 1.19445e-05 0.133961 0.983386 0.931429 -0.0132917 4.92862e-06 0.514712 -2.00243e-20 7.42511e-24 -2.00169e-20 0.00139638 0.997815 8.60176e-05 0.152722 2.85273 0.00139638 0.997815 0.784899 0.0010664 0.00188129 0.000860176 0.455401 0.00188129 0.444116 0.000131082 1.02 0.888691 0.534397 0.287453 1.71927e-07 3.08266e-09 2371.96 3134.86 -0.0577711 0.482203 0.277294 0.254512 -0.593123 -0.169569 0.488996 -0.265937 -0.223068 2.59 1 0 295.733 0 2.22515 2.588 0.000299201 0.865099 0.697271 0.31863 0.432665 2.22533 138.647 83.6923 18.7077 60.7563 0.00403472 0 -40 10
1.689 4.88643e-08 2.53982e-06 0.144981 0.144981 0.0120273 2.22111e-05 0.00115446 0.181227 0.000658776 0.181881 0.945394 101.485 0.235722 0.845539 4.51532 0.0642778 0.0425974 0.957403 0.019472 0.00456856 0.0187298 0.00436067 0.00552801 0.00627016 0.22112 0.250806 58.0452 -87.8989 126.172 15.9374 145.035 0.00014211 0.267303 192.737 0.310219 0.0673284 0.00409829 0.000562336 0.00138496 0.986961 0.991717 -2.98917e-06 -85.6576 0.0930797 31170.4 309.382 0.983499 0.319146 0.737197 0.737193 9.99958 2.98614e-06 1.19445e-05 0.133965 0.983387 0.931428 -0.0132917 4.92865e-06 0.514731 -2.00259e-20 7.42572e-24 -2.00185e-20 0.00139638 0.997815 8.60176e-05 0.152722 2.85273 0.00139638 0.997815 0.784974 0.00106641 0.0018813 0.000860176 0.455401 0.00188129 0.444121 0.000131084 1.02 0.888692 0.534397 0.287454 1.71927e-07 3.08268e-09 2371.94 3134.91 -0.057776 0.482203 0.277294 0.254515 -0.593122 -0.169569 0.488981 -0.265935 -0.223055 2.591 1 0 295.729 0 2.22529 2.589 0.0002992 0.865126 0.697314 0.318587 0.432688 2.22547 138.654 83.6917 18.7076 60.756 0.00403475 0 -40 10
1.69 4.88932e-08 2.53982e-06 0.145016 0.145016 0.0120273 2.22242e-05 0.00115446 0.18127 0.000658777 0.181924 0.945483 101.484 0.235712 0.845671 4.51592 0.0642884 0.042603 0.957397 0.0194714 0.004569 0.0187293 0.00436105 0.00552855 0.00627071 0.221142 0.250829 58.0452 -87.8989 126.171 15.9374 145.035 0.000142113 0.267303 192.737 0.310219 0.0673283 0.00409829 0.000562337 0.00138496 0.986961 0.991717 -2.98918e-06 -85.6576 0.0930798 31170.4 309.394 0.983499 0.319146 0.737209 0.737204 9.99958 2.98615e-06 1.19445e-05 0.13397 0.983387 0.931427 -0.0132917 4.92867e-06 0.51475 -2.00274e-20 7.42634e-24 -2.002e-20 0.00139638 0.997815 8.60177e-05 0.152722 2.85273 0.00139638 0.997815 0.785048 0.00106643 0.0018813 0.000860177 0.455401 0.0018813 0.444127 0.000131087 1.02 0.888693 0.534397 0.287456 1.71928e-07 3.08271e-09 2371.93 3134.96 -0.0577809 0.482203 0.277293 0.254518 -0.593121 -0.169569 0.488965 -0.265933 -0.223041 2.592 1 0 295.724 0 2.22543 2.59 0.000299199 0.865154 0.697357 0.318544 0.43271 2.22561 138.662 83.6911 18.7076 60.7558 0.00403477 0 -40 10
1.691 4.8922e-08 2.53982e-06 0.145051 0.14505 0.0120273 2.22373e-05 0.00115446 0.181314 0.000658778 0.181968 0.945572 101.483 0.235701 0.845803 4.51651 0.0642991 0.0426086 0.957391 0.0194709 0.00456944 0.0187287 0.00436143 0.00552909 0.00627127 0.221164 0.250851 58.0453 -87.8989 126.171 15.9374 145.035 0.000142115 0.267303 192.737 0.310219 0.0673283 0.0040983 0.000562337 0.00138496 0.986961 0.991717 -2.9892e-06 -85.6576 0.0930799 31170.4 309.406 0.983499 0.319146 0.73722 0.737216 9.99958 2.98615e-06 1.19445e-05 0.133974 0.983388 0.931426 -0.0132917 4.9287e-06 0.51477 -2.00289e-20 7.42695e-24 -2.00215e-20 0.00139639 0.997815 8.60178e-05 0.152722 2.85273 0.00139639 0.997815 0.785123 0.00106645 0.0018813 0.000860178 0.455401 0.0018813 0.444132 0.000131089 1.02 0.888694 0.534396 0.287458 1.71928e-07 3.08273e-09 2371.91 3135.01 -0.0577859 0.482203 0.277293 0.254521 -0.593121 -0.169569 0.488949 -0.265931 -0.223028 2.593 1 0 295.72 0 2.22556 2.591 0.000299198 0.865182 0.6974 0.318501 0.432732 2.22575 138.669 83.6906 18.7076 60.7555 0.00403479 0 -40 10
1.692 4.89509e-08 2.53982e-06 0.145086 0.145085 0.0120273 2.22504e-05 0.00115447 0.181357 0.000658778 0.182011 0.945661 101.483 0.23569 0.845934 4.51711 0.0643097 0.0426142 0.957386 0.0194704 0.00456988 0.0187282 0.00436181 0.00552964 0.00627183 0.221185 0.250873 58.0453 -87.8989 126.171 15.9373 145.035 0.000142117 0.267304 192.737 0.310218 0.0673282 0.0040983 0.000562338 0.00138496 0.986961 0.991717 -2.98921e-06 -85.6576 0.09308 31170.4 309.418 0.983499 0.319146 0.737232 0.737228 9.99958 2.98616e-06 1.19445e-05 0.133979 0.983388 0.931425 -0.0132917 4.92873e-06 0.514789 -2.00305e-20 7.42756e-24 -2.0023e-20 0.00139639 0.997815 8.60179e-05 0.152723 2.85273 0.00139639 0.997815 0.785197 0.00106646 0.0018813 0.000860179 0.455401 0.0018813 0.444137 0.000131092 1.02 0.888695 0.534396 0.287459 1.71928e-07 3.08275e-09 2371.89 3135.05 -0.0577908 0.482203 0.277293 0.254525 -0.59312 -0.169569 0.488934 -0.265929 -0.223014 2.594 1 0 295.715 0 2.2257 2.592 0.000299196 0.865209 0.697443 0.318458 0.432755 2.22588 138.677 83.69 18.7075 60.7552 0.00403482 0 -40 10
1.693 4.89797e-08 2.53983e-06 0.14512 0.14512 0.0120273 2.22635e-05 0.00115447 0.181401 0.000658779 0.182055 0.94575 101.482 0.23568 0.846066 4.5177 0.0643204 0.0426199 0.95738 0.0194698 0.00457032 0.0187276 0.00436219 0.00553018 0.00627239 0.221207 0.250895 58.0454 -87.8989 126.171 15.9373 145.035 0.000142119 0.267304 192.737 0.310218 0.0673281 0.0040983 0.000562339 0.00138496 0.986961 0.991717 -2.98923e-06 -85.6576 0.0930801 31170.4 309.429 0.983499 0.319146 0.737244 0.737239 9.99958 2.98616e-06 1.19445e-05 0.133983 0.983388 0.931424 -0.0132917 4.92876e-06 0.514808 -2.0032e-20 7.42818e-24 -2.00246e-20 0.00139639 0.997815 8.6018e-05 0.152723 2.85273 0.00139639 0.997815 0.785272 0.00106648 0.0018813 0.00086018 0.4554 0.0018813 0.444143 0.000131094 1.02 0.888696 0.534396 0.287461 1.71929e-07 3.08278e-09 2371.88 3135.1 -0.0577957 0.482203 0.277293 0.254528 -0.59312 -0.16957 0.488918 -0.265927 -0.223 2.595 1 0 295.711 0 2.22584 2.593 0.000299195 0.865237 0.697487 0.318415 0.432777 2.22602 138.684 83.6894 18.7075 60.7549 0.00403484 0 -40 10
1.694 4.90086e-08 2.53983e-06 0.145155 0.145155 0.0120273 2.22766e-05 0.00115447 0.181444 0.000658779 0.182098 0.945839 101.482 0.235669 0.846198 4.5183 0.064331 0.0426255 0.957375 0.0194693 0.00457076 0.0187271 0.00436257 0.00553072 0.00627294 0.221229 0.250918 58.0455 -87.8989 126.171 15.9372 145.035 0.000142122 0.267304 192.737 0.310217 0.0673281 0.00409831 0.000562339 0.00138497 0.986961 0.991717 -2.98924e-06 -85.6576 0.0930802 31170.3 309.441 0.983499 0.319146 0.737255 0.737251 9.99958 2.98617e-06 1.19446e-05 0.133988 0.983389 0.931423 -0.0132917 4.92879e-06 0.514827 -2.00335e-20 7.42879e-24 -2.00261e-20 0.00139639 0.997815 8.6018e-05 0.152723 2.85273 0.00139639 0.997815 0.785346 0.0010665 0.0018813 0.00086018 0.4554 0.0018813 0.444148 0.000131096 1.02 0.888698 0.534396 0.287462 1.71929e-07 3.0828e-09 2371.86 3135.15 -0.0578007 0.482203 0.277292 0.254531 -0.593119 -0.16957 0.488902 -0.265925 -0.222987 2.596 1 0 295.706 0 2.22598 2.594 0.000299194 0.865265 0.69753 0.318372 0.432799 2.22616 138.691 83.6888 18.7075 60.7547 0.00403486 0 -40 10
1.695 4.90374e-08 2.53983e-06 0.14519 0.145189 0.0120272 2.22897e-05 0.00115447 0.181487 0.00065878 0.182141 0.945928 101.481 0.235658 0.846329 4.5189 0.0643417 0.0426311 0.957369 0.0194687 0.0045712 0.0187265 0.00436295 0.00553127 0.0062735 0.221251 0.25094 58.0455 -87.8989 126.17 15.9372 145.035 0.000142124 0.267304 192.736 0.310217 0.067328 0.00409831 0.00056234 0.00138497 0.986961 0.991717 -2.98926e-06 -85.6576 0.0930803 31170.3 309.453 0.983499 0.319146 0.737267 0.737263 9.99958 2.98617e-06 1.19446e-05 0.133992 0.983389 0.931422 -0.0132917 4.92882e-06 0.514846 -2.00351e-20 7.4294e-24 -2.00276e-20 0.00139639 0.997815 8.60181e-05 0.152723 2.85273 0.00139639 0.997815 0.785421 0.00106651 0.0018813 0.000860181 0.4554 0.0018813 0.444154 0.000131099 1.02 0.888699 0.534395 0.287464 1.71929e-07 3.08282e-09 2371.84 3135.2 -0.0578056 0.482203 0.277292 0.254534 -0.593118 -0.16957 0.488886 -0.265923 -0.222973 2.597 1 0 295.702 0 2.22612 2.595 0.000299193 0.865292 0.697573 0.318329 0.432822 2.2263 138.699 83.6883 18.7074 60.7544 0.00403489 0 -40 10
1.696 4.90663e-08 2.53983e-06 0.145224 0.145224 0.0120272 2.23029e-05 0.00115447 0.181531 0.00065878 0.182185 0.946018 101.481 0.235648 0.846461 4.5195 0.0643523 0.0426368 0.957363 0.0194682 0.00457164 0.0187259 0.00436333 0.00553181 0.00627406 0.221272 0.250962 58.0456 -87.8989 126.17 15.9372 145.035 0.000142126 0.267304 192.736 0.310216 0.067328 0.00409831 0.000562341 0.00138497 0.986961 0.991717 -2.98927e-06 -85.6576 0.0930803 31170.3 309.465 0.983499 0.319146 0.737279 0.737274 9.99958 2.98618e-06 1.19446e-05 0.133997 0.983389 0.931421 -0.0132917 4.92885e-06 0.514865 -2.00366e-20 7.43002e-24 -2.00292e-20 0.00139639 0.997815 8.60182e-05 0.152723 2.85274 0.00139639 0.997815 0.785495 0.00106653 0.00188131 0.000860182 0.4554 0.0018813 0.444159 0.000131101 1.02 0.8887 0.534395 0.287465 1.71929e-07 3.08284e-09 2371.83 3135.25 -0.0578105 0.482203 0.277292 0.254537 -0.593118 -0.16957 0.488871 -0.265921 -0.22296 2.598 1 0 295.697 0 2.22625 2.596 0.000299192 0.86532 0.697616 0.318286 0.432844 2.22643 138.706 83.6877 18.7074 60.7541 0.00403491 0 -40 10
1.697 4.90951e-08 2.53983e-06 0.145259 0.145258 0.0120272 2.2316e-05 0.00115447 0.181574 0.000658781 0.182228 0.946107 101.48 0.235637 0.846593 4.52009 0.064363 0.0426424 0.957358 0.0194676 0.00457208 0.0187254 0.00436371 0.00553235 0.00627462 0.221294 0.250985 58.0457 -87.8989 126.17 15.9371 145.035 0.000142128 0.267305 192.736 0.310216 0.0673279 0.00409831 0.000562341 0.00138497 0.986961 0.991717 -2.98929e-06 -85.6576 0.0930804 31170.3 309.477 0.983499 0.319146 0.73729 0.737286 9.99958 2.98618e-06 1.19446e-05 0.134001 0.98339 0.93142 -0.0132917 4.92888e-06 0.514884 -2.00381e-20 7.43063e-24 -2.00307e-20 0.00139639 0.997815 8.60183e-05 0.152723 2.85274 0.00139639 0.997815 0.78557 0.00106654 0.00188131 0.000860183 0.455399 0.00188131 0.444164 0.000131104 1.02 0.888701 0.534395 0.287467 1.7193e-07 3.08287e-09 2371.81 3135.3 -0.0578155 0.482203 0.277291 0.25454 -0.593117 -0.16957 0.488855 -0.265919 -0.222946 2.599 1 0 295.693 0 2.22639 2.597 0.000299191 0.865348 0.697659 0.318243 0.432867 2.22657 138.713 83.6871 18.7074 60.7538 0.00403494 0 -40 10
1.698 4.9124e-08 2.53983e-06 0.145294 0.145293 0.0120272 2.23291e-05 0.00115447 0.181617 0.000658782 0.182271 0.946196 101.479 0.235626 0.846724 4.52069 0.0643737 0.042648 0.957352 0.0194671 0.00457252 0.0187248 0.00436409 0.0055329 0.00627518 0.221316 0.251007 58.0457 -87.8989 126.17 15.9371 145.035 0.00014213 0.267305 192.736 0.310216 0.0673279 0.00409832 0.000562342 0.00138497 0.986961 0.991717 -2.9893e-06 -85.6575 0.0930805 31170.2 309.489 0.983499 0.319146 0.737302 0.737297 9.99958 2.98619e-06 1.19446e-05 0.134006 0.98339 0.931419 -0.0132917 4.92891e-06 0.514903 -2.00397e-20 7.43125e-24 -2.00322e-20 0.00139639 0.997815 8.60184e-05 0.152723 2.85274 0.00139639 0.997815 0.785644 0.00106656 0.00188131 0.000860184 0.455399 0.00188131 0.44417 0.000131106 1.02 0.888702 0.534394 0.287468 1.7193e-07 3.08289e-09 2371.79 3135.35 -0.0578204 0.482203 0.277291 0.254543 -0.593116 -0.16957 0.488839 -0.265916 -0.222932 2.6 1 0 295.688 0 2.22653 2.598 0.000299189 0.865375 0.697702 0.3182 0.432889 2.22671 138.721 83.6866 18.7073 60.7536 0.00403496 0 -40 10
1.699 4.91528e-08 2.53984e-06 0.145328 0.145328 0.0120272 2.23422e-05 0.00115447 0.18166 0.000658782 0.182314 0.946285 101.479 0.235616 0.846856 4.52129 0.0643843 0.0426537 0.957346 0.0194666 0.00457297 0.0187243 0.00436447 0.00553344 0.00627574 0.221338 0.251029 58.0458 -87.8989 126.17 15.9371 145.035 0.000142133 0.267305 192.736 0.310215 0.0673278 0.00409832 0.000562343 0.00138498 0.986961 0.991717 -2.98932e-06 -85.6575 0.0930806 31170.2 309.501 0.983499 0.319146 0.737313 0.737309 9.99958 2.98619e-06 1.19447e-05 0.13401 0.98339 0.931418 -0.0132917 4.92894e-06 0.514923 -2.00412e-20 7.43186e-24 -2.00338e-20 0.00139639 0.997815 8.60184e-05 0.152724 2.85274 0.00139639 0.997815 0.785718 0.00106658 0.00188131 0.000860184 0.455399 0.00188131 0.444175 0.000131109 1.02 0.888703 0.534394 0.28747 1.7193e-07 3.08291e-09 2371.78 3135.4 -0.0578253 0.482203 0.277291 0.254546 -0.593116 -0.16957 0.488824 -0.265914 -0.222919 2.601 1 0 295.684 0 2.22667 2.599 0.000299188 0.865403 0.697746 0.318158 0.432911 2.22685 138.728 83.686 18.7073 60.7533 0.00403498 0 -40 10
1.7 4.91817e-08 2.53984e-06 0.145363 0.145362 0.0120272 2.23553e-05 0.00115447 0.181703 0.000658783 0.182358 0.946375 101.478 0.235605 0.846988 4.52189 0.064395 0.0426593 0.957341 0.019466 0.00457341 0.0187237 0.00436485 0.00553399 0.0062763 0.221359 0.251052 58.0458 -87.8989 126.169 15.937 145.035 0.000142135 0.267305 192.736 0.310215 0.0673278 0.00409832 0.000562343 0.00138498 0.986961 0.991717 -2.98933e-06 -85.6575 0.0930807 31170.2 309.513 0.983499 0.319146 0.737325 0.737321 9.99958 2.9862e-06 1.19447e-05 0.134015 0.983391 0.931417 -0.0132917 4.92897e-06 0.514942 -2.00427e-20 7.43248e-24 -2.00353e-20 0.0013964 0.997815 8.60185e-05 0.152724 2.85274 0.0013964 0.997815 0.785793 0.00106659 0.00188131 0.000860185 0.455399 0.00188131 0.44418 0.000131111 1.02 0.888704 0.534394 0.287471 1.7193e-07 3.08294e-09 2371.76 3135.44 -0.0578303 0.482204 0.277291 0.25455 -0.593115 -0.16957 0.488808 -0.265912 -0.222905 2.602 1 0 295.68 0 2.2268 2.6 0.000299187 0.865431 0.697789 0.318115 0.432934 2.22699 138.736 83.6854 18.7073 60.753 0.00403501 0 -40 10
1.701 4.92105e-08 2.53984e-06 0.145397 0.145397 0.0120272 2.23684e-05 0.00115447 0.181746 0.000658783 0.182401 0.946464 101.478 0.235594 0.84712 4.52249 0.0644057 0.042665 0.957335 0.0194655 0.00457385 0.0187231 0.00436524 0.00553453 0.00627686 0.221381 0.251074 58.0459 -87.8989 126.169 15.937 145.035 0.000142137 0.267305 192.735 0.310214 0.0673277 0.00409833 0.000562344 0.00138498 0.986961 0.991717 -2.98935e-06 -85.6575 0.0930808 31170.2 309.525 0.983499 0.319146 0.737337 0.737332 9.99958 2.9862e-06 1.19447e-05 0.134019 0.983391 0.931416 -0.0132917 4.929e-06 0.514961 -2.00443e-20 7.43309e-24 -2.00368e-20 0.0013964 0.997815 8.60186e-05 0.152724 2.85274 0.0013964 0.997815 0.785867 0.00106661 0.00188131 0.000860186 0.455399 0.00188131 0.444186 0.000131114 1.02 0.888705 0.534393 0.287473 1.71931e-07 3.08296e-09 2371.75 3135.49 -0.0578352 0.482204 0.27729 0.254553 -0.593115 -0.16957 0.488792 -0.26591 -0.222891 2.603 1 0 295.675 0 2.22694 2.601 0.000299186 0.865459 0.697832 0.318072 0.432956 2.22712 138.743 83.6848 18.7072 60.7527 0.00403503 0 -40 10
1.702 4.92394e-08 2.53984e-06 0.145432 0.145431 0.0120271 2.23815e-05 0.00115447 0.18179 0.000658784 0.182444 0.946553 101.477 0.235584 0.847252 4.52309 0.0644163 0.0426707 0.957329 0.0194649 0.00457429 0.0187226 0.00436562 0.00553508 0.00627742 0.221403 0.251097 58.046 -87.899 126.169 15.9369 145.035 0.000142139 0.267305 192.735 0.310214 0.0673277 0.00409833 0.000562345 0.00138498 0.986961 0.991717 -2.98936e-06 -85.6575 0.0930809 31170.2 309.537 0.983499 0.319146 0.737348 0.737344 9.99958 2.98621e-06 1.19447e-05 0.134024 0.983391 0.931415 -0.0132917 4.92903e-06 0.51498 -2.00458e-20 7.43371e-24 -2.00384e-20 0.0013964 0.997815 8.60187e-05 0.152724 2.85274 0.0013964 0.997815 0.785941 0.00106663 0.00188132 0.000860187 0.455398 0.00188131 0.444191 0.000131116 1.02 0.888706 0.534393 0.287474 1.71931e-07 3.08298e-09 2371.73 3135.54 -0.0578402 0.482204 0.27729 0.254556 -0.593114 -0.16957 0.488776 -0.265908 -0.222878 2.604 1 0 295.671 0 2.22708 2.602 0.000299185 0.865487 0.697875 0.318029 0.432978 2.22726 138.75 83.6843 18.7072 60.7525 0.00403505 0 -40 10
1.703 4.92682e-08 2.53984e-06 0.145466 0.145466 0.0120271 2.23947e-05 0.00115447 0.181833 0.000658784 0.182487 0.946642 101.476 0.235573 0.847383 4.52369 0.064427 0.0426763 0.957324 0.0194644 0.00457474 0.018722 0.004366 0.00553562 0.00627798 0.221425 0.251119 58.046 -87.899 126.169 15.9369 145.035 0.000142142 0.267306 192.735 0.310213 0.0673276 0.00409833 0.000562345 0.00138499 0.986961 0.991717 -2.98938e-06 -85.6575 0.093081 31170.1 309.549 0.983499 0.319146 0.73736 0.737356 9.99958 2.98621e-06 1.19447e-05 0.134028 0.983392 0.931414 -0.0132917 4.92906e-06 0.514999 -2.00474e-20 7.43433e-24 -2.00399e-20 0.0013964 0.997815 8.60188e-05 0.152724 2.85274 0.0013964 0.997815 0.786016 0.00106664 0.00188132 0.000860188 0.455398 0.00188132 0.444196 0.000131118 1.02 0.888707 0.534393 0.287476 1.71931e-07 3.08301e-09 2371.71 3135.59 -0.0578451 0.482204 0.27729 0.254559 -0.593113 -0.16957 0.488761 -0.265906 -0.222864 2.605 1 0 295.666 0 2.22722 2.603 0.000299184 0.865514 0.697918 0.317987 0.433001 2.2274 138.758 83.6837 18.7072 60.7522 0.00403508 0 -40 10
1.704 4.92971e-08 2.53984e-06 0.1455 0.1455 0.0120271 2.24078e-05 0.00115447 0.181876 0.000658785 0.18253 0.946732 101.476 0.235562 0.847515 4.52429 0.0644377 0.042682 0.957318 0.0194638 0.00457518 0.0187215 0.00436638 0.00553617 0.00627854 0.221447 0.251142 58.0461 -87.899 126.168 15.9369 145.035 0.000142144 0.267306 192.735 0.310213 0.0673276 0.00409834 0.000562346 0.00138499 0.986961 0.991717 -2.98939e-06 -85.6575 0.093081 31170.1 309.562 0.983499 0.319146 0.737372 0.737367 9.99958 2.98622e-06 1.19448e-05 0.134033 0.983392 0.931413 -0.0132917 4.92909e-06 0.515018 -2.00489e-20 7.43494e-24 -2.00415e-20 0.0013964 0.997815 8.60189e-05 0.152724 2.85274 0.0013964 0.997815 0.78609 0.00106666 0.00188132 0.000860189 0.455398 0.00188132 0.444202 0.000131121 1.02 0.888709 0.534392 0.287477 1.71932e-07 3.08303e-09 2371.7 3135.64 -0.0578501 0.482204 0.277289 0.254562 -0.593113 -0.16957 0.488745 -0.265904 -0.22285 2.606 1 0 295.662 0 2.22735 2.604 0.000299183 0.865542 0.697961 0.317944 0.433023 2.22754 138.765 83.6831 18.7071 60.7519 0.0040351 0 -40 10
1.705 4.93259e-08 2.53984e-06 0.145535 0.145534 0.0120271 2.24209e-05 0.00115447 0.181919 0.000658785 0.182573 0.946821 101.475 0.235552 0.847647 4.52489 0.0644483 0.0426877 0.957312 0.0194633 0.00457562 0.0187209 0.00436676 0.00553671 0.0062791 0.221469 0.251164 58.0462 -87.899 126.168 15.9368 145.035 0.000142146 0.267306 192.735 0.310213 0.0673275 0.00409834 0.000562347 0.00138499 0.986961 0.991717 -2.98941e-06 -85.6575 0.0930811 31170.1 309.574 0.983498 0.319146 0.737383 0.737379 9.99958 2.98622e-06 1.19448e-05 0.134037 0.983392 0.931412 -0.0132917 4.92912e-06 0.515038 -2.00504e-20 7.43556e-24 -2.0043e-20 0.0013964 0.997815 8.60189e-05 0.152725 2.85274 0.0013964 0.997815 0.786164 0.00106668 0.00188132 0.000860189 0.455398 0.00188132 0.444207 0.000131123 1.02 0.88871 0.534392 0.287479 1.71932e-07 3.08305e-09 2371.68 3135.69 -0.057855 0.482204 0.277289 0.254565 -0.593112 -0.16957 0.488729 -0.265902 -0.222837 2.607 1 0 295.657 0 2.22749 2.605 0.000299181 0.86557 0.698004 0.317902 0.433045 2.22767 138.773 83.6825 18.7071 60.7516 0.00403513 0 -40 10
1.706 4.93548e-08 2.53985e-06 0.145569 0.145569 0.0120271 2.2434e-05 0.00115448 0.181962 0.000658786 0.182616 0.94691 101.475 0.235541 0.847779 4.5255 0.064459 0.0426934 0.957307 0.0194627 0.00457606 0.0187203 0.00436715 0.00553726 0.00627966 0.22149 0.251186 58.0462 -87.899 126.168 15.9368 145.035 0.000142148 0.267306 192.735 0.310212 0.0673275 0.00409834 0.000562347 0.00138499 0.986961 0.991717 -2.98943e-06 -85.6575 0.0930812 31170.1 309.586 0.983498 0.319146 0.737395 0.737391 9.99958 2.98623e-06 1.19448e-05 0.134042 0.983393 0.931411 -0.0132917 4.92915e-06 0.515057 -2.0052e-20 7.43618e-24 -2.00445e-20 0.0013964 0.997815 8.6019e-05 0.152725 2.85274 0.0013964 0.997815 0.786238 0.00106669 0.00188132 0.00086019 0.455397 0.00188132 0.444212 0.000131126 1.02 0.888711 0.534392 0.28748 1.71932e-07 3.08307e-09 2371.66 3135.74 -0.0578599 0.482204 0.277289 0.254568 -0.593111 -0.16957 0.488713 -0.2659 -0.222823 2.608 1 0 295.653 0 2.22763 2.606 0.00029918 0.865598 0.698048 0.317859 0.433068 2.22781 138.78 83.682 18.7071 60.7513 0.00403515 0 -40 10
1.707 4.93836e-08 2.53985e-06 0.145604 0.145603 0.0120271 2.24471e-05 0.00115448 0.182004 0.000658787 0.182659 0.947 101.474 0.23553 0.847911 4.5261 0.0644697 0.042699 0.957301 0.0194622 0.00457651 0.0187198 0.00436753 0.00553781 0.00628022 0.221512 0.251209 58.0463 -87.899 126.168 15.9368 145.035 0.000142151 0.267306 192.735 0.310212 0.0673274 0.00409835 0.000562348 0.00138499 0.986961 0.991717 -2.98944e-06 -85.6575 0.0930813 31170 309.598 0.983498 0.319146 0.737407 0.737402 9.99958 2.98623e-06 1.19448e-05 0.134046 0.983393 0.93141 -0.0132917 4.92918e-06 0.515076 -2.00535e-20 7.43679e-24 -2.00461e-20 0.0013964 0.997815 8.60191e-05 0.152725 2.85275 0.0013964 0.997815 0.786312 0.00106671 0.00188132 0.000860191 0.455397 0.00188132 0.444218 0.000131128 1.02 0.888712 0.534392 0.287482 1.71932e-07 3.0831e-09 2371.65 3135.79 -0.0578649 0.482204 0.277289 0.254572 -0.593111 -0.16957 0.488698 -0.265898 -0.22281 2.609 1 0 295.648 0 2.22777 2.607 0.000299179 0.865626 0.698091 0.317817 0.43309 2.22795 138.787 83.6814 18.707 60.7511 0.00403517 0 -40 10
1.708 4.94125e-08 2.53985e-06 0.145638 0.145637 0.0120271 2.24602e-05 0.00115448 0.182047 0.000658787 0.182701 0.947089 101.473 0.23552 0.848043 4.5267 0.0644804 0.0427047 0.957295 0.0194616 0.00457695 0.0187192 0.00436791 0.00553835 0.00628079 0.221534 0.251231 58.0463 -87.899 126.168 15.9367 145.035 0.000142153 0.267307 192.734 0.310211 0.0673274 0.00409835 0.000562349 0.001385 0.986961 0.991717 -2.98946e-06 -85.6575 0.0930814 31170 309.61 0.983498 0.319146 0.737418 0.737414 9.99958 2.98624e-06 1.19448e-05 0.134051 0.983393 0.93141 -0.0132917 4.92921e-06 0.515095 -2.00551e-20 7.43741e-24 -2.00476e-20 0.00139641 0.997815 8.60192e-05 0.152725 2.85275 0.00139641 0.997815 0.786386 0.00106672 0.00188132 0.000860192 0.455397 0.00188132 0.444223 0.000131131 1.02 0.888713 0.534391 0.287483 1.71933e-07 3.08312e-09 2371.63 3135.84 -0.0578698 0.482204 0.277288 0.254575 -0.59311 -0.16957 0.488682 -0.265895 -0.222796 2.61 1 0 295.644 0 2.22791 2.608 0.000299178 0.865654 0.698134 0.317774 0.433112 2.22809 138.795 83.6808 18.707 60.7508 0.0040352 0 -40 10
1.709 4.94413e-08 2.53985e-06 0.145672 0.145672 0.012027 2.24733e-05 0.00115448 0.18209 0.000658788 0.182744 0.947178 101.473 0.235509 0.848175 4.52731 0.064491 0.0427104 0.95729 0.0194611 0.0045774 0.0187187 0.00436829 0.0055389 0.00628135 0.221556 0.251254 58.0464 -87.899 126.167 15.9367 145.035 0.000142155 0.267307 192.734 0.310211 0.0673273 0.00409835 0.00056235 0.001385 0.986961 0.991717 -2.98947e-06 -85.6574 0.0930815 31170 309.622 0.983498 0.319146 0.73743 0.737426 9.99958 2.98624e-06 1.19449e-05 0.134055 0.983394 0.931409 -0.0132917 4.92924e-06 0.515115 -2.00566e-20 7.43803e-24 -2.00492e-20 0.00139641 0.997815 8.60193e-05 0.152725 2.85275 0.00139641 0.997815 0.786461 0.00106674 0.00188133 0.000860193 0.455397 0.00188132 0.444228 0.000131133 1.02 0.888714 0.534391 0.287485 1.71933e-07 3.08314e-09 2371.61 3135.88 -0.0578748 0.482204 0.277288 0.254578 -0.59311 -0.169571 0.488666 -0.265893 -0.222782 2.611 1 0 295.639 0 2.22804 2.609 0.000299177 0.865681 0.698177 0.317732 0.433135 2.22822 138.802 83.6802 18.707 60.7505 0.00403522 0 -40 10
1.71 4.94702e-08 2.53985e-06 0.145706 0.145706 0.012027 2.24864e-05 0.00115448 0.182133 0.000658788 0.182787 0.947268 101.472 0.235498 0.848307 4.52791 0.0645017 0.0427161 0.957284 0.0194606 0.00457784 0.0187181 0.00436868 0.00553945 0.00628191 0.221578 0.251276 58.0465 -87.899 126.167 15.9366 145.035 0.000142157 0.267307 192.734 0.31021 0.0673272 0.00409835 0.00056235 0.001385 0.986961 0.991717 -2.98949e-06 -85.6574 0.0930816 31170 309.634 0.983498 0.319146 0.737442 0.737437 9.99958 2.98625e-06 1.19449e-05 0.13406 0.983394 0.931408 -0.0132917 4.92927e-06 0.515134 -2.00582e-20 7.43865e-24 -2.00507e-20 0.00139641 0.997815 8.60193e-05 0.152725 2.85275 0.00139641 0.997815 0.786535 0.00106676 0.00188133 0.000860193 0.455396 0.00188133 0.444234 0.000131136 1.02 0.888715 0.534391 0.287486 1.71933e-07 3.08317e-09 2371.6 3135.93 -0.0578798 0.482204 0.277288 0.254581 -0.593109 -0.169571 0.48865 -0.265891 -0.222769 2.612 1 0 295.635 0 2.22818 2.61 0.000299176 0.865709 0.69822 0.31769 0.433157 2.22836 138.81 83.6797 18.7069 60.7502 0.00403524 0 -40 10
1.711 4.9499e-08 2.53985e-06 0.145741 0.14574 0.012027 2.24996e-05 0.00115448 0.182176 0.000658789 0.18283 0.947357 101.471 0.235488 0.848439 4.52851 0.0645124 0.0427218 0.957278 0.01946 0.00457828 0.0187175 0.00436906 0.00554 0.00628247 0.2216 0.251299 58.0465 -87.899 126.167 15.9366 145.035 0.00014216 0.267307 192.734 0.31021 0.0673272 0.00409836 0.000562351 0.001385 0.986961 0.991717 -2.9895e-06 -85.6574 0.0930817 31169.9 309.646 0.983498 0.319146 0.737453 0.737449 9.99958 2.98625e-06 1.19449e-05 0.134064 0.983394 0.931407 -0.0132917 4.9293e-06 0.515153 -2.00597e-20 7.43927e-24 -2.00523e-20 0.00139641 0.997815 8.60194e-05 0.152725 2.85275 0.00139641 0.997815 0.786609 0.00106677 0.00188133 0.000860194 0.455396 0.00188133 0.444239 0.000131138 1.02 0.888716 0.53439 0.287488 1.71933e-07 3.08319e-09 2371.58 3135.98 -0.0578847 0.482204 0.277287 0.254584 -0.593108 -0.169571 0.488635 -0.265889 -0.222755 2.613 1 0 295.631 0 2.22832 2.611 0.000299174 0.865737 0.698263 0.317647 0.433179 2.2285 138.817 83.6791 18.7069 60.75 0.00403527 0 -40 10
1.712 4.95279e-08 2.53986e-06 0.145775 0.145774 0.012027 2.25127e-05 0.00115448 0.182218 0.000658789 0.182873 0.947447 101.471 0.235477 0.848571 4.52912 0.0645231 0.0427275 0.957272 0.0194595 0.00457873 0.018717 0.00436944 0.00554054 0.00628304 0.221622 0.251321 58.0466 -87.899 126.167 15.9366 145.035 0.000142162 0.267307 192.734 0.31021 0.0673271 0.00409836 0.000562352 0.00138501 0.986961 0.991717 -2.98952e-06 -85.6574 0.0930817 31169.9 309.658 0.983498 0.319146 0.737465 0.737461 9.99958 2.98626e-06 1.19449e-05 0.134069 0.983395 0.931406 -0.0132917 4.92933e-06 0.515172 -2.00612e-20 7.43988e-24 -2.00538e-20 0.00139641 0.997815 8.60195e-05 0.152726 2.85275 0.00139641 0.997815 0.786683 0.00106679 0.00188133 0.000860195 0.455396 0.00188133 0.444244 0.00013114 1.02 0.888717 0.53439 0.287489 1.71934e-07 3.08321e-09 2371.57 3136.03 -0.0578897 0.482204 0.277287 0.254587 -0.593108 -0.169571 0.488619 -0.265887 -0.222741 2.614 1 0 295.626 0 2.22846 2.612 0.000299173 0.865765 0.698306 0.317605 0.433201 2.22864 138.824 83.6785 18.7069 60.7497 0.00403529 0 -40 10
1.713 4.95567e-08 2.53986e-06 0.145809 0.145808 0.012027 2.25258e-05 0.00115448 0.182261 0.00065879 0.182915 0.947536 101.47 0.235466 0.848703 4.52972 0.0645338 0.0427332 0.957267 0.0194589 0.00457917 0.0187164 0.00436983 0.00554109 0.0062836 0.221644 0.251344 58.0467 -87.899 126.167 15.9365 145.035 0.000142164 0.267308 192.734 0.310209 0.0673271 0.00409836 0.000562352 0.00138501 0.986961 0.991717 -2.98953e-06 -85.6574 0.0930818 31169.9 309.67 0.983498 0.319146 0.737477 0.737472 9.99958 2.98626e-06 1.19449e-05 0.134073 0.983395 0.931405 -0.0132917 4.92936e-06 0.515192 -2.00628e-20 7.4405e-24 -2.00553e-20 0.00139641 0.997815 8.60196e-05 0.152726 2.85275 0.00139641 0.997815 0.786757 0.00106681 0.00188133 0.000860196 0.455396 0.00188133 0.444249 0.000131143 1.02 0.888718 0.53439 0.287491 1.71934e-07 3.08323e-09 2371.55 3136.08 -0.0578946 0.482205 0.277287 0.25459 -0.593107 -0.169571 0.488603 -0.265885 -0.222728 2.615 1 0 295.622 0 2.22859 2.613 0.000299172 0.865793 0.698349 0.317563 0.433224 2.22877 138.832 83.6779 18.7068 60.7494 0.00403532 0 -40 10
1.714 4.95856e-08 2.53986e-06 0.145843 0.145842 0.012027 2.25389e-05 0.00115448 0.182304 0.00065879 0.182958 0.947626 101.47 0.235456 0.848835 4.53033 0.0645444 0.042739 0.957261 0.0194584 0.00457962 0.0187158 0.00437021 0.00554164 0.00628416 0.221666 0.251367 58.0467 -87.899 126.166 15.9365 145.035 0.000142166 0.267308 192.733 0.310209 0.067327 0.00409837 0.000562353 0.00138501 0.986961 0.991717 -2.98955e-06 -85.6574 0.0930819 31169.9 309.682 0.983498 0.319146 0.737488 0.737484 9.99958 2.98627e-06 1.1945e-05 0.134078 0.983395 0.931404 -0.0132917 4.92939e-06 0.515211 -2.00643e-20 7.44112e-24 -2.00569e-20 0.00139641 0.997815 8.60197e-05 0.152726 2.85275 0.00139641 0.997815 0.786831 0.00106682 0.00188133 0.000860197 0.455396 0.00188133 0.444255 0.000131145 1.02 0.88872 0.534389 0.287492 1.71934e-07 3.08326e-09 2371.53 3136.13 -0.0578996 0.482205 0.277287 0.254594 -0.593107 -0.169571 0.488587 -0.265883 -0.222714 2.616 1 0 295.617 0 2.22873 2.614 0.000299171 0.865821 0.698392 0.317521 0.433246 2.22891 138.839 83.6774 18.7068 60.7491 0.00403534 0 -40 10
1.715 4.96144e-08 2.53986e-06 0.145877 0.145877 0.012027 2.2552e-05 0.00115448 0.182346 0.000658791 0.183001 0.947715 101.469 0.235445 0.848967 4.53094 0.0645551 0.0427447 0.957255 0.0194578 0.00458006 0.0187153 0.0043706 0.00554219 0.00628473 0.221688 0.251389 58.0468 -87.899 126.166 15.9365 145.035 0.000142169 0.267308 192.733 0.310208 0.067327 0.00409837 0.000562354 0.00138501 0.986961 0.991717 -2.98956e-06 -85.6574 0.093082 31169.9 309.694 0.983498 0.319146 0.7375 0.737496 9.99958 2.98627e-06 1.1945e-05 0.134083 0.983396 0.931403 -0.0132917 4.92942e-06 0.51523 -2.00659e-20 7.44174e-24 -2.00584e-20 0.00139641 0.997815 8.60197e-05 0.152726 2.85275 0.00139641 0.997815 0.786905 0.00106684 0.00188133 0.000860197 0.455395 0.00188133 0.44426 0.000131148 1.02 0.888721 0.534389 0.287494 1.71934e-07 3.08328e-09 2371.52 3136.18 -0.0579045 0.482205 0.277286 0.254597 -0.593106 -0.169571 0.488571 -0.265881 -0.2227 2.617 1 0 295.613 0 2.22887 2.615 0.00029917 0.865849 0.698436 0.317479 0.433268 2.22905 138.846 83.6768 18.7068 60.7488 0.00403536 0 -40 10
1.716 4.96433e-08 2.53986e-06 0.145911 0.145911 0.012027 2.25651e-05 0.00115448 0.182389 0.000658792 0.183043 0.947805 101.468 0.235434 0.849099 4.53154 0.0645658 0.0427504 0.95725 0.0194573 0.00458051 0.0187147 0.00437098 0.00554274 0.00628529 0.221709 0.251412 58.0468 -87.899 126.166 15.9364 145.035 0.000142171 0.267308 192.733 0.310208 0.0673269 0.00409837 0.000562354 0.00138501 0.986961 0.991717 -2.98958e-06 -85.6574 0.0930821 31169.8 309.706 0.983498 0.319146 0.737512 0.737507 9.99958 2.98628e-06 1.1945e-05 0.134087 0.983396 0.931402 -0.0132917 4.92945e-06 0.51525 -2.00674e-20 7.44236e-24 -2.006e-20 0.00139641 0.997815 8.60198e-05 0.152726 2.85275 0.00139641 0.997815 0.786979 0.00106686 0.00188134 0.000860198 0.455395 0.00188133 0.444265 0.00013115 1.02 0.888722 0.534389 0.287496 1.71935e-07 3.0833e-09 2371.5 3136.23 -0.0579095 0.482205 0.277286 0.2546 -0.593105 -0.169571 0.488556 -0.265879 -0.222686 2.618 1 0 295.608 0 2.22901 2.616 0.000299168 0.865877 0.698479 0.317436 0.433291 2.22919 138.854 83.6762 18.7067 60.7486 0.00403539 0 -40 10
1.717 4.96721e-08 2.53986e-06 0.145945 0.145945 0.0120269 2.25782e-05 0.00115448 0.182432 0.000658792 0.183086 0.947894 101.468 0.235423 0.849231 4.53215 0.0645765 0.0427561 0.957244 0.0194567 0.00458095 0.0187141 0.00437137 0.00554329 0.00628586 0.221731 0.251434 58.0469 -87.899 126.166 15.9364 145.035 0.000142173 0.267308 192.733 0.310207 0.0673269 0.00409838 0.000562355 0.00138502 0.986961 0.991717 -2.98959e-06 -85.6574 0.0930822 31169.8 309.718 0.983498 0.319146 0.737524 0.737519 9.99958 2.98628e-06 1.1945e-05 0.134092 0.983396 0.931401 -0.0132917 4.92948e-06 0.515269 -2.0069e-20 7.44298e-24 -2.00615e-20 0.00139642 0.997815 8.60199e-05 0.152726 2.85275 0.00139642 0.997815 0.787052 0.00106687 0.00188134 0.000860199 0.455395 0.00188134 0.444271 0.000131153 1.02 0.888723 0.534388 0.287497 1.71935e-07 3.08333e-09 2371.48 3136.28 -0.0579145 0.482205 0.277286 0.254603 -0.593105 -0.169571 0.48854 -0.265877 -0.222673 2.619 1 0 295.604 0 2.22914 2.617 0.000299167 0.865905 0.698522 0.317394 0.433313 2.22932 138.861 83.6756 18.7067 60.7483 0.00403541 0 -40 10
1.718 4.97009e-08 2.53987e-06 0.145979 0.145979 0.0120269 2.25913e-05 0.00115448 0.182474 0.000658793 0.183128 0.947984 101.467 0.235413 0.849363 4.53276 0.0645872 0.0427619 0.957238 0.0194562 0.0045814 0.0187136 0.00437175 0.00554384 0.00628642 0.221753 0.251457 58.047 -87.899 126.166 15.9364 145.035 0.000142175 0.267309 192.733 0.310207 0.0673268 0.00409838 0.000562356 0.00138502 0.986961 0.991717 -2.98961e-06 -85.6574 0.0930823 31169.8 309.731 0.983498 0.319146 0.737535 0.737531 9.99958 2.98629e-06 1.1945e-05 0.134096 0.983397 0.9314 -0.0132917 4.92951e-06 0.515288 -2.00705e-20 7.4436e-24 -2.00631e-20 0.00139642 0.997815 8.602e-05 0.152727 2.85276 0.00139642 0.997815 0.787126 0.00106689 0.00188134 0.0008602 0.455395 0.00188134 0.444276 0.000131155 1.02 0.888724 0.534388 0.287499 1.71935e-07 3.08335e-09 2371.47 3136.33 -0.0579194 0.482205 0.277286 0.254606 -0.593104 -0.169571 0.488524 -0.265874 -0.222659 2.62 1 0 295.599 0 2.22928 2.618 0.000299166 0.865933 0.698565 0.317352 0.433335 2.22946 138.869 83.675 18.7067 60.748 0.00403543 0 -40 10
1.719 4.97298e-08 2.53987e-06 0.146013 0.146013 0.0120269 2.26045e-05 0.00115448 0.182517 0.000658793 0.183171 0.948073 101.467 0.235402 0.849495 4.53336 0.0645979 0.0427676 0.957232 0.0194556 0.00458185 0.018713 0.00437214 0.00554439 0.00628699 0.221775 0.251479 58.047 -87.899 126.165 15.9363 145.035 0.000142178 0.267309 192.733 0.310207 0.0673268 0.00409838 0.000562356 0.00138502 0.986961 0.991717 -2.98962e-06 -85.6574 0.0930824 31169.8 309.743 0.983498 0.319146 0.737547 0.737543 9.99958 2.98629e-06 1.19451e-05 0.134101 0.983397 0.931399 -0.0132917 4.92953e-06 0.515308 -2.00721e-20 7.44422e-24 -2.00646e-20 0.00139642 0.997815 8.60201e-05 0.152727 2.85276 0.00139642 0.997815 0.7872 0.0010669 0.00188134 0.000860201 0.455394 0.00188134 0.444281 0.000131158 1.02 0.888725 0.534388 0.2875 1.71936e-07 3.08337e-09 2371.45 3136.37 -0.0579244 0.482205 0.277285 0.254609 -0.593103 -0.169571 0.488508 -0.265872 -0.222645 2.621 1 0 295.595 0 2.22942 2.619 0.000299165 0.865961 0.698608 0.31731 0.433358 2.2296 138.876 83.6745 18.7066 60.7477 0.00403546 0 -40 10
1.72 4.97586e-08 2.53987e-06 0.146047 0.146047 0.0120269 2.26176e-05 0.00115449 0.182559 0.000658794 0.183213 0.948163 101.466 0.235391 0.849627 4.53397 0.0646086 0.0427733 0.957227 0.0194551 0.00458229 0.0187124 0.00437252 0.00554493 0.00628755 0.221797 0.251502 58.0471 -87.899 126.165 15.9363 145.035 0.00014218 0.267309 192.732 0.310206 0.0673267 0.00409838 0.000562357 0.00138502 0.986961 0.991717 -2.98964e-06 -85.6573 0.0930824 31169.7 309.755 0.983498 0.319146 0.737559 0.737554 9.99958 2.9863e-06 1.19451e-05 0.134105 0.983397 0.931398 -0.0132916 4.92956e-06 0.515327 -2.00736e-20 7.44484e-24 -2.00662e-20 0.00139642 0.997815 8.60201e-05 0.152727 2.85276 0.00139642 0.997815 0.787274 0.00106692 0.00188134 0.000860201 0.455394 0.00188134 0.444287 0.00013116 1.02 0.888726 0.534388 0.287502 1.71936e-07 3.08339e-09 2371.43 3136.42 -0.0579294 0.482205 0.277285 0.254612 -0.593103 -0.169571 0.488493 -0.26587 -0.222632 2.622 1 0 295.59 0 2.22956 2.62 0.000299164 0.865989 0.698651 0.317268 0.43338 2.22974 138.883 83.6739 18.7066 60.7475 0.00403548 0 -40 10
1.721 4.97875e-08 2.53987e-06 0.146081 0.146081 0.0120269 2.26307e-05 0.00115449 0.182601 0.000658794 0.183256 0.948252 101.465 0.235381 0.849759 4.53458 0.0646193 0.0427791 0.957221 0.0194545 0.00458274 0.0187119 0.00437291 0.00554549 0.00628812 0.221819 0.251525 58.0472 -87.899 126.165 15.9362 145.035 0.000142182 0.267309 192.732 0.310206 0.0673267 0.00409839 0.000562358 0.00138502 0.986961 0.991717 -2.98965e-06 -85.6573 0.0930825 31169.7 309.767 0.983498 0.319146 0.73757 0.737566 9.99958 2.9863e-06 1.19451e-05 0.13411 0.983397 0.931397 -0.0132916 4.92959e-06 0.515347 -2.00752e-20 7.44547e-24 -2.00677e-20 0.00139642 0.997815 8.60202e-05 0.152727 2.85276 0.00139642 0.997815 0.787348 0.00106694 0.00188134 0.000860202 0.455394 0.00188134 0.444292 0.000131162 1.02 0.888727 0.534387 0.287503 1.71936e-07 3.08342e-09 2371.42 3136.47 -0.0579343 0.482205 0.277285 0.254616 -0.593102 -0.169571 0.488477 -0.265868 -0.222618 2.623 1 0 295.586 0 2.22969 2.621 0.000299163 0.866017 0.698694 0.317226 0.433402 2.22987 138.891 83.6733 18.7066 60.7472 0.00403551 0 -40 10
1.722 4.98163e-08 2.53987e-06 0.146115 0.146115 0.0120269 2.26438e-05 0.00115449 0.182644 0.000658795 0.183298 0.948342 101.465 0.23537 0.849891 4.53519 0.06463 0.0427848 0.957215 0.019454 0.00458318 0.0187113 0.00437329 0.00554604 0.00628868 0.221841 0.251547 58.0472 -87.899 126.165 15.9362 145.035 0.000142185 0.267309 192.732 0.310205 0.0673266 0.00409839 0.000562358 0.00138503 0.98696 0.991717 -2.98967e-06 -85.6573 0.0930826 31169.7 309.779 0.983498 0.319146 0.737582 0.737578 9.99958 2.98631e-06 1.19451e-05 0.134114 0.983398 0.931396 -0.0132916 4.92962e-06 0.515366 -2.00767e-20 7.44609e-24 -2.00693e-20 0.00139642 0.997815 8.60203e-05 0.152727 2.85276 0.00139642 0.997815 0.787422 0.00106695 0.00188134 0.000860203 0.455394 0.00188134 0.444297 0.000131165 1.02 0.888728 0.534387 0.287505 1.71936e-07 3.08344e-09 2371.4 3136.52 -0.0579393 0.482205 0.277284 0.254619 -0.593102 -0.169571 0.488461 -0.265866 -0.222604 2.624 1 0 295.581 0 2.22983 2.622 0.000299161 0.866045 0.698737 0.317184 0.433424 2.23001 138.898 83.6727 18.7065 60.7469 0.00403553 0 -40 10
1.723 4.98452e-08 2.53987e-06 0.146149 0.146148 0.0120269 2.26569e-05 0.00115449 0.182686 0.000658795 0.18334 0.948432 101.464 0.235359 0.850024 4.5358 0.0646407 0.0427906 0.957209 0.0194534 0.00458363 0.0187107 0.00437368 0.00554659 0.00628925 0.221863 0.25157 58.0473 -87.899 126.164 15.9362 145.035 0.000142187 0.267309 192.732 0.310205 0.0673266 0.00409839 0.000562359 0.00138503 0.98696 0.991717 -2.98968e-06 -85.6573 0.0930827 31169.7 309.791 0.983498 0.319146 0.737594 0.73759 9.99958 2.98631e-06 1.19451e-05 0.134119 0.983398 0.931395 -0.0132916 4.92965e-06 0.515385 -2.00783e-20 7.44671e-24 -2.00708e-20 0.00139642 0.997815 8.60204e-05 0.152727 2.85276 0.00139642 0.997815 0.787495 0.00106697 0.00188135 0.000860204 0.455394 0.00188135 0.444302 0.000131167 1.02 0.888729 0.534387 0.287506 1.71937e-07 3.08346e-09 2371.39 3136.57 -0.0579443 0.482205 0.277284 0.254622 -0.593101 -0.169571 0.488445 -0.265864 -0.222591 2.625 1 0 295.577 0 2.22997 2.623 0.00029916 0.866073 0.69878 0.317142 0.433447 2.23015 138.906 83.6722 18.7065 60.7466 0.00403555 0 -40 10
1.724 4.9874e-08 2.53987e-06 0.146183 0.146182 0.0120268 2.267e-05 0.00115449 0.182729 0.000658796 0.183383 0.948521 101.464 0.235349 0.850156 4.53641 0.0646514 0.0427963 0.957204 0.0194529 0.00458408 0.0187102 0.00437406 0.00554714 0.00628982 0.221885 0.251593 58.0473 -87.899 126.164 15.9361 145.035 0.000142189 0.26731 192.732 0.310204 0.0673265 0.0040984 0.00056236 0.00138503 0.98696 0.991717 -2.9897e-06 -85.6573 0.0930828 31169.7 309.803 0.983498 0.319146 0.737606 0.737601 9.99958 2.98632e-06 1.19452e-05 0.134123 0.983398 0.931394 -0.0132916 4.92968e-06 0.515405 -2.00798e-20 7.44733e-24 -2.00724e-20 0.00139642 0.997815 8.60205e-05 0.152727 2.85276 0.00139642 0.997815 0.787569 0.00106699 0.00188135 0.000860205 0.455393 0.00188135 0.444308 0.00013117 1.02 0.888731 0.534386 0.287508 1.71937e-07 3.08349e-09 2371.37 3136.62 -0.0579492 0.482205 0.277284 0.254625 -0.5931 -0.169571 0.488429 -0.265862 -0.222577 2.626 1 0 295.572 0 2.23011 2.624 0.000299159 0.866101 0.698823 0.317101 0.433469 2.23029 138.913 83.6716 18.7065 60.7463 0.00403558 0 -40 10
1.725 4.99029e-08 2.53988e-06 0.146217 0.146216 0.0120268 2.26831e-05 0.00115449 0.182771 0.000658797 0.183425 0.948611 101.463 0.235338 0.850288 4.53702 0.0646621 0.0428021 0.957198 0.0194523 0.00458453 0.0187096 0.00437445 0.00554769 0.00629038 0.221908 0.251615 58.0474 -87.899 126.164 15.9361 145.035 0.000142191 0.26731 192.732 0.310204 0.0673265 0.0040984 0.00056236 0.00138503 0.98696 0.991717 -2.98971e-06 -85.6573 0.0930829 31169.6 309.816 0.983498 0.319146 0.737617 0.737613 9.99958 2.98632e-06 1.19452e-05 0.134128 0.983399 0.931393 -0.0132916 4.92971e-06 0.515424 -2.00814e-20 7.44795e-24 -2.0074e-20 0.00139642 0.997815 8.60205e-05 0.152728 2.85276 0.00139642 0.997815 0.787643 0.001067 0.00188135 0.000860205 0.455393 0.00188135 0.444313 0.000131172 1.02 0.888732 0.534386 0.287509 1.71937e-07 3.08351e-09 2371.35 3136.67 -0.0579542 0.482205 0.277284 0.254628 -0.5931 -0.169572 0.488413 -0.26586 -0.222563 2.627 1 0 295.568 0 2.23024 2.625 0.000299158 0.866129 0.698866 0.317059 0.433491 2.23042 138.92 83.671 18.7064 60.7461 0.0040356 0 -40 10
1.726 4.99317e-08 2.53988e-06 0.14625 0.14625 0.0120268 2.26962e-05 0.00115449 0.182813 0.000658797 0.183467 0.9487 101.462 0.235327 0.85042 4.53763 0.0646728 0.0428079 0.957192 0.0194518 0.00458497 0.018709 0.00437484 0.00554824 0.00629095 0.22193 0.251638 58.0475 -87.899 126.164 15.9361 145.035 0.000142194 0.26731 192.731 0.310204 0.0673264 0.0040984 0.000562361 0.00138504 0.98696 0.991717 -2.98973e-06 -85.6573 0.093083 31169.6 309.828 0.983498 0.319146 0.737629 0.737625 9.99958 2.98633e-06 1.19452e-05 0.134133 0.983399 0.931392 -0.0132916 4.92974e-06 0.515444 -2.0083e-20 7.44858e-24 -2.00755e-20 0.00139643 0.997815 8.60206e-05 0.152728 2.85276 0.00139643 0.997815 0.787716 0.00106702 0.00188135 0.000860206 0.455393 0.00188135 0.444318 0.000131175 1.02 0.888733 0.534386 0.287511 1.71937e-07 3.08353e-09 2371.34 3136.72 -0.0579592 0.482206 0.277283 0.254631 -0.593099 -0.169572 0.488398 -0.265858 -0.222549 2.628 1 0 295.563 0 2.23038 2.626 0.000299157 0.866157 0.698909 0.317017 0.433514 2.23056 138.928 83.6704 18.7064 60.7458 0.00403563 0 -40 10
1.727 4.99606e-08 2.53988e-06 0.146284 0.146284 0.0120268 2.27093e-05 0.00115449 0.182855 0.000658798 0.183509 0.94879 101.462 0.235317 0.850552 4.53824 0.0646835 0.0428136 0.957186 0.0194512 0.00458542 0.0187085 0.00437522 0.00554879 0.00629152 0.221952 0.251661 58.0475 -87.899 126.164 15.936 145.035 0.000142196 0.26731 192.731 0.310203 0.0673264 0.00409841 0.000562362 0.00138504 0.98696 0.991717 -2.98974e-06 -85.6573 0.0930831 31169.6 309.84 0.983498 0.319146 0.737641 0.737636 9.99958 2.98633e-06 1.19452e-05 0.134137 0.983399 0.931391 -0.0132916 4.92977e-06 0.515463 -2.00845e-20 7.4492e-24 -2.00771e-20 0.00139643 0.997815 8.60207e-05 0.152728 2.85276 0.00139643 0.997815 0.78779 0.00106704 0.00188135 0.000860207 0.455393 0.00188135 0.444324 0.000131177 1.02 0.888734 0.534385 0.287512 1.71938e-07 3.08356e-09 2371.32 3136.77 -0.0579642 0.482206 0.277283 0.254634 -0.593098 -0.169572 0.488382 -0.265856 -0.222536 2.629 1 0 295.559 0 2.23052 2.627 0.000299155 0.866185 0.698952 0.316975 0.433536 2.2307 138.935 83.6698 18.7064 60.7455 0.00403565 0 -40 10
1.728 4.99894e-08 2.53988e-06 0.146318 0.146317 0.0120268 2.27225e-05 0.00115449 0.182897 0.000658798 0.183552 0.94888 101.461 0.235306 0.850684 4.53886 0.0646942 0.0428194 0.957181 0.0194507 0.00458587 0.0187079 0.00437561 0.00554934 0.00629209 0.221974 0.251683 58.0476 -87.899 126.163 15.936 145.035 0.000142198 0.26731 192.731 0.310203 0.0673263 0.00409841 0.000562362 0.00138504 0.98696 0.991717 -2.98976e-06 -85.6573 0.0930831 31169.6 309.852 0.983498 0.319146 0.737653 0.737648 9.99958 2.98634e-06 1.19452e-05 0.134142 0.9834 0.93139 -0.0132916 4.9298e-06 0.515482 -2.00861e-20 7.44982e-24 -2.00786e-20 0.00139643 0.997815 8.60208e-05 0.152728 2.85276 0.00139643 0.997815 0.787864 0.00106705 0.00188135 0.000860208 0.455392 0.00188135 0.444329 0.000131179 1.02 0.888735 0.534385 0.287514 1.71938e-07 3.08358e-09 2371.3 3136.82 -0.0579691 0.482206 0.277283 0.254638 -0.593098 -0.169572 0.488366 -0.265853 -0.222522 2.63 1 0 295.554 0 2.23066 2.628 0.000299154 0.866214 0.698995 0.316934 0.433558 2.23084 138.942 83.6693 18.7063 60.7452 0.00403567 0 -40 10
1.729 5.00183e-08 2.53988e-06 0.146352 0.146351 0.0120268 2.27356e-05 0.00115449 0.18294 0.000658799 0.183594 0.948969 101.461 0.235295 0.850817 4.53947 0.0647049 0.0428252 0.957175 0.0194501 0.00458632 0.0187073 0.004376 0.0055499 0.00629266 0.221996 0.251706 58.0477 -87.8991 126.163 15.9359 145.035 0.0001422 0.267311 192.731 0.310202 0.0673262 0.00409841 0.000562363 0.00138504 0.98696 0.991717 -2.98977e-06 -85.6573 0.0930832 31169.5 309.864 0.983498 0.319146 0.737664 0.73766 9.99958 2.98634e-06 1.19453e-05 0.134146 0.9834 0.931389 -0.0132916 4.92983e-06 0.515502 -2.00876e-20 7.45045e-24 -2.00802e-20 0.00139643 0.997815 8.60209e-05 0.152728 2.85277 0.00139643 0.997815 0.787937 0.00106707 0.00188136 0.000860209 0.455392 0.00188135 0.444334 0.000131182 1.02 0.888736 0.534385 0.287515 1.71938e-07 3.0836e-09 2371.29 3136.87 -0.0579741 0.482206 0.277282 0.254641 -0.593097 -0.169572 0.48835 -0.265851 -0.222508 2.631 1 0 295.55 0 2.23079 2.629 0.000299153 0.866242 0.699038 0.316892 0.43358 2.23097 138.95 83.6687 18.7063 60.7449 0.0040357 0 -40 10
1.73 5.00471e-08 2.53988e-06 0.146385 0.146385 0.0120268 2.27487e-05 0.00115449 0.182982 0.000658799 0.183636 0.949059 101.46 0.235284 0.850949 4.54008 0.0647156 0.042831 0.957169 0.0194496 0.00458677 0.0187068 0.00437638 0.00555045 0.00629322 0.222018 0.251729 58.0477 -87.8991 126.163 15.9359 145.035 0.000142203 0.267311 192.731 0.310202 0.0673262 0.00409842 0.000562364 0.00138504 0.98696 0.991717 -2.98979e-06 -85.6572 0.0930833 31169.5 309.876 0.983498 0.319146 0.737676 0.737672 9.99958 2.98635e-06 1.19453e-05 0.134151 0.9834 0.931388 -0.0132916 4.92986e-06 0.515521 -2.00892e-20 7.45107e-24 -2.00817e-20 0.00139643 0.997815 8.60209e-05 0.152728 2.85277 0.00139643 0.997815 0.788011 0.00106708 0.00188136 0.000860209 0.455392 0.00188136 0.444339 0.000131184 1.02 0.888737 0.534384 0.287517 1.71939e-07 3.08362e-09 2371.27 3136.92 -0.0579791 0.482206 0.277282 0.254644 -0.593097 -0.169572 0.488334 -0.265849 -0.222494 2.632 1 0 295.545 0 2.23093 2.63 0.000299152 0.86627 0.699082 0.31685 0.433603 2.23111 138.957 83.6681 18.7063 60.7447 0.00403572 0 -40 10
1.731 5.00759e-08 2.53989e-06 0.146419 0.146419 0.0120267 2.27618e-05 0.00115449 0.183024 0.0006588 0.183678 0.949149 101.459 0.235274 0.851081 4.5407 0.0647263 0.0428368 0.957163 0.019449 0.00458721 0.0187062 0.00437677 0.005551 0.00629379 0.22204 0.251752 58.0478 -87.8991 126.163 15.9359 145.035 0.000142205 0.267311 192.731 0.310201 0.0673261 0.00409842 0.000562364 0.00138505 0.98696 0.991717 -2.9898e-06 -85.6572 0.0930834 31169.5 309.889 0.983498 0.319146 0.737688 0.737684 9.99958 2.98635e-06 1.19453e-05 0.134155 0.983401 0.931387 -0.0132916 4.92989e-06 0.515541 -2.00907e-20 7.45169e-24 -2.00833e-20 0.00139643 0.997815 8.6021e-05 0.152729 2.85277 0.00139643 0.997815 0.788084 0.0010671 0.00188136 0.00086021 0.455392 0.00188136 0.444345 0.000131187 1.02 0.888738 0.534384 0.287518 1.71939e-07 3.08365e-09 2371.25 3136.97 -0.0579841 0.482206 0.277282 0.254647 -0.593096 -0.169572 0.488318 -0.265847 -0.222481 2.633 1 0 295.541 0 2.23107 2.631 0.000299151 0.866298 0.699125 0.316809 0.433625 2.23125 138.965 83.6675 18.7062 60.7444 0.00403575 0 -40 10
1.732 5.01048e-08 2.53989e-06 0.146453 0.146452 0.0120267 2.27749e-05 0.00115449 0.183066 0.0006588 0.18372 0.949239 101.459 0.235263 0.851214 4.54131 0.064737 0.0428425 0.957157 0.0194484 0.00458766 0.0187056 0.00437716 0.00555155 0.00629436 0.222062 0.251774 58.0478 -87.8991 126.163 15.9358 145.035 0.000142207 0.267311 192.73 0.310201 0.0673261 0.00409842 0.000562365 0.00138505 0.98696 0.991717 -2.98982e-06 -85.6572 0.0930835 31169.5 309.901 0.983498 0.319146 0.7377 0.737695 9.99958 2.98636e-06 1.19453e-05 0.13416 0.983401 0.931386 -0.0132916 4.92992e-06 0.51556 -2.00923e-20 7.45232e-24 -2.00849e-20 0.00139643 0.997815 8.60211e-05 0.152729 2.85277 0.00139643 0.997815 0.788158 0.00106712 0.00188136 0.000860211 0.455391 0.00188136 0.44435 0.000131189 1.02 0.888739 0.534384 0.28752 1.71939e-07 3.08367e-09 2371.24 3137.01 -0.0579891 0.482206 0.277282 0.25465 -0.593095 -0.169572 0.488303 -0.265845 -0.222467 2.634 1 0 295.536 0 2.23121 2.632 0.00029915 0.866326 0.699168 0.316767 0.433647 2.23139 138.972 83.667 18.7062 60.7441 0.00403577 0 -40 10
1.733 5.01336e-08 2.53989e-06 0.146486 0.146486 0.0120267 2.2788e-05 0.00115449 0.183108 0.000658801 0.183762 0.949328 101.458 0.235252 0.851346 4.54192 0.0647478 0.0428483 0.957152 0.0194479 0.00458811 0.0187051 0.00437755 0.00555211 0.00629493 0.222084 0.251797 58.0479 -87.8991 126.162 15.9358 145.035 0.000142209 0.267311 192.73 0.310201 0.067326 0.00409842 0.000562366 0.00138505 0.98696 0.991717 -2.98983e-06 -85.6572 0.0930836 31169.5 309.913 0.983498 0.319146 0.737711 0.737707 9.99958 2.98636e-06 1.19453e-05 0.134165 0.983401 0.931385 -0.0132916 4.92995e-06 0.51558 -2.00939e-20 7.45294e-24 -2.00864e-20 0.00139643 0.997815 8.60212e-05 0.152729 2.85277 0.00139643 0.997815 0.788231 0.00106713 0.00188136 0.000860212 0.455391 0.00188136 0.444355 0.000131192 1.02 0.88874 0.534384 0.287521 1.71939e-07 3.08369e-09 2371.22 3137.06 -0.057994 0.482206 0.277281 0.254653 -0.593095 -0.169572 0.488287 -0.265843 -0.222453 2.635 1 0 295.532 0 2.23134 2.633 0.000299148 0.866354 0.699211 0.316726 0.433669 2.23152 138.979 83.6664 18.7062 60.7438 0.00403579 0 -40 10
1.734 5.01625e-08 2.53989e-06 0.14652 0.146519 0.0120267 2.28011e-05 0.0011545 0.18315 0.000658801 0.183804 0.949418 101.457 0.235242 0.851478 4.54254 0.0647585 0.0428541 0.957146 0.0194473 0.00458856 0.0187045 0.00437793 0.00555266 0.0062955 0.222106 0.25182 58.048 -87.8991 126.162 15.9358 145.035 0.000142212 0.267312 192.73 0.3102 0.067326 0.00409843 0.000562366 0.00138505 0.98696 0.991717 -2.98985e-06 -85.6572 0.0930837 31169.4 309.925 0.983498 0.319146 0.737723 0.737719 9.99958 2.98637e-06 1.19454e-05 0.134169 0.983401 0.931384 -0.0132916 4.92998e-06 0.515599 -2.00954e-20 7.45357e-24 -2.0088e-20 0.00139644 0.997815 8.60213e-05 0.152729 2.85277 0.00139643 0.997815 0.788305 0.00106715 0.00188136 0.000860213 0.455391 0.00188136 0.44436 0.000131194 1.02 0.888742 0.534383 0.287523 1.7194e-07 3.08372e-09 2371.21 3137.11 -0.057999 0.482206 0.277281 0.254657 -0.593094 -0.169572 0.488271 -0.265841 -0.222439 2.636 1 0 295.527 0 2.23148 2.634 0.000299147 0.866383 0.699254 0.316684 0.433692 2.23166 138.987 83.6658 18.7061 60.7436 0.00403582 0 -40 10
1.735 5.01913e-08 2.53989e-06 0.146553 0.146553 0.0120267 2.28142e-05 0.0011545 0.183192 0.000658802 0.183846 0.949508 101.457 0.235231 0.85161 4.54315 0.0647692 0.0428599 0.95714 0.0194468 0.00458901 0.0187039 0.00437832 0.00555321 0.00629607 0.222129 0.251843 58.048 -87.8991 126.162 15.9357 145.035 0.000142214 0.267312 192.73 0.3102 0.0673259 0.00409843 0.000562367 0.00138506 0.98696 0.991717 -2.98986e-06 -85.6572 0.0930838 31169.4 309.937 0.983498 0.319146 0.737735 0.737731 9.99958 2.98637e-06 1.19454e-05 0.134174 0.983402 0.931383 -0.0132916 4.93001e-06 0.515619 -2.0097e-20 7.45419e-24 -2.00895e-20 0.00139644 0.997815 8.60214e-05 0.152729 2.85277 0.00139644 0.997815 0.788378 0.00106717 0.00188136 0.000860214 0.455391 0.00188136 0.444366 0.000131196 1.02 0.888743 0.534383 0.287524 1.7194e-07 3.08374e-09 2371.19 3137.16 -0.058004 0.482206 0.277281 0.25466 -0.593093 -0.169572 0.488255 -0.265839 -0.222426 2.637 1 0 295.523 0 2.23162 2.635 0.000299146 0.866411 0.699297 0.316643 0.433714 2.2318 138.994 83.6652 18.7061 60.7433 0.00403584 0 -40 10
1.736 5.02202e-08 2.53989e-06 0.146587 0.146586 0.0120267 2.28274e-05 0.0011545 0.183234 0.000658802 0.183888 0.949598 101.456 0.23522 0.851743 4.54377 0.0647799 0.0428658 0.957134 0.0194462 0.00458946 0.0187034 0.00437871 0.00555377 0.00629664 0.222151 0.251866 58.0481 -87.8991 126.162 15.9357 145.036 0.000142216 0.267312 192.73 0.310199 0.0673259 0.00409843 0.000562368 0.00138506 0.98696 0.991717 -2.98988e-06 -85.6572 0.0930838 31169.4 309.95 0.983498 0.319146 0.737747 0.737742 9.99958 2.98638e-06 1.19454e-05 0.134178 0.983402 0.931382 -0.0132916 4.93004e-06 0.515638 -2.00986e-20 7.45482e-24 -2.00911e-20 0.00139644 0.997815 8.60214e-05 0.152729 2.85277 0.00139644 0.997815 0.788452 0.00106718 0.00188137 0.000860214 0.455391 0.00188136 0.444371 0.000131199 1.02 0.888744 0.534383 0.287526 1.7194e-07 3.08376e-09 2371.17 3137.21 -0.058009 0.482206 0.27728 0.254663 -0.593093 -0.169572 0.488239 -0.265837 -0.222412 2.638 1 0 295.518 0 2.23175 2.636 0.000299145 0.866439 0.69934 0.316601 0.433736 2.23194 139.001 83.6646 18.7061 60.743 0.00403587 0 -40 10
1.737 5.0249e-08 2.5399e-06 0.146621 0.14662 0.0120267 2.28405e-05 0.0011545 0.183276 0.000658803 0.18393 0.949688 101.456 0.235209 0.851875 4.54439 0.0647906 0.0428716 0.957128 0.0194457 0.00458991 0.0187028 0.0043791 0.00555432 0.00629721 0.222173 0.251888 58.0482 -87.8991 126.161 15.9356 145.036 0.000142219 0.267312 192.73 0.310199 0.0673258 0.00409844 0.000562368 0.00138506 0.98696 0.991716 -2.98989e-06 -85.6572 0.0930839 31169.4 309.962 0.983498 0.319146 0.737759 0.737754 9.99958 2.98638e-06 1.19454e-05 0.134183 0.983402 0.931382 -0.0132916 4.93007e-06 0.515658 -2.01001e-20 7.45544e-24 -2.00927e-20 0.00139644 0.997815 8.60215e-05 0.152729 2.85277 0.00139644 0.997815 0.788525 0.0010672 0.00188137 0.000860215 0.45539 0.00188137 0.444376 0.000131201 1.02 0.888745 0.534382 0.287527 1.7194e-07 3.08378e-09 2371.16 3137.26 -0.058014 0.482206 0.27728 0.254666 -0.593092 -0.169572 0.488223 -0.265835 -0.222398 2.639 1 0 295.514 0 2.23189 2.637 0.000299144 0.866467 0.699383 0.31656 0.433758 2.23207 139.009 83.6641 18.706 60.7427 0.00403589 0 -40 10
1.738 5.02779e-08 2.5399e-06 0.146654 0.146653 0.0120266 2.28536e-05 0.0011545 0.183317 0.000658804 0.183972 0.949777 101.455 0.235199 0.852008 4.545 0.0648013 0.0428774 0.957123 0.0194451 0.00459036 0.0187022 0.00437949 0.00555488 0.00629778 0.222195 0.251911 58.0482 -87.8991 126.161 15.9356 145.036 0.000142221 0.267312 192.729 0.310198 0.0673258 0.00409844 0.000562369 0.00138506 0.98696 0.991716 -2.98991e-06 -85.6572 0.093084 31169.3 309.974 0.983498 0.319146 0.73777 0.737766 9.99958 2.98639e-06 1.19454e-05 0.134187 0.983403 0.931381 -0.0132916 4.9301e-06 0.515677 -2.01017e-20 7.45607e-24 -2.00942e-20 0.00139644 0.997815 8.60216e-05 0.15273 2.85277 0.00139644 0.997815 0.788598 0.00106721 0.00188137 0.000860216 0.45539 0.00188137 0.444381 0.000131204 1.02 0.888746 0.534382 0.287529 1.71941e-07 3.08381e-09 2371.14 3137.31 -0.058019 0.482206 0.27728 0.254669 -0.593092 -0.169572 0.488207 -0.265832 -0.222384 2.64 1 0 295.509 0 2.23203 2.638 0.000299142 0.866495 0.699426 0.316518 0.433781 2.23221 139.016 83.6635 18.706 60.7424 0.00403591 0 -40 10
1.739 5.03067e-08 2.5399e-06 0.146687 0.146687 0.0120266 2.28667e-05 0.0011545 0.183359 0.000658804 0.184014 0.949867 101.454 0.235188 0.85214 4.54562 0.0648121 0.0428832 0.957117 0.0194446 0.00459081 0.0187016 0.00437988 0.00555543 0.00629835 0.222217 0.251934 58.0483 -87.8991 126.161 15.9356 145.036 0.000142223 0.267313 192.729 0.310198 0.0673257 0.00409844 0.00056237 0.00138506 0.98696 0.991716 -2.98992e-06 -85.6572 0.0930841 31169.3 309.986 0.983498 0.319146 0.737782 0.737778 9.99958 2.98639e-06 1.19455e-05 0.134192 0.983403 0.93138 -0.0132916 4.93013e-06 0.515697 -2.01033e-20 7.4567e-24 -2.00958e-20 0.00139644 0.997815 8.60217e-05 0.15273 2.85277 0.00139644 0.997815 0.788672 0.00106723 0.00188137 0.000860217 0.45539 0.00188137 0.444387 0.000131206 1.02 0.888747 0.534382 0.28753 1.71941e-07 3.08383e-09 2371.12 3137.36 -0.058024 0.482206 0.27728 0.254672 -0.593091 -0.169572 0.488192 -0.26583 -0.222371 2.641 1 0 295.505 0 2.23217 2.639 0.000299141 0.866524 0.699469 0.316477 0.433803 2.23235 139.024 83.6629 18.706 60.7422 0.00403594 0 -40 10
1.74 5.03356e-08 2.5399e-06 0.146721 0.14672 0.0120266 2.28798e-05 0.0011545 0.183401 0.000658805 0.184055 0.949957 101.454 0.235177 0.852272 4.54624 0.0648228 0.042889 0.957111 0.019444 0.00459126 0.0187011 0.00438027 0.00555599 0.00629892 0.22224 0.251957 58.0483 -87.8991 126.161 15.9355 145.036 0.000142225 0.267313 192.729 0.310198 0.0673257 0.00409845 0.00056237 0.00138507 0.98696 0.991716 -2.98994e-06 -85.6572 0.0930842 31169.3 309.999 0.983498 0.319146 0.737794 0.73779 9.99958 2.9864e-06 1.19455e-05 0.134197 0.983403 0.931379 -0.0132916 4.93016e-06 0.515717 -2.01048e-20 7.45732e-24 -2.00974e-20 0.00139644 0.997815 8.60218e-05 0.15273 2.85278 0.00139644 0.997815 0.788745 0.00106725 0.00188137 0.000860218 0.45539 0.00188137 0.444392 0.000131209 1.02 0.888748 0.534381 0.287532 1.71941e-07 3.08385e-09 2371.11 3137.41 -0.058029 0.482207 0.277279 0.254676 -0.59309 -0.169572 0.488176 -0.265828 -0.222357 2.642 1 0 295.5 0 2.2323 2.64 0.00029914 0.866552 0.699512 0.316436 0.433825 2.23248 139.031 83.6623 18.7059 60.7419 0.00403596 0 -40 10
1.741 5.03644e-08 2.5399e-06 0.146754 0.146754 0.0120266 2.28929e-05 0.0011545 0.183443 0.000658805 0.184097 0.950047 101.453 0.235166 0.852405 4.54686 0.0648335 0.0428949 0.957105 0.0194435 0.00459171 0.0187005 0.00438065 0.00555654 0.00629949 0.222262 0.25198 58.0484 -87.8991 126.161 15.9355 145.036 0.000142228 0.267313 192.729 0.310197 0.0673256 0.00409845 0.000562371 0.00138507 0.98696 0.991716 -2.98995e-06 -85.6571 0.0930843 31169.3 310.011 0.983498 0.319146 0.737806 0.737801 9.99958 2.9864e-06 1.19455e-05 0.134201 0.983404 0.931378 -0.0132916 4.93019e-06 0.515736 -2.01064e-20 7.45795e-24 -2.00989e-20 0.00139644 0.997815 8.60218e-05 0.15273 2.85278 0.00139644 0.997815 0.788818 0.00106726 0.00188137 0.000860218 0.455389 0.00188137 0.444397 0.000131211 1.02 0.888749 0.534381 0.287533 1.71942e-07 3.08388e-09 2371.09 3137.46 -0.0580339 0.482207 0.277279 0.254679 -0.59309 -0.169573 0.48816 -0.265826 -0.222343 2.643 1 0 295.496 0 2.23244 2.641 0.000299139 0.86658 0.699555 0.316394 0.433847 2.23262 139.038 83.6617 18.7059 60.7416 0.00403599 0 -40 10
1.742 5.03932e-08 2.5399e-06 0.146788 0.146787 0.0120266 2.2906e-05 0.0011545 0.183485 0.000658806 0.184139 0.950137 101.453 0.235156 0.852537 4.54747 0.0648442 0.0429007 0.957099 0.0194429 0.00459216 0.0186999 0.00438104 0.0055571 0.00630007 0.222284 0.252003 58.0485 -87.8991 126.16 15.9355 145.036 0.00014223 0.267313 192.729 0.310197 0.0673256 0.00409845 0.000562372 0.00138507 0.98696 0.991716 -2.98997e-06 -85.6571 0.0930844 31169.2 310.023 0.983498 0.319146 0.737818 0.737813 9.99958 2.98641e-06 1.19455e-05 0.134206 0.983404 0.931377 -0.0132916 4.93022e-06 0.515756 -2.0108e-20 7.45858e-24 -2.01005e-20 0.00139644 0.997815 8.60219e-05 0.15273 2.85278 0.00139644 0.997815 0.788891 0.00106728 0.00188137 0.000860219 0.455389 0.00188137 0.444402 0.000131213 1.02 0.88875 0.534381 0.287535 1.71942e-07 3.0839e-09 2371.07 3137.51 -0.0580389 0.482207 0.277279 0.254682 -0.593089 -0.169573 0.488144 -0.265824 -0.222329 2.644 1 0 295.491 0 2.23258 2.642 0.000299138 0.866608 0.699598 0.316353 0.43387 2.23276 139.046 83.6611 18.7059 60.7413 0.00403601 0 -40 10
1.743 5.04221e-08 2.5399e-06 0.146821 0.14682 0.0120266 2.29191e-05 0.0011545 0.183526 0.000658806 0.18418 0.950227 101.452 0.235145 0.85267 4.54809 0.064855 0.0429065 0.957093 0.0194423 0.00459261 0.0186994 0.00438143 0.00555765 0.00630064 0.222306 0.252026 58.0485 -87.8991 126.16 15.9354 145.036 0.000142232 0.267313 192.729 0.310196 0.0673255 0.00409845 0.000562372 0.00138507 0.98696 0.991716 -2.98998e-06 -85.6571 0.0930845 31169.2 310.035 0.983498 0.319146 0.737829 0.737825 9.99958 2.98641e-06 1.19455e-05 0.13421 0.983404 0.931376 -0.0132916 4.93025e-06 0.515775 -2.01095e-20 7.4592e-24 -2.01021e-20 0.00139645 0.997815 8.6022e-05 0.15273 2.85278 0.00139645 0.997815 0.788965 0.0010673 0.00188138 0.00086022 0.455389 0.00188137 0.444408 0.000131216 1.02 0.888751 0.53438 0.287537 1.71942e-07 3.08392e-09 2371.06 3137.56 -0.0580439 0.482207 0.277278 0.254685 -0.593088 -0.169573 0.488128 -0.265822 -0.222315 2.645 1 0 295.487 0 2.23272 2.643 0.000299136 0.866637 0.699641 0.316312 0.433892 2.2329 139.053 83.6606 18.7058 60.741 0.00403603 0 -40 10
1.744 5.04509e-08 2.53991e-06 0.146854 0.146854 0.0120266 2.29322e-05 0.0011545 0.183568 0.000658807 0.184222 0.950317 101.451 0.235134 0.852802 4.54871 0.0648657 0.0429124 0.957088 0.0194418 0.00459306 0.0186988 0.00438182 0.00555821 0.00630121 0.222328 0.252048 58.0486 -87.8991 126.16 15.9354 145.036 0.000142234 0.267314 192.728 0.310196 0.0673255 0.00409846 0.000562373 0.00138507 0.98696 0.991716 -2.99e-06 -85.6571 0.0930845 31169.2 310.048 0.983498 0.319146 0.737841 0.737837 9.99958 2.98642e-06 1.19456e-05 0.134215 0.983404 0.931375 -0.0132916 4.93028e-06 0.515795 -2.01111e-20 7.45983e-24 -2.01036e-20 0.00139645 0.997815 8.60221e-05 0.152731 2.85278 0.00139645 0.997815 0.789038 0.00106731 0.00188138 0.000860221 0.455389 0.00188138 0.444413 0.000131218 1.02 0.888752 0.53438 0.287538 1.71942e-07 3.08394e-09 2371.04 3137.61 -0.0580489 0.482207 0.277278 0.254688 -0.593088 -0.169573 0.488112 -0.26582 -0.222302 2.646 1 0 295.482 0 2.23285 2.644 0.000299135 0.866665 0.699684 0.316271 0.433914 2.23303 139.06 83.66 18.7058 60.7407 0.00403606 0 -40 10
1.745 5.04798e-08 2.53991e-06 0.146888 0.146887 0.0120266 2.29454e-05 0.0011545 0.183609 0.000658807 0.184264 0.950407 101.451 0.235124 0.852935 4.54933 0.0648764 0.0429182 0.957082 0.0194412 0.00459351 0.0186982 0.00438221 0.00555877 0.00630178 0.222351 0.252071 58.0487 -87.8991 126.16 15.9353 145.036 0.000142237 0.267314 192.728 0.310195 0.0673254 0.00409846 0.000562374 0.00138508 0.98696 0.991716 -2.99001e-06 -85.6571 0.0930846 31169.2 310.06 0.983498 0.319146 0.737853 0.737849 9.99958 2.98642e-06 1.19456e-05 0.13422 0.983405 0.931374 -0.0132916 4.93031e-06 0.515814 -2.01127e-20 7.46046e-24 -2.01052e-20 0.00139645 0.997815 8.60222e-05 0.152731 2.85278 0.00139645 0.997815 0.789111 0.00106733 0.00188138 0.000860222 0.455389 0.00188138 0.444418 0.000131221 1.02 0.888754 0.53438 0.28754 1.71943e-07 3.08397e-09 2371.03 3137.66 -0.0580539 0.482207 0.277278 0.254692 -0.593087 -0.169573 0.488096 -0.265818 -0.222288 2.647 1 0 295.478 0 2.23299 2.645 0.000299134 0.866693 0.699727 0.31623 0.433936 2.23317 139.068 83.6594 18.7058 60.7405 0.00403608 0 -40 10
1.746 5.05086e-08 2.53991e-06 0.146921 0.14692 0.0120265 2.29585e-05 0.0011545 0.183651 0.000658808 0.184305 0.950497 101.45 0.235113 0.853067 4.54995 0.0648872 0.0429241 0.957076 0.0194407 0.00459397 0.0186976 0.0043826 0.00555932 0.00630236 0.222373 0.252094 58.0487 -87.8991 126.16 15.9353 145.036 0.000142239 0.267314 192.728 0.310195 0.0673254 0.00409846 0.000562374 0.00138508 0.98696 0.991716 -2.99003e-06 -85.6571 0.0930847 31169.2 310.072 0.983498 0.319146 0.737865 0.73786 9.99958 2.98643e-06 1.19456e-05 0.134224 0.983405 0.931373 -0.0132916 4.93034e-06 0.515834 -2.01142e-20 7.46109e-24 -2.01068e-20 0.00139645 0.997815 8.60222e-05 0.152731 2.85278 0.00139645 0.997815 0.789184 0.00106734 0.00188138 0.000860222 0.455388 0.00188138 0.444423 0.000131223 1.02 0.888755 0.53438 0.287541 1.71943e-07 3.08399e-09 2371.01 3137.71 -0.0580589 0.482207 0.277278 0.254695 -0.593087 -0.169573 0.48808 -0.265816 -0.222274 2.648 1 0 295.473 0 2.23313 2.646 0.000299133 0.866722 0.69977 0.316189 0.433959 2.23331 139.075 83.6588 18.7057 60.7402 0.00403611 0 -40 10
1.747 5.05375e-08 2.53991e-06 0.146954 0.146954 0.0120265 2.29716e-05 0.00115451 0.183693 0.000658808 0.184347 0.950586 101.449 0.235102 0.8532 4.55057 0.0648979 0.0429299 0.95707 0.0194401 0.00459442 0.0186971 0.00438299 0.00555988 0.00630293 0.222395 0.252117 58.0488 -87.8991 126.159 15.9353 145.036 0.000142241 0.267314 192.728 0.310195 0.0673253 0.00409847 0.000562375 0.00138508 0.98696 0.991716 -2.99004e-06 -85.6571 0.0930848 31169.1 310.084 0.983498 0.319146 0.737877 0.737872 9.99958 2.98643e-06 1.19456e-05 0.134229 0.983405 0.931372 -0.0132916 4.93036e-06 0.515854 -2.01158e-20 7.46172e-24 -2.01083e-20 0.00139645 0.997815 8.60223e-05 0.152731 2.85278 0.00139645 0.997815 0.789257 0.00106736 0.00188138 0.000860223 0.455388 0.00188138 0.444428 0.000131225 1.02 0.888756 0.534379 0.287543 1.71943e-07 3.08401e-09 2370.99 3137.76 -0.0580639 0.482207 0.277277 0.254698 -0.593086 -0.169573 0.488064 -0.265814 -0.22226 2.649 1 0 295.469 0 2.23326 2.647 0.000299132 0.86675 0.699813 0.316148 0.433981 2.23344 139.082 83.6582 18.7057 60.7399 0.00403613 0 -40 10
1.748 5.05663e-08 2.53991e-06 0.146987 0.146987 0.0120265 2.29847e-05 0.00115451 0.183734 0.000658809 0.184388 0.950676 101.449 0.235091 0.853332 4.55119 0.0649086 0.0429358 0.957064 0.0194396 0.00459487 0.0186965 0.00438338 0.00556044 0.0063035 0.222418 0.25214 58.0489 -87.8991 126.159 15.9352 145.036 0.000142244 0.267314 192.728 0.310194 0.0673252 0.00409847 0.000562376 0.00138508 0.98696 0.991716 -2.99006e-06 -85.6571 0.0930849 31169.1 310.097 0.983498 0.319146 0.737889 0.737884 9.99958 2.98644e-06 1.19456e-05 0.134233 0.983406 0.931371 -0.0132916 4.93039e-06 0.515873 -2.01174e-20 7.46235e-24 -2.01099e-20 0.00139645 0.997815 8.60224e-05 0.152731 2.85278 0.00139645 0.997815 0.78933 0.00106738 0.00188138 0.000860224 0.455388 0.00188138 0.444434 0.000131228 1.02 0.888757 0.534379 0.287544 1.71943e-07 3.08404e-09 2370.98 3137.81 -0.0580689 0.482207 0.277277 0.254701 -0.593085 -0.169573 0.488049 -0.265811 -0.222246 2.65 1 0 295.464 0 2.2334 2.648 0.00029913 0.866778 0.699856 0.316106 0.434003 2.23358 139.09 83.6577 18.7057 60.7396 0.00403615 0 -40 10
1.749 5.05952e-08 2.53991e-06 0.14702 0.14702 0.0120265 2.29978e-05 0.00115451 0.183776 0.000658809 0.18443 0.950766 101.448 0.235081 0.853465 4.55182 0.0649194 0.0429417 0.957058 0.019439 0.00459532 0.0186959 0.00438377 0.005561 0.00630408 0.22244 0.252163 58.0489 -87.8991 126.159 15.9352 145.036 0.000142246 0.267314 192.728 0.310194 0.0673252 0.00409847 0.000562376 0.00138509 0.98696 0.991716 -2.99007e-06 -85.6571 0.093085 31169.1 310.109 0.983498 0.319146 0.7379 0.737896 9.99958 2.98644e-06 1.19457e-05 0.134238 0.983406 0.93137 -0.0132916 4.93042e-06 0.515893 -2.01189e-20 7.46297e-24 -2.01115e-20 0.00139645 0.997815 8.60225e-05 0.152731 2.85278 0.00139645 0.997815 0.789403 0.00106739 0.00188139 0.000860225 0.455388 0.00188138 0.444439 0.00013123 1.02 0.888758 0.534379 0.287546 1.71944e-07 3.08406e-09 2370.96 3137.86 -0.0580739 0.482207 0.277277 0.254704 -0.593085 -0.169573 0.488033 -0.265809 -0.222233 2.651 1 0 295.46 0 2.23354 2.649 0.000299129 0.866807 0.699899 0.316065 0.434025 2.23372 139.097 83.6571 18.7056 60.7393 0.00403618 0 -40 10
1.75 5.0624e-08 2.53992e-06 0.147054 0.147053 0.0120265 2.30109e-05 0.00115451 0.183817 0.00065881 0.184471 0.950856 101.448 0.23507 0.853597 4.55244 0.0649301 0.0429475 0.957052 0.0194384 0.00459577 0.0186954 0.00438417 0.00556155 0.00630465 0.222462 0.252186 58.049 -87.8991 126.159 15.9352 145.036 0.000142248 0.267315 192.727 0.310193 0.0673251 0.00409848 0.000562377 0.00138509 0.98696 0.991716 -2.99009e-06 -85.6571 0.0930851 31169.1 310.121 0.983498 0.319146 0.737912 0.737908 9.99958 2.98645e-06 1.19457e-05 0.134243 0.983406 0.931369 -0.0132916 4.93045e-06 0.515913 -2.01205e-20 7.4636e-24 -2.01131e-20 0.00139645 0.997815 8.60226e-05 0.152731 2.85278 0.00139645 0.997815 0.789476 0.00106741 0.00188139 0.000860226 0.455387 0.00188139 0.444444 0.000131233 1.02 0.888759 0.534378 0.287547 1.71944e-07 3.08408e-09 2370.94 3137.91 -0.0580789 0.482207 0.277277 0.254707 -0.593084 -0.169573 0.488017 -0.265807 -0.222219 2.652 1 0 295.455 0 2.23368 2.65 0.000299128 0.866835 0.699942 0.316025 0.434047 2.23386 139.105 83.6565 18.7056 60.7391 0.0040362 0 -40 10
1.751 5.06528e-08 2.53992e-06 0.147087 0.147086 0.0120265 2.3024e-05 0.00115451 0.183858 0.00065881 0.184513 0.950946 101.447 0.235059 0.85373 4.55306 0.0649408 0.0429534 0.957047 0.0194379 0.00459623 0.0186948 0.00438456 0.00556211 0.00630522 0.222484 0.252209 58.049 -87.8991 126.158 15.9351 145.036 0.00014225 0.267315 192.727 0.310193 0.0673251 0.00409848 0.000562378 0.00138509 0.98696 0.991716 -2.9901e-06 -85.6571 0.0930852 31169 310.134 0.983498 0.319146 0.737924 0.73792 9.99958 2.98645e-06 1.19457e-05 0.134247 0.983406 0.931368 -0.0132916 4.93048e-06 0.515932 -2.01221e-20 7.46423e-24 -2.01146e-20 0.00139645 0.997815 8.60226e-05 0.152732 2.85279 0.00139645 0.997815 0.789549 0.00106743 0.00188139 0.000860226 0.455387 0.00188139 0.444449 0.000131235 1.02 0.88876 0.534378 0.287549 1.71944e-07 3.08411e-09 2370.93 3137.95 -0.0580839 0.482207 0.277276 0.254711 -0.593083 -0.169573 0.488001 -0.265805 -0.222205 2.653 1 0 295.451 0 2.23381 2.651 0.000299127 0.866864 0.699985 0.315984 0.43407 2.23399 139.112 83.6559 18.7056 60.7388 0.00403623 0 -40 10
1.752 5.06817e-08 2.53992e-06 0.14712 0.147119 0.0120265 2.30371e-05 0.00115451 0.1839 0.000658811 0.184554 0.951036 101.446 0.235048 0.853862 4.55368 0.0649516 0.0429593 0.957041 0.0194373 0.00459668 0.0186942 0.00438495 0.00556267 0.0063058 0.222507 0.252232 58.0491 -87.8991 126.158 15.9351 145.036 0.000142253 0.267315 192.727 0.310192 0.067325 0.00409848 0.000562378 0.00138509 0.98696 0.991716 -2.99012e-06 -85.657 0.0930852 31169 310.146 0.983498 0.319146 0.737936 0.737931 9.99958 2.98646e-06 1.19457e-05 0.134252 0.983407 0.931367 -0.0132916 4.93051e-06 0.515952 -2.01237e-20 7.46486e-24 -2.01162e-20 0.00139646 0.997815 8.60227e-05 0.152732 2.85279 0.00139646 0.997815 0.789622 0.00106744 0.00188139 0.000860227 0.455387 0.00188139 0.444454 0.000131237 1.02 0.888761 0.534378 0.28755 1.71944e-07 3.08413e-09 2370.91 3138 -0.0580889 0.482207 0.277276 0.254714 -0.593083 -0.169573 0.487985 -0.265803 -0.222191 2.654 1 0 295.446 0 2.23395 2.652 0.000299126 0.866892 0.700028 0.315943 0.434092 2.23413 139.119 83.6553 18.7055 60.7385 0.00403625 0 -40 10
1.753 5.07105e-08 2.53992e-06 0.147153 0.147152 0.0120264 2.30502e-05 0.00115451 0.183941 0.000658812 0.184595 0.951127 101.446 0.235038 0.853995 4.55431 0.0649623 0.0429652 0.957035 0.0194368 0.00459713 0.0186936 0.00438534 0.00556323 0.00630637 0.222529 0.252255 58.0492 -87.8991 126.158 15.935 145.036 0.000142255 0.267315 192.727 0.310192 0.067325 0.00409849 0.000562379 0.00138509 0.98696 0.991716 -2.99013e-06 -85.657 0.0930853 31169 310.158 0.983498 0.319146 0.737948 0.737943 9.99958 2.98646e-06 1.19457e-05 0.134256 0.983407 0.931366 -0.0132916 4.93054e-06 0.515972 -2.01252e-20 7.46549e-24 -2.01178e-20 0.00139646 0.997815 8.60228e-05 0.152732 2.85279 0.00139646 0.997815 0.789695 0.00106746 0.00188139 0.000860228 0.455387 0.00188139 0.44446 0.00013124 1.02 0.888762 0.534377 0.287552 1.71945e-07 3.08415e-09 2370.89 3138.05 -0.0580939 0.482208 0.277276 0.254717 -0.593082 -0.169573 0.487969 -0.265801 -0.222177 2.655 1 0 295.442 0 2.23409 2.653 0.000299124 0.86692 0.700071 0.315902 0.434114 2.23427 139.127 83.6547 18.7055 60.7382 0.00403628 0 -40 10
1.754 5.07394e-08 2.53992e-06 0.147186 0.147185 0.0120264 2.30634e-05 0.00115451 0.183982 0.000658812 0.184637 0.951217 101.445 0.235027 0.854128 4.55493 0.0649731 0.042971 0.957029 0.0194362 0.00459759 0.0186931 0.00438573 0.00556379 0.00630695 0.222551 0.252278 58.0492 -87.8991 126.158 15.935 145.036 0.000142257 0.267315 192.727 0.310192 0.0673249 0.00409849 0.00056238 0.0013851 0.98696 0.991716 -2.99015e-06 -85.657 0.0930854 31169 310.17 0.983497 0.319146 0.73796 0.737955 9.99958 2.98647e-06 1.19458e-05 0.134261 0.983407 0.931365 -0.0132916 4.93057e-06 0.515991 -2.01268e-20 7.46612e-24 -2.01194e-20 0.00139646 0.997815 8.60229e-05 0.152732 2.85279 0.00139646 0.997815 0.789768 0.00106747 0.00188139 0.000860229 0.455387 0.00188139 0.444465 0.000131242 1.02 0.888763 0.534377 0.287553 1.71945e-07 3.08417e-09 2370.88 3138.1 -0.0580989 0.482208 0.277275 0.25472 -0.593082 -0.169573 0.487953 -0.265799 -0.222164 2.656 1 0 295.437 0 2.23422 2.654 0.000299123 0.866949 0.700113 0.315861 0.434136 2.2344 139.134 83.6542 18.7055 60.7379 0.0040363 0 -40 10
1.755 5.07682e-08 2.53992e-06 0.147219 0.147218 0.0120264 2.30765e-05 0.00115451 0.184024 0.000658813 0.184678 0.951307 101.444 0.235016 0.85426 4.55555 0.0649838 0.0429769 0.957023 0.0194357 0.00459804 0.0186925 0.00438612 0.00556435 0.00630752 0.222574 0.252301 58.0493 -87.8991 126.158 15.935 145.036 0.00014226 0.267316 192.727 0.310191 0.0673249 0.00409849 0.00056238 0.0013851 0.98696 0.991716 -2.99016e-06 -85.657 0.0930855 31169 310.183 0.983497 0.319146 0.737971 0.737967 9.99958 2.98647e-06 1.19458e-05 0.134266 0.983408 0.931364 -0.0132916 4.9306e-06 0.516011 -2.01284e-20 7.46675e-24 -2.01209e-20 0.00139646 0.997815 8.6023e-05 0.152732 2.85279 0.00139646 0.997815 0.789841 0.00106749 0.00188139 0.00086023 0.455386 0.00188139 0.44447 0.000131245 1.02 0.888765 0.534377 0.287555 1.71945e-07 3.0842e-09 2370.86 3138.15 -0.0581039 0.482208 0.277275 0.254723 -0.593081 -0.169573 0.487937 -0.265797 -0.22215 2.657 1 0 295.433 0 2.23436 2.655 0.000299122 0.866977 0.700156 0.31582 0.434158 2.23454 139.141 83.6536 18.7054 60.7377 0.00403632 0 -40 10
1.756 5.07971e-08 2.53993e-06 0.147252 0.147251 0.0120264 2.30896e-05 0.00115451 0.184065 0.000658813 0.184719 0.951397 101.444 0.235005 0.854393 4.55618 0.0649946 0.0429828 0.957017 0.0194351 0.00459849 0.0186919 0.00438652 0.0055649 0.0063081 0.222596 0.252324 58.0494 -87.8992 126.157 15.9349 145.036 0.000142262 0.267316 192.726 0.310191 0.0673248 0.00409849 0.000562381 0.0013851 0.98696 0.991716 -2.99018e-06 -85.657 0.0930856 31168.9 310.195 0.983497 0.319146 0.737983 0.737979 9.99958 2.98648e-06 1.19458e-05 0.13427 0.983408 0.931363 -0.0132916 4.93063e-06 0.516031 -2.013e-20 7.46739e-24 -2.01225e-20 0.00139646 0.997815 8.6023e-05 0.152732 2.85279 0.00139646 0.997815 0.789914 0.00106751 0.0018814 0.00086023 0.455386 0.00188139 0.444475 0.000131247 1.02 0.888766 0.534376 0.287556 1.71946e-07 3.08422e-09 2370.85 3138.2 -0.058109 0.482208 0.277275 0.254727 -0.59308 -0.169573 0.487921 -0.265795 -0.222136 2.658 1 0 295.428 0 2.2345 2.656 0.000299121 0.867006 0.700199 0.315779 0.434181 2.23468 139.149 83.653 18.7054 60.7374 0.00403635 0 -40 10
1.757 5.08259e-08 2.53993e-06 0.147285 0.147284 0.0120264 2.31027e-05 0.00115451 0.184106 0.000658814 0.18476 0.951487 101.443 0.234995 0.854526 4.5568 0.0650053 0.0429887 0.957011 0.0194345 0.00459895 0.0186913 0.00438691 0.00556546 0.00630868 0.222619 0.252347 58.0494 -87.8992 126.157 15.9349 145.036 0.000142264 0.267316 192.726 0.31019 0.0673248 0.0040985 0.000562382 0.0013851 0.98696 0.991716 -2.99019e-06 -85.657 0.0930857 31168.9 310.207 0.983497 0.319146 0.737995 0.737991 9.99958 2.98648e-06 1.19458e-05 0.134275 0.983408 0.931362 -0.0132916 4.93066e-06 0.516051 -2.01316e-20 7.46802e-24 -2.01241e-20 0.00139646 0.997815 8.60231e-05 0.152733 2.85279 0.00139646 0.997815 0.789987 0.00106752 0.0018814 0.000860231 0.455386 0.0018814 0.44448 0.00013125 1.02 0.888767 0.534376 0.287558 1.71946e-07 3.08424e-09 2370.83 3138.25 -0.058114 0.482208 0.277275 0.25473 -0.59308 -0.169574 0.487905 -0.265793 -0.222122 2.659 1 0 295.424 0 2.23464 2.657 0.00029912 0.867034 0.700242 0.315739 0.434203 2.23482 139.156 83.6524 18.7053 60.7371 0.00403637 0 -40 10
1.758 5.08547e-08 2.53993e-06 0.147318 0.147317 0.0120264 2.31158e-05 0.00115451 0.184147 0.000658814 0.184802 0.951577 101.443 0.234984 0.854658 4.55743 0.0650161 0.0429946 0.957005 0.019434 0.0045994 0.0186907 0.0043873 0.00556602 0.00630925 0.222641 0.25237 58.0495 -87.8992 126.157 15.9349 145.036 0.000142266 0.267316 192.726 0.31019 0.0673247 0.0040985 0.000562382 0.00138511 0.98696 0.991716 -2.99021e-06 -85.657 0.0930858 31168.9 310.22 0.983497 0.319146 0.738007 0.738003 9.99958 2.98649e-06 1.19458e-05 0.134279 0.983408 0.931361 -0.0132916 4.93069e-06 0.51607 -2.01331e-20 7.46865e-24 -2.01257e-20 0.00139646 0.997815 8.60232e-05 0.152733 2.85279 0.00139646 0.997815 0.79006 0.00106754 0.0018814 0.000860232 0.455386 0.0018814 0.444486 0.000131252 1.02 0.888768 0.534376 0.287559 1.71946e-07 3.08427e-09 2370.81 3138.3 -0.058119 0.482208 0.277274 0.254733 -0.593079 -0.169574 0.487889 -0.26579 -0.222108 2.66 1 0 295.419 0 2.23477 2.658 0.000299118 0.867063 0.700285 0.315698 0.434225 2.23495 139.163 83.6518 18.7053 60.7368 0.0040364 0 -40 10
1.759 5.08836e-08 2.53993e-06 0.147351 0.14735 0.0120264 2.31289e-05 0.00115451 0.184189 0.000658815 0.184843 0.951667 101.442 0.234973 0.854791 4.55806 0.0650268 0.0430005 0.956999 0.0194334 0.00459986 0.0186902 0.00438769 0.00556658 0.00630983 0.222663 0.252393 58.0495 -87.8992 126.157 15.9348 145.036 0.000142269 0.267316 192.726 0.310189 0.0673247 0.0040985 0.000562383 0.00138511 0.986959 0.991716 -2.99022e-06 -85.657 0.0930859 31168.9 310.232 0.983497 0.319146 0.738019 0.738014 9.99958 2.98649e-06 1.19459e-05 0.134284 0.983409 0.93136 -0.0132916 4.93072e-06 0.51609 -2.01347e-20 7.46928e-24 -2.01272e-20 0.00139646 0.997815 8.60233e-05 0.152733 2.85279 0.00139646 0.997815 0.790133 0.00106756 0.0018814 0.000860233 0.455385 0.0018814 0.444491 0.000131254 1.02 0.888769 0.534376 0.287561 1.71946e-07 3.08429e-09 2370.8 3138.35 -0.058124 0.482208 0.277274 0.254736 -0.593078 -0.169574 0.487873 -0.265788 -0.222094 2.661 1 0 295.415 0 2.23491 2.659 0.000299117 0.867091 0.700328 0.315657 0.434247 2.23509 139.171 83.6512 18.7053 60.7365 0.00403642 0 -40 10
1.76 5.09124e-08 2.53993e-06 0.147384 0.147383 0.0120263 2.3142e-05 0.00115451 0.18423 0.000658815 0.184884 0.951757 101.441 0.234962 0.854924 4.55868 0.0650376 0.0430064 0.956994 0.0194329 0.00460031 0.0186896 0.00438809 0.00556714 0.0063104 0.222686 0.252416 58.0496 -87.8992 126.157 15.9348 145.036 0.000142271 0.267317 192.726 0.310189 0.0673246 0.00409851 0.000562384 0.00138511 0.986959 0.991716 -2.99024e-06 -85.657 0.0930859 31168.8 310.244 0.983497 0.319146 0.738031 0.738026 9.99958 2.9865e-06 1.19459e-05 0.134289 0.983409 0.931359 -0.0132916 4.93075e-06 0.51611 -2.01363e-20 7.46991e-24 -2.01288e-20 0.00139646 0.997815 8.60234e-05 0.152733 2.85279 0.00139646 0.997815 0.790205 0.00106757 0.0018814 0.000860234 0.455385 0.0018814 0.444496 0.000131257 1.02 0.88877 0.534375 0.287562 1.71947e-07 3.08431e-09 2370.78 3138.4 -0.058129 0.482208 0.277274 0.254739 -0.593078 -0.169574 0.487857 -0.265786 -0.222081 2.662 1 0 295.41 0 2.23505 2.66 0.000299116 0.86712 0.700371 0.315617 0.434269 2.23523 139.178 83.6507 18.7052 60.7362 0.00403644 0 -40 10
1.761 5.09413e-08 2.53993e-06 0.147417 0.147416 0.0120263 2.31551e-05 0.00115452 0.184271 0.000658816 0.184925 0.951847 101.441 0.234952 0.855056 4.55931 0.0650483 0.0430124 0.956988 0.0194323 0.00460077 0.018689 0.00438848 0.0055677 0.00631098 0.222708 0.252439 58.0497 -87.8992 126.156 15.9347 145.036 0.000142273 0.267317 192.726 0.310189 0.0673246 0.00409851 0.000562384 0.00138511 0.986959 0.991716 -2.99025e-06 -85.657 0.093086 31168.8 310.257 0.983497 0.319146 0.738043 0.738038 9.99958 2.9865e-06 1.19459e-05 0.134293 0.983409 0.931358 -0.0132916 4.93078e-06 0.51613 -2.01379e-20 7.47054e-24 -2.01304e-20 0.00139647 0.997815 8.60235e-05 0.152733 2.8528 0.00139647 0.997815 0.790278 0.00106759 0.0018814 0.000860235 0.455385 0.0018814 0.444501 0.000131259 1.02 0.888771 0.534375 0.287564 1.71947e-07 3.08433e-09 2370.76 3138.45 -0.058134 0.482208 0.277273 0.254742 -0.593077 -0.169574 0.487842 -0.265784 -0.222067 2.663 1 0 295.406 0 2.23518 2.661 0.000299115 0.867148 0.700414 0.315576 0.434292 2.23536 139.186 83.6501 18.7052 60.736 0.00403647 0 -40 10
1.762 5.09701e-08 2.53994e-06 0.147449 0.147449 0.0120263 2.31682e-05 0.00115452 0.184312 0.000658816 0.184966 0.951938 101.44 0.234941 0.855189 4.55994 0.0650591 0.0430183 0.956982 0.0194317 0.00460122 0.0186884 0.00438887 0.00556826 0.00631156 0.222731 0.252462 58.0497 -87.8992 126.156 15.9347 145.036 0.000142276 0.267317 192.725 0.310188 0.0673245 0.00409851 0.000562385 0.00138511 0.986959 0.991716 -2.99027e-06 -85.6569 0.0930861 31168.8 310.269 0.983497 0.319146 0.738055 0.73805 9.99958 2.98651e-06 1.19459e-05 0.134298 0.98341 0.931357 -0.0132916 4.93081e-06 0.516149 -2.01395e-20 7.47118e-24 -2.0132e-20 0.00139647 0.997815 8.60235e-05 0.152733 2.8528 0.00139647 0.997815 0.790351 0.0010676 0.0018814 0.000860235 0.455385 0.0018814 0.444506 0.000131262 1.02 0.888772 0.534375 0.287565 1.71947e-07 3.08436e-09 2370.75 3138.5 -0.058139 0.482208 0.277273 0.254746 -0.593077 -0.169574 0.487826 -0.265782 -0.222053 2.664 1 0 295.401 0 2.23532 2.662 0.000299113 0.867177 0.700457 0.315535 0.434314 2.2355 139.193 83.6495 18.7052 60.7357 0.00403649 0 -40 10
1.763 5.0999e-08 2.53994e-06 0.147482 0.147482 0.0120263 2.31813e-05 0.00115452 0.184353 0.000658817 0.185007 0.952028 101.439 0.23493 0.855322 4.56057 0.0650698 0.0430242 0.956976 0.0194312 0.00460168 0.0186879 0.00438926 0.00556883 0.00631214 0.222753 0.252485 58.0498 -87.8992 126.156 15.9347 145.036 0.000142278 0.267317 192.725 0.310188 0.0673245 0.00409852 0.000562386 0.00138512 0.986959 0.991716 -2.99028e-06 -85.6569 0.0930862 31168.8 310.282 0.983497 0.319146 0.738066 0.738062 9.99958 2.98651e-06 1.19459e-05 0.134303 0.98341 0.931356 -0.0132916 4.93084e-06 0.516169 -2.0141e-20 7.47181e-24 -2.01336e-20 0.00139647 0.997815 8.60236e-05 0.152733 2.8528 0.00139647 0.997815 0.790424 0.00106762 0.00188141 0.000860236 0.455384 0.0018814 0.444512 0.000131264 1.02 0.888773 0.534374 0.287567 1.71947e-07 3.08438e-09 2370.73 3138.55 -0.058144 0.482208 0.277273 0.254749 -0.593076 -0.169574 0.48781 -0.26578 -0.222039 2.665 1 0 295.397 0 2.23546 2.663 0.000299112 0.867205 0.7005 0.315495 0.434336 2.23564 139.2 83.6489 18.7051 60.7354 0.00403652 0 -40 10
1.764 5.10278e-08 2.53994e-06 0.147515 0.147515 0.0120263 2.31945e-05 0.00115452 0.184394 0.000658817 0.185048 0.952118 101.439 0.234919 0.855455 4.56119 0.0650806 0.0430301 0.95697 0.0194306 0.00460213 0.0186873 0.00438966 0.00556939 0.00631271 0.222775 0.252509 58.0499 -87.8992 126.156 15.9346 145.036 0.00014228 0.267317 192.725 0.310187 0.0673244 0.00409852 0.000562386 0.00138512 0.986959 0.991716 -2.9903e-06 -85.6569 0.0930863 31168.8 310.294 0.983497 0.319146 0.738078 0.738074 9.99958 2.98652e-06 1.1946e-05 0.134307 0.98341 0.931355 -0.0132916 4.93087e-06 0.516189 -2.01426e-20 7.47244e-24 -2.01351e-20 0.00139647 0.997815 8.60237e-05 0.152734 2.8528 0.00139647 0.997815 0.790496 0.00106764 0.00188141 0.000860237 0.455384 0.00188141 0.444517 0.000131266 1.02 0.888774 0.534374 0.287568 1.71948e-07 3.0844e-09 2370.71 3138.6 -0.0581491 0.482208 0.277273 0.254752 -0.593075 -0.169574 0.487794 -0.265778 -0.222025 2.666 1 0 295.392 0 2.2356 2.664 0.000299111 0.867234 0.700543 0.315454 0.434358 2.23578 139.208 83.6483 18.7051 60.7351 0.00403654 0 -40 10
1.765 5.10566e-08 2.53994e-06 0.147548 0.147547 0.0120263 2.32076e-05 0.00115452 0.184435 0.000658818 0.185089 0.952208 101.438 0.234909 0.855587 4.56182 0.0650913 0.0430361 0.956964 0.0194301 0.00460259 0.0186867 0.00439005 0.00556995 0.00631329 0.222798 0.252532 58.0499 -87.8992 126.155 15.9346 145.036 0.000142282 0.267318 192.725 0.310187 0.0673244 0.00409852 0.000562387 0.00138512 0.986959 0.991716 -2.99031e-06 -85.6569 0.0930864 31168.7 310.306 0.983497 0.319146 0.73809 0.738086 9.99958 2.98652e-06 1.1946e-05 0.134312 0.98341 0.931354 -0.0132916 4.9309e-06 0.516209 -2.01442e-20 7.47308e-24 -2.01367e-20 0.00139647 0.997815 8.60238e-05 0.152734 2.8528 0.00139647 0.997815 0.790569 0.00106765 0.00188141 0.000860238 0.455384 0.00188141 0.444522 0.000131269 1.02 0.888776 0.534374 0.28757 1.71948e-07 3.08443e-09 2370.7 3138.65 -0.0581541 0.482208 0.277272 0.254755 -0.593075 -0.169574 0.487778 -0.265776 -0.222011 2.667 1 0 295.388 0 2.23573 2.665 0.00029911 0.867262 0.700586 0.315414 0.43438 2.23591 139.215 83.6477 18.7051 60.7348 0.00403657 0 -40 10
1.766 5.10855e-08 2.53994e-06 0.147581 0.14758 0.0120263 2.32207e-05 0.00115452 0.184476 0.000658818 0.18513 0.952298 101.438 0.234898 0.85572 4.56245 0.0651021 0.043042 0.956958 0.0194295 0.00460304 0.0186861 0.00439045 0.00557051 0.00631387 0.22282 0.252555 58.05 -87.8992 126.155 15.9346 145.036 0.000142285 0.267318 192.725 0.310186 0.0673243 0.00409852 0.000562388 0.00138512 0.986959 0.991716 -2.99033e-06 -85.6569 0.0930865 31168.7 310.319 0.983497 0.319146 0.738102 0.738098 9.99958 2.98653e-06 1.1946e-05 0.134317 0.983411 0.931353 -0.0132916 4.93093e-06 0.516228 -2.01458e-20 7.47371e-24 -2.01383e-20 0.00139647 0.997815 8.60239e-05 0.152734 2.8528 0.00139647 0.997815 0.790642 0.00106767 0.00188141 0.000860239 0.455384 0.00188141 0.444527 0.000131271 1.02 0.888777 0.534373 0.287571 1.71948e-07 3.08445e-09 2370.68 3138.7 -0.0581591 0.482209 0.277272 0.254758 -0.593074 -0.169574 0.487762 -0.265774 -0.221997 2.668 1 0 295.383 0 2.23587 2.666 0.000299109 0.867291 0.700629 0.315373 0.434403 2.23605 139.222 83.6471 18.705 60.7346 0.00403659 0 -40 10
1.767 5.11143e-08 2.53994e-06 0.147613 0.147613 0.0120262 2.32338e-05 0.00115452 0.184517 0.000658819 0.185171 0.952389 101.437 0.234887 0.855853 4.56308 0.0651129 0.0430479 0.956952 0.0194289 0.0046035 0.0186856 0.00439084 0.00557107 0.00631445 0.222843 0.252578 58.05 -87.8992 126.155 15.9345 145.036 0.000142287 0.267318 192.725 0.310186 0.0673242 0.00409853 0.000562388 0.00138512 0.986959 0.991716 -2.99034e-06 -85.6569 0.0930866 31168.7 310.331 0.983497 0.319146 0.738114 0.73811 9.99958 2.98653e-06 1.1946e-05 0.134321 0.983411 0.931352 -0.0132916 4.93096e-06 0.516248 -2.01474e-20 7.47434e-24 -2.01399e-20 0.00139647 0.997815 8.60239e-05 0.152734 2.8528 0.00139647 0.997815 0.790714 0.00106769 0.00188141 0.000860239 0.455384 0.00188141 0.444532 0.000131274 1.02 0.888778 0.534373 0.287573 1.71949e-07 3.08447e-09 2370.67 3138.75 -0.0581641 0.482209 0.277272 0.254762 -0.593073 -0.169574 0.487746 -0.265772 -0.221984 2.669 1 0 295.379 0 2.23601 2.667 0.000299107 0.867319 0.700672 0.315333 0.434425 2.23619 139.23 83.6466 18.705 60.7343 0.00403661 0 -40 10
1.768 5.11432e-08 2.53995e-06 0.147646 0.147645 0.0120262 2.32469e-05 0.00115452 0.184557 0.000658819 0.185212 0.952479 101.436 0.234876 0.855986 4.56371 0.0651236 0.0430539 0.956946 0.0194284 0.00460395 0.018685 0.00439123 0.00557163 0.00631503 0.222865 0.252601 58.0501 -87.8992 126.155 15.9345 145.036 0.000142289 0.267318 192.724 0.310186 0.0673242 0.00409853 0.000562389 0.00138513 0.986959 0.991716 -2.99036e-06 -85.6569 0.0930866 31168.7 310.343 0.983497 0.319146 0.738126 0.738121 9.99958 2.98654e-06 1.1946e-05 0.134326 0.983411 0.931351 -0.0132916 4.93099e-06 0.516268 -2.0149e-20 7.47498e-24 -2.01415e-20 0.00139647 0.997815 8.6024e-05 0.152734 2.8528 0.00139647 0.997815 0.790787 0.0010677 0.00188141 0.00086024 0.455383 0.00188141 0.444537 0.000131276 1.02 0.888779 0.534373 0.287575 1.71949e-07 3.08449e-09 2370.65 3138.8 -0.0581691 0.482209 0.277271 0.254765 -0.593073 -0.169574 0.48773 -0.26577 -0.22197 2.67 1 0 295.374 0 2.23614 2.668 0.000299106 0.867348 0.700715 0.315293 0.434447 2.23632 139.237 83.646 18.705 60.734 0.00403664 0 -40 10
1.769 5.1172e-08 2.53995e-06 0.147679 0.147678 0.0120262 2.326e-05 0.00115452 0.184598 0.00065882 0.185252 0.952569 101.436 0.234866 0.856119 4.56434 0.0651344 0.0430598 0.95694 0.0194278 0.00460441 0.0186844 0.00439163 0.0055722 0.00631561 0.222888 0.252624 58.0502 -87.8992 126.155 15.9344 145.036 0.000142292 0.267318 192.724 0.310185 0.0673241 0.00409853 0.00056239 0.00138513 0.986959 0.991716 -2.99037e-06 -85.6569 0.0930867 31168.6 310.356 0.983497 0.319146 0.738138 0.738133 9.99958 2.98654e-06 1.19461e-05 0.13433 0.983411 0.93135 -0.0132916 4.93102e-06 0.516288 -2.01505e-20 7.47561e-24 -2.01431e-20 0.00139648 0.997815 8.60241e-05 0.152734 2.8528 0.00139648 0.997815 0.790859 0.00106772 0.00188142 0.000860241 0.455383 0.00188141 0.444543 0.000131278 1.02 0.88878 0.534372 0.287576 1.71949e-07 3.08452e-09 2370.63 3138.85 -0.0581742 0.482209 0.277271 0.254768 -0.593072 -0.169574 0.487714 -0.265767 -0.221956 2.671 1 0 295.369 0 2.23628 2.669 0.000299105 0.867376 0.700758 0.315252 0.434469 2.23646 139.244 83.6454 18.7049 60.7337 0.00403666 0 -40 10
1.77 5.12009e-08 2.53995e-06 0.147711 0.147711 0.0120262 2.32731e-05 0.00115452 0.184639 0.00065882 0.185293 0.95266 101.435 0.234855 0.856251 4.56497 0.0651451 0.0430658 0.956934 0.0194272 0.00460487 0.0186838 0.00439202 0.00557276 0.00631619 0.22291 0.252647 58.0502 -87.8992 126.154 15.9344 145.036 0.000142294 0.267318 192.724 0.310185 0.0673241 0.00409854 0.00056239 0.00138513 0.986959 0.991716 -2.99039e-06 -85.6569 0.0930868 31168.6 310.368 0.983497 0.319146 0.73815 0.738145 9.99958 2.98655e-06 1.19461e-05 0.134335 0.983412 0.931349 -0.0132916 4.93105e-06 0.516308 -2.01521e-20 7.47625e-24 -2.01447e-20 0.00139648 0.997815 8.60242e-05 0.152735 2.8528 0.00139648 0.997815 0.790932 0.00106773 0.00188142 0.000860242 0.455383 0.00188142 0.444548 0.000131281 1.02 0.888781 0.534372 0.287578 1.71949e-07 3.08454e-09 2370.62 3138.9 -0.0581792 0.482209 0.277271 0.254771 -0.593072 -0.169574 0.487698 -0.265765 -0.221942 2.672 1 0 295.365 0 2.23642 2.67 0.000299104 0.867405 0.7008 0.315212 0.434491 2.2366 139.252 83.6448 18.7049 60.7334 0.00403669 0 -40 10
1.771 5.12297e-08 2.53995e-06 0.147744 0.147743 0.0120262 2.32862e-05 0.00115452 0.18468 0.000658821 0.185334 0.95275 101.434 0.234844 0.856384 4.56561 0.0651559 0.0430718 0.956928 0.0194267 0.00460532 0.0186832 0.00439242 0.00557332 0.00631677 0.222933 0.252671 58.0503 -87.8992 126.154 15.9344 145.036 0.000142296 0.267319 192.724 0.310184 0.067324 0.00409854 0.000562391 0.00138513 0.986959 0.991716 -2.9904e-06 -85.6569 0.0930869 31168.6 310.381 0.983497 0.319146 0.738162 0.738157 9.99958 2.98655e-06 1.19461e-05 0.13434 0.983412 0.931348 -0.0132916 4.93108e-06 0.516328 -2.01537e-20 7.47688e-24 -2.01462e-20 0.00139648 0.997815 8.60243e-05 0.152735 2.8528 0.00139648 0.997815 0.791004 0.00106775 0.00188142 0.000860243 0.455383 0.00188142 0.444553 0.000131283 1.02 0.888782 0.534372 0.287579 1.7195e-07 3.08456e-09 2370.6 3138.95 -0.0581842 0.482209 0.277271 0.254774 -0.593071 -0.169574 0.487682 -0.265763 -0.221928 2.673 1 0 295.36 0 2.23655 2.671 0.000299102 0.867434 0.700843 0.315172 0.434513 2.23673 139.259 83.6442 18.7049 60.7331 0.00403671 0 -40 10
1.772 5.12585e-08 2.53995e-06 0.147776 0.147776 0.0120262 2.32993e-05 0.00115452 0.18472 0.000658821 0.185375 0.95284 101.434 0.234833 0.856517 4.56624 0.0651667 0.0430777 0.956922 0.0194261 0.00460578 0.0186827 0.00439281 0.00557389 0.00631735 0.222955 0.252694 58.0504 -87.8992 126.154 15.9343 145.036 0.000142298 0.267319 192.724 0.310184 0.067324 0.00409854 0.000562392 0.00138514 0.986959 0.991716 -2.99042e-06 -85.6569 0.093087 31168.6 310.393 0.983497 0.319146 0.738173 0.738169 9.99958 2.98656e-06 1.19461e-05 0.134344 0.983412 0.931347 -0.0132916 4.93111e-06 0.516348 -2.01553e-20 7.47752e-24 -2.01478e-20 0.00139648 0.997815 8.60243e-05 0.152735 2.85281 0.00139648 0.997815 0.791077 0.00106777 0.00188142 0.000860243 0.455382 0.00188142 0.444558 0.000131286 1.02 0.888783 0.534372 0.287581 1.7195e-07 3.08459e-09 2370.58 3139 -0.0581892 0.482209 0.27727 0.254778 -0.59307 -0.169575 0.487666 -0.265761 -0.221914 2.674 1 0 295.356 0 2.23669 2.672 0.000299101 0.867462 0.700886 0.315131 0.434536 2.23687 139.266 83.6436 18.7048 60.7329 0.00403674 0 -40 10
1.773 5.12874e-08 2.53995e-06 0.147809 0.147808 0.0120262 2.33124e-05 0.00115452 0.184761 0.000658822 0.185415 0.952931 101.433 0.234823 0.85665 4.56687 0.0651774 0.0430837 0.956916 0.0194256 0.00460624 0.0186821 0.00439321 0.00557445 0.00631793 0.222978 0.252717 58.0504 -87.8992 126.154 15.9343 145.036 0.000142301 0.267319 192.724 0.310183 0.0673239 0.00409855 0.000562392 0.00138514 0.986959 0.991716 -2.99043e-06 -85.6568 0.0930871 31168.6 310.406 0.983497 0.319146 0.738185 0.738181 9.99958 2.98656e-06 1.19461e-05 0.134349 0.983413 0.931346 -0.0132916 4.93114e-06 0.516367 -2.01569e-20 7.47815e-24 -2.01494e-20 0.00139648 0.997815 8.60244e-05 0.152735 2.85281 0.00139648 0.997815 0.791149 0.00106778 0.00188142 0.000860244 0.455382 0.00188142 0.444563 0.000131288 1.02 0.888784 0.534371 0.287582 1.7195e-07 3.08461e-09 2370.57 3139.05 -0.0581943 0.482209 0.27727 0.254781 -0.59307 -0.169575 0.48765 -0.265759 -0.2219 2.675 1 0 295.351 0 2.23683 2.673 0.0002991 0.867491 0.700929 0.315091 0.434558 2.23701 139.274 83.643 18.7048 60.7326 0.00403676 0 -40 10
1.774 5.13162e-08 2.53996e-06 0.147841 0.147841 0.0120261 2.33256e-05 0.00115453 0.184802 0.000658822 0.185456 0.953021 101.432 0.234812 0.856783 4.5675 0.0651882 0.0430897 0.95691 0.019425 0.00460669 0.0186815 0.0043936 0.00557501 0.00631851 0.223 0.25274 58.0505 -87.8992 126.154 15.9343 145.036 0.000142303 0.267319 192.723 0.310183 0.0673239 0.00409855 0.000562393 0.00138514 0.986959 0.991716 -2.99045e-06 -85.6568 0.0930872 31168.5 310.418 0.983497 0.319146 0.738197 0.738193 9.99958 2.98657e-06 1.19462e-05 0.134354 0.983413 0.931345 -0.0132916 4.93117e-06 0.516387 -2.01585e-20 7.47879e-24 -2.0151e-20 0.00139648 0.997815 8.60245e-05 0.152735 2.85281 0.00139648 0.997815 0.791222 0.0010678 0.00188142 0.000860245 0.455382 0.00188142 0.444568 0.00013129 1.02 0.888785 0.534371 0.287584 1.7195e-07 3.08463e-09 2370.55 3139.1 -0.0581993 0.482209 0.27727 0.254784 -0.593069 -0.169575 0.487634 -0.265757 -0.221886 2.676 1 0 295.347 0 2.23697 2.674 0.000299099 0.867519 0.700972 0.315051 0.43458 2.23714 139.281 83.6425 18.7048 60.7323 0.00403678 0 -40 10
1.775 5.13451e-08 2.53996e-06 0.147874 0.147873 0.0120261 2.33387e-05 0.00115453 0.184842 0.000658823 0.185497 0.953111 101.432 0.234801 0.856916 4.56814 0.065199 0.0430956 0.956904 0.0194244 0.00460715 0.0186809 0.004394 0.00557558 0.00631909 0.223023 0.252764 58.0505 -87.8992 126.153 15.9342 145.036 0.000142305 0.267319 192.723 0.310183 0.0673238 0.00409855 0.000562394 0.00138514 0.986959 0.991716 -2.99046e-06 -85.6568 0.0930873 31168.5 310.43 0.983497 0.319146 0.738209 0.738205 9.99958 2.98657e-06 1.19462e-05 0.134358 0.983413 0.931344 -0.0132916 4.93119e-06 0.516407 -2.01601e-20 7.47943e-24 -2.01526e-20 0.00139648 0.997815 8.60246e-05 0.152735 2.85281 0.00139648 0.997815 0.791294 0.00106782 0.00188142 0.000860246 0.455382 0.00188142 0.444574 0.000131293 1.02 0.888787 0.534371 0.287585 1.71951e-07 3.08465e-09 2370.53 3139.15 -0.0582043 0.482209 0.27727 0.254787 -0.593068 -0.169575 0.487618 -0.265755 -0.221873 2.677 1 0 295.342 0 2.2371 2.675 0.000299098 0.867548 0.701015 0.315011 0.434602 2.23728 139.288 83.6419 18.7047 60.732 0.00403681 0 -40 10
1.776 5.13739e-08 2.53996e-06 0.147906 0.147906 0.0120261 2.33518e-05 0.00115453 0.184883 0.000658823 0.185537 0.953202 101.431 0.23479 0.857049 4.56877 0.0652098 0.0431016 0.956898 0.0194239 0.00460761 0.0186803 0.0043944 0.00557614 0.00631967 0.223046 0.252787 58.0506 -87.8992 126.153 15.9342 145.036 0.000142308 0.26732 192.723 0.310182 0.0673238 0.00409856 0.000562394 0.00138514 0.986959 0.991716 -2.99048e-06 -85.6568 0.0930873 31168.5 310.443 0.983497 0.319146 0.738221 0.738217 9.99958 2.98658e-06 1.19462e-05 0.134363 0.983413 0.931343 -0.0132916 4.93122e-06 0.516427 -2.01617e-20 7.48006e-24 -2.01542e-20 0.00139648 0.997815 8.60247e-05 0.152735 2.85281 0.00139648 0.997815 0.791367 0.00106783 0.00188143 0.000860247 0.455382 0.00188142 0.444579 0.000131295 1.02 0.888788 0.53437 0.287587 1.71951e-07 3.08468e-09 2370.52 3139.2 -0.0582093 0.482209 0.277269 0.25479 -0.593068 -0.169575 0.487602 -0.265753 -0.221859 2.678 1 0 295.338 0 2.23724 2.676 0.000299096 0.867577 0.701058 0.314971 0.434624 2.23742 139.296 83.6413 18.7047 60.7317 0.00403683 0 -40 10
1.777 5.14027e-08 2.53996e-06 0.147939 0.147938 0.0120261 2.33649e-05 0.00115453 0.184924 0.000658824 0.185578 0.953292 101.431 0.234779 0.857182 4.5694 0.0652205 0.0431076 0.956892 0.0194233 0.00460807 0.0186797 0.00439479 0.0055767 0.00632025 0.223068 0.25281 58.0507 -87.8992 126.153 15.9341 145.036 0.00014231 0.26732 192.723 0.310182 0.0673237 0.00409856 0.000562395 0.00138515 0.986959 0.991716 -2.99049e-06 -85.6568 0.0930874 31168.5 310.455 0.983497 0.319146 0.738233 0.738229 9.99958 2.98658e-06 1.19462e-05 0.134368 0.983414 0.931342 -0.0132916 4.93125e-06 0.516447 -2.01633e-20 7.4807e-24 -2.01558e-20 0.00139648 0.997815 8.60247e-05 0.152736 2.85281 0.00139648 0.997815 0.791439 0.00106785 0.00188143 0.000860247 0.455381 0.00188143 0.444584 0.000131298 1.02 0.888789 0.53437 0.287588 1.71951e-07 3.0847e-09 2370.5 3139.25 -0.0582144 0.482209 0.277269 0.254794 -0.593067 -0.169575 0.487586 -0.265751 -0.221845 2.679 1 0 295.333 0 2.23738 2.677 0.000299095 0.867605 0.701101 0.31493 0.434646 2.23756 139.303 83.6407 18.7047 60.7314 0.00403686 0 -40 10
1.778 5.14316e-08 2.53996e-06 0.147971 0.147971 0.0120261 2.3378e-05 0.00115453 0.184964 0.000658824 0.185618 0.953382 101.43 0.234769 0.857315 4.57004 0.0652313 0.0431136 0.956886 0.0194227 0.00460853 0.0186792 0.00439519 0.00557727 0.00632083 0.223091 0.252833 58.0507 -87.8992 126.153 15.9341 145.036 0.000142312 0.26732 192.723 0.310181 0.0673237 0.00409856 0.000562396 0.00138515 0.986959 0.991716 -2.99051e-06 -85.6568 0.0930875 31168.4 310.468 0.983497 0.319146 0.738245 0.738241 9.99958 2.98659e-06 1.19462e-05 0.134372 0.983414 0.931341 -0.0132916 4.93128e-06 0.516467 -2.01649e-20 7.48134e-24 -2.01574e-20 0.00139649 0.997815 8.60248e-05 0.152736 2.85281 0.00139649 0.997815 0.791511 0.00106786 0.00188143 0.000860248 0.455381 0.00188143 0.444589 0.0001313 1.02 0.88879 0.53437 0.28759 1.71952e-07 3.08472e-09 2370.49 3139.3 -0.0582194 0.482209 0.277269 0.254797 -0.593067 -0.169575 0.48757 -0.265749 -0.221831 2.68 1 0 295.329 0 2.23751 2.678 0.000299094 0.867634 0.701144 0.31489 0.434668 2.23769 139.31 83.6401 18.7046 60.7312 0.00403688 0 -40 10
1.779 5.14604e-08 2.53996e-06 0.148004 0.148003 0.0120261 2.33911e-05 0.00115453 0.185005 0.000658825 0.185659 0.953473 101.429 0.234758 0.857448 4.57067 0.0652421 0.0431196 0.95688 0.0194222 0.00460898 0.0186786 0.00439558 0.00557783 0.00632142 0.223113 0.252857 58.0508 -87.8992 126.152 15.9341 145.036 0.000142315 0.26732 192.723 0.310181 0.0673236 0.00409856 0.000562396 0.00138515 0.986959 0.991716 -2.99052e-06 -85.6568 0.0930876 31168.4 310.48 0.983497 0.319146 0.738257 0.738253 9.99958 2.98659e-06 1.19463e-05 0.134377 0.983414 0.93134 -0.0132916 4.93131e-06 0.516487 -2.01665e-20 7.48197e-24 -2.0159e-20 0.00139649 0.997815 8.60249e-05 0.152736 2.85281 0.00139649 0.997815 0.791584 0.00106788 0.00188143 0.000860249 0.455381 0.00188143 0.444594 0.000131302 1.02 0.888791 0.534369 0.287591 1.71952e-07 3.08475e-09 2370.47 3139.35 -0.0582244 0.48221 0.277268 0.2548 -0.593066 -0.169575 0.487554 -0.265746 -0.221817 2.681 1 0 295.324 0 2.23765 2.679 0.000299093 0.867663 0.701186 0.31485 0.434691 2.23783 139.318 83.6395 18.7046 60.7309 0.00403691 0 -40 10
1.78 5.14893e-08 2.53997e-06 0.148036 0.148036 0.0120261 2.34042e-05 0.00115453 0.185045 0.000658825 0.185699 0.953563 101.429 0.234747 0.85758 4.57131 0.0652529 0.0431256 0.956874 0.0194216 0.00460944 0.018678 0.00439598 0.0055784 0.006322 0.223136 0.25288 58.0509 -87.8992 126.152 15.934 145.036 0.000142317 0.26732 192.722 0.31018 0.0673236 0.00409857 0.000562397 0.00138515 0.986959 0.991716 -2.99054e-06 -85.6568 0.0930877 31168.4 310.493 0.983497 0.319146 0.738269 0.738264 9.99958 2.9866e-06 1.19463e-05 0.134382 0.983414 0.931339 -0.0132916 4.93134e-06 0.516507 -2.01681e-20 7.48261e-24 -2.01606e-20 0.00139649 0.997815 8.6025e-05 0.152736 2.85281 0.00139649 0.997815 0.791656 0.0010679 0.00188143 0.00086025 0.455381 0.00188143 0.444599 0.000131305 1.02 0.888792 0.534369 0.287593 1.71952e-07 3.08477e-09 2370.45 3139.4 -0.0582295 0.48221 0.277268 0.254803 -0.593065 -0.169575 0.487538 -0.265744 -0.221803 2.682 1 0 295.32 0 2.23779 2.68 0.000299091 0.867692 0.701229 0.31481 0.434713 2.23797 139.325 83.6389 18.7046 60.7306 0.00403693 0 -40 10
1.781 5.15181e-08 2.53997e-06 0.148068 0.148068 0.0120261 2.34173e-05 0.00115453 0.185085 0.000658826 0.18574 0.953654 101.428 0.234736 0.857713 4.57195 0.0652636 0.0431316 0.956868 0.019421 0.0046099 0.0186774 0.00439638 0.00557897 0.00632258 0.223159 0.252903 58.0509 -87.8992 126.152 15.934 145.036 0.000142319 0.267321 192.722 0.31018 0.0673235 0.00409857 0.000562398 0.00138516 0.986959 0.991716 -2.99055e-06 -85.6568 0.0930878 31168.4 310.505 0.983497 0.319146 0.738281 0.738276 9.99958 2.9866e-06 1.19463e-05 0.134386 0.983415 0.931338 -0.0132916 4.93137e-06 0.516527 -2.01696e-20 7.48325e-24 -2.01622e-20 0.00139649 0.997815 8.60251e-05 0.152736 2.85281 0.00139649 0.997815 0.791728 0.00106791 0.00188143 0.000860251 0.45538 0.00188143 0.444604 0.000131307 1.02 0.888793 0.534369 0.287594 1.71952e-07 3.08479e-09 2370.44 3139.45 -0.0582345 0.48221 0.277268 0.254806 -0.593065 -0.169575 0.487522 -0.265742 -0.221789 2.683 1 0 295.315 0 2.23792 2.681 0.00029909 0.86772 0.701272 0.31477 0.434735 2.2381 139.333 83.6383 18.7045 60.7303 0.00403695 0 -40 10
1.782 5.1547e-08 2.53997e-06 0.148101 0.1481 0.012026 2.34304e-05 0.00115453 0.185126 0.000658826 0.18578 0.953744 101.427 0.234726 0.857846 4.57258 0.0652744 0.0431376 0.956862 0.0194205 0.00461036 0.0186768 0.00439677 0.00557953 0.00632316 0.223181 0.252927 58.051 -87.8992 126.152 15.934 145.036 0.000142321 0.267321 192.722 0.31018 0.0673235 0.00409857 0.000562398 0.00138516 0.986959 0.991716 -2.99057e-06 -85.6568 0.0930879 31168.3 310.518 0.983497 0.319146 0.738293 0.738288 9.99958 2.98661e-06 1.19463e-05 0.134391 0.983415 0.931337 -0.0132916 4.9314e-06 0.516547 -2.01712e-20 7.48389e-24 -2.01638e-20 0.00139649 0.997815 8.60251e-05 0.152736 2.85281 0.00139649 0.997815 0.7918 0.00106793 0.00188143 0.000860251 0.45538 0.00188143 0.44461 0.000131309 1.02 0.888794 0.534368 0.287596 1.71953e-07 3.08482e-09 2370.42 3139.5 -0.0582395 0.48221 0.277268 0.25481 -0.593064 -0.169575 0.487506 -0.26574 -0.221775 2.684 1 0 295.31 0 2.23806 2.682 0.000299089 0.867749 0.701315 0.31473 0.434757 2.23824 139.34 83.6378 18.7045 60.73 0.00403698 0 -40 10
1.783 5.15758e-08 2.53997e-06 0.148133 0.148132 0.012026 2.34435e-05 0.00115453 0.185166 0.000658827 0.18582 0.953835 101.427 0.234715 0.857979 4.57322 0.0652852 0.0431436 0.956856 0.0194199 0.00461082 0.0186763 0.00439717 0.0055801 0.00632375 0.223204 0.25295 58.051 -87.8993 126.152 15.9339 145.036 0.000142324 0.267321 192.722 0.310179 0.0673234 0.00409858 0.000562399 0.00138516 0.986959 0.991716 -2.99058e-06 -85.6568 0.093088 31168.3 310.53 0.983497 0.319146 0.738305 0.7383 9.99958 2.98661e-06 1.19463e-05 0.134396 0.983415 0.931336 -0.0132916 4.93143e-06 0.516567 -2.01728e-20 7.48452e-24 -2.01654e-20 0.00139649 0.997815 8.60252e-05 0.152737 2.85282 0.00139649 0.997815 0.791873 0.00106794 0.00188144 0.000860252 0.45538 0.00188143 0.444615 0.000131312 1.02 0.888795 0.534368 0.287597 1.71953e-07 3.08484e-09 2370.4 3139.55 -0.0582446 0.48221 0.277267 0.254813 -0.593063 -0.169575 0.48749 -0.265738 -0.221761 2.685 1 0 295.306 0 2.2382 2.683 0.000299088 0.867778 0.701358 0.31469 0.434779 2.23838 139.347 83.6372 18.7045 60.7297 0.004037 0 -40 10
1.784 5.16046e-08 2.53997e-06 0.148165 0.148165 0.012026 2.34567e-05 0.00115453 0.185207 0.000658828 0.185861 0.953925 101.426 0.234704 0.858113 4.57386 0.065296 0.0431496 0.95685 0.0194193 0.00461128 0.0186757 0.00439757 0.00558066 0.00632433 0.223227 0.252973 58.0511 -87.8993 126.151 15.9339 145.036 0.000142326 0.267321 192.722 0.310179 0.0673233 0.00409858 0.0005624 0.00138516 0.986959 0.991716 -2.9906e-06 -85.6567 0.093088 31168.3 310.543 0.983497 0.319146 0.738317 0.738312 9.99958 2.98662e-06 1.19464e-05 0.1344 0.983415 0.931335 -0.0132916 4.93146e-06 0.516587 -2.01744e-20 7.48516e-24 -2.0167e-20 0.00139649 0.997815 8.60253e-05 0.152737 2.85282 0.00139649 0.997815 0.791945 0.00106796 0.00188144 0.000860253 0.45538 0.00188144 0.44462 0.000131314 1.02 0.888796 0.534368 0.287599 1.71953e-07 3.08486e-09 2370.39 3139.6 -0.0582496 0.48221 0.277267 0.254816 -0.593063 -0.169575 0.487474 -0.265736 -0.221747 2.686 1 0 295.301 0 2.23833 2.684 0.000299087 0.867806 0.701401 0.314651 0.434801 2.23851 139.355 83.6366 18.7044 60.7295 0.00403703 0 -40 10
1.785 5.16335e-08 2.53997e-06 0.148197 0.148197 0.012026 2.34698e-05 0.00115453 0.185247 0.000658828 0.185901 0.954016 101.426 0.234693 0.858246 4.5745 0.0653068 0.0431556 0.956844 0.0194188 0.00461174 0.0186751 0.00439797 0.00558123 0.00632491 0.223249 0.252997 58.0512 -87.8993 126.151 15.9339 145.037 0.000142328 0.267321 192.722 0.310178 0.0673233 0.00409858 0.0005624 0.00138516 0.986959 0.991716 -2.99061e-06 -85.6567 0.0930881 31168.3 310.555 0.983497 0.319146 0.738329 0.738324 9.99958 2.98662e-06 1.19464e-05 0.134405 0.983416 0.931334 -0.0132916 4.93149e-06 0.516607 -2.0176e-20 7.4858e-24 -2.01685e-20 0.00139649 0.997815 8.60254e-05 0.152737 2.85282 0.00139649 0.997815 0.792017 0.00106798 0.00188144 0.000860254 0.45538 0.00188144 0.444625 0.000131317 1.02 0.888797 0.534368 0.2876 1.71953e-07 3.08488e-09 2370.37 3139.65 -0.0582546 0.48221 0.277267 0.254819 -0.593062 -0.169575 0.487458 -0.265734 -0.221734 2.687 1 0 295.297 0 2.23847 2.685 0.000299085 0.867835 0.701444 0.314611 0.434823 2.23865 139.362 83.636 18.7044 60.7292 0.00403705 0 -40 10
1.786 5.16623e-08 2.53998e-06 0.14823 0.148229 0.012026 2.34829e-05 0.00115453 0.185287 0.000658829 0.185941 0.954106 101.425 0.234682 0.858379 4.57513 0.0653176 0.0431616 0.956838 0.0194182 0.0046122 0.0186745 0.00439836 0.0055818 0.0063255 0.223272 0.25302 58.0512 -87.8993 126.151 15.9338 145.037 0.000142331 0.267322 192.721 0.310178 0.0673232 0.00409859 0.000562401 0.00138517 0.986959 0.991716 -2.99063e-06 -85.6567 0.0930882 31168.3 310.568 0.983497 0.319146 0.738341 0.738336 9.99958 2.98663e-06 1.19464e-05 0.13441 0.983416 0.931333 -0.0132916 4.93152e-06 0.516627 -2.01776e-20 7.48644e-24 -2.01701e-20 0.00139649 0.997815 8.60255e-05 0.152737 2.85282 0.00139649 0.997815 0.792089 0.00106799 0.00188144 0.000860255 0.455379 0.00188144 0.44463 0.000131319 1.02 0.888799 0.534367 0.287602 1.71954e-07 3.08491e-09 2370.35 3139.7 -0.0582597 0.48221 0.277266 0.254822 -0.593061 -0.169575 0.487442 -0.265732 -0.22172 2.688 1 0 295.292 0 2.23861 2.686 0.000299084 0.867864 0.701486 0.314571 0.434846 2.23879 139.369 83.6354 18.7044 60.7289 0.00403708 0 -40 10
1.787 5.16912e-08 2.53998e-06 0.148262 0.148261 0.012026 2.3496e-05 0.00115454 0.185327 0.000658829 0.185982 0.954197 101.424 0.234672 0.858512 4.57577 0.0653283 0.0431677 0.956832 0.0194176 0.00461266 0.0186739 0.00439876 0.00558236 0.00632608 0.223295 0.253043 58.0513 -87.8993 126.151 15.9338 145.037 0.000142333 0.267322 192.721 0.310177 0.0673232 0.00409859 0.000562402 0.00138517 0.986959 0.991716 -2.99064e-06 -85.6567 0.0930883 31168.2 310.58 0.983497 0.319146 0.738352 0.738348 9.99958 2.98663e-06 1.19464e-05 0.134414 0.983416 0.931332 -0.0132916 4.93155e-06 0.516647 -2.01792e-20 7.48708e-24 -2.01717e-20 0.0013965 0.997815 8.60255e-05 0.152737 2.85282 0.0013965 0.997815 0.792161 0.00106801 0.00188144 0.000860255 0.455379 0.00188144 0.444635 0.000131321 1.02 0.8888 0.534367 0.287603 1.71954e-07 3.08493e-09 2370.34 3139.75 -0.0582647 0.48221 0.277266 0.254826 -0.593061 -0.169575 0.487426 -0.26573 -0.221706 2.689 1 0 295.288 0 2.23874 2.687 0.000299083 0.867893 0.701529 0.314531 0.434868 2.23892 139.377 83.6348 18.7043 60.7286 0.0040371 0 -40 10
1.788 5.172e-08 2.53998e-06 0.148294 0.148293 0.012026 2.35091e-05 0.00115454 0.185367 0.00065883 0.186022 0.954287 101.424 0.234661 0.858645 4.57641 0.0653391 0.0431737 0.956826 0.0194171 0.00461312 0.0186733 0.00439916 0.00558293 0.00632667 0.223317 0.253067 58.0513 -87.8993 126.151 15.9337 145.037 0.000142335 0.267322 192.721 0.310177 0.0673231 0.00409859 0.000562403 0.00138517 0.986959 0.991716 -2.99066e-06 -85.6567 0.0930884 31168.2 310.593 0.983497 0.319146 0.738364 0.73836 9.99958 2.98664e-06 1.19464e-05 0.134419 0.983416 0.931331 -0.0132916 4.93158e-06 0.516667 -2.01808e-20 7.48772e-24 -2.01733e-20 0.0013965 0.997815 8.60256e-05 0.152737 2.85282 0.0013965 0.997815 0.792233 0.00106803 0.00188144 0.000860256 0.455379 0.00188144 0.44464 0.000131324 1.02 0.888801 0.534367 0.287605 1.71954e-07 3.08495e-09 2370.32 3139.8 -0.0582698 0.48221 0.277266 0.254829 -0.59306 -0.169576 0.48741 -0.265728 -0.221692 2.69 1 0 295.283 0 2.23888 2.688 0.000299082 0.867921 0.701572 0.314491 0.43489 2.23906 139.384 83.6342 18.7043 60.7283 0.00403712 0 -40 10
1.789 5.17488e-08 2.53998e-06 0.148326 0.148326 0.0120259 2.35222e-05 0.00115454 0.185408 0.00065883 0.186062 0.954378 101.423 0.23465 0.858778 4.57705 0.0653499 0.0431797 0.95682 0.0194165 0.00461358 0.0186727 0.00439956 0.0055835 0.00632725 0.22334 0.25309 58.0514 -87.8993 126.15 15.9337 145.037 0.000142338 0.267322 192.721 0.310177 0.0673231 0.00409859 0.000562403 0.00138517 0.986959 0.991716 -2.99067e-06 -85.6567 0.0930885 31168.2 310.605 0.983497 0.319146 0.738376 0.738372 9.99958 2.98664e-06 1.19465e-05 0.134424 0.983417 0.93133 -0.0132916 4.93161e-06 0.516687 -2.01824e-20 7.48836e-24 -2.01749e-20 0.0013965 0.997815 8.60257e-05 0.152737 2.85282 0.0013965 0.997815 0.792305 0.00106804 0.00188144 0.000860257 0.455379 0.00188144 0.444645 0.000131326 1.02 0.888802 0.534366 0.287606 1.71954e-07 3.08498e-09 2370.31 3139.85 -0.0582748 0.48221 0.277266 0.254832 -0.59306 -0.169576 0.487394 -0.265725 -0.221678 2.691 1 0 295.279 0 2.23902 2.689 0.00029908 0.86795 0.701615 0.314451 0.434912 2.2392 139.391 83.6336 18.7043 60.728 0.00403715 0 -40 10
1.79 5.17777e-08 2.53998e-06 0.148358 0.148358 0.0120259 2.35353e-05 0.00115454 0.185448 0.000658831 0.186102 0.954468 101.422 0.234639 0.858911 4.57769 0.0653607 0.0431858 0.956814 0.0194159 0.00461404 0.0186722 0.00439996 0.00558407 0.00632784 0.223363 0.253113 58.0515 -87.8993 126.15 15.9337 145.037 0.00014234 0.267322 192.721 0.310176 0.067323 0.0040986 0.000562404 0.00138517 0.986959 0.991716 -2.99069e-06 -85.6567 0.0930886 31168.2 310.618 0.983497 0.319146 0.738388 0.738384 9.99958 2.98665e-06 1.19465e-05 0.134429 0.983417 0.931329 -0.0132915 4.93164e-06 0.516707 -2.0184e-20 7.489e-24 -2.01765e-20 0.0013965 0.997815 8.60258e-05 0.152738 2.85282 0.0013965 0.997815 0.792377 0.00106806 0.00188145 0.000860258 0.455378 0.00188145 0.44465 0.000131329 1.02 0.888803 0.534366 0.287608 1.71955e-07 3.085e-09 2370.29 3139.9 -0.0582798 0.48221 0.277265 0.254835 -0.593059 -0.169576 0.487378 -0.265723 -0.221664 2.692 1 0 295.274 0 2.23915 2.69 0.000299079 0.867979 0.701658 0.314412 0.434934 2.23933 139.399 83.633 18.7042 60.7278 0.00403717 0 -40 10
1.791 5.18065e-08 2.53998e-06 0.14839 0.14839 0.0120259 2.35484e-05 0.00115454 0.185488 0.000658831 0.186142 0.954559 101.422 0.234628 0.859044 4.57833 0.0653715 0.0431918 0.956808 0.0194154 0.0046145 0.0186716 0.00440035 0.00558463 0.00632842 0.223385 0.253137 58.0515 -87.8993 126.15 15.9336 145.037 0.000142342 0.267323 192.721 0.310176 0.067323 0.0040986 0.000562405 0.00138518 0.986959 0.991716 -2.9907e-06 -85.6567 0.0930886 31168.1 310.63 0.983497 0.319146 0.7384 0.738396 9.99958 2.98665e-06 1.19465e-05 0.134433 0.983417 0.931328 -0.0132915 4.93167e-06 0.516727 -2.01856e-20 7.48964e-24 -2.01781e-20 0.0013965 0.997815 8.60259e-05 0.152738 2.85282 0.0013965 0.997815 0.792449 0.00106807 0.00188145 0.000860259 0.455378 0.00188145 0.444656 0.000131331 1.02 0.888804 0.534366 0.287609 1.71955e-07 3.08502e-09 2370.27 3139.95 -0.0582849 0.48221 0.277265 0.254839 -0.593058 -0.169576 0.487362 -0.265721 -0.22165 2.693 1 0 295.27 0 2.23929 2.691 0.000299078 0.868008 0.701701 0.314372 0.434956 2.23947 139.406 83.6325 18.7042 60.7275 0.0040372 0 -40 10
1.792 5.18354e-08 2.53999e-06 0.148422 0.148422 0.0120259 2.35615e-05 0.00115454 0.185528 0.000658832 0.186182 0.95465 101.421 0.234618 0.859177 4.57897 0.0653823 0.0431979 0.956802 0.0194148 0.00461496 0.018671 0.00440075 0.0055852 0.00632901 0.223408 0.25316 58.0516 -87.8993 126.15 15.9336 145.037 0.000142345 0.267323 192.721 0.310175 0.0673229 0.0040986 0.000562405 0.00138518 0.986959 0.991716 -2.99072e-06 -85.6567 0.0930887 31168.1 310.643 0.983497 0.319146 0.738412 0.738408 9.99958 2.98666e-06 1.19465e-05 0.134438 0.983417 0.931327 -0.0132915 4.9317e-06 0.516747 -2.01872e-20 7.49028e-24 -2.01798e-20 0.0013965 0.997815 8.6026e-05 0.152738 2.85282 0.0013965 0.997815 0.792521 0.00106809 0.00188145 0.00086026 0.455378 0.00188145 0.444661 0.000131333 1.02 0.888805 0.534365 0.287611 1.71955e-07 3.08504e-09 2370.26 3140 -0.0582899 0.48221 0.277265 0.254842 -0.593058 -0.169576 0.487346 -0.265719 -0.221636 2.694 1 0 295.265 0 2.23943 2.692 0.000299077 0.868037 0.701744 0.314332 0.434978 2.23961 139.413 83.6319 18.7042 60.7272 0.00403722 0 -40 10
1.793 5.18642e-08 2.53999e-06 0.148454 0.148454 0.0120259 2.35746e-05 0.00115454 0.185568 0.000658832 0.186222 0.95474 101.42 0.234607 0.85931 4.57962 0.0653931 0.0432039 0.956796 0.0194142 0.00461542 0.0186704 0.00440115 0.00558577 0.00632959 0.223431 0.253184 58.0517 -87.8993 126.149 15.9336 145.037 0.000142347 0.267323 192.72 0.310175 0.0673229 0.00409861 0.000562406 0.00138518 0.986959 0.991716 -2.99073e-06 -85.6567 0.0930888 31168.1 310.655 0.983497 0.319146 0.738424 0.73842 9.99958 2.98666e-06 1.19465e-05 0.134443 0.983418 0.931326 -0.0132915 4.93173e-06 0.516767 -2.01888e-20 7.49092e-24 -2.01814e-20 0.0013965 0.997815 8.6026e-05 0.152738 2.85282 0.0013965 0.997815 0.792593 0.00106811 0.00188145 0.00086026 0.455378 0.00188145 0.444666 0.000131336 1.02 0.888806 0.534365 0.287612 1.71956e-07 3.08507e-09 2370.24 3140.05 -0.058295 0.482211 0.277265 0.254845 -0.593057 -0.169576 0.48733 -0.265717 -0.221622 2.695 1 0 295.26 0 2.23956 2.693 0.000299075 0.868066 0.701786 0.314293 0.435 2.23974 139.421 83.6313 18.7041 60.7269 0.00403725 0 -40 10
1.794 5.1893e-08 2.53999e-06 0.148486 0.148486 0.0120259 2.35877e-05 0.00115454 0.185608 0.000658833 0.186262 0.954831 101.42 0.234596 0.859444 4.58026 0.0654039 0.04321 0.95679 0.0194137 0.00461588 0.0186698 0.00440155 0.00558634 0.00633018 0.223454 0.253207 58.0517 -87.8993 126.149 15.9335 145.037 0.000142349 0.267323 192.72 0.310174 0.0673228 0.00409861 0.000562407 0.00138518 0.986959 0.991716 -2.99075e-06 -85.6566 0.0930889 31168.1 310.668 0.983497 0.319146 0.738436 0.738432 9.99958 2.98667e-06 1.19466e-05 0.134447 0.983418 0.931325 -0.0132915 4.93176e-06 0.516787 -2.01905e-20 7.49156e-24 -2.0183e-20 0.0013965 0.997815 8.60261e-05 0.152738 2.85283 0.0013965 0.997815 0.792665 0.00106812 0.00188145 0.000860261 0.455377 0.00188145 0.444671 0.000131338 1.02 0.888807 0.534365 0.287614 1.71956e-07 3.08509e-09 2370.22 3140.1 -0.0583 0.482211 0.277264 0.254848 -0.593056 -0.169576 0.487314 -0.265715 -0.221608 2.696 1 0 295.256 0 2.2397 2.694 0.000299074 0.868094 0.701829 0.314253 0.435023 2.23988 139.428 83.6307 18.7041 60.7266 0.00403727 0 -40 10
1.795 5.19219e-08 2.53999e-06 0.148518 0.148518 0.0120259 2.36009e-05 0.00115454 0.185648 0.000658833 0.186302 0.954921 101.419 0.234585 0.859577 4.5809 0.0654147 0.043216 0.956784 0.0194131 0.00461634 0.0186692 0.00440195 0.00558691 0.00633076 0.223476 0.253231 58.0518 -87.8993 126.149 15.9335 145.037 0.000142351 0.267323 192.72 0.310174 0.0673228 0.00409861 0.000562407 0.00138519 0.986959 0.991716 -2.99076e-06 -85.6566 0.093089 31168.1 310.68 0.983497 0.319146 0.738448 0.738444 9.99958 2.98667e-06 1.19466e-05 0.134452 0.983418 0.931324 -0.0132915 4.93179e-06 0.516807 -2.01921e-20 7.4922e-24 -2.01846e-20 0.0013965 0.997815 8.60262e-05 0.152738 2.85283 0.0013965 0.997815 0.792737 0.00106814 0.00188145 0.000860262 0.455377 0.00188145 0.444676 0.00013134 1.02 0.888808 0.534364 0.287616 1.71956e-07 3.08511e-09 2370.21 3140.15 -0.0583051 0.482211 0.277264 0.254851 -0.593056 -0.169576 0.487298 -0.265713 -0.221594 2.697 1 0 295.251 0 2.23984 2.695 0.000299073 0.868123 0.701872 0.314214 0.435045 2.24002 139.435 83.6301 18.7041 60.7263 0.0040373 0 -40 10
1.796 5.19507e-08 2.53999e-06 0.14855 0.14855 0.0120258 2.3614e-05 0.00115454 0.185688 0.000658834 0.186342 0.955012 101.418 0.234575 0.85971 4.58154 0.0654255 0.0432221 0.956778 0.0194125 0.0046168 0.0186686 0.00440235 0.00558748 0.00633135 0.223499 0.253254 58.0518 -87.8993 126.149 15.9334 145.037 0.000142354 0.267323 192.72 0.310174 0.0673227 0.00409862 0.000562408 0.00138519 0.986958 0.991716 -2.99078e-06 -85.6566 0.0930891 31168 310.693 0.983497 0.319146 0.73846 0.738456 9.99958 2.98668e-06 1.19466e-05 0.134457 0.983418 0.931323 -0.0132915 4.93182e-06 0.516827 -2.01937e-20 7.49285e-24 -2.01862e-20 0.00139651 0.997815 8.60263e-05 0.152739 2.85283 0.00139651 0.997815 0.792809 0.00106815 0.00188146 0.000860263 0.455377 0.00188145 0.444681 0.000131343 1.02 0.88881 0.534364 0.287617 1.71956e-07 3.08514e-09 2370.19 3140.2 -0.0583101 0.482211 0.277264 0.254855 -0.593055 -0.169576 0.487282 -0.265711 -0.22158 2.698 1 0 295.247 0 2.23997 2.696 0.000299072 0.868152 0.701915 0.314174 0.435067 2.24015 139.443 83.6295 18.704 60.7261 0.00403732 0 -40 10
1.797 5.19796e-08 2.53999e-06 0.148582 0.148582 0.0120258 2.36271e-05 0.00115454 0.185728 0.000658834 0.186382 0.955103 101.418 0.234564 0.859843 4.58219 0.0654363 0.0432282 0.956772 0.019412 0.00461727 0.0186681 0.00440275 0.00558805 0.00633194 0.223522 0.253278 58.0519 -87.8993 126.149 15.9334 145.037 0.000142356 0.267324 192.72 0.310173 0.0673227 0.00409862 0.000562409 0.00138519 0.986958 0.991716 -2.99079e-06 -85.6566 0.0930892 31168 310.705 0.983497 0.319146 0.738472 0.738468 9.99958 2.98668e-06 1.19466e-05 0.134461 0.983419 0.931322 -0.0132915 4.93185e-06 0.516847 -2.01953e-20 7.49349e-24 -2.01878e-20 0.00139651 0.997815 8.60264e-05 0.152739 2.85283 0.00139651 0.997815 0.792881 0.00106817 0.00188146 0.000860264 0.455377 0.00188146 0.444686 0.000131345 1.02 0.888811 0.534364 0.287619 1.71957e-07 3.08516e-09 2370.18 3140.25 -0.0583152 0.482211 0.277263 0.254858 -0.593055 -0.169576 0.487266 -0.265709 -0.221566 2.699 1 0 295.242 0 2.24011 2.697 0.00029907 0.868181 0.701958 0.314135 0.435089 2.24029 139.45 83.6289 18.704 60.7258 0.00403734 0 -40 10
1.798 5.20084e-08 2.54e-06 0.148614 0.148614 0.0120258 2.36402e-05 0.00115454 0.185768 0.000658835 0.186422 0.955193 101.417 0.234553 0.859976 4.58283 0.0654471 0.0432342 0.956766 0.0194114 0.00461773 0.0186675 0.00440315 0.00558862 0.00633252 0.223545 0.253301 58.052 -87.8993 126.148 15.9334 145.037 0.000142358 0.267324 192.72 0.310173 0.0673226 0.00409862 0.000562409 0.00138519 0.986958 0.991716 -2.99081e-06 -85.6566 0.0930893 31168 310.718 0.983497 0.319146 0.738484 0.73848 9.99958 2.98669e-06 1.19466e-05 0.134466 0.983419 0.931321 -0.0132915 4.93188e-06 0.516867 -2.01969e-20 7.49413e-24 -2.01894e-20 0.00139651 0.997815 8.60264e-05 0.152739 2.85283 0.00139651 0.997815 0.792953 0.00106819 0.00188146 0.000860264 0.455377 0.00188146 0.444691 0.000131348 1.02 0.888812 0.534364 0.28762 1.71957e-07 3.08518e-09 2370.16 3140.3 -0.0583202 0.482211 0.277263 0.254861 -0.593054 -0.169576 0.48725 -0.265707 -0.221552 2.7 1 0 295.238 0 2.24025 2.698 0.000299069 0.86821 0.702001 0.314095 0.435111 2.24043 139.457 83.6283 18.704 60.7255 0.00403737 0 -40 10
1.799 5.20372e-08 2.54e-06 0.148646 0.148646 0.0120258 2.36533e-05 0.00115454 0.185808 0.000658835 0.186462 0.955284 101.417 0.234542 0.86011 4.58347 0.0654579 0.0432403 0.95676 0.0194108 0.00461819 0.0186669 0.00440355 0.00558919 0.00633311 0.223567 0.253324 58.052 -87.8993 126.148 15.9333 145.037 0.000142361 0.267324 192.719 0.310172 0.0673226 0.00409863 0.00056241 0.00138519 0.986958 0.991715 -2.99082e-06 -85.6566 0.0930893 31168 310.73 0.983497 0.319146 0.738496 0.738492 9.99958 2.98669e-06 1.19467e-05 0.134471 0.983419 0.93132 -0.0132915 4.93191e-06 0.516887 -2.01985e-20 7.49477e-24 -2.0191e-20 0.00139651 0.997815 8.60265e-05 0.152739 2.85283 0.00139651 0.997815 0.793024 0.0010682 0.00188146 0.000860265 0.455376 0.00188146 0.444696 0.00013135 1.02 0.888813 0.534363 0.287622 1.71957e-07 3.0852e-09 2370.14 3140.35 -0.0583252 0.482211 0.277263 0.254864 -0.593053 -0.169576 0.487234 -0.265705 -0.221538 2.701 1 0 295.233 0 2.24038 2.699 0.000299068 0.868239 0.702043 0.314056 0.435133 2.24056 139.465 83.6277 18.7039 60.7252 0.00403739 0 -40 10
1.8 5.20661e-08 2.54e-06 0.148678 0.148677 0.0120258 2.36664e-05 0.00115455 0.185847 0.000658836 0.186502 0.955375 101.416 0.234531 0.860243 4.58412 0.0654687 0.0432464 0.956754 0.0194102 0.00461865 0.0186663 0.00440395 0.00558976 0.0063337 0.22359 0.253348 58.0521 -87.8993 126.148 15.9333 145.037 0.000142363 0.267324 192.719 0.310172 0.0673225 0.00409863 0.000562411 0.0013852 0.986958 0.991715 -2.99084e-06 -85.6566 0.0930894 31167.9 310.743 0.983497 0.319146 0.738508 0.738504 9.99958 2.9867e-06 1.19467e-05 0.134475 0.983419 0.931319 -0.0132915 4.93194e-06 0.516908 -2.02001e-20 7.49542e-24 -2.01926e-20 0.00139651 0.997815 8.60266e-05 0.152739 2.85283 0.00139651 0.997815 0.793096 0.00106822 0.00188146 0.000860266 0.455376 0.00188146 0.444701 0.000131352 1.02 0.888814 0.534363 0.287623 1.71957e-07 3.08523e-09 2370.13 3140.4 -0.0583303 0.482211 0.277263 0.254868 -0.593053 -0.169576 0.487217 -0.265702 -0.221524 2.702 1 0 295.229 0 2.24052 2.7 0.000299067 0.868268 0.702086 0.314016 0.435155 2.2407 139.472 83.6272 18.7039 60.7249 0.00403742 0 -40 10
1.801 5.20949e-08 2.54e-06 0.14871 0.148709 0.0120258 2.36795e-05 0.00115455 0.185887 0.000658836 0.186541 0.955466 101.415 0.23452 0.860376 4.58476 0.0654795 0.0432525 0.956748 0.0194097 0.00461912 0.0186657 0.00440435 0.00559033 0.00633429 0.223613 0.253372 58.0522 -87.8993 126.148 15.9333 145.037 0.000142365 0.267324 192.719 0.310171 0.0673225 0.00409863 0.000562411 0.0013852 0.986958 0.991715 -2.99085e-06 -85.6566 0.0930895 31167.9 310.756 0.983497 0.319146 0.73852 0.738516 9.99958 2.9867e-06 1.19467e-05 0.13448 0.98342 0.931318 -0.0132915 4.93197e-06 0.516928 -2.02017e-20 7.49606e-24 -2.01942e-20 0.00139651 0.997815 8.60267e-05 0.152739 2.85283 0.00139651 0.997815 0.793168 0.00106823 0.00188146 0.000860267 0.455376 0.00188146 0.444706 0.000131355 1.02 0.888815 0.534363 0.287625 1.71958e-07 3.08525e-09 2370.11 3140.45 -0.0583353 0.482211 0.277262 0.254871 -0.593052 -0.169576 0.487201 -0.2657 -0.221511 2.703 1 0 295.224 0 2.24066 2.701 0.000299065 0.868297 0.702129 0.313977 0.435177 2.24084 139.479 83.6266 18.7038 60.7246 0.00403744 0 -40 10
1.802 5.21237e-08 2.54e-06 0.148741 0.148741 0.0120258 2.36926e-05 0.00115455 0.185927 0.000658837 0.186581 0.955556 101.415 0.23451 0.860509 4.58541 0.0654903 0.0432586 0.956741 0.0194091 0.00461958 0.0186651 0.00440475 0.0055909 0.00633488 0.223636 0.253395 58.0522 -87.8993 126.147 15.9332 145.037 0.000142368 0.267325 192.719 0.310171 0.0673224 0.00409863 0.000562412 0.0013852 0.986958 0.991715 -2.99087e-06 -85.6566 0.0930896 31167.9 310.768 0.983497 0.319146 0.738532 0.738528 9.99958 2.98671e-06 1.19467e-05 0.134485 0.98342 0.931317 -0.0132915 4.932e-06 0.516948 -2.02033e-20 7.4967e-24 -2.01958e-20 0.00139651 0.997815 8.60268e-05 0.152739 2.85283 0.00139651 0.997815 0.79324 0.00106825 0.00188146 0.000860268 0.455376 0.00188146 0.444712 0.000131357 1.02 0.888816 0.534362 0.287626 1.71958e-07 3.08527e-09 2370.09 3140.5 -0.0583404 0.482211 0.277262 0.254874 -0.593051 -0.169576 0.487185 -0.265698 -0.221497 2.704 1 0 295.219 0 2.24079 2.702 0.000299064 0.868325 0.702172 0.313938 0.435199 2.24097 139.487 83.626 18.7038 60.7243 0.00403747 0 -40 10
1.803 5.21526e-08 2.54e-06 0.148773 0.148773 0.0120257 2.37057e-05 0.00115455 0.185967 0.000658837 0.186621 0.955647 101.414 0.234499 0.860643 4.58606 0.0655011 0.0432647 0.956735 0.0194085 0.00462004 0.0186645 0.00440515 0.00559147 0.00633546 0.223659 0.253419 58.0523 -87.8993 126.147 15.9332 145.037 0.00014237 0.267325 192.719 0.310171 0.0673223 0.00409864 0.000562413 0.0013852 0.986958 0.991715 -2.99088e-06 -85.6566 0.0930897 31167.9 310.781 0.983497 0.319146 0.738544 0.73854 9.99958 2.98671e-06 1.19467e-05 0.13449 0.98342 0.931316 -0.0132915 4.93202e-06 0.516968 -2.02049e-20 7.49735e-24 -2.01974e-20 0.00139651 0.997815 8.60268e-05 0.15274 2.85283 0.00139651 0.997815 0.793311 0.00106827 0.00188147 0.000860268 0.455375 0.00188146 0.444717 0.000131359 1.02 0.888817 0.534362 0.287628 1.71958e-07 3.0853e-09 2370.08 3140.55 -0.0583455 0.482211 0.277262 0.254877 -0.593051 -0.169576 0.487169 -0.265696 -0.221483 2.705 1 0 295.215 0 2.24093 2.703 0.000299063 0.868354 0.702215 0.313898 0.435221 2.24111 139.494 83.6254 18.7038 60.7241 0.00403749 0 -40 10
1.804 5.21814e-08 2.54001e-06 0.148805 0.148805 0.0120257 2.37188e-05 0.00115455 0.186006 0.000658838 0.18666 0.955738 101.413 0.234488 0.860776 4.5867 0.0655119 0.0432708 0.956729 0.019408 0.00462051 0.0186639 0.00440555 0.00559204 0.00633605 0.223682 0.253442 58.0523 -87.8993 126.147 15.9331 145.037 0.000142372 0.267325 192.719 0.31017 0.0673223 0.00409864 0.000562413 0.00138521 0.986958 0.991715 -2.9909e-06 -85.6566 0.0930898 31167.9 310.793 0.983496 0.319146 0.738556 0.738552 9.99958 2.98672e-06 1.19468e-05 0.134494 0.98342 0.931315 -0.0132915 4.93205e-06 0.516988 -2.02065e-20 7.49799e-24 -2.0199e-20 0.00139652 0.997815 8.60269e-05 0.15274 2.85283 0.00139652 0.997815 0.793383 0.00106828 0.00188147 0.000860269 0.455375 0.00188147 0.444722 0.000131362 1.02 0.888818 0.534362 0.287629 1.71959e-07 3.08532e-09 2370.06 3140.6 -0.0583505 0.482211 0.277261 0.25488 -0.59305 -0.169577 0.487153 -0.265694 -0.221469 2.706 1 0 295.21 0 2.24107 2.704 0.000299062 0.868383 0.702257 0.313859 0.435243 2.24125 139.501 83.6248 18.7037 60.7238 0.00403751 0 -40 10
1.805 5.22103e-08 2.54001e-06 0.148837 0.148836 0.0120257 2.37319e-05 0.00115455 0.186046 0.000658838 0.1867 0.955829 101.413 0.234477 0.860909 4.58735 0.0655227 0.0432769 0.956723 0.0194074 0.00462097 0.0186634 0.00440595 0.00559261 0.00633664 0.223704 0.253466 58.0524 -87.8993 126.147 15.9331 145.037 0.000142375 0.267325 192.718 0.31017 0.0673222 0.00409864 0.000562414 0.00138521 0.986958 0.991715 -2.99091e-06 -85.6565 0.0930899 31167.8 310.806 0.983496 0.319146 0.738568 0.738564 9.99958 2.98672e-06 1.19468e-05 0.134499 0.983421 0.931314 -0.0132915 4.93208e-06 0.517008 -2.02081e-20 7.49863e-24 -2.02006e-20 0.00139652 0.997815 8.6027e-05 0.15274 2.85284 0.00139652 0.997815 0.793455 0.0010683 0.00188147 0.00086027 0.455375 0.00188147 0.444727 0.000131364 1.02 0.888819 0.534361 0.287631 1.71959e-07 3.08534e-09 2370.04 3140.66 -0.0583556 0.482211 0.277261 0.254884 -0.593049 -0.169577 0.487137 -0.265692 -0.221455 2.707 1 0 295.206 0 2.2412 2.705 0.00029906 0.868412 0.7023 0.31382 0.435266 2.24138 139.509 83.6242 18.7037 60.7235 0.00403754 0 -40 10
1.806 5.22391e-08 2.54001e-06 0.148868 0.148868 0.0120257 2.3745e-05 0.00115455 0.186086 0.000658838 0.18674 0.955919 101.412 0.234466 0.861042 4.588 0.0655335 0.043283 0.956717 0.0194068 0.00462143 0.0186628 0.00440635 0.00559318 0.00633723 0.223727 0.253489 58.0525 -87.8993 126.147 15.9331 145.037 0.000142377 0.267325 192.718 0.310169 0.0673222 0.00409865 0.000562415 0.00138521 0.986958 0.991715 -2.99093e-06 -85.6565 0.09309 31167.8 310.819 0.983496 0.319146 0.73858 0.738576 9.99958 2.98673e-06 1.19468e-05 0.134504 0.983421 0.931313 -0.0132915 4.93211e-06 0.517028 -2.02098e-20 7.49928e-24 -2.02023e-20 0.00139652 0.997815 8.60271e-05 0.15274 2.85284 0.00139652 0.997815 0.793526 0.00106832 0.00188147 0.000860271 0.455375 0.00188147 0.444732 0.000131367 1.02 0.888821 0.534361 0.287632 1.71959e-07 3.08537e-09 2370.03 3140.71 -0.0583606 0.482212 0.277261 0.254887 -0.593049 -0.169577 0.487121 -0.26569 -0.221441 2.708 1 0 295.201 0 2.24134 2.706 0.000299059 0.868441 0.702343 0.31378 0.435288 2.24152 139.516 83.6236 18.7037 60.7232 0.00403756 0 -40 10
1.807 5.22679e-08 2.54001e-06 0.1489 0.1489 0.0120257 2.37582e-05 0.00115455 0.186125 0.000658839 0.186779 0.95601 101.411 0.234456 0.861176 4.58864 0.0655444 0.0432891 0.956711 0.0194062 0.0046219 0.0186622 0.00440676 0.00559375 0.00633782 0.22375 0.253513 58.0525 -87.8993 126.146 15.933 145.037 0.000142379 0.267326 192.718 0.310169 0.0673221 0.00409865 0.000562415 0.00138521 0.986958 0.991715 -2.99094e-06 -85.6565 0.09309 31167.8 310.831 0.983496 0.319146 0.738592 0.738588 9.99958 2.98673e-06 1.19468e-05 0.134508 0.983421 0.931312 -0.0132915 4.93214e-06 0.517049 -2.02114e-20 7.49992e-24 -2.02039e-20 0.00139652 0.997815 8.60272e-05 0.15274 2.85284 0.00139652 0.997815 0.793598 0.00106833 0.00188147 0.000860272 0.455375 0.00188147 0.444737 0.000131369 1.02 0.888822 0.534361 0.287634 1.71959e-07 3.08539e-09 2370.01 3140.76 -0.0583657 0.482212 0.277261 0.25489 -0.593048 -0.169577 0.487105 -0.265688 -0.221427 2.709 1 0 295.197 0 2.24148 2.707 0.000299058 0.86847 0.702386 0.313741 0.43531 2.24166 139.523 83.623 18.7036 60.7229 0.00403759 0 -40 10
1.808 5.22968e-08 2.54001e-06 0.148932 0.148931 0.0120257 2.37713e-05 0.00115455 0.186165 0.000658839 0.186819 0.956101 101.411 0.234445 0.861309 4.58929 0.0655552 0.0432952 0.956705 0.0194057 0.00462236 0.0186616 0.00440716 0.00559432 0.00633841 0.223773 0.253536 58.0526 -87.8993 126.146 15.933 145.037 0.000142382 0.267326 192.718 0.310168 0.0673221 0.00409865 0.000562416 0.00138521 0.986958 0.991715 -2.99096e-06 -85.6565 0.0930901 31167.8 310.844 0.983496 0.319146 0.738604 0.7386 9.99958 2.98674e-06 1.19468e-05 0.134513 0.983421 0.931311 -0.0132915 4.93217e-06 0.517069 -2.0213e-20 7.50057e-24 -2.02055e-20 0.00139652 0.997815 8.60272e-05 0.15274 2.85284 0.00139652 0.997815 0.793669 0.00106835 0.00188147 0.000860272 0.455374 0.00188147 0.444742 0.000131371 1.02 0.888823 0.53436 0.287635 1.7196e-07 3.08541e-09 2370 3140.81 -0.0583707 0.482212 0.27726 0.254893 -0.593048 -0.169577 0.487089 -0.265686 -0.221413 2.71 1 0 295.192 0 2.24161 2.708 0.000299057 0.868499 0.702428 0.313702 0.435332 2.24179 139.531 83.6224 18.7036 60.7226 0.00403761 0 -40 10
1.809 5.23256e-08 2.54001e-06 0.148963 0.148963 0.0120257 2.37844e-05 0.00115455 0.186204 0.00065884 0.186858 0.956192 101.41 0.234434 0.861442 4.58994 0.065566 0.0433013 0.956699 0.0194051 0.00462282 0.018661 0.00440756 0.0055949 0.006339 0.223796 0.25356 58.0527 -87.8994 126.146 15.933 145.037 0.000142384 0.267326 192.718 0.310168 0.067322 0.00409866 0.000562417 0.00138522 0.986958 0.991715 -2.99097e-06 -85.6565 0.0930902 31167.7 310.856 0.983496 0.319146 0.738616 0.738612 9.99958 2.98674e-06 1.19469e-05 0.134518 0.983422 0.93131 -0.0132915 4.9322e-06 0.517089 -2.02146e-20 7.50121e-24 -2.02071e-20 0.00139652 0.997815 8.60273e-05 0.152741 2.85284 0.00139652 0.997815 0.793741 0.00106836 0.00188147 0.000860273 0.455374 0.00188147 0.444747 0.000131374 1.02 0.888824 0.53436 0.287637 1.7196e-07 3.08543e-09 2369.98 3140.86 -0.0583758 0.482212 0.27726 0.254897 -0.593047 -0.169577 0.487073 -0.265684 -0.221399 2.711 1 0 295.188 0 2.24175 2.709 0.000299055 0.868528 0.702471 0.313663 0.435354 2.24193 139.538 83.6218 18.7036 60.7224 0.00403764 0 -40 10
1.81 5.23545e-08 2.54002e-06 0.148995 0.148994 0.0120256 2.37975e-05 0.00115455 0.186244 0.00065884 0.186898 0.956283 101.409 0.234423 0.861576 4.59059 0.0655768 0.0433075 0.956693 0.0194045 0.00462329 0.0186604 0.00440796 0.00559547 0.00633959 0.223819 0.253584 58.0527 -87.8994 126.146 15.9329 145.037 0.000142386 0.267326 192.718 0.310168 0.067322 0.00409866 0.000562417 0.00138522 0.986958 0.991715 -2.99099e-06 -85.6565 0.0930903 31167.7 310.869 0.983496 0.319146 0.738628 0.738624 9.99958 2.98674e-06 1.19469e-05 0.134523 0.983422 0.931309 -0.0132915 4.93223e-06 0.517109 -2.02162e-20 7.50186e-24 -2.02087e-20 0.00139652 0.997815 8.60274e-05 0.152741 2.85284 0.00139652 0.997815 0.793812 0.00106838 0.00188148 0.000860274 0.455374 0.00188147 0.444752 0.000131376 1.02 0.888825 0.53436 0.287638 1.7196e-07 3.08546e-09 2369.96 3140.91 -0.0583808 0.482212 0.27726 0.2549 -0.593046 -0.169577 0.487057 -0.265681 -0.221385 2.712 1 0 295.183 0 2.24189 2.71 0.000299054 0.868557 0.702514 0.313624 0.435376 2.24207 139.545 83.6212 18.7035 60.7221 0.00403766 0 -40 10
1.811 5.23833e-08 2.54002e-06 0.149027 0.149026 0.0120256 2.38106e-05 0.00115455 0.186283 0.000658841 0.186937 0.956374 101.409 0.234412 0.861709 4.59124 0.0655876 0.0433136 0.956686 0.019404 0.00462375 0.0186598 0.00440836 0.00559604 0.00634018 0.223842 0.253607 58.0528 -87.8994 126.146 15.9329 145.037 0.000142388 0.267326 192.717 0.310167 0.0673219 0.00409866 0.000562418 0.00138522 0.986958 0.991715 -2.991e-06 -85.6565 0.0930904 31167.7 310.882 0.983496 0.319146 0.73864 0.738636 9.99958 2.98675e-06 1.19469e-05 0.134527 0.983422 0.931308 -0.0132915 4.93226e-06 0.51713 -2.02178e-20 7.5025e-24 -2.02103e-20 0.00139652 0.997815 8.60275e-05 0.152741 2.85284 0.00139652 0.997815 0.793884 0.0010684 0.00188148 0.000860275 0.455374 0.00188148 0.444757 0.000131378 1.02 0.888826 0.53436 0.28764 1.7196e-07 3.08548e-09 2369.95 3140.96 -0.0583859 0.482212 0.277259 0.254903 -0.593046 -0.169577 0.487041 -0.265679 -0.221371 2.713 1 0 295.178 0 2.24202 2.711 0.000299053 0.868586 0.702557 0.313585 0.435398 2.2422 139.553 83.6207 18.7035 60.7218 0.00403769 0 -40 10
1.812 5.24121e-08 2.54002e-06 0.149058 0.149058 0.0120256 2.38237e-05 0.00115455 0.186323 0.000658841 0.186977 0.956465 101.408 0.234402 0.861843 4.59189 0.0655984 0.0433197 0.95668 0.0194034 0.00462422 0.0186592 0.00440877 0.00559662 0.00634077 0.223865 0.253631 58.0528 -87.8994 126.145 15.9328 145.037 0.000142391 0.267327 192.717 0.310167 0.0673219 0.00409866 0.000562419 0.00138522 0.986958 0.991715 -2.99102e-06 -85.6565 0.0930905 31167.7 310.894 0.983496 0.319146 0.738652 0.738648 9.99958 2.98675e-06 1.19469e-05 0.134532 0.983422 0.931307 -0.0132915 4.93229e-06 0.51715 -2.02195e-20 7.50315e-24 -2.0212e-20 0.00139652 0.997815 8.60276e-05 0.152741 2.85284 0.00139652 0.997815 0.793955 0.00106841 0.00188148 0.000860276 0.455373 0.00188148 0.444762 0.000131381 1.02 0.888827 0.534359 0.287641 1.71961e-07 3.0855e-09 2369.93 3141.01 -0.058391 0.482212 0.277259 0.254906 -0.593045 -0.169577 0.487025 -0.265677 -0.221357 2.714 1 0 295.174 0 2.24216 2.712 0.000299052 0.868615 0.7026 0.313545 0.43542 2.24234 139.56 83.6201 18.7035 60.7215 0.00403771 0 -40 10
1.813 5.2441e-08 2.54002e-06 0.14909 0.149089 0.0120256 2.38368e-05 0.00115456 0.186362 0.000658842 0.187016 0.956555 101.407 0.234391 0.861976 4.59254 0.0656093 0.0433259 0.956674 0.0194028 0.00462468 0.0186586 0.00440917 0.00559719 0.00634136 0.223888 0.253655 58.0529 -87.8994 126.145 15.9328 145.037 0.000142393 0.267327 192.717 0.310166 0.0673218 0.00409867 0.000562419 0.00138522 0.986958 0.991715 -2.99103e-06 -85.6565 0.0930906 31167.7 310.907 0.983496 0.319146 0.738664 0.73866 9.99958 2.98676e-06 1.19469e-05 0.134537 0.983422 0.931306 -0.0132915 4.93232e-06 0.51717 -2.02211e-20 7.5038e-24 -2.02136e-20 0.00139653 0.997815 8.60276e-05 0.152741 2.85284 0.00139653 0.997815 0.794027 0.00106843 0.00188148 0.000860276 0.455373 0.00188148 0.444767 0.000131383 1.02 0.888828 0.534359 0.287643 1.71961e-07 3.08553e-09 2369.91 3141.06 -0.058396 0.482212 0.277259 0.254909 -0.593044 -0.169577 0.487009 -0.265675 -0.221343 2.715 1 0 295.169 0 2.2423 2.713 0.00029905 0.868644 0.702642 0.313506 0.435442 2.24248 139.567 83.6195 18.7034 60.7212 0.00403774 0 -40 10
1.814 5.24698e-08 2.54002e-06 0.149121 0.149121 0.0120256 2.38499e-05 0.00115456 0.186401 0.000658842 0.187056 0.956646 101.407 0.23438 0.862109 4.59319 0.0656201 0.043332 0.956668 0.0194022 0.00462515 0.018658 0.00440957 0.00559776 0.00634196 0.22391 0.253678 58.053 -87.8994 126.145 15.9328 145.037 0.000142395 0.267327 192.717 0.310166 0.0673218 0.00409867 0.00056242 0.00138523 0.986958 0.991715 -2.99105e-06 -85.6565 0.0930907 31167.6 310.92 0.983496 0.319146 0.738676 0.738672 9.99958 2.98676e-06 1.1947e-05 0.134542 0.983423 0.931305 -0.0132915 4.93235e-06 0.51719 -2.02227e-20 7.50444e-24 -2.02152e-20 0.00139653 0.997815 8.60277e-05 0.152741 2.85284 0.00139653 0.997815 0.794098 0.00106844 0.00188148 0.000860277 0.455373 0.00188148 0.444772 0.000131385 1.02 0.888829 0.534359 0.287644 1.71961e-07 3.08555e-09 2369.9 3141.11 -0.0584011 0.482212 0.277259 0.254913 -0.593044 -0.169577 0.486993 -0.265673 -0.221329 2.716 1 0 295.165 0 2.24243 2.714 0.000299049 0.868673 0.702685 0.313467 0.435464 2.24261 139.575 83.6189 18.7034 60.7209 0.00403776 0 -40 10
1.815 5.24986e-08 2.54002e-06 0.149153 0.149152 0.0120256 2.3863e-05 0.00115456 0.186441 0.000658843 0.187095 0.956737 101.406 0.234369 0.862243 4.59384 0.0656309 0.0433381 0.956662 0.0194017 0.00462561 0.0186575 0.00440997 0.00559834 0.00634255 0.223933 0.253702 58.053 -87.8994 126.145 15.9327 145.037 0.000142398 0.267327 192.717 0.310165 0.0673217 0.00409867 0.000562421 0.00138523 0.986958 0.991715 -2.99106e-06 -85.6565 0.0930907 31167.6 310.932 0.983496 0.319146 0.738688 0.738684 9.99958 2.98677e-06 1.1947e-05 0.134546 0.983423 0.931304 -0.0132915 4.93238e-06 0.517211 -2.02243e-20 7.50509e-24 -2.02168e-20 0.00139653 0.997815 8.60278e-05 0.152741 2.85284 0.00139653 0.997815 0.79417 0.00106846 0.00188148 0.000860278 0.455373 0.00188148 0.444777 0.000131388 1.02 0.88883 0.534358 0.287646 1.71962e-07 3.08557e-09 2369.88 3141.16 -0.0584061 0.482212 0.277258 0.254916 -0.593043 -0.169577 0.486976 -0.265671 -0.221315 2.717 1 0 295.16 0 2.24257 2.715 0.000299048 0.868702 0.702728 0.313428 0.435486 2.24275 139.582 83.6183 18.7034 60.7206 0.00403778 0 -40 10
1.816 5.25275e-08 2.54003e-06 0.149184 0.149183 0.0120256 2.38761e-05 0.00115456 0.18648 0.000658843 0.187134 0.956828 101.406 0.234358 0.862376 4.5945 0.0656417 0.0433443 0.956656 0.0194011 0.00462608 0.0186569 0.00441038 0.00559891 0.00634314 0.223956 0.253726 58.0531 -87.8994 126.144 15.9327 145.037 0.0001424 0.267327 192.717 0.310165 0.0673217 0.00409868 0.000562421 0.00138523 0.986958 0.991715 -2.99108e-06 -85.6564 0.0930908 31167.6 310.945 0.983496 0.319146 0.7387 0.738696 9.99958 2.98677e-06 1.1947e-05 0.134551 0.983423 0.931303 -0.0132915 4.93241e-06 0.517231 -2.02259e-20 7.50574e-24 -2.02184e-20 0.00139653 0.997815 8.60279e-05 0.152742 2.85285 0.00139653 0.997815 0.794241 0.00106848 0.00188149 0.000860279 0.455372 0.00188148 0.444782 0.00013139 1.02 0.888831 0.534358 0.287647 1.71962e-07 3.08559e-09 2369.87 3141.21 -0.0584112 0.482212 0.277258 0.254919 -0.593042 -0.169577 0.48696 -0.265669 -0.221301 2.718 1 0 295.156 0 2.24271 2.716 0.000299047 0.868731 0.702771 0.313389 0.435508 2.24289 139.589 83.6177 18.7033 60.7204 0.00403781 0 -40 10
1.817 5.25563e-08 2.54003e-06 0.149215 0.149215 0.0120256 2.38892e-05 0.00115456 0.186519 0.000658844 0.187173 0.956919 101.405 0.234347 0.86251 4.59515 0.0656526 0.0433505 0.95665 0.0194005 0.00462654 0.0186563 0.00441078 0.00559948 0.00634373 0.223979 0.253749 58.0532 -87.8994 126.144 15.9327 145.037 0.000142402 0.267327 192.716 0.310165 0.0673216 0.00409868 0.000562422 0.00138523 0.986958 0.991715 -2.99109e-06 -85.6564 0.0930909 31167.6 310.958 0.983496 0.319146 0.738712 0.738708 9.99958 2.98678e-06 1.1947e-05 0.134556 0.983423 0.931302 -0.0132915 4.93244e-06 0.517251 -2.02276e-20 7.50638e-24 -2.022e-20 0.00139653 0.997815 8.6028e-05 0.152742 2.85285 0.00139653 0.997815 0.794312 0.00106849 0.00188149 0.00086028 0.455372 0.00188149 0.444787 0.000131393 1.02 0.888833 0.534358 0.287649 1.71962e-07 3.08562e-09 2369.85 3141.26 -0.0584163 0.482212 0.277258 0.254922 -0.593042 -0.169577 0.486944 -0.265667 -0.221287 2.719 1 0 295.151 0 2.24284 2.717 0.000299045 0.86876 0.702813 0.313351 0.43553 2.24302 139.597 83.6171 18.7033 60.7201 0.00403783 0 -40 10
1.818 5.25852e-08 2.54003e-06 0.149247 0.149246 0.0120255 2.39023e-05 0.00115456 0.186558 0.000658844 0.187213 0.95701 101.404 0.234337 0.862643 4.5958 0.0656634 0.0433566 0.956643 0.0193999 0.00462701 0.0186557 0.00441118 0.00560006 0.00634432 0.224002 0.253773 58.0532 -87.8994 126.144 15.9326 145.037 0.000142405 0.267328 192.716 0.310164 0.0673216 0.00409868 0.000562423 0.00138524 0.986958 0.991715 -2.99111e-06 -85.6564 0.093091 31167.5 310.97 0.983496 0.319146 0.738725 0.73872 9.99958 2.98678e-06 1.1947e-05 0.134561 0.983424 0.931301 -0.0132915 4.93247e-06 0.517271 -2.02292e-20 7.50703e-24 -2.02217e-20 0.00139653 0.997815 8.6028e-05 0.152742 2.85285 0.00139653 0.997815 0.794384 0.00106851 0.00188149 0.00086028 0.455372 0.00188149 0.444793 0.000131395 1.02 0.888834 0.534357 0.28765 1.71962e-07 3.08564e-09 2369.83 3141.31 -0.0584213 0.482212 0.277258 0.254926 -0.593041 -0.169577 0.486928 -0.265665 -0.221273 2.72 1 0 295.146 0 2.24298 2.718 0.000299044 0.86879 0.702856 0.313312 0.435552 2.24316 139.604 83.6165 18.7033 60.7198 0.00403786 0 -40 10
1.819 5.2614e-08 2.54003e-06 0.149278 0.149278 0.0120255 2.39155e-05 0.00115456 0.186598 0.000658845 0.187252 0.957101 101.404 0.234326 0.862777 4.59645 0.0656742 0.0433628 0.956637 0.0193994 0.00462748 0.0186551 0.00441159 0.00560063 0.00634492 0.224025 0.253797 58.0533 -87.8994 126.144 15.9326 145.037 0.000142407 0.267328 192.716 0.310164 0.0673215 0.00409869 0.000562423 0.00138524 0.986958 0.991715 -2.99112e-06 -85.6564 0.0930911 31167.5 310.983 0.983496 0.319146 0.738737 0.738732 9.99958 2.98679e-06 1.19471e-05 0.134565 0.983424 0.9313 -0.0132915 4.9325e-06 0.517292 -2.02308e-20 7.50768e-24 -2.02233e-20 0.00139653 0.997815 8.60281e-05 0.152742 2.85285 0.00139653 0.997815 0.794455 0.00106852 0.00188149 0.000860281 0.455372 0.00188149 0.444798 0.000131397 1.02 0.888835 0.534357 0.287652 1.71963e-07 3.08566e-09 2369.82 3141.36 -0.0584264 0.482213 0.277257 0.254929 -0.593041 -0.169577 0.486912 -0.265663 -0.221259 2.721 1 0 295.142 0 2.24312 2.719 0.000299043 0.868819 0.702899 0.313273 0.435574 2.24329 139.611 83.6159 18.7032 60.7195 0.00403788 0 -40 10
1.82 5.26428e-08 2.54003e-06 0.149309 0.149309 0.0120255 2.39286e-05 0.00115456 0.186637 0.000658845 0.187291 0.957192 101.403 0.234315 0.86291 4.59711 0.065685 0.0433689 0.956631 0.0193988 0.00462794 0.0186545 0.00441199 0.00560121 0.00634551 0.224048 0.25382 58.0533 -87.8994 126.144 15.9325 145.037 0.000142409 0.267328 192.716 0.310163 0.0673215 0.00409869 0.000562424 0.00138524 0.986958 0.991715 -2.99114e-06 -85.6564 0.0930912 31167.5 310.996 0.983496 0.319146 0.738749 0.738744 9.99958 2.98679e-06 1.19471e-05 0.13457 0.983424 0.931299 -0.0132915 4.93253e-06 0.517312 -2.02324e-20 7.50833e-24 -2.02249e-20 0.00139653 0.997815 8.60282e-05 0.152742 2.85285 0.00139653 0.997815 0.794526 0.00106854 0.00188149 0.000860282 0.455372 0.00188149 0.444803 0.0001314 1.02 0.888836 0.534357 0.287653 1.71963e-07 3.08569e-09 2369.8 3141.41 -0.0584315 0.482213 0.277257 0.254932 -0.59304 -0.169578 0.486896 -0.26566 -0.221245 2.722 1 0 295.137 0 2.24325 2.72 0.000299041 0.868848 0.702942 0.313234 0.435596 2.24343 139.619 83.6153 18.7032 60.7192 0.00403791 0 -40 10
1.821 5.26717e-08 2.54003e-06 0.149341 0.14934 0.0120255 2.39417e-05 0.00115456 0.186676 0.000658846 0.18733 0.957283 101.402 0.234304 0.863044 4.59776 0.0656959 0.0433751 0.956625 0.0193982 0.00462841 0.0186539 0.00441239 0.00560178 0.0063461 0.224071 0.253844 58.0534 -87.8994 126.143 15.9325 145.037 0.000142412 0.267328 192.716 0.310163 0.0673214 0.00409869 0.000562425 0.00138524 0.986958 0.991715 -2.99115e-06 -85.6564 0.0930913 31167.5 311.008 0.983496 0.319146 0.738761 0.738756 9.99958 2.9868e-06 1.19471e-05 0.134575 0.983424 0.931298 -0.0132915 4.93256e-06 0.517332 -2.0234e-20 7.50898e-24 -2.02265e-20 0.00139653 0.997815 8.60283e-05 0.152742 2.85285 0.00139653 0.997815 0.794598 0.00106856 0.00188149 0.000860283 0.455371 0.00188149 0.444808 0.000131402 1.02 0.888837 0.534356 0.287655 1.71963e-07 3.08571e-09 2369.78 3141.46 -0.0584365 0.482213 0.277257 0.254935 -0.593039 -0.169578 0.48688 -0.265658 -0.221231 2.723 1 0 295.133 0 2.24339 2.721 0.00029904 0.868877 0.702984 0.313195 0.435619 2.24357 139.626 83.6147 18.7032 60.7189 0.00403793 0 -40 10
1.822 5.27005e-08 2.54004e-06 0.149372 0.149372 0.0120255 2.39548e-05 0.00115456 0.186715 0.000658846 0.187369 0.957374 101.402 0.234293 0.863177 4.59842 0.0657067 0.0433813 0.956619 0.0193976 0.00462888 0.0186533 0.0044128 0.00560236 0.0063467 0.224094 0.253868 58.0535 -87.8994 126.143 15.9325 145.037 0.000142414 0.267328 192.716 0.310162 0.0673213 0.0040987 0.000562425 0.00138524 0.986958 0.991715 -2.99117e-06 -85.6564 0.0930914 31167.4 311.021 0.983496 0.319146 0.738773 0.738768 9.99958 2.9868e-06 1.19471e-05 0.13458 0.983424 0.931297 -0.0132915 4.93259e-06 0.517353 -2.02357e-20 7.50962e-24 -2.02282e-20 0.00139654 0.997815 8.60284e-05 0.152743 2.85285 0.00139654 0.997815 0.794669 0.00106857 0.00188149 0.000860284 0.455371 0.00188149 0.444813 0.000131404 1.02 0.888838 0.534356 0.287657 1.71963e-07 3.08573e-09 2369.77 3141.51 -0.0584416 0.482213 0.277256 0.254939 -0.593039 -0.169578 0.486864 -0.265656 -0.221217 2.724 1 0 295.128 0 2.24353 2.722 0.000299039 0.868906 0.703027 0.313156 0.435641 2.2437 139.633 83.6141 18.7031 60.7186 0.00403796 0 -40 10
1.823 5.27293e-08 2.54004e-06 0.149403 0.149403 0.0120255 2.39679e-05 0.00115456 0.186754 0.000658847 0.187408 0.957465 101.401 0.234282 0.863311 4.59907 0.0657175 0.0433875 0.956613 0.0193971 0.00462934 0.0186527 0.0044132 0.00560293 0.00634729 0.224117 0.253892 58.0535 -87.8994 126.143 15.9324 145.037 0.000142416 0.267329 192.715 0.310162 0.0673213 0.0040987 0.000562426 0.00138525 0.986958 0.991715 -2.99118e-06 -85.6564 0.0930914 31167.4 311.034 0.983496 0.319146 0.738785 0.73878 9.99958 2.98681e-06 1.19471e-05 0.134584 0.983425 0.931296 -0.0132915 4.93262e-06 0.517373 -2.02373e-20 7.51027e-24 -2.02298e-20 0.00139654 0.997815 8.60285e-05 0.152743 2.85285 0.00139654 0.997815 0.79474 0.00106859 0.0018815 0.000860285 0.455371 0.00188149 0.444818 0.000131407 1.02 0.888839 0.534356 0.287658 1.71964e-07 3.08575e-09 2369.75 3141.56 -0.0584467 0.482213 0.277256 0.254942 -0.593038 -0.169578 0.486848 -0.265654 -0.221203 2.725 1 0 295.124 0 2.24366 2.723 0.000299038 0.868935 0.70307 0.313118 0.435663 2.24384 139.641 83.6135 18.7031 60.7184 0.00403798 0 -40 10
1.824 5.27582e-08 2.54004e-06 0.149435 0.149434 0.0120255 2.3981e-05 0.00115456 0.186793 0.000658847 0.187447 0.957556 101.4 0.234272 0.863444 4.59973 0.0657284 0.0433937 0.956606 0.0193965 0.00462981 0.0186521 0.00441361 0.00560351 0.00634788 0.22414 0.253915 58.0536 -87.8994 126.143 15.9324 145.037 0.000142419 0.267329 192.715 0.310162 0.0673212 0.0040987 0.000562427 0.00138525 0.986958 0.991715 -2.9912e-06 -85.6564 0.0930915 31167.4 311.046 0.983496 0.319146 0.738797 0.738792 9.99958 2.98681e-06 1.19472e-05 0.134589 0.983425 0.931295 -0.0132915 4.93265e-06 0.517393 -2.02389e-20 7.51092e-24 -2.02314e-20 0.00139654 0.997815 8.60285e-05 0.152743 2.85285 0.00139654 0.997815 0.794811 0.0010686 0.0018815 0.000860285 0.455371 0.0018815 0.444823 0.000131409 1.02 0.88884 0.534356 0.28766 1.71964e-07 3.08578e-09 2369.73 3141.61 -0.0584517 0.482213 0.277256 0.254945 -0.593037 -0.169578 0.486832 -0.265652 -0.221189 2.726 1 0 295.119 0 2.2438 2.724 0.000299036 0.868964 0.703113 0.313079 0.435685 2.24398 139.648 83.6129 18.7031 60.7181 0.00403801 0 -40 10
1.825 5.2787e-08 2.54004e-06 0.149466 0.149465 0.0120254 2.39941e-05 0.00115456 0.186832 0.000658848 0.187486 0.957647 101.4 0.234261 0.863578 4.60038 0.0657392 0.0433998 0.9566 0.0193959 0.00463028 0.0186515 0.00441401 0.00560409 0.00634848 0.224163 0.253939 58.0537 -87.8994 126.142 15.9324 145.037 0.000142421 0.267329 192.715 0.310161 0.0673212 0.0040987 0.000562427 0.00138525 0.986958 0.991715 -2.99121e-06 -85.6564 0.0930916 31167.4 311.059 0.983496 0.319146 0.738809 0.738804 9.99958 2.98682e-06 1.19472e-05 0.134594 0.983425 0.931294 -0.0132915 4.93268e-06 0.517414 -2.02405e-20 7.51157e-24 -2.0233e-20 0.00139654 0.997815 8.60286e-05 0.152743 2.85285 0.00139654 0.997815 0.794882 0.00106862 0.0018815 0.000860286 0.45537 0.0018815 0.444828 0.000131411 1.02 0.888841 0.534355 0.287661 1.71964e-07 3.0858e-09 2369.72 3141.66 -0.0584568 0.482213 0.277256 0.254948 -0.593037 -0.169578 0.486815 -0.26565 -0.221175 2.727 1 0 295.114 0 2.24393 2.725 0.000299035 0.868993 0.703155 0.31304 0.435707 2.24411 139.655 83.6124 18.703 60.7178 0.00403803 0 -40 10
1.826 5.28158e-08 2.54004e-06 0.149497 0.149496 0.0120254 2.40072e-05 0.00115457 0.186871 0.000658848 0.187525 0.957738 101.399 0.23425 0.863711 4.60104 0.06575 0.043406 0.956594 0.0193953 0.00463075 0.0186509 0.00441442 0.00560466 0.00634907 0.224187 0.253963 58.0537 -87.8994 126.142 15.9323 145.037 0.000142423 0.267329 192.715 0.310161 0.0673211 0.00409871 0.000562428 0.00138525 0.986958 0.991715 -2.99123e-06 -85.6563 0.0930917 31167.4 311.072 0.983496 0.319146 0.738821 0.738816 9.99958 2.98682e-06 1.19472e-05 0.134599 0.983425 0.931293 -0.0132915 4.93271e-06 0.517434 -2.02422e-20 7.51222e-24 -2.02347e-20 0.00139654 0.997815 8.60287e-05 0.152743 2.85285 0.00139654 0.997815 0.794953 0.00106864 0.0018815 0.000860287 0.45537 0.0018815 0.444833 0.000131414 1.02 0.888842 0.534355 0.287663 1.71964e-07 3.08582e-09 2369.7 3141.71 -0.0584619 0.482213 0.277255 0.254952 -0.593036 -0.169578 0.486799 -0.265648 -0.221161 2.728 1 0 295.11 0 2.24407 2.726 0.000299034 0.869022 0.703198 0.313001 0.435729 2.24425 139.663 83.6118 18.703 60.7175 0.00403805 0 -40 10
1.827 5.28447e-08 2.54005e-06 0.149528 0.149528 0.0120254 2.40203e-05 0.00115457 0.18691 0.000658849 0.187564 0.957829 101.398 0.234239 0.863845 4.6017 0.0657609 0.0434122 0.956588 0.0193948 0.00463121 0.0186503 0.00441482 0.00560524 0.00634967 0.22421 0.253987 58.0538 -87.8994 126.142 15.9323 145.037 0.000142426 0.267329 192.715 0.31016 0.0673211 0.00409871 0.000562429 0.00138525 0.986958 0.991715 -2.99124e-06 -85.6563 0.0930918 31167.3 311.084 0.983496 0.319146 0.738833 0.738829 9.99958 2.98683e-06 1.19472e-05 0.134603 0.983426 0.931292 -0.0132915 4.93274e-06 0.517454 -2.02438e-20 7.51287e-24 -2.02363e-20 0.00139654 0.997815 8.60288e-05 0.152743 2.85286 0.00139654 0.997815 0.795024 0.00106865 0.0018815 0.000860288 0.45537 0.0018815 0.444838 0.000131416 1.02 0.888844 0.534355 0.287664 1.71965e-07 3.08585e-09 2369.69 3141.77 -0.0584669 0.482213 0.277255 0.254955 -0.593035 -0.169578 0.486783 -0.265646 -0.221147 2.729 1 0 295.105 0 2.24421 2.727 0.000299033 0.869052 0.703241 0.312963 0.435751 2.24439 139.67 83.6112 18.703 60.7172 0.00403808 0 -40 10
1.828 5.28735e-08 2.54005e-06 0.149559 0.149559 0.0120254 2.40334e-05 0.00115457 0.186949 0.000658849 0.187603 0.95792 101.398 0.234228 0.863979 4.60235 0.0657717 0.0434184 0.956582 0.0193942 0.00463168 0.0186497 0.00441523 0.00560582 0.00635026 0.224233 0.254011 58.0538 -87.8994 126.142 15.9323 145.037 0.000142428 0.26733 192.715 0.31016 0.067321 0.00409871 0.000562429 0.00138526 0.986958 0.991715 -2.99126e-06 -85.6563 0.0930919 31167.3 311.097 0.983496 0.319146 0.738845 0.738841 9.99958 2.98683e-06 1.19472e-05 0.134608 0.983426 0.931291 -0.0132915 4.93277e-06 0.517475 -2.02454e-20 7.51352e-24 -2.02379e-20 0.00139654 0.997815 8.60289e-05 0.152743 2.85286 0.00139654 0.997815 0.795096 0.00106867 0.0018815 0.000860289 0.45537 0.0018815 0.444843 0.000131419 1.02 0.888845 0.534354 0.287666 1.71965e-07 3.08587e-09 2369.67 3141.82 -0.058472 0.482213 0.277255 0.254958 -0.593035 -0.169578 0.486767 -0.265644 -0.221133 2.73 1 0 295.101 0 2.24434 2.728 0.000299031 0.869081 0.703284 0.312924 0.435773 2.24452 139.677 83.6106 18.7029 60.7169 0.0040381 0 -40 10
1.829 5.29024e-08 2.54005e-06 0.14959 0.14959 0.0120254 2.40465e-05 0.00115457 0.186988 0.00065885 0.187642 0.958012 101.397 0.234217 0.864112 4.60301 0.0657825 0.0434246 0.956575 0.0193936 0.00463215 0.0186491 0.00441563 0.00560639 0.00635086 0.224256 0.254034 58.0539 -87.8994 126.142 15.9322 145.037 0.00014243 0.26733 192.714 0.310159 0.067321 0.00409872 0.00056243 0.00138526 0.986958 0.991715 -2.99127e-06 -85.6563 0.093092 31167.3 311.11 0.983496 0.319146 0.738857 0.738853 9.99958 2.98684e-06 1.19472e-05 0.134613 0.983426 0.93129 -0.0132915 4.9328e-06 0.517495 -2.02471e-20 7.51417e-24 -2.02395e-20 0.00139654 0.997814 8.60289e-05 0.152744 2.85286 0.00139654 0.997815 0.795167 0.00106868 0.0018815 0.000860289 0.45537 0.0018815 0.444848 0.000131421 1.02 0.888846 0.534354 0.287667 1.71965e-07 3.08589e-09 2369.65 3141.87 -0.0584771 0.482213 0.277254 0.254961 -0.593034 -0.169578 0.486751 -0.265642 -0.221119 2.731 1 0 295.096 0 2.24448 2.729 0.00029903 0.86911 0.703326 0.312886 0.435795 2.24466 139.685 83.61 18.7029 60.7166 0.00403813 0 -40 10
1.83 5.29312e-08 2.54005e-06 0.149621 0.149621 0.0120254 2.40596e-05 0.00115457 0.187027 0.00065885 0.187681 0.958103 101.396 0.234207 0.864246 4.60367 0.0657934 0.0434308 0.956569 0.019393 0.00463262 0.0186485 0.00441604 0.00560697 0.00635145 0.224279 0.254058 58.054 -87.8994 126.141 15.9322 145.037 0.000142433 0.26733 192.714 0.310159 0.0673209 0.00409872 0.000562431 0.00138526 0.986958 0.991715 -2.99129e-06 -85.6563 0.0930921 31167.3 311.123 0.983496 0.319146 0.738869 0.738865 9.99958 2.98684e-06 1.19473e-05 0.134618 0.983426 0.931289 -0.0132915 4.93282e-06 0.517516 -2.02487e-20 7.51482e-24 -2.02412e-20 0.00139655 0.997814 8.6029e-05 0.152744 2.85286 0.00139655 0.997815 0.795238 0.0010687 0.00188151 0.00086029 0.455369 0.0018815 0.444853 0.000131423 1.02 0.888847 0.534354 0.287669 1.71966e-07 3.08591e-09 2369.64 3141.92 -0.0584822 0.482213 0.277254 0.254964 -0.593034 -0.169578 0.486735 -0.26564 -0.221105 2.732 1 0 295.092 0 2.24462 2.73 0.000299029 0.869139 0.703369 0.312847 0.435817 2.24479 139.692 83.6094 18.7029 60.7163 0.00403815 0 -40 10
1.831 5.296e-08 2.54005e-06 0.149653 0.149652 0.0120254 2.40727e-05 0.00115457 0.187066 0.000658851 0.18772 0.958194 101.396 0.234196 0.864379 4.60433 0.0658042 0.0434371 0.956563 0.0193925 0.00463309 0.018648 0.00441644 0.00560755 0.00635205 0.224302 0.254082 58.054 -87.8994 126.141 15.9321 145.037 0.000142435 0.26733 192.714 0.310159 0.0673209 0.00409872 0.000562431 0.00138526 0.986958 0.991715 -2.9913e-06 -85.6563 0.0930921 31167.2 311.135 0.983496 0.319146 0.738881 0.738877 9.99958 2.98685e-06 1.19473e-05 0.134622 0.983426 0.931288 -0.0132915 4.93285e-06 0.517536 -2.02503e-20 7.51547e-24 -2.02428e-20 0.00139655 0.997814 8.60291e-05 0.152744 2.85286 0.00139655 0.997815 0.795309 0.00106872 0.00188151 0.000860291 0.455369 0.00188151 0.444858 0.000131426 1.02 0.888848 0.534353 0.28767 1.71966e-07 3.08594e-09 2369.62 3141.97 -0.0584872 0.482213 0.277254 0.254968 -0.593033 -0.169578 0.486719 -0.265637 -0.221091 2.733 1 0 295.087 0 2.24475 2.731 0.000299027 0.869168 0.703412 0.312808 0.435839 2.24493 139.699 83.6088 18.7028 60.7161 0.00403818 0 -40 10
1.832 5.29889e-08 2.54005e-06 0.149684 0.149683 0.0120253 2.40858e-05 0.00115457 0.187104 0.000658851 0.187759 0.958285 101.395 0.234185 0.864513 4.60499 0.0658151 0.0434433 0.956557 0.0193919 0.00463355 0.0186474 0.00441685 0.00560813 0.00635265 0.224325 0.254106 58.0541 -87.8994 126.141 15.9321 145.037 0.000142437 0.26733 192.714 0.310158 0.0673208 0.00409873 0.000562432 0.00138527 0.986957 0.991715 -2.99132e-06 -85.6563 0.0930922 31167.2 311.148 0.983496 0.319146 0.738893 0.738889 9.99958 2.98685e-06 1.19473e-05 0.134627 0.983427 0.931287 -0.0132915 4.93288e-06 0.517556 -2.02519e-20 7.51612e-24 -2.02444e-20 0.00139655 0.997814 8.60292e-05 0.152744 2.85286 0.00139655 0.997815 0.79538 0.00106873 0.00188151 0.000860292 0.455369 0.00188151 0.444863 0.000131428 1.02 0.888849 0.534353 0.287672 1.71966e-07 3.08596e-09 2369.6 3142.02 -0.0584923 0.482213 0.277254 0.254971 -0.593032 -0.169578 0.486703 -0.265635 -0.221077 2.734 1 0 295.082 0 2.24489 2.732 0.000299026 0.869198 0.703454 0.31277 0.435861 2.24507 139.706 83.6082 18.7028 60.7158 0.0040382 0 -40 10
1.833 5.30177e-08 2.54006e-06 0.149715 0.149714 0.0120253 2.4099e-05 0.00115457 0.187143 0.000658852 0.187797 0.958376 101.394 0.234174 0.864647 4.60565 0.0658259 0.0434495 0.95655 0.0193913 0.00463402 0.0186468 0.00441726 0.0056087 0.00635324 0.224348 0.25413 58.0542 -87.8994 126.141 15.9321 145.037 0.00014244 0.267331 192.714 0.310158 0.0673208 0.00409873 0.000562433 0.00138527 0.986957 0.991715 -2.99133e-06 -85.6563 0.0930923 31167.2 311.161 0.983496 0.319146 0.738905 0.738901 9.99958 2.98686e-06 1.19473e-05 0.134632 0.983427 0.931286 -0.0132915 4.93291e-06 0.517577 -2.02536e-20 7.51678e-24 -2.02461e-20 0.00139655 0.997814 8.60293e-05 0.152744 2.85286 0.00139655 0.997815 0.795451 0.00106875 0.00188151 0.000860293 0.455369 0.00188151 0.444868 0.00013143 1.02 0.88885 0.534353 0.287673 1.71966e-07 3.08598e-09 2369.59 3142.07 -0.0584974 0.482214 0.277253 0.254974 -0.593032 -0.169578 0.486686 -0.265633 -0.221063 2.735 1 0 295.078 0 2.24503 2.733 0.000299025 0.869227 0.703497 0.312731 0.435883 2.2452 139.714 83.6076 18.7027 60.7155 0.00403823 0 -40 10
1.834 5.30465e-08 2.54006e-06 0.149746 0.149745 0.0120253 2.41121e-05 0.00115457 0.187182 0.000658852 0.187836 0.958467 101.394 0.234163 0.86478 4.60631 0.0658368 0.0434557 0.956544 0.0193907 0.00463449 0.0186462 0.00441766 0.00560928 0.00635384 0.224371 0.254154 58.0542 -87.8994 126.141 15.932 145.037 0.000142442 0.267331 192.714 0.310157 0.0673207 0.00409873 0.000562433 0.00138527 0.986957 0.991715 -2.99135e-06 -85.6563 0.0930924 31167.2 311.174 0.983496 0.319146 0.738917 0.738913 9.99958 2.98686e-06 1.19473e-05 0.134637 0.983427 0.931285 -0.0132915 4.93294e-06 0.517597 -2.02552e-20 7.51743e-24 -2.02477e-20 0.00139655 0.997814 8.60293e-05 0.152744 2.85286 0.00139655 0.997815 0.795521 0.00106876 0.00188151 0.000860293 0.455368 0.00188151 0.444873 0.000131433 1.02 0.888851 0.534352 0.287675 1.71967e-07 3.08601e-09 2369.57 3142.12 -0.0585025 0.482214 0.277253 0.254977 -0.593031 -0.169578 0.48667 -0.265631 -0.221049 2.736 1 0 295.073 0 2.24516 2.734 0.000299024 0.869256 0.70354 0.312693 0.435905 2.24534 139.721 83.607 18.7027 60.7152 0.00403825 0 -40 10
1.835 5.30754e-08 2.54006e-06 0.149777 0.149776 0.0120253 2.41252e-05 0.00115457 0.187221 0.000658853 0.187875 0.958558 101.393 0.234152 0.864914 4.60697 0.0658476 0.043462 0.956538 0.0193901 0.00463496 0.0186456 0.00441807 0.00560986 0.00635444 0.224394 0.254177 58.0543 -87.8994 126.14 15.932 145.038 0.000142444 0.267331 192.713 0.310157 0.0673207 0.00409873 0.000562434 0.00138527 0.986957 0.991715 -2.99136e-06 -85.6563 0.0930925 31167.2 311.186 0.983496 0.319146 0.73893 0.738925 9.99958 2.98687e-06 1.19474e-05 0.134641 0.983427 0.931284 -0.0132915 4.93297e-06 0.517618 -2.02568e-20 7.51808e-24 -2.02493e-20 0.00139655 0.997814 8.60294e-05 0.152745 2.85286 0.00139655 0.997815 0.795592 0.00106878 0.00188151 0.000860294 0.455368 0.00188151 0.444878 0.000131435 1.02 0.888852 0.534352 0.287676 1.71967e-07 3.08603e-09 2369.56 3142.17 -0.0585075 0.482214 0.277253 0.254981 -0.59303 -0.169578 0.486654 -0.265629 -0.221035 2.737 1 0 295.069 0 2.2453 2.735 0.000299022 0.869285 0.703582 0.312655 0.435927 2.24548 139.728 83.6064 18.7027 60.7149 0.00403828 0 -40 10
1.836 5.31042e-08 2.54006e-06 0.149807 0.149807 0.0120253 2.41383e-05 0.00115457 0.187259 0.000658853 0.187914 0.95865 101.392 0.234142 0.865048 4.60763 0.0658585 0.0434682 0.956532 0.0193896 0.00463543 0.018645 0.00441847 0.00561044 0.00635503 0.224418 0.254201 58.0543 -87.8995 126.14 15.932 145.038 0.000142447 0.267331 192.713 0.310156 0.0673206 0.00409874 0.000562435 0.00138527 0.986957 0.991715 -2.99138e-06 -85.6563 0.0930926 31167.1 311.199 0.983496 0.319146 0.738942 0.738937 9.99958 2.98687e-06 1.19474e-05 0.134646 0.983428 0.931283 -0.0132915 4.933e-06 0.517638 -2.02585e-20 7.51873e-24 -2.0251e-20 0.00139655 0.997814 8.60295e-05 0.152745 2.85286 0.00139655 0.997815 0.795663 0.0010688 0.00188152 0.000860295 0.455368 0.00188151 0.444883 0.000131437 1.02 0.888853 0.534352 0.287678 1.71967e-07 3.08605e-09 2369.54 3142.22 -0.0585126 0.482214 0.277252 0.254984 -0.59303 -0.169579 0.486638 -0.265627 -0.221021 2.738 1 0 295.064 0 2.24543 2.736 0.000299021 0.869314 0.703625 0.312616 0.435949 2.24561 139.736 83.6058 18.7026 60.7146 0.0040383 0 -40 10
1.837 5.3133e-08 2.54006e-06 0.149838 0.149838 0.0120253 2.41514e-05 0.00115457 0.187298 0.000658853 0.187952 0.958741 101.392 0.234131 0.865181 4.60829 0.0658693 0.0434744 0.956526 0.019389 0.0046359 0.0186444 0.00441888 0.00561102 0.00635563 0.224441 0.254225 58.0544 -87.8995 126.14 15.9319 145.038 0.000142449 0.267331 192.713 0.310156 0.0673206 0.00409874 0.000562435 0.00138528 0.986957 0.991715 -2.99139e-06 -85.6562 0.0930927 31167.1 311.212 0.983496 0.319146 0.738954 0.738949 9.99958 2.98688e-06 1.19474e-05 0.134651 0.983428 0.931282 -0.0132915 4.93303e-06 0.517659 -2.02601e-20 7.51939e-24 -2.02526e-20 0.00139655 0.997814 8.60296e-05 0.152745 2.85287 0.00139655 0.997815 0.795734 0.00106881 0.00188152 0.000860296 0.455368 0.00188152 0.444888 0.00013144 1.02 0.888855 0.534352 0.287679 1.71967e-07 3.08608e-09 2369.52 3142.27 -0.0585177 0.482214 0.277252 0.254987 -0.593029 -0.169579 0.486622 -0.265625 -0.221006 2.739 1 0 295.06 0 2.24557 2.737 0.00029902 0.869344 0.703668 0.312578 0.435971 2.24575 139.743 83.6052 18.7026 60.7143 0.00403833 0 -40 10
1.838 5.31619e-08 2.54006e-06 0.149869 0.149869 0.0120253 2.41645e-05 0.00115457 0.187337 0.000658854 0.187991 0.958832 101.391 0.23412 0.865315 4.60895 0.0658802 0.0434807 0.956519 0.0193884 0.00463637 0.0186438 0.00441929 0.0056116 0.00635623 0.224464 0.254249 58.0545 -87.8995 126.14 15.9319 145.038 0.000142451 0.267331 192.713 0.310156 0.0673205 0.00409874 0.000562436 0.00138528 0.986957 0.991715 -2.99141e-06 -85.6562 0.0930928 31167.1 311.225 0.983496 0.319146 0.738966 0.738961 9.99958 2.98688e-06 1.19474e-05 0.134656 0.983428 0.931281 -0.0132915 4.93306e-06 0.517679 -2.02617e-20 7.52004e-24 -2.02542e-20 0.00139655 0.997814 8.60297e-05 0.152745 2.85287 0.00139655 0.997815 0.795805 0.00106883 0.00188152 0.000860297 0.455368 0.00188152 0.444893 0.000131442 1.02 0.888856 0.534351 0.287681 1.71968e-07 3.0861e-09 2369.51 3142.32 -0.0585228 0.482214 0.277252 0.25499 -0.593028 -0.169579 0.486606 -0.265623 -0.220992 2.74 1 0 295.055 0 2.24571 2.738 0.000299019 0.869373 0.703711 0.312539 0.435993 2.24588 139.75 83.6046 18.7026 60.7141 0.00403835 0 -40 10
1.839 5.31907e-08 2.54007e-06 0.1499 0.1499 0.0120252 2.41776e-05 0.00115458 0.187375 0.000658854 0.188029 0.958923 101.39 0.234109 0.865449 4.60961 0.065891 0.0434869 0.956513 0.0193878 0.00463684 0.0186432 0.0044197 0.00561218 0.00635683 0.224487 0.254273 58.0545 -87.8995 126.139 15.9318 145.038 0.000142454 0.267332 192.713 0.310155 0.0673205 0.00409875 0.000562437 0.00138528 0.986957 0.991715 -2.99142e-06 -85.6562 0.0930928 31167.1 311.237 0.983496 0.319146 0.738978 0.738973 9.99958 2.98689e-06 1.19474e-05 0.134661 0.983428 0.93128 -0.0132915 4.93309e-06 0.5177 -2.02634e-20 7.52069e-24 -2.02559e-20 0.00139656 0.997814 8.60297e-05 0.152745 2.85287 0.00139656 0.997815 0.795876 0.00106884 0.00188152 0.000860297 0.455367 0.00188152 0.444898 0.000131444 1.02 0.888857 0.534351 0.287682 1.71968e-07 3.08612e-09 2369.49 3142.37 -0.0585279 0.482214 0.277252 0.254994 -0.593028 -0.169579 0.48659 -0.265621 -0.220978 2.741 1 0 295.05 0 2.24584 2.739 0.000299017 0.869402 0.703753 0.312501 0.436015 2.24602 139.758 83.604 18.7025 60.7138 0.00403837 0 -40 10
1.84 5.32195e-08 2.54007e-06 0.149931 0.14993 0.0120252 2.41907e-05 0.00115458 0.187414 0.000658855 0.188068 0.959015 101.39 0.234098 0.865582 4.61028 0.0659019 0.0434932 0.956507 0.0193872 0.00463731 0.0186426 0.0044201 0.00561276 0.00635742 0.22451 0.254297 58.0546 -87.8995 126.139 15.9318 145.038 0.000142456 0.267332 192.713 0.310155 0.0673204 0.00409875 0.000562437 0.00138528 0.986957 0.991715 -2.99144e-06 -85.6562 0.0930929 31167 311.25 0.983496 0.319146 0.73899 0.738986 9.99958 2.98689e-06 1.19475e-05 0.134665 0.983428 0.931279 -0.0132915 4.93312e-06 0.51772 -2.0265e-20 7.52134e-24 -2.02575e-20 0.00139656 0.997814 8.60298e-05 0.152745 2.85287 0.00139656 0.997815 0.795946 0.00106886 0.00188152 0.000860298 0.455367 0.00188152 0.444903 0.000131447 1.02 0.888858 0.534351 0.287684 1.71968e-07 3.08614e-09 2369.47 3142.42 -0.0585329 0.482214 0.277251 0.254997 -0.593027 -0.169579 0.486574 -0.265619 -0.220964 2.742 1 0 295.046 0 2.24598 2.74 0.000299016 0.869431 0.703796 0.312463 0.436037 2.24616 139.765 83.6034 18.7025 60.7135 0.0040384 0 -40 10
1.841 5.32484e-08 2.54007e-06 0.149962 0.149961 0.0120252 2.42038e-05 0.00115458 0.187452 0.000658855 0.188106 0.959106 101.389 0.234087 0.865716 4.61094 0.0659127 0.0434994 0.956501 0.0193867 0.00463778 0.018642 0.00442051 0.00561334 0.00635802 0.224533 0.254321 58.0547 -87.8995 126.139 15.9318 145.038 0.000142458 0.267332 192.712 0.310154 0.0673203 0.00409875 0.000562438 0.00138529 0.986957 0.991715 -2.99145e-06 -85.6562 0.093093 31167 311.263 0.983496 0.319146 0.739002 0.738998 9.99958 2.9869e-06 1.19475e-05 0.13467 0.983429 0.931278 -0.0132915 4.93315e-06 0.51774 -2.02667e-20 7.522e-24 -2.02591e-20 0.00139656 0.997814 8.60299e-05 0.152745 2.85287 0.00139656 0.997815 0.796017 0.00106888 0.00188152 0.000860299 0.455367 0.00188152 0.444908 0.000131449 1.02 0.888859 0.53435 0.287685 1.71969e-07 3.08617e-09 2369.46 3142.47 -0.058538 0.482214 0.277251 0.255 -0.593027 -0.169579 0.486557 -0.265616 -0.22095 2.743 1 0 295.041 0 2.24612 2.741 0.000299015 0.869461 0.703839 0.312425 0.436059 2.24629 139.772 83.6029 18.7025 60.7132 0.00403842 0 -40 10
1.842 5.32772e-08 2.54007e-06 0.149993 0.149992 0.0120252 2.42169e-05 0.00115458 0.187491 0.000658856 0.188145 0.959197 101.388 0.234076 0.86585 4.6116 0.0659236 0.0435057 0.956494 0.0193861 0.00463825 0.0186414 0.00442092 0.00561392 0.00635862 0.224557 0.254345 58.0547 -87.8995 126.139 15.9317 145.038 0.000142461 0.267332 192.712 0.310154 0.0673203 0.00409876 0.000562439 0.00138529 0.986957 0.991715 -2.99147e-06 -85.6562 0.0930931 31167 311.276 0.983496 0.319146 0.739014 0.73901 9.99958 2.9869e-06 1.19475e-05 0.134675 0.983429 0.931277 -0.0132915 4.93318e-06 0.517761 -2.02683e-20 7.52265e-24 -2.02608e-20 0.00139656 0.997814 8.603e-05 0.152746 2.85287 0.00139656 0.997815 0.796088 0.00106889 0.00188152 0.0008603 0.455367 0.00188152 0.444913 0.000131451 1.02 0.88886 0.53435 0.287687 1.71969e-07 3.08619e-09 2369.44 3142.53 -0.0585431 0.482214 0.277251 0.255003 -0.593026 -0.169579 0.486541 -0.265614 -0.220936 2.744 1 0 295.037 0 2.24625 2.742 0.000299013 0.86949 0.703881 0.312386 0.436081 2.24643 139.78 83.6023 18.7024 60.7129 0.00403845 0 -40 10
1.843 5.33061e-08 2.54007e-06 0.150023 0.150023 0.0120252 2.423e-05 0.00115458 0.187529 0.000658856 0.188183 0.959288 101.388 0.234066 0.865984 4.61227 0.0659344 0.043512 0.956488 0.0193855 0.00463872 0.0186408 0.00442133 0.0056145 0.00635922 0.22458 0.254369 58.0548 -87.8995 126.139 15.9317 145.038 0.000142463 0.267332 192.712 0.310153 0.0673202 0.00409876 0.000562439 0.00138529 0.986957 0.991715 -2.99148e-06 -85.6562 0.0930932 31167 311.289 0.983496 0.319146 0.739026 0.739022 9.99958 2.98691e-06 1.19475e-05 0.13468 0.983429 0.931276 -0.0132915 4.93321e-06 0.517782 -2.02699e-20 7.52331e-24 -2.02624e-20 0.00139656 0.997814 8.60301e-05 0.152746 2.85287 0.00139656 0.997815 0.796159 0.00106891 0.00188153 0.000860301 0.455366 0.00188152 0.444918 0.000131454 1.02 0.888861 0.53435 0.287688 1.71969e-07 3.08621e-09 2369.42 3142.58 -0.0585482 0.482214 0.277251 0.255007 -0.593025 -0.169579 0.486525 -0.265612 -0.220922 2.745 1 0 295.032 0 2.24639 2.743 0.000299012 0.869519 0.703924 0.312348 0.436103 2.24657 139.787 83.6017 18.7024 60.7126 0.00403847 0 -40 10
1.844 5.33349e-08 2.54007e-06 0.150054 0.150054 0.0120252 2.42431e-05 0.00115458 0.187568 0.000658857 0.188222 0.95938 101.387 0.234055 0.866117 4.61293 0.0659453 0.0435182 0.956482 0.0193849 0.00463919 0.0186402 0.00442173 0.00561508 0.00635982 0.224603 0.254393 58.0548 -87.8995 126.138 15.9317 145.038 0.000142465 0.267333 192.712 0.310153 0.0673202 0.00409876 0.00056244 0.00138529 0.986957 0.991715 -2.9915e-06 -85.6562 0.0930933 31167 311.301 0.983496 0.319146 0.739038 0.739034 9.99958 2.98691e-06 1.19475e-05 0.134685 0.983429 0.931275 -0.0132915 4.93324e-06 0.517802 -2.02716e-20 7.52396e-24 -2.0264e-20 0.00139656 0.997814 8.60301e-05 0.152746 2.85287 0.00139656 0.997815 0.796229 0.00106892 0.00188153 0.000860301 0.455366 0.00188153 0.444923 0.000131456 1.02 0.888862 0.534349 0.28769 1.71969e-07 3.08624e-09 2369.41 3142.63 -0.0585533 0.482214 0.27725 0.25501 -0.593025 -0.169579 0.486509 -0.26561 -0.220908 2.746 1 0 295.027 0 2.24652 2.744 0.000299011 0.869549 0.703967 0.31231 0.436125 2.2467 139.794 83.6011 18.7024 60.7123 0.0040385 0 -40 10
1.845 5.33637e-08 2.54008e-06 0.150085 0.150084 0.0120252 2.42562e-05 0.00115458 0.187606 0.000658857 0.18826 0.959471 101.386 0.234044 0.866251 4.6136 0.0659561 0.0435245 0.956475 0.0193843 0.00463966 0.0186396 0.00442214 0.00561566 0.00636042 0.224626 0.254417 58.0549 -87.8995 126.138 15.9316 145.038 0.000142468 0.267333 192.712 0.310153 0.0673201 0.00409877 0.000562441 0.00138529 0.986957 0.991715 -2.99151e-06 -85.6562 0.0930934 31166.9 311.314 0.983496 0.319146 0.73905 0.739046 9.99958 2.98692e-06 1.19476e-05 0.134689 0.983429 0.931274 -0.0132915 4.93327e-06 0.517823 -2.02732e-20 7.52462e-24 -2.02657e-20 0.00139656 0.997814 8.60302e-05 0.152746 2.85287 0.00139656 0.997815 0.7963 0.00106894 0.00188153 0.000860302 0.455366 0.00188153 0.444928 0.000131458 1.02 0.888863 0.534349 0.287691 1.7197e-07 3.08626e-09 2369.39 3142.68 -0.0585583 0.482214 0.27725 0.255013 -0.593024 -0.169579 0.486493 -0.265608 -0.220894 2.747 1 0 295.023 0 2.24666 2.745 0.00029901 0.869578 0.704009 0.312272 0.436147 2.24684 139.802 83.6005 18.7023 60.712 0.00403852 0 -40 10
1.846 5.33926e-08 2.54008e-06 0.150115 0.150115 0.0120251 2.42693e-05 0.00115458 0.187644 0.000658858 0.188299 0.959562 101.386 0.234033 0.866385 4.61426 0.065967 0.0435308 0.956469 0.0193838 0.00464013 0.018639 0.00442255 0.00561624 0.00636102 0.22465 0.254441 58.055 -87.8995 126.138 15.9316 145.038 0.00014247 0.267333 192.712 0.310152 0.0673201 0.00409877 0.000562441 0.0013853 0.986957 0.991715 -2.99153e-06 -85.6562 0.0930935 31166.9 311.327 0.983496 0.319146 0.739063 0.739058 9.99958 2.98692e-06 1.19476e-05 0.134694 0.98343 0.931273 -0.0132915 4.9333e-06 0.517843 -2.02748e-20 7.52527e-24 -2.02673e-20 0.00139656 0.997814 8.60303e-05 0.152746 2.85287 0.00139656 0.997815 0.796371 0.00106896 0.00188153 0.000860303 0.455366 0.00188153 0.444933 0.000131461 1.02 0.888864 0.534349 0.287693 1.7197e-07 3.08628e-09 2369.38 3142.73 -0.0585634 0.482215 0.27725 0.255016 -0.593023 -0.169579 0.486477 -0.265606 -0.22088 2.748 1 0 295.018 0 2.2468 2.746 0.000299008 0.869607 0.704052 0.312234 0.436169 2.24697 139.809 83.5999 18.7023 60.7118 0.00403855 0 -40 10
1.847 5.34214e-08 2.54008e-06 0.150146 0.150146 0.0120251 2.42825e-05 0.00115458 0.187683 0.000658858 0.188337 0.959654 101.385 0.234022 0.866519 4.61493 0.0659779 0.0435371 0.956463 0.0193832 0.00464061 0.0186384 0.00442296 0.00561682 0.00636162 0.224673 0.254465 58.055 -87.8995 126.138 15.9315 145.038 0.000142472 0.267333 192.711 0.310152 0.06732 0.00409877 0.000562442 0.0013853 0.986957 0.991715 -2.99154e-06 -85.6561 0.0930935 31166.9 311.34 0.983496 0.319146 0.739075 0.73907 9.99958 2.98693e-06 1.19476e-05 0.134699 0.98343 0.931272 -0.0132915 4.93333e-06 0.517864 -2.02765e-20 7.52593e-24 -2.0269e-20 0.00139656 0.997814 8.60304e-05 0.152746 2.85287 0.00139656 0.997815 0.796441 0.00106897 0.00188153 0.000860304 0.455365 0.00188153 0.444938 0.000131463 1.02 0.888866 0.534348 0.287694 1.7197e-07 3.0863e-09 2369.36 3142.78 -0.0585685 0.482215 0.277249 0.25502 -0.593023 -0.169579 0.486461 -0.265604 -0.220866 2.749 1 0 295.014 0 2.24693 2.747 0.000299007 0.869637 0.704095 0.312195 0.436191 2.24711 139.816 83.5993 18.7023 60.7115 0.00403857 0 -40 10
1.848 5.34502e-08 2.54008e-06 0.150177 0.150176 0.0120251 2.42956e-05 0.00115458 0.187721 0.000658859 0.188375 0.959745 101.384 0.234011 0.866653 4.6156 0.0659887 0.0435434 0.956457 0.0193826 0.00464108 0.0186378 0.00442337 0.0056174 0.00636222 0.224696 0.254489 58.0551 -87.8995 126.137 15.9315 145.038 0.000142475 0.267333 192.711 0.310151 0.06732 0.00409877 0.000562443 0.0013853 0.986957 0.991715 -2.99156e-06 -85.6561 0.0930936 31166.9 311.353 0.983496 0.319146 0.739087 0.739082 9.99958 2.98693e-06 1.19476e-05 0.134704 0.98343 0.931271 -0.0132915 4.93336e-06 0.517884 -2.02781e-20 7.52658e-24 -2.02706e-20 0.00139657 0.997814 8.60305e-05 0.152747 2.85288 0.00139657 0.997815 0.796512 0.00106899 0.00188153 0.000860305 0.455365 0.00188153 0.444943 0.000131465 1.02 0.888867 0.534348 0.287696 1.7197e-07 3.08633e-09 2369.34 3142.83 -0.0585736 0.482215 0.277249 0.255023 -0.593022 -0.169579 0.486444 -0.265602 -0.220852 2.75 1 0 295.009 0 2.24707 2.748 0.000299006 0.869666 0.704137 0.312157 0.436213 2.24725 139.824 83.5987 18.7022 60.7112 0.0040386 0 -40 10
1.849 5.34791e-08 2.54008e-06 0.150207 0.150207 0.0120251 2.43087e-05 0.00115458 0.187759 0.000658859 0.188414 0.959836 101.384 0.234 0.866787 4.61626 0.0659996 0.0435496 0.95645 0.019382 0.00464155 0.0186372 0.00442378 0.00561798 0.00636282 0.224719 0.254513 58.0552 -87.8995 126.137 15.9315 145.038 0.000142477 0.267334 192.711 0.310151 0.0673199 0.00409878 0.000562443 0.0013853 0.986957 0.991715 -2.99157e-06 -85.6561 0.0930937 31166.8 311.365 0.983496 0.319146 0.739099 0.739094 9.99958 2.98694e-06 1.19476e-05 0.134709 0.98343 0.93127 -0.0132915 4.93339e-06 0.517905 -2.02798e-20 7.52724e-24 -2.02722e-20 0.00139657 0.997814 8.60305e-05 0.152747 2.85288 0.00139657 0.997815 0.796582 0.001069 0.00188153 0.000860305 0.455365 0.00188153 0.444947 0.000131468 1.02 0.888868 0.534348 0.287698 1.71971e-07 3.08635e-09 2369.33 3142.88 -0.0585787 0.482215 0.277249 0.255026 -0.593021 -0.169579 0.486428 -0.2656 -0.220838 2.751 1 0 295.005 0 2.24721 2.749 0.000299004 0.869695 0.70418 0.312119 0.436235 2.24738 139.831 83.5981 18.7022 60.7109 0.00403862 0 -40 10
1.85 5.35079e-08 2.54009e-06 0.150238 0.150238 0.0120251 2.43218e-05 0.00115458 0.187797 0.00065886 0.188452 0.959928 101.383 0.23399 0.86692 4.61693 0.0660104 0.0435559 0.956444 0.0193814 0.00464202 0.0186366 0.00442419 0.00561857 0.00636342 0.224743 0.254537 58.0552 -87.8995 126.137 15.9314 145.038 0.000142479 0.267334 192.711 0.31015 0.0673199 0.00409878 0.000562444 0.0013853 0.986957 0.991715 -2.99159e-06 -85.6561 0.0930938 31166.8 311.378 0.983496 0.319146 0.739111 0.739107 9.99958 2.98694e-06 1.19477e-05 0.134713 0.98343 0.931269 -0.0132915 4.93342e-06 0.517925 -2.02814e-20 7.52789e-24 -2.02739e-20 0.00139657 0.997814 8.60306e-05 0.152747 2.85288 0.00139657 0.997815 0.796653 0.00106902 0.00188154 0.000860306 0.455365 0.00188153 0.444952 0.00013147 1.02 0.888869 0.534348 0.287699 1.71971e-07 3.08637e-09 2369.31 3142.93 -0.0585838 0.482215 0.277249 0.255029 -0.593021 -0.169579 0.486412 -0.265598 -0.220824 2.752 1 0 295 0 2.24734 2.75 0.000299003 0.869725 0.704223 0.312081 0.436257 2.24752 139.838 83.5975 18.7022 60.7106 0.00403865 0 -40 10
1.851 5.35367e-08 2.54009e-06 0.150269 0.150268 0.0120251 2.43349e-05 0.00115459 0.187836 0.00065886 0.18849 0.960019 101.382 0.233979 0.867054 4.6176 0.0660213 0.0435622 0.956438 0.0193809 0.00464249 0.018636 0.00442459 0.00561915 0.00636402 0.224766 0.254561 58.0553 -87.8995 126.137 15.9314 145.038 0.000142482 0.267334 192.711 0.31015 0.0673198 0.00409878 0.000562445 0.00138531 0.986957 0.991715 -2.9916e-06 -85.6561 0.0930939 31166.8 311.391 0.983496 0.319146 0.739123 0.739119 9.99958 2.98695e-06 1.19477e-05 0.134718 0.983431 0.931268 -0.0132915 4.93345e-06 0.517946 -2.02831e-20 7.52855e-24 -2.02755e-20 0.00139657 0.997814 8.60307e-05 0.152747 2.85288 0.00139657 0.997815 0.796723 0.00106904 0.00188154 0.000860307 0.455365 0.00188154 0.444957 0.000131472 1.02 0.88887 0.534347 0.287701 1.71971e-07 3.0864e-09 2369.29 3142.98 -0.0585888 0.482215 0.277248 0.255033 -0.59302 -0.169579 0.486396 -0.265596 -0.22081 2.753 1 0 294.995 0 2.24748 2.751 0.000299002 0.869754 0.704265 0.312043 0.436279 2.24766 139.845 83.5969 18.7021 60.7103 0.00403867 0 -40 10
1.852 5.35656e-08 2.54009e-06 0.150299 0.150299 0.0120251 2.4348e-05 0.00115459 0.187874 0.000658861 0.188528 0.960111 101.382 0.233968 0.867188 4.61827 0.0660322 0.0435685 0.956431 0.0193803 0.00464297 0.0186354 0.004425 0.00561973 0.00636462 0.224789 0.254585 58.0553 -87.8995 126.137 15.9314 145.038 0.000142484 0.267334 192.711 0.31015 0.0673198 0.00409879 0.000562445 0.00138531 0.986957 0.991715 -2.99162e-06 -85.6561 0.093094 31166.8 311.404 0.983496 0.319146 0.739135 0.739131 9.99958 2.98695e-06 1.19477e-05 0.134723 0.983431 0.931267 -0.0132915 4.93348e-06 0.517967 -2.02847e-20 7.52921e-24 -2.02772e-20 0.00139657 0.997814 8.60308e-05 0.152747 2.85288 0.00139657 0.997815 0.796794 0.00106905 0.00188154 0.000860308 0.455364 0.00188154 0.444962 0.000131475 1.02 0.888871 0.534347 0.287702 1.71971e-07 3.08642e-09 2369.28 3143.03 -0.0585939 0.482215 0.277248 0.255036 -0.593019 -0.16958 0.48638 -0.265593 -0.220796 2.754 1 0 294.991 0 2.24761 2.752 0.000299001 0.869783 0.704308 0.312005 0.436301 2.24779 139.853 83.5963 18.7021 60.71 0.0040387 0 -40 10
1.853 5.35944e-08 2.54009e-06 0.15033 0.150329 0.0120251 2.43611e-05 0.00115459 0.187912 0.000658861 0.188566 0.960202 101.381 0.233957 0.867322 4.61893 0.066043 0.0435749 0.956425 0.0193797 0.00464344 0.0186348 0.00442541 0.00562031 0.00636522 0.224813 0.254609 58.0554 -87.8995 126.136 15.9313 145.038 0.000142486 0.267334 192.71 0.310149 0.0673197 0.00409879 0.000562446 0.00138531 0.986957 0.991715 -2.99163e-06 -85.6561 0.0930941 31166.8 311.417 0.983495 0.319146 0.739147 0.739143 9.99958 2.98696e-06 1.19477e-05 0.134728 0.983431 0.931265 -0.0132915 4.93351e-06 0.517987 -2.02864e-20 7.52986e-24 -2.02788e-20 0.00139657 0.997814 8.60309e-05 0.152747 2.85288 0.00139657 0.997815 0.796864 0.00106907 0.00188154 0.000860309 0.455364 0.00188154 0.444967 0.000131477 1.02 0.888872 0.534347 0.287704 1.71972e-07 3.08644e-09 2369.26 3143.08 -0.058599 0.482215 0.277248 0.255039 -0.593019 -0.16958 0.486364 -0.265591 -0.220782 2.755 1 0 294.986 0 2.24775 2.753 0.000298999 0.869813 0.704351 0.311967 0.436323 2.24793 139.86 83.5957 18.7021 60.7097 0.00403872 0 -40 10
1.854 5.36232e-08 2.54009e-06 0.15036 0.15036 0.012025 2.43742e-05 0.00115459 0.18795 0.000658861 0.188604 0.960293 101.38 0.233946 0.867456 4.6196 0.0660539 0.0435812 0.956419 0.0193791 0.00464391 0.0186342 0.00442582 0.0056209 0.00636583 0.224836 0.254633 58.0555 -87.8995 126.136 15.9313 145.038 0.000142489 0.267335 192.71 0.310149 0.0673197 0.00409879 0.000562447 0.00138531 0.986957 0.991715 -2.99165e-06 -85.6561 0.0930942 31166.7 311.43 0.983495 0.319146 0.739159 0.739155 9.99958 2.98696e-06 1.19477e-05 0.134733 0.983431 0.931264 -0.0132915 4.93354e-06 0.518008 -2.0288e-20 7.53052e-24 -2.02805e-20 0.00139657 0.997814 8.6031e-05 0.152747 2.85288 0.00139657 0.997815 0.796935 0.00106908 0.00188154 0.00086031 0.455364 0.00188154 0.444972 0.000131479 1.02 0.888873 0.534346 0.287705 1.71972e-07 3.08646e-09 2369.25 3143.13 -0.0586041 0.482215 0.277247 0.255042 -0.593018 -0.16958 0.486347 -0.265589 -0.220768 2.756 1 0 294.982 0 2.24789 2.754 0.000298998 0.869842 0.704393 0.311929 0.436345 2.24806 139.867 83.5951 18.702 60.7095 0.00403874 0 -40 10
1.855 5.36521e-08 2.54009e-06 0.150391 0.15039 0.012025 2.43873e-05 0.00115459 0.187988 0.000658862 0.188642 0.960385 101.38 0.233935 0.86759 4.62027 0.0660648 0.0435875 0.956413 0.0193785 0.00464438 0.0186336 0.00442623 0.00562148 0.00636643 0.224859 0.254657 58.0555 -87.8995 126.136 15.9312 145.038 0.000142491 0.267335 192.71 0.310148 0.0673196 0.0040988 0.000562447 0.00138532 0.986957 0.991715 -2.99167e-06 -85.6561 0.0930942 31166.7 311.442 0.983495 0.319146 0.739172 0.739167 9.99958 2.98697e-06 1.19478e-05 0.134737 0.983431 0.931263 -0.0132915 4.93357e-06 0.518028 -2.02896e-20 7.53118e-24 -2.02821e-20 0.00139657 0.997814 8.6031e-05 0.152748 2.85288 0.00139657 0.997815 0.797005 0.0010691 0.00188154 0.00086031 0.455364 0.00188154 0.444977 0.000131482 1.02 0.888874 0.534346 0.287707 1.71972e-07 3.08649e-09 2369.23 3143.19 -0.0586092 0.482215 0.277247 0.255046 -0.593018 -0.16958 0.486331 -0.265587 -0.220753 2.757 1 0 294.977 0 2.24802 2.755 0.000298997 0.869872 0.704436 0.311892 0.436367 2.2482 139.875 83.5945 18.702 60.7092 0.00403877 0 -40 10
1.856 5.36809e-08 2.5401e-06 0.150421 0.150421 0.012025 2.44004e-05 0.00115459 0.188026 0.000658862 0.188681 0.960476 101.379 0.233924 0.867724 4.62094 0.0660756 0.0435938 0.956406 0.0193779 0.00464486 0.018633 0.00442664 0.00562206 0.00636703 0.224883 0.254681 58.0556 -87.8995 126.136 15.9312 145.038 0.000142493 0.267335 192.71 0.310148 0.0673196 0.0040988 0.000562448 0.00138532 0.986957 0.991715 -2.99168e-06 -85.6561 0.0930943 31166.7 311.455 0.983495 0.319146 0.739184 0.739179 9.99958 2.98697e-06 1.19478e-05 0.134742 0.983432 0.931262 -0.0132915 4.9336e-06 0.518049 -2.02913e-20 7.53183e-24 -2.02838e-20 0.00139657 0.997814 8.60311e-05 0.152748 2.85288 0.00139657 0.997815 0.797075 0.00106912 0.00188154 0.000860311 0.455363 0.00188154 0.444982 0.000131484 1.02 0.888875 0.534346 0.287708 1.71973e-07 3.08651e-09 2369.21 3143.24 -0.0586143 0.482215 0.277247 0.255049 -0.593017 -0.16958 0.486315 -0.265585 -0.220739 2.758 1 0 294.972 0 2.24816 2.756 0.000298995 0.869901 0.704478 0.311854 0.436389 2.24834 139.882 83.5939 18.702 60.7089 0.00403879 0 -40 10
1.857 5.37097e-08 2.5401e-06 0.150451 0.150451 0.012025 2.44135e-05 0.00115459 0.188064 0.000658863 0.188719 0.960568 101.378 0.233913 0.867858 4.62161 0.0660865 0.0436001 0.9564 0.0193774 0.00464533 0.0186324 0.00442705 0.00562265 0.00636763 0.224906 0.254705 58.0557 -87.8995 126.135 15.9312 145.038 0.000142496 0.267335 192.71 0.310147 0.0673195 0.0040988 0.000562449 0.00138532 0.986957 0.991715 -2.9917e-06 -85.6561 0.0930944 31166.7 311.468 0.983495 0.319146 0.739196 0.739191 9.99958 2.98698e-06 1.19478e-05 0.134747 0.983432 0.931261 -0.0132915 4.93362e-06 0.51807 -2.02929e-20 7.53249e-24 -2.02854e-20 0.00139658 0.997814 8.60312e-05 0.152748 2.85288 0.00139658 0.997815 0.797146 0.00106913 0.00188155 0.000860312 0.455363 0.00188155 0.444987 0.000131486 1.02 0.888876 0.534345 0.28771 1.71973e-07 3.08653e-09 2369.2 3143.29 -0.0586194 0.482215 0.277247 0.255052 -0.593016 -0.16958 0.486299 -0.265583 -0.220725 2.759 1 0 294.968 0 2.24829 2.757 0.000298994 0.86993 0.704521 0.311816 0.436411 2.24847 139.889 83.5933 18.7019 60.7086 0.00403882 0 -40 10
1.858 5.37386e-08 2.5401e-06 0.150482 0.150481 0.012025 2.44266e-05 0.00115459 0.188102 0.000658863 0.188757 0.960659 101.378 0.233903 0.867991 4.62228 0.0660974 0.0436065 0.956394 0.0193768 0.0046458 0.0186318 0.00442746 0.00562323 0.00636824 0.224929 0.254729 58.0557 -87.8995 126.135 15.9311 145.038 0.000142498 0.267335 192.71 0.310147 0.0673195 0.0040988 0.000562449 0.00138532 0.986957 0.991715 -2.99171e-06 -85.656 0.0930945 31166.6 311.481 0.983495 0.319146 0.739208 0.739204 9.99958 2.98698e-06 1.19478e-05 0.134752 0.983432 0.93126 -0.0132915 4.93365e-06 0.51809 -2.02946e-20 7.53315e-24 -2.02871e-20 0.00139658 0.997814 8.60313e-05 0.152748 2.85288 0.00139658 0.997815 0.797216 0.00106915 0.00188155 0.000860313 0.455363 0.00188155 0.444992 0.000131489 1.02 0.888878 0.534345 0.287711 1.71973e-07 3.08656e-09 2369.18 3143.34 -0.0586245 0.482215 0.277246 0.255055 -0.593016 -0.16958 0.486283 -0.265581 -0.220711 2.76 1 0 294.963 0 2.24843 2.758 0.000298993 0.86996 0.704564 0.311778 0.436433 2.24861 139.897 83.5927 18.7019 60.7083 0.00403884 0 -40 10
1.859 5.37674e-08 2.5401e-06 0.150512 0.150512 0.012025 2.44397e-05 0.00115459 0.18814 0.000658864 0.188795 0.960751 101.377 0.233892 0.868125 4.62296 0.0661083 0.0436128 0.956387 0.0193762 0.00464628 0.0186312 0.00442787 0.00562381 0.00636884 0.224953 0.254754 58.0558 -87.8995 126.135 15.9311 145.038 0.0001425 0.267336 192.709 0.310147 0.0673194 0.00409881 0.00056245 0.00138532 0.986957 0.991715 -2.99173e-06 -85.656 0.0930946 31166.6 311.494 0.983495 0.319146 0.73922 0.739216 9.99958 2.98699e-06 1.19478e-05 0.134757 0.983432 0.931259 -0.0132914 4.93368e-06 0.518111 -2.02962e-20 7.53381e-24 -2.02887e-20 0.00139658 0.997814 8.60314e-05 0.152748 2.85289 0.00139658 0.997815 0.797286 0.00106916 0.00188155 0.000860314 0.455363 0.00188155 0.444997 0.000131491 1.02 0.888879 0.534345 0.287713 1.71973e-07 3.08658e-09 2369.16 3143.39 -0.0586296 0.482216 0.277246 0.255059 -0.593015 -0.16958 0.486267 -0.265579 -0.220697 2.761 1 0 294.959 0 2.24857 2.759 0.000298991 0.869989 0.704606 0.31174 0.436454 2.24874 139.904 83.5921 18.7018 60.708 0.00403887 0 -40 10
1.86 5.37962e-08 2.5401e-06 0.150543 0.150542 0.012025 2.44528e-05 0.00115459 0.188178 0.000658864 0.188832 0.960842 101.376 0.233881 0.868259 4.62363 0.0661191 0.0436191 0.956381 0.0193756 0.00464675 0.0186306 0.00442829 0.0056244 0.00636944 0.224976 0.254778 58.0558 -87.8995 126.135 15.9311 145.038 0.000142503 0.267336 192.709 0.310146 0.0673193 0.00409881 0.000562451 0.00138533 0.986957 0.991715 -2.99174e-06 -85.656 0.0930947 31166.6 311.507 0.983495 0.319146 0.739232 0.739228 9.99958 2.98699e-06 1.19479e-05 0.134761 0.983432 0.931258 -0.0132914 4.93371e-06 0.518132 -2.02979e-20 7.53447e-24 -2.02904e-20 0.00139658 0.997814 8.60314e-05 0.152748 2.85289 0.00139658 0.997815 0.797357 0.00106918 0.00188155 0.000860314 0.455363 0.00188155 0.445002 0.000131493 1.02 0.88888 0.534344 0.287714 1.71974e-07 3.0866e-09 2369.15 3143.44 -0.0586347 0.482216 0.277246 0.255062 -0.593014 -0.16958 0.48625 -0.265577 -0.220683 2.762 1 0 294.954 0 2.2487 2.76 0.00029899 0.870019 0.704649 0.311702 0.436476 2.24888 139.911 83.5915 18.7018 60.7077 0.00403889 0 -40 10
1.861 5.38251e-08 2.5401e-06 0.150573 0.150572 0.0120249 2.44659e-05 0.00115459 0.188216 0.000658865 0.18887 0.960934 101.376 0.23387 0.868393 4.6243 0.06613 0.0436255 0.956375 0.019375 0.00464723 0.01863 0.0044287 0.00562498 0.00637005 0.224999 0.254802 58.0559 -87.8995 126.135 15.931 145.038 0.000142505 0.267336 192.709 0.310146 0.0673193 0.00409881 0.000562451 0.00138533 0.986957 0.991714 -2.99176e-06 -85.656 0.0930948 31166.6 311.52 0.983495 0.319146 0.739244 0.73924 9.99958 2.987e-06 1.19479e-05 0.134766 0.983433 0.931257 -0.0132914 4.93374e-06 0.518152 -2.02995e-20 7.53512e-24 -2.0292e-20 0.00139658 0.997814 8.60315e-05 0.152749 2.85289 0.00139658 0.997815 0.797427 0.00106919 0.00188155 0.000860315 0.455362 0.00188155 0.445007 0.000131496 1.02 0.888881 0.534344 0.287716 1.71974e-07 3.08662e-09 2369.13 3143.49 -0.0586397 0.482216 0.277246 0.255065 -0.593014 -0.16958 0.486234 -0.265575 -0.220669 2.763 1 0 294.949 0 2.24884 2.761 0.000298989 0.870048 0.704692 0.311665 0.436498 2.24902 139.919 83.5909 18.7018 60.7074 0.00403892 0 -40 10
1.862 5.38539e-08 2.54011e-06 0.150603 0.150603 0.0120249 2.4479e-05 0.00115459 0.188254 0.000658865 0.188908 0.961025 101.375 0.233859 0.868527 4.62497 0.0661409 0.0436318 0.956368 0.0193744 0.0046477 0.0186293 0.00442911 0.00562557 0.00637065 0.225023 0.254826 58.056 -87.8995 126.134 15.931 145.038 0.000142507 0.267336 192.709 0.310145 0.0673192 0.00409882 0.000562452 0.00138533 0.986957 0.991714 -2.99177e-06 -85.656 0.0930949 31166.5 311.533 0.983495 0.319146 0.739257 0.739252 9.99958 2.987e-06 1.19479e-05 0.134771 0.983433 0.931256 -0.0132914 4.93377e-06 0.518173 -2.03012e-20 7.53578e-24 -2.02937e-20 0.00139658 0.997814 8.60316e-05 0.152749 2.85289 0.00139658 0.997815 0.797497 0.00106921 0.00188155 0.000860316 0.455362 0.00188155 0.445012 0.000131498 1.02 0.888882 0.534344 0.287717 1.71974e-07 3.08665e-09 2369.12 3143.54 -0.0586448 0.482216 0.277245 0.255069 -0.593013 -0.16958 0.486218 -0.265573 -0.220655 2.764 1 0 294.945 0 2.24897 2.762 0.000298988 0.870078 0.704734 0.311627 0.43652 2.24915 139.926 83.5903 18.7017 60.7072 0.00403894 0 -40 10
1.863 5.38827e-08 2.54011e-06 0.150633 0.150633 0.0120249 2.44922e-05 0.00115459 0.188292 0.000658866 0.188946 0.961117 101.374 0.233848 0.868661 4.62565 0.0661518 0.0436382 0.956362 0.0193738 0.00464817 0.0186287 0.00442952 0.00562615 0.00637125 0.225046 0.25485 58.056 -87.8996 126.134 15.9309 145.038 0.00014251 0.267336 192.709 0.310145 0.0673192 0.00409882 0.000562453 0.00138533 0.986957 0.991714 -2.99179e-06 -85.656 0.0930949 31166.5 311.546 0.983495 0.319146 0.739269 0.739264 9.99958 2.98701e-06 1.19479e-05 0.134776 0.983433 0.931255 -0.0132914 4.9338e-06 0.518194 -2.03028e-20 7.53644e-24 -2.02953e-20 0.00139658 0.997814 8.60317e-05 0.152749 2.85289 0.00139658 0.997815 0.797567 0.00106923 0.00188156 0.000860317 0.455362 0.00188155 0.445017 0.0001315 1.02 0.888883 0.534344 0.287719 1.71974e-07 3.08667e-09 2369.1 3143.59 -0.0586499 0.482216 0.277245 0.255072 -0.593012 -0.16958 0.486202 -0.26557 -0.220641 2.765 1 0 294.94 0 2.24911 2.763 0.000298986 0.870107 0.704777 0.311589 0.436542 2.24929 139.933 83.5897 18.7017 60.7069 0.00403897 0 -40 10
1.864 5.39116e-08 2.54011e-06 0.150664 0.150663 0.0120249 2.45053e-05 0.0011546 0.18833 0.000658866 0.188984 0.961209 101.374 0.233837 0.868795 4.62632 0.0661626 0.0436445 0.956355 0.0193733 0.00464865 0.0186281 0.00442993 0.00562674 0.00637186 0.22507 0.254874 58.0561 -87.8996 126.134 15.9309 145.038 0.000142512 0.267336 192.709 0.310144 0.0673191 0.00409882 0.000562453 0.00138534 0.986957 0.991714 -2.9918e-06 -85.656 0.093095 31166.5 311.558 0.983495 0.319146 0.739281 0.739276 9.99958 2.98701e-06 1.19479e-05 0.134781 0.983433 0.931254 -0.0132914 4.93383e-06 0.518214 -2.03045e-20 7.5371e-24 -2.0297e-20 0.00139658 0.997814 8.60318e-05 0.152749 2.85289 0.00139658 0.997815 0.797638 0.00106924 0.00188156 0.000860318 0.455362 0.00188156 0.445022 0.000131503 1.02 0.888884 0.534343 0.28772 1.71975e-07 3.08669e-09 2369.08 3143.64 -0.058655 0.482216 0.277245 0.255075 -0.593012 -0.16958 0.486186 -0.265568 -0.220627 2.766 1 0 294.936 0 2.24925 2.764 0.000298985 0.870137 0.704819 0.311552 0.436564 2.24942 139.94 83.5891 18.7017 60.7066 0.00403899 0 -40 10
1.865 5.39404e-08 2.54011e-06 0.150694 0.150693 0.0120249 2.45184e-05 0.0011546 0.188367 0.000658867 0.189022 0.9613 101.373 0.233826 0.868929 4.62699 0.0661735 0.0436509 0.956349 0.0193727 0.00464912 0.0186275 0.00443034 0.00562732 0.00637246 0.225093 0.254899 58.0562 -87.8996 126.134 15.9309 145.038 0.000142514 0.267337 192.709 0.310144 0.0673191 0.00409883 0.000562454 0.00138534 0.986957 0.991714 -2.99182e-06 -85.656 0.0930951 31166.5 311.571 0.983495 0.319146 0.739293 0.739289 9.99958 2.98702e-06 1.1948e-05 0.134786 0.983433 0.931253 -0.0132914 4.93386e-06 0.518235 -2.03061e-20 7.53776e-24 -2.02986e-20 0.00139659 0.997814 8.60318e-05 0.152749 2.85289 0.00139659 0.997815 0.797708 0.00106926 0.00188156 0.000860318 0.455361 0.00188156 0.445027 0.000131505 1.02 0.888885 0.534343 0.287722 1.71975e-07 3.08672e-09 2369.07 3143.69 -0.0586601 0.482216 0.277244 0.255078 -0.593011 -0.16958 0.486169 -0.265566 -0.220613 2.767 1 0 294.931 0 2.24938 2.765 0.000298984 0.870166 0.704862 0.311514 0.436586 2.24956 139.948 83.5885 18.7016 60.7063 0.00403902 0 -40 10
1.866 5.39692e-08 2.54011e-06 0.150724 0.150724 0.0120249 2.45315e-05 0.0011546 0.188405 0.000658867 0.189059 0.961392 101.372 0.233816 0.869063 4.62767 0.0661844 0.0436572 0.956343 0.0193721 0.0046496 0.0186269 0.00443075 0.00562791 0.00637307 0.225116 0.254923 58.0562 -87.8996 126.134 15.9308 145.038 0.000142517 0.267337 192.708 0.310144 0.067319 0.00409883 0.000562455 0.00138534 0.986957 0.991714 -2.99183e-06 -85.656 0.0930952 31166.5 311.584 0.983495 0.319146 0.739305 0.739301 9.99958 2.98702e-06 1.1948e-05 0.13479 0.983434 0.931252 -0.0132914 4.93389e-06 0.518256 -2.03078e-20 7.53842e-24 -2.03003e-20 0.00139659 0.997814 8.60319e-05 0.152749 2.85289 0.00139659 0.997815 0.797778 0.00106927 0.00188156 0.000860319 0.455361 0.00188156 0.445031 0.000131507 1.02 0.888886 0.534343 0.287723 1.71975e-07 3.08674e-09 2369.05 3143.74 -0.0586652 0.482216 0.277244 0.255082 -0.593011 -0.16958 0.486153 -0.265564 -0.220599 2.768 1 0 294.927 0 2.24952 2.766 0.000298982 0.870195 0.704905 0.311476 0.436608 2.2497 139.955 83.5879 18.7016 60.706 0.00403904 0 -40 10
1.867 5.39981e-08 2.54012e-06 0.150754 0.150754 0.0120249 2.45446e-05 0.0011546 0.188443 0.000658867 0.189097 0.961483 101.372 0.233805 0.869197 4.62834 0.0661953 0.0436636 0.956336 0.0193715 0.00465007 0.0186263 0.00443117 0.0056285 0.00637367 0.22514 0.254947 58.0563 -87.8996 126.133 15.9308 145.038 0.000142519 0.267337 192.708 0.310143 0.067319 0.00409883 0.000562455 0.00138534 0.986957 0.991714 -2.99185e-06 -85.656 0.0930953 31166.4 311.597 0.983495 0.319146 0.739317 0.739313 9.99958 2.98703e-06 1.1948e-05 0.134795 0.983434 0.931251 -0.0132914 4.93392e-06 0.518276 -2.03095e-20 7.53908e-24 -2.03019e-20 0.00139659 0.997814 8.6032e-05 0.152749 2.85289 0.00139659 0.997815 0.797848 0.00106929 0.00188156 0.00086032 0.455361 0.00188156 0.445036 0.00013151 1.02 0.888887 0.534342 0.287725 1.71976e-07 3.08676e-09 2369.03 3143.8 -0.0586703 0.482216 0.277244 0.255085 -0.59301 -0.16958 0.486137 -0.265562 -0.220584 2.769 1 0 294.922 0 2.24965 2.767 0.000298981 0.870225 0.704947 0.311439 0.43663 2.24983 139.962 83.5874 18.7016 60.7057 0.00403907 0 -40 10
1.868 5.40269e-08 2.54012e-06 0.150784 0.150784 0.0120248 2.45577e-05 0.0011546 0.188481 0.000658868 0.189135 0.961575 101.371 0.233794 0.869331 4.62902 0.0662062 0.04367 0.95633 0.0193709 0.00465055 0.0186257 0.00443158 0.00562908 0.00637428 0.225163 0.254971 58.0563 -87.8996 126.133 15.9308 145.038 0.000142521 0.267337 192.708 0.310143 0.0673189 0.00409883 0.000562456 0.00138534 0.986957 0.991714 -2.99186e-06 -85.656 0.0930954 31166.4 311.61 0.983495 0.319146 0.739329 0.739325 9.99958 2.98703e-06 1.1948e-05 0.1348 0.983434 0.93125 -0.0132914 4.93395e-06 0.518297 -2.03111e-20 7.53974e-24 -2.03036e-20 0.00139659 0.997814 8.60321e-05 0.15275 2.85289 0.00139659 0.997815 0.797918 0.00106931 0.00188156 0.000860321 0.455361 0.00188156 0.445041 0.000131512 1.02 0.888889 0.534342 0.287726 1.71976e-07 3.08678e-09 2369.02 3143.85 -0.0586754 0.482216 0.277244 0.255088 -0.593009 -0.169581 0.486121 -0.26556 -0.22057 2.77 1 0 294.917 0 2.24979 2.768 0.00029898 0.870254 0.70499 0.311401 0.436652 2.24997 139.97 83.5868 18.7015 60.7054 0.00403909 0 -40 10
1.869 5.40557e-08 2.54012e-06 0.150815 0.150814 0.0120248 2.45708e-05 0.0011546 0.188518 0.000658868 0.189172 0.961666 101.37 0.233783 0.869465 4.62969 0.0662171 0.0436764 0.956324 0.0193703 0.00465102 0.0186251 0.00443199 0.00562967 0.00637488 0.225187 0.254995 58.0564 -87.8996 126.133 15.9307 145.038 0.000142524 0.267337 192.708 0.310142 0.0673189 0.00409884 0.000562457 0.00138535 0.986956 0.991714 -2.99188e-06 -85.6559 0.0930955 31166.4 311.623 0.983495 0.319146 0.739342 0.739337 9.99958 2.98704e-06 1.1948e-05 0.134805 0.983434 0.931249 -0.0132914 4.93398e-06 0.518318 -2.03128e-20 7.5404e-24 -2.03052e-20 0.00139659 0.997814 8.60322e-05 0.15275 2.85289 0.00139659 0.997815 0.797988 0.00106932 0.00188156 0.000860322 0.455361 0.00188156 0.445046 0.000131514 1.02 0.88889 0.534342 0.287728 1.71976e-07 3.08681e-09 2369 3143.9 -0.0586805 0.482216 0.277243 0.255091 -0.593009 -0.169581 0.486105 -0.265558 -0.220556 2.771 1 0 294.913 0 2.24993 2.769 0.000298978 0.870284 0.705032 0.311364 0.436674 2.2501 139.977 83.5862 18.7015 60.7051 0.00403912 0 -40 10
1.87 5.40846e-08 2.54012e-06 0.150845 0.150844 0.0120248 2.45839e-05 0.0011546 0.188556 0.000658869 0.18921 0.961758 101.37 0.233772 0.869599 4.63037 0.0662279 0.0436827 0.956317 0.0193697 0.0046515 0.0186245 0.0044324 0.00563025 0.00637549 0.22521 0.25502 58.0565 -87.8996 126.133 15.9307 145.038 0.000142526 0.267338 192.708 0.310142 0.0673188 0.00409884 0.000562458 0.00138535 0.986956 0.991714 -2.99189e-06 -85.6559 0.0930956 31166.4 311.636 0.983495 0.319146 0.739354 0.739349 9.99958 2.98704e-06 1.19481e-05 0.13481 0.983434 0.931248 -0.0132914 4.93401e-06 0.518339 -2.03144e-20 7.54107e-24 -2.03069e-20 0.00139659 0.997814 8.60322e-05 0.15275 2.8529 0.00139659 0.997815 0.798058 0.00106934 0.00188157 0.000860322 0.45536 0.00188156 0.445051 0.000131517 1.02 0.888891 0.534341 0.287729 1.71976e-07 3.08683e-09 2368.98 3143.95 -0.0586856 0.482216 0.277243 0.255095 -0.593008 -0.169581 0.486089 -0.265556 -0.220542 2.772 1 0 294.908 0 2.25006 2.77 0.000298977 0.870314 0.705075 0.311326 0.436696 2.25024 139.984 83.5856 18.7015 60.7049 0.00403914 0 -40 10
1.871 5.41134e-08 2.54012e-06 0.150875 0.150874 0.0120248 2.4597e-05 0.0011546 0.188593 0.000658869 0.189248 0.96185 101.369 0.233761 0.869734 4.63105 0.0662388 0.0436891 0.956311 0.0193692 0.00465198 0.0186239 0.00443282 0.00563084 0.0063761 0.225234 0.255044 58.0565 -87.8996 126.132 15.9307 145.038 0.000142528 0.267338 192.708 0.310141 0.0673188 0.00409884 0.000562458 0.00138535 0.986956 0.991714 -2.99191e-06 -85.6559 0.0930956 31166.3 311.649 0.983495 0.319146 0.739366 0.739361 9.99958 2.98705e-06 1.19481e-05 0.134815 0.983435 0.931247 -0.0132914 4.93404e-06 0.518359 -2.03161e-20 7.54173e-24 -2.03085e-20 0.00139659 0.997814 8.60323e-05 0.15275 2.8529 0.00139659 0.997815 0.798128 0.00106935 0.00188157 0.000860323 0.45536 0.00188157 0.445056 0.000131519 1.02 0.888892 0.534341 0.287731 1.71977e-07 3.08685e-09 2368.97 3144 -0.0586907 0.482216 0.277243 0.255098 -0.593007 -0.169581 0.486072 -0.265554 -0.220528 2.773 1 0 294.904 0 2.2502 2.771 0.000298976 0.870343 0.705118 0.311289 0.436718 2.25038 139.992 83.585 18.7014 60.7046 0.00403917 0 -40 10
1.872 5.41422e-08 2.54012e-06 0.150905 0.150904 0.0120248 2.46101e-05 0.0011546 0.188631 0.00065887 0.189285 0.961941 101.368 0.23375 0.869868 4.63172 0.0662497 0.0436955 0.956304 0.0193686 0.00465245 0.0186233 0.00443323 0.00563143 0.0063767 0.225257 0.255068 58.0566 -87.8996 126.132 15.9306 145.038 0.000142531 0.267338 192.707 0.310141 0.0673187 0.00409885 0.000562459 0.00138535 0.986956 0.991714 -2.99192e-06 -85.6559 0.0930957 31166.3 311.662 0.983495 0.319146 0.739378 0.739374 9.99958 2.98705e-06 1.19481e-05 0.134819 0.983435 0.931246 -0.0132914 4.93407e-06 0.51838 -2.03177e-20 7.54239e-24 -2.03102e-20 0.00139659 0.997814 8.60324e-05 0.15275 2.8529 0.00139659 0.997815 0.798198 0.00106937 0.00188157 0.000860324 0.45536 0.00188157 0.445061 0.000131521 1.02 0.888893 0.534341 0.287732 1.71977e-07 3.08688e-09 2368.95 3144.05 -0.0586958 0.482216 0.277242 0.255101 -0.593007 -0.169581 0.486056 -0.265552 -0.220514 2.774 1 0 294.899 0 2.25033 2.772 0.000298974 0.870373 0.70516 0.311251 0.43674 2.25051 139.999 83.5844 18.7014 60.7043 0.00403919 0 -40 10
1.873 5.41711e-08 2.54013e-06 0.150935 0.150934 0.0120248 2.46232e-05 0.0011546 0.188669 0.00065887 0.189323 0.962033 101.368 0.233739 0.870002 4.6324 0.0662606 0.0437019 0.956298 0.019368 0.00465293 0.0186227 0.00443364 0.00563202 0.00637731 0.225281 0.255092 58.0567 -87.8996 126.132 15.9306 145.038 0.000142533 0.267338 192.707 0.310141 0.0673187 0.00409885 0.00056246 0.00138535 0.986956 0.991714 -2.99194e-06 -85.6559 0.0930958 31166.3 311.675 0.983495 0.319146 0.73939 0.739386 9.99958 2.98706e-06 1.19481e-05 0.134824 0.983435 0.931245 -0.0132914 4.9341e-06 0.518401 -2.03194e-20 7.54305e-24 -2.03119e-20 0.00139659 0.997814 8.60325e-05 0.15275 2.8529 0.00139659 0.997815 0.798268 0.00106939 0.00188157 0.000860325 0.45536 0.00188157 0.445066 0.000131524 1.02 0.888894 0.534341 0.287734 1.71977e-07 3.0869e-09 2368.94 3144.1 -0.0587009 0.482217 0.277242 0.255104 -0.593006 -0.169581 0.48604 -0.265549 -0.2205 2.775 1 0 294.894 0 2.25047 2.773 0.000298973 0.870402 0.705203 0.311214 0.436762 2.25065 140.006 83.5838 18.7014 60.704 0.00403921 0 -40 10
1.874 5.41999e-08 2.54013e-06 0.150965 0.150964 0.0120248 2.46363e-05 0.0011546 0.188706 0.000658871 0.18936 0.962125 101.367 0.233729 0.870136 4.63308 0.0662715 0.0437083 0.956292 0.0193674 0.0046534 0.0186221 0.00443405 0.0056326 0.00637792 0.225304 0.255117 58.0567 -87.8996 126.132 15.9305 145.038 0.000142535 0.267338 192.707 0.31014 0.0673186 0.00409885 0.00056246 0.00138536 0.986956 0.991714 -2.99195e-06 -85.6559 0.0930959 31166.3 311.688 0.983495 0.319146 0.739402 0.739398 9.99958 2.98706e-06 1.19481e-05 0.134829 0.983435 0.931244 -0.0132914 4.93413e-06 0.518422 -2.03211e-20 7.54371e-24 -2.03135e-20 0.0013966 0.997814 8.60326e-05 0.152751 2.8529 0.0013966 0.997815 0.798338 0.0010694 0.00188157 0.000860326 0.455359 0.00188157 0.445071 0.000131526 1.02 0.888895 0.53434 0.287735 1.71977e-07 3.08692e-09 2368.92 3144.15 -0.058706 0.482217 0.277242 0.255108 -0.593005 -0.169581 0.486024 -0.265547 -0.220486 2.776 1 0 294.89 0 2.25061 2.774 0.000298972 0.870432 0.705245 0.311176 0.436784 2.25078 140.013 83.5832 18.7013 60.7037 0.00403924 0 -40 10
1.875 5.42287e-08 2.54013e-06 0.150995 0.150994 0.0120247 2.46494e-05 0.0011546 0.188743 0.000658871 0.189398 0.962217 101.366 0.233718 0.87027 4.63376 0.0662824 0.0437147 0.956285 0.0193668 0.00465388 0.0186215 0.00443447 0.00563319 0.00637852 0.225328 0.255141 58.0568 -87.8996 126.132 15.9305 145.038 0.000142538 0.267339 192.707 0.31014 0.0673186 0.00409886 0.000562461 0.00138536 0.986956 0.991714 -2.99197e-06 -85.6559 0.093096 31166.3 311.701 0.983495 0.319146 0.739414 0.73941 9.99958 2.98707e-06 1.19482e-05 0.134834 0.983435 0.931243 -0.0132914 4.93416e-06 0.518443 -2.03227e-20 7.54438e-24 -2.03152e-20 0.0013966 0.997814 8.60326e-05 0.152751 2.8529 0.0013966 0.997815 0.798408 0.00106942 0.00188157 0.000860326 0.455359 0.00188157 0.445076 0.000131528 1.02 0.888896 0.53434 0.287737 1.71978e-07 3.08695e-09 2368.9 3144.2 -0.0587111 0.482217 0.277242 0.255111 -0.593005 -0.169581 0.486008 -0.265545 -0.220472 2.777 1 0 294.885 0 2.25074 2.775 0.00029897 0.870461 0.705288 0.311139 0.436805 2.25092 140.021 83.5826 18.7013 60.7034 0.00403926 0 -40 10
1.876 5.42576e-08 2.54013e-06 0.151025 0.151024 0.0120247 2.46625e-05 0.00115461 0.188781 0.000658872 0.189435 0.962308 101.366 0.233707 0.870404 4.63444 0.0662933 0.0437211 0.956279 0.0193662 0.00465436 0.0186209 0.00443488 0.00563378 0.00637913 0.225351 0.255165 58.0568 -87.8996 126.131 15.9305 145.038 0.00014254 0.267339 192.707 0.310139 0.0673185 0.00409886 0.000562462 0.00138536 0.986956 0.991714 -2.99198e-06 -85.6559 0.0930961 31166.2 311.714 0.983495 0.319146 0.739427 0.739422 9.99958 2.98707e-06 1.19482e-05 0.134839 0.983436 0.931242 -0.0132914 4.93419e-06 0.518463 -2.03244e-20 7.54504e-24 -2.03168e-20 0.0013966 0.997814 8.60327e-05 0.152751 2.8529 0.0013966 0.997815 0.798478 0.00106943 0.00188157 0.000860327 0.455359 0.00188157 0.445081 0.000131531 1.02 0.888897 0.53434 0.287738 1.71978e-07 3.08697e-09 2368.89 3144.25 -0.0587162 0.482217 0.277241 0.255114 -0.593004 -0.169581 0.485991 -0.265543 -0.220458 2.778 1 0 294.881 0 2.25088 2.776 0.000298969 0.870491 0.705331 0.311102 0.436827 2.25106 140.028 83.582 18.7013 60.7031 0.00403929 0 -40 10
1.877 5.42864e-08 2.54013e-06 0.151055 0.151054 0.0120247 2.46756e-05 0.00115461 0.188818 0.000658872 0.189473 0.9624 101.365 0.233696 0.870538 4.63512 0.0663042 0.0437275 0.956272 0.0193656 0.00465484 0.0186203 0.00443529 0.00563437 0.00637974 0.225375 0.25519 58.0569 -87.8996 126.131 15.9304 145.038 0.000142542 0.267339 192.707 0.310139 0.0673185 0.00409886 0.000562462 0.00138536 0.986956 0.991714 -2.992e-06 -85.6559 0.0930962 31166.2 311.727 0.983495 0.319146 0.739439 0.739434 9.99958 2.98708e-06 1.19482e-05 0.134844 0.983436 0.931241 -0.0132914 4.93422e-06 0.518484 -2.0326e-20 7.5457e-24 -2.03185e-20 0.0013966 0.997814 8.60328e-05 0.152751 2.8529 0.0013966 0.997815 0.798548 0.00106945 0.00188158 0.000860328 0.455359 0.00188157 0.445085 0.000131533 1.02 0.888898 0.534339 0.28774 1.71978e-07 3.08699e-09 2368.87 3144.31 -0.0587213 0.482217 0.277241 0.255117 -0.593003 -0.169581 0.485975 -0.265541 -0.220443 2.779 1 0 294.876 0 2.25101 2.777 0.000298968 0.87052 0.705373 0.311064 0.436849 2.25119 140.035 83.5814 18.7012 60.7028 0.00403931 0 -40 10
1.878 5.43152e-08 2.54014e-06 0.151085 0.151084 0.0120247 2.46887e-05 0.00115461 0.188856 0.000658872 0.18951 0.962492 101.364 0.233685 0.870672 4.6358 0.0663151 0.0437339 0.956266 0.019365 0.00465531 0.0186197 0.00443571 0.00563496 0.00638035 0.225398 0.255214 58.057 -87.8996 126.131 15.9304 145.038 0.000142545 0.267339 192.706 0.310138 0.0673184 0.00409887 0.000562463 0.00138537 0.986956 0.991714 -2.99201e-06 -85.6559 0.0930963 31166.2 311.74 0.983495 0.319146 0.739451 0.739447 9.99958 2.98708e-06 1.19482e-05 0.134849 0.983436 0.93124 -0.0132914 4.93425e-06 0.518505 -2.03277e-20 7.54636e-24 -2.03202e-20 0.0013966 0.997814 8.60329e-05 0.152751 2.8529 0.0013966 0.997815 0.798617 0.00106946 0.00188158 0.000860329 0.455358 0.00188158 0.44509 0.000131535 1.02 0.8889 0.534339 0.287742 1.71979e-07 3.08701e-09 2368.85 3144.36 -0.0587264 0.482217 0.277241 0.255121 -0.593003 -0.169581 0.485959 -0.265539 -0.220429 2.78 1 0 294.871 0 2.25115 2.778 0.000298967 0.87055 0.705416 0.311027 0.436871 2.25133 140.043 83.5808 18.7012 60.7025 0.00403934 0 -40 10
1.879 5.4344e-08 2.54014e-06 0.151114 0.151114 0.0120247 2.47018e-05 0.00115461 0.188893 0.000658873 0.189547 0.962583 101.364 0.233674 0.870806 4.63648 0.066326 0.0437404 0.95626 0.0193645 0.00465579 0.018619 0.00443612 0.00563554 0.00638096 0.225422 0.255238 58.057 -87.8996 126.131 15.9304 145.038 0.000142547 0.267339 192.706 0.310138 0.0673183 0.00409887 0.000562464 0.00138537 0.986956 0.991714 -2.99203e-06 -85.6558 0.0930963 31166.2 311.753 0.983495 0.319146 0.739463 0.739459 9.99958 2.98709e-06 1.19482e-05 0.134853 0.983436 0.931239 -0.0132914 4.93428e-06 0.518526 -2.03294e-20 7.54703e-24 -2.03218e-20 0.0013966 0.997814 8.6033e-05 0.152751 2.8529 0.0013966 0.997815 0.798687 0.00106948 0.00188158 0.00086033 0.455358 0.00188158 0.445095 0.000131538 1.02 0.888901 0.534339 0.287743 1.71979e-07 3.08704e-09 2368.84 3144.41 -0.0587315 0.482217 0.27724 0.255124 -0.593002 -0.169581 0.485943 -0.265537 -0.220415 2.781 1 0 294.867 0 2.25129 2.779 0.000298965 0.87058 0.705458 0.31099 0.436893 2.25146 140.05 83.5802 18.7012 60.7023 0.00403936 0 -40 10
1.88 5.43729e-08 2.54014e-06 0.151144 0.151144 0.0120247 2.47149e-05 0.00115461 0.18893 0.000658873 0.189585 0.962675 101.363 0.233663 0.870941 4.63716 0.0663369 0.0437468 0.956253 0.0193639 0.00465627 0.0186184 0.00443654 0.00563613 0.00638156 0.225445 0.255263 58.0571 -87.8996 126.13 15.9303 145.038 0.000142549 0.26734 192.706 0.310138 0.0673183 0.00409887 0.000562464 0.00138537 0.986956 0.991714 -2.99204e-06 -85.6558 0.0930964 31166.1 311.766 0.983495 0.319146 0.739475 0.739471 9.99958 2.98709e-06 1.19483e-05 0.134858 0.983436 0.931238 -0.0132914 4.93431e-06 0.518547 -2.0331e-20 7.54769e-24 -2.03235e-20 0.0013966 0.997814 8.6033e-05 0.152751 2.8529 0.0013966 0.997815 0.798757 0.0010695 0.00188158 0.00086033 0.455358 0.00188158 0.4451 0.00013154 1.02 0.888902 0.534338 0.287745 1.71979e-07 3.08706e-09 2368.82 3144.46 -0.0587366 0.482217 0.27724 0.255127 -0.593002 -0.169581 0.485927 -0.265535 -0.220401 2.782 1 0 294.862 0 2.25142 2.78 0.000298964 0.870609 0.705501 0.310952 0.436915 2.2516 140.057 83.5796 18.7011 60.702 0.00403939 0 -40 10
1.881 5.44017e-08 2.54014e-06 0.151174 0.151174 0.0120247 2.4728e-05 0.00115461 0.188968 0.000658874 0.189622 0.962767 101.362 0.233652 0.871075 4.63784 0.0663478 0.0437532 0.956247 0.0193633 0.00465674 0.0186178 0.00443695 0.00563672 0.00638217 0.225469 0.255287 58.0572 -87.8996 126.13 15.9303 145.038 0.000142552 0.26734 192.706 0.310137 0.0673182 0.00409887 0.000562465 0.00138537 0.986956 0.991714 -2.99206e-06 -85.6558 0.0930965 31166.1 311.779 0.983495 0.319146 0.739487 0.739483 9.99958 2.9871e-06 1.19483e-05 0.134863 0.983436 0.931237 -0.0132914 4.93434e-06 0.518568 -2.03327e-20 7.54835e-24 -2.03251e-20 0.0013966 0.997814 8.60331e-05 0.152752 2.85291 0.0013966 0.997815 0.798827 0.00106951 0.00188158 0.000860331 0.455358 0.00188158 0.445105 0.000131542 1.02 0.888903 0.534338 0.287746 1.71979e-07 3.08708e-09 2368.81 3144.51 -0.0587417 0.482217 0.27724 0.255131 -0.593001 -0.169581 0.48591 -0.265533 -0.220387 2.783 1 0 294.858 0 2.25156 2.781 0.000298963 0.870639 0.705543 0.310915 0.436937 2.25173 140.065 83.579 18.7011 60.7017 0.00403941 0 -40 10
1.882 5.44305e-08 2.54014e-06 0.151204 0.151204 0.0120246 2.47412e-05 0.00115461 0.189005 0.000658874 0.189659 0.962859 101.361 0.233641 0.871209 4.63852 0.0663587 0.0437596 0.95624 0.0193627 0.00465722 0.0186172 0.00443737 0.00563731 0.00638278 0.225492 0.255311 58.0572 -87.8996 126.13 15.9302 145.038 0.000142554 0.26734 192.706 0.310137 0.0673182 0.00409888 0.000562466 0.00138537 0.986956 0.991714 -2.99207e-06 -85.6558 0.0930966 31166.1 311.792 0.983495 0.319146 0.7395 0.739495 9.99958 2.9871e-06 1.19483e-05 0.134868 0.983437 0.931236 -0.0132914 4.93437e-06 0.518588 -2.03344e-20 7.54902e-24 -2.03268e-20 0.0013966 0.997814 8.60332e-05 0.152752 2.85291 0.0013966 0.997815 0.798897 0.00106953 0.00188158 0.000860332 0.455358 0.00188158 0.44511 0.000131545 1.02 0.888904 0.534338 0.287748 1.7198e-07 3.08711e-09 2368.79 3144.56 -0.0587468 0.482217 0.27724 0.255134 -0.593 -0.169581 0.485894 -0.265531 -0.220373 2.784 1 0 294.853 0 2.25169 2.782 0.000298961 0.870668 0.705586 0.310878 0.436959 2.25187 140.072 83.5784 18.701 60.7014 0.00403944 0 -40 10
1.883 5.44594e-08 2.54014e-06 0.151234 0.151233 0.0120246 2.47543e-05 0.00115461 0.189042 0.000658875 0.189696 0.962951 101.361 0.23363 0.871343 4.6392 0.0663696 0.0437661 0.956234 0.0193621 0.0046577 0.0186166 0.00443778 0.0056379 0.00638339 0.225516 0.255336 58.0573 -87.8996 126.13 15.9302 145.038 0.000142556 0.26734 192.706 0.310136 0.0673181 0.00409888 0.000562466 0.00138538 0.986956 0.991714 -2.99209e-06 -85.6558 0.0930967 31166.1 311.805 0.983495 0.319146 0.739512 0.739507 9.99958 2.98711e-06 1.19483e-05 0.134873 0.983437 0.931235 -0.0132914 4.93439e-06 0.518609 -2.0336e-20 7.54968e-24 -2.03285e-20 0.00139661 0.997814 8.60333e-05 0.152752 2.85291 0.00139661 0.997815 0.798966 0.00106954 0.00188159 0.000860333 0.455357 0.00188158 0.445115 0.000131547 1.02 0.888905 0.534337 0.287749 1.7198e-07 3.08713e-09 2368.77 3144.61 -0.0587519 0.482217 0.277239 0.255137 -0.593 -0.169581 0.485878 -0.265529 -0.220359 2.785 1 0 294.848 0 2.25183 2.783 0.00029896 0.870698 0.705629 0.310841 0.436981 2.25201 140.079 83.5778 18.701 60.7011 0.00403946 0 -40 10
1.884 5.44882e-08 2.54015e-06 0.151264 0.151263 0.0120246 2.47674e-05 0.00115461 0.189079 0.000658875 0.189734 0.963042 101.36 0.23362 0.871477 4.63989 0.0663805 0.0437725 0.956227 0.0193615 0.00465818 0.018616 0.0044382 0.00563849 0.006384 0.22554 0.25536 58.0573 -87.8996 126.13 15.9302 145.039 0.000142559 0.26734 192.705 0.310136 0.0673181 0.00409888 0.000562467 0.00138538 0.986956 0.991714 -2.9921e-06 -85.6558 0.0930968 31166.1 311.818 0.983495 0.319146 0.739524 0.73952 9.99958 2.98711e-06 1.19483e-05 0.134878 0.983437 0.931234 -0.0132914 4.93442e-06 0.51863 -2.03377e-20 7.55035e-24 -2.03301e-20 0.00139661 0.997814 8.60334e-05 0.152752 2.85291 0.00139661 0.997815 0.799036 0.00106956 0.00188159 0.000860334 0.455357 0.00188159 0.44512 0.000131549 1.02 0.888906 0.534337 0.287751 1.7198e-07 3.08715e-09 2368.76 3144.66 -0.058757 0.482217 0.277239 0.25514 -0.592999 -0.169582 0.485862 -0.265526 -0.220345 2.786 1 0 294.844 0 2.25196 2.784 0.000298959 0.870728 0.705671 0.310803 0.437003 2.25214 140.086 83.5772 18.701 60.7008 0.00403949 0 -40 10
1.885 5.4517e-08 2.54015e-06 0.151293 0.151293 0.0120246 2.47805e-05 0.00115461 0.189117 0.000658876 0.189771 0.963134 101.359 0.233609 0.871612 4.64057 0.0663914 0.043779 0.956221 0.0193609 0.00465866 0.0186154 0.00443861 0.00563908 0.00638461 0.225563 0.255384 58.0574 -87.8996 126.129 15.9301 145.039 0.000142561 0.26734 192.705 0.310135 0.067318 0.00409889 0.000562468 0.00138538 0.986956 0.991714 -2.99212e-06 -85.6558 0.0930969 31166 311.831 0.983495 0.319146 0.739536 0.739532 9.99958 2.98712e-06 1.19484e-05 0.134883 0.983437 0.931233 -0.0132914 4.93445e-06 0.518651 -2.03394e-20 7.55101e-24 -2.03318e-20 0.00139661 0.997814 8.60335e-05 0.152752 2.85291 0.00139661 0.997815 0.799106 0.00106958 0.00188159 0.000860335 0.455357 0.00188159 0.445124 0.000131552 1.02 0.888907 0.534337 0.287752 1.7198e-07 3.08717e-09 2368.74 3144.71 -0.0587621 0.482217 0.277239 0.255144 -0.592998 -0.169582 0.485845 -0.265524 -0.220331 2.787 1 0 294.839 0 2.2521 2.785 0.000298957 0.870757 0.705714 0.310766 0.437025 2.25228 140.094 83.5766 18.7009 60.7005 0.00403951 0 -40 10
1.886 5.45459e-08 2.54015e-06 0.151323 0.151323 0.0120246 2.47936e-05 0.00115461 0.189154 0.000658876 0.189808 0.963226 101.359 0.233598 0.871746 4.64125 0.0664023 0.0437854 0.956215 0.0193603 0.00465914 0.0186148 0.00443903 0.00563967 0.00638522 0.225587 0.255409 58.0575 -87.8996 126.129 15.9301 145.039 0.000142564 0.267341 192.705 0.310135 0.067318 0.00409889 0.000562468 0.00138538 0.986956 0.991714 -2.99213e-06 -85.6558 0.093097 31166 311.844 0.983495 0.319146 0.739548 0.739544 9.99958 2.98712e-06 1.19484e-05 0.134887 0.983437 0.931232 -0.0132914 4.93448e-06 0.518672 -2.0341e-20 7.55168e-24 -2.03335e-20 0.00139661 0.997814 8.60335e-05 0.152752 2.85291 0.00139661 0.997815 0.799175 0.00106959 0.00188159 0.000860335 0.455357 0.00188159 0.445129 0.000131554 1.02 0.888908 0.534337 0.287754 1.71981e-07 3.0872e-09 2368.72 3144.76 -0.0587672 0.482218 0.277239 0.255147 -0.592998 -0.169582 0.485829 -0.265522 -0.220316 2.788 1 0 294.835 0 2.25224 2.786 0.000298956 0.870787 0.705756 0.310729 0.437046 2.25241 140.101 83.576 18.7009 60.7002 0.00403954 0 -40 10
1.887 5.45747e-08 2.54015e-06 0.151353 0.151352 0.0120246 2.48067e-05 0.00115461 0.189191 0.000658876 0.189845 0.963318 101.358 0.233587 0.87188 4.64194 0.0664132 0.0437919 0.956208 0.0193597 0.00465961 0.0186142 0.00443944 0.00564026 0.00638583 0.22561 0.255433 58.0575 -87.8996 126.129 15.9301 145.039 0.000142566 0.267341 192.705 0.310135 0.0673179 0.00409889 0.000562469 0.00138539 0.986956 0.991714 -2.99215e-06 -85.6558 0.093097 31166 311.857 0.983495 0.319146 0.73956 0.739556 9.99958 2.98713e-06 1.19484e-05 0.134892 0.983438 0.931231 -0.0132914 4.93451e-06 0.518693 -2.03427e-20 7.55234e-24 -2.03351e-20 0.00139661 0.997814 8.60336e-05 0.152753 2.85291 0.00139661 0.997815 0.799245 0.00106961 0.00188159 0.000860336 0.455356 0.00188159 0.445134 0.000131556 1.02 0.888909 0.534336 0.287755 1.71981e-07 3.08722e-09 2368.71 3144.82 -0.0587723 0.482218 0.277238 0.25515 -0.592997 -0.169582 0.485813 -0.26552 -0.220302 2.789 1 0 294.83 0 2.25237 2.787 0.000298955 0.870817 0.705799 0.310692 0.437068 2.25255 140.108 83.5754 18.7009 60.6999 0.00403956 0 -40 10
1.888 5.46035e-08 2.54015e-06 0.151382 0.151382 0.0120246 2.48198e-05 0.00115462 0.189228 0.000658877 0.189882 0.96341 101.357 0.233576 0.872014 4.64262 0.0664241 0.0437983 0.956202 0.0193591 0.00466009 0.0186136 0.00443986 0.00564085 0.00638644 0.225634 0.255458 58.0576 -87.8996 126.129 15.93 145.039 0.000142568 0.267341 192.705 0.310134 0.0673179 0.0040989 0.00056247 0.00138539 0.986956 0.991714 -2.99216e-06 -85.6558 0.0930971 31166 311.87 0.983495 0.319146 0.739573 0.739568 9.99958 2.98713e-06 1.19484e-05 0.134897 0.983438 0.93123 -0.0132914 4.93454e-06 0.518714 -2.03444e-20 7.55301e-24 -2.03368e-20 0.00139661 0.997814 8.60337e-05 0.152753 2.85291 0.00139661 0.997815 0.799314 0.00106962 0.00188159 0.000860337 0.455356 0.00188159 0.445139 0.000131558 1.02 0.88891 0.534336 0.287757 1.71981e-07 3.08724e-09 2368.69 3144.87 -0.0587774 0.482218 0.277238 0.255153 -0.592996 -0.169582 0.485797 -0.265518 -0.220288 2.79 1 0 294.825 0 2.25251 2.788 0.000298953 0.870846 0.705841 0.310655 0.43709 2.25268 140.116 83.5748 18.7008 60.6997 0.00403959 0 -40 10
1.889 5.46324e-08 2.54015e-06 0.151412 0.151412 0.0120246 2.48329e-05 0.00115462 0.189265 0.000658877 0.189919 0.963502 101.357 0.233565 0.872149 4.64331 0.066435 0.0438048 0.956195 0.0193586 0.00466057 0.0186129 0.00444027 0.00564144 0.00638705 0.225658 0.255482 58.0576 -87.8996 126.128 15.93 145.039 0.000142571 0.267341 192.705 0.310134 0.0673178 0.0040989 0.00056247 0.00138539 0.986956 0.991714 -2.99218e-06 -85.6558 0.0930972 31165.9 311.883 0.983495 0.319146 0.739585 0.73958 9.99958 2.98714e-06 1.19484e-05 0.134902 0.983438 0.931229 -0.0132914 4.93457e-06 0.518735 -2.0346e-20 7.55368e-24 -2.03385e-20 0.00139661 0.997814 8.60338e-05 0.152753 2.85291 0.00139661 0.997815 0.799384 0.00106964 0.00188159 0.000860338 0.455356 0.00188159 0.445144 0.000131561 1.02 0.888912 0.534336 0.287758 1.71981e-07 3.08727e-09 2368.68 3144.92 -0.0587826 0.482218 0.277238 0.255157 -0.592996 -0.169582 0.485781 -0.265516 -0.220274 2.791 1 0 294.821 0 2.25264 2.789 0.000298952 0.870876 0.705884 0.310618 0.437112 2.25282 140.123 83.5742 18.7008 60.6994 0.00403961 0 -40 10
1.89 5.46612e-08 2.54016e-06 0.151442 0.151441 0.0120245 2.4846e-05 0.00115462 0.189302 0.000658878 0.189956 0.963594 101.356 0.233554 0.872283 4.64399 0.0664459 0.0438112 0.956189 0.019358 0.00466105 0.0186123 0.00444069 0.00564203 0.00638766 0.225681 0.255506 58.0577 -87.8997 126.128 15.9299 145.039 0.000142573 0.267341 192.704 0.310133 0.0673178 0.0040989 0.000562471 0.00138539 0.986956 0.991714 -2.99219e-06 -85.6557 0.0930973 31165.9 311.896 0.983495 0.319146 0.739597 0.739593 9.99958 2.98714e-06 1.19485e-05 0.134907 0.983438 0.931227 -0.0132914 4.9346e-06 0.518756 -2.03477e-20 7.55434e-24 -2.03401e-20 0.00139661 0.997814 8.60339e-05 0.152753 2.85291 0.00139661 0.997815 0.799454 0.00106965 0.0018816 0.000860339 0.455356 0.00188159 0.445149 0.000131563 1.02 0.888913 0.534335 0.28776 1.71982e-07 3.08729e-09 2368.66 3144.97 -0.0587877 0.482218 0.277237 0.25516 -0.592995 -0.169582 0.485764 -0.265514 -0.22026 2.792 1 0 294.816 0 2.25278 2.79 0.000298951 0.870906 0.705926 0.310581 0.437134 2.25296 140.13 83.5736 18.7008 60.6991 0.00403964 0 -40 10
1.891 5.469e-08 2.54016e-06 0.151471 0.151471 0.0120245 2.48591e-05 0.00115462 0.189339 0.000658878 0.189993 0.963685 101.355 0.233543 0.872417 4.64468 0.0664568 0.0438177 0.956182 0.0193574 0.00466153 0.0186117 0.0044411 0.00564263 0.00638827 0.225705 0.255531 58.0578 -87.8997 126.128 15.9299 145.039 0.000142575 0.267342 192.704 0.310133 0.0673177 0.0040989 0.000562472 0.00138539 0.986956 0.991714 -2.99221e-06 -85.6557 0.0930974 31165.9 311.909 0.983495 0.319146 0.739609 0.739605 9.99958 2.98715e-06 1.19485e-05 0.134912 0.983438 0.931226 -0.0132914 4.93463e-06 0.518776 -2.03494e-20 7.55501e-24 -2.03418e-20 0.00139662 0.997814 8.60339e-05 0.152753 2.85291 0.00139661 0.997815 0.799523 0.00106967 0.0018816 0.000860339 0.455356 0.0018816 0.445154 0.000131565 1.02 0.888914 0.534335 0.287761 1.71982e-07 3.08731e-09 2368.64 3145.02 -0.0587928 0.482218 0.277237 0.255163 -0.592994 -0.169582 0.485748 -0.265512 -0.220246 2.793 1 0 294.811 0 2.25292 2.791 0.000298949 0.870935 0.705969 0.310544 0.437156 2.25309 140.137 83.573 18.7007 60.6988 0.00403966 0 -40 10
1.892 5.47188e-08 2.54016e-06 0.151501 0.1515 0.0120245 2.48722e-05 0.00115462 0.189376 0.000658879 0.19003 0.963777 101.355 0.233532 0.872551 4.64536 0.0664677 0.0438242 0.956176 0.0193568 0.00466201 0.0186111 0.00444152 0.00564322 0.00638888 0.225729 0.255555 58.0578 -87.8997 126.128 15.9299 145.039 0.000142578 0.267342 192.704 0.310132 0.0673177 0.00409891 0.000562472 0.0013854 0.986956 0.991714 -2.99222e-06 -85.6557 0.0930975 31165.9 311.922 0.983495 0.319146 0.739621 0.739617 9.99958 2.98715e-06 1.19485e-05 0.134917 0.983438 0.931225 -0.0132914 4.93466e-06 0.518797 -2.0351e-20 7.55567e-24 -2.03435e-20 0.00139662 0.997814 8.6034e-05 0.152753 2.85292 0.00139662 0.997815 0.799593 0.00106969 0.0018816 0.00086034 0.455355 0.0018816 0.445159 0.000131568 1.02 0.888915 0.534335 0.287763 1.71982e-07 3.08733e-09 2368.63 3145.07 -0.0587979 0.482218 0.277237 0.255166 -0.592994 -0.169582 0.485732 -0.26551 -0.220232 2.794 1 0 294.807 0 2.25305 2.792 0.000298948 0.870965 0.706011 0.310507 0.437178 2.25323 140.145 83.5724 18.7007 60.6985 0.00403969 0 -40 10
1.893 5.47477e-08 2.54016e-06 0.15153 0.15153 0.0120245 2.48853e-05 0.00115462 0.189413 0.000658879 0.190067 0.963869 101.354 0.233521 0.872686 4.64605 0.0664786 0.0438307 0.956169 0.0193562 0.00466249 0.0186105 0.00444194 0.00564381 0.0063895 0.225752 0.25558 58.0579 -87.8997 126.128 15.9298 145.039 0.00014258 0.267342 192.704 0.310132 0.0673176 0.00409891 0.000562473 0.0013854 0.986956 0.991714 -2.99224e-06 -85.6557 0.0930976 31165.9 311.935 0.983495 0.319146 0.739634 0.739629 9.99958 2.98716e-06 1.19485e-05 0.134922 0.983439 0.931224 -0.0132914 4.93469e-06 0.518818 -2.03527e-20 7.55634e-24 -2.03452e-20 0.00139662 0.997814 8.60341e-05 0.152753 2.85292 0.00139662 0.997815 0.799662 0.0010697 0.0018816 0.000860341 0.455355 0.0018816 0.445163 0.00013157 1.02 0.888916 0.534334 0.287764 1.71983e-07 3.08736e-09 2368.61 3145.12 -0.058803 0.482218 0.277237 0.25517 -0.592993 -0.169582 0.485716 -0.265508 -0.220218 2.795 1 0 294.802 0 2.25319 2.793 0.000298947 0.870995 0.706054 0.31047 0.4372 2.25336 140.152 83.5718 18.7007 60.6982 0.00403971 0 -40 10
1.894 5.47765e-08 2.54016e-06 0.15156 0.151559 0.0120245 2.48984e-05 0.00115462 0.18945 0.00065888 0.190104 0.963961 101.353 0.23351 0.87282 4.64674 0.0664895 0.0438371 0.956163 0.0193556 0.00466297 0.0186099 0.00444235 0.0056444 0.00639011 0.225776 0.255604 58.058 -87.8997 126.127 15.9298 145.039 0.000142582 0.267342 192.704 0.310132 0.0673176 0.00409891 0.000562474 0.0013854 0.986956 0.991714 -2.99225e-06 -85.6557 0.0930976 31165.8 311.948 0.983495 0.319146 0.739646 0.739641 9.99958 2.98716e-06 1.19485e-05 0.134926 0.983439 0.931223 -0.0132914 4.93472e-06 0.518839 -2.03544e-20 7.55701e-24 -2.03468e-20 0.00139662 0.997814 8.60342e-05 0.152754 2.85292 0.00139662 0.997815 0.799731 0.00106972 0.0018816 0.000860342 0.455355 0.0018816 0.445168 0.000131572 1.02 0.888917 0.534334 0.287766 1.71983e-07 3.08738e-09 2368.59 3145.17 -0.0588081 0.482218 0.277236 0.255173 -0.592993 -0.169582 0.4857 -0.265506 -0.220203 2.796 1 0 294.798 0 2.25332 2.794 0.000298945 0.871024 0.706096 0.310433 0.437222 2.2535 140.159 83.5712 18.7006 60.6979 0.00403974 0 -40 10
1.895 5.48053e-08 2.54017e-06 0.151589 0.151589 0.0120245 2.49115e-05 0.00115462 0.189487 0.00065888 0.190141 0.964053 101.353 0.2335 0.872954 4.64742 0.0665004 0.0438436 0.956156 0.019355 0.00466345 0.0186093 0.00444277 0.00564499 0.00639072 0.2258 0.255629 58.058 -87.8997 126.127 15.9298 145.039 0.000142585 0.267342 192.704 0.310131 0.0673175 0.00409892 0.000562474 0.0013854 0.986956 0.991714 -2.99227e-06 -85.6557 0.0930977 31165.8 311.961 0.983495 0.319146 0.739658 0.739654 9.99958 2.98717e-06 1.19486e-05 0.134931 0.983439 0.931222 -0.0132914 4.93475e-06 0.51886 -2.03561e-20 7.55768e-24 -2.03485e-20 0.00139662 0.997814 8.60343e-05 0.152754 2.85292 0.00139662 0.997815 0.799801 0.00106973 0.0018816 0.000860343 0.455355 0.0018816 0.445173 0.000131575 1.02 0.888918 0.534334 0.287767 1.71983e-07 3.0874e-09 2368.58 3145.22 -0.0588132 0.482218 0.277236 0.255176 -0.592992 -0.169582 0.485683 -0.265503 -0.220189 2.797 1 0 294.793 0 2.25346 2.795 0.000298944 0.871054 0.706139 0.310396 0.437243 2.25364 140.167 83.5706 18.7006 60.6976 0.00403976 0 -40 10
1.896 5.48342e-08 2.54017e-06 0.151619 0.151618 0.0120245 2.49246e-05 0.00115462 0.189524 0.00065888 0.190178 0.964145 101.352 0.233489 0.873089 4.64811 0.0665113 0.0438501 0.95615 0.0193544 0.00466393 0.0186087 0.00444319 0.00564559 0.00639133 0.225823 0.255653 58.0581 -87.8997 126.127 15.9297 145.039 0.000142587 0.267343 192.703 0.310131 0.0673175 0.00409892 0.000562475 0.0013854 0.986956 0.991714 -2.99228e-06 -85.6557 0.0930978 31165.8 311.974 0.983495 0.319146 0.73967 0.739666 9.99958 2.98717e-06 1.19486e-05 0.134936 0.983439 0.931221 -0.0132914 4.93478e-06 0.518881 -2.03577e-20 7.55834e-24 -2.03502e-20 0.00139662 0.997814 8.60343e-05 0.152754 2.85292 0.00139662 0.997815 0.79987 0.00106975 0.0018816 0.000860343 0.455354 0.0018816 0.445178 0.000131577 1.02 0.888919 0.534333 0.287769 1.71983e-07 3.08743e-09 2368.56 3145.28 -0.0588183 0.482218 0.277236 0.25518 -0.592991 -0.169582 0.485667 -0.265501 -0.220175 2.798 1 0 294.788 0 2.25359 2.796 0.000298943 0.871084 0.706181 0.310359 0.437265 2.25377 140.174 83.57 18.7006 60.6973 0.00403979 0 -40 10
1.897 5.4863e-08 2.54017e-06 0.151648 0.151648 0.0120244 2.49377e-05 0.00115462 0.18956 0.000658881 0.190215 0.964237 101.351 0.233478 0.873223 4.6488 0.0665223 0.0438566 0.956143 0.0193538 0.00466441 0.0186081 0.0044436 0.00564618 0.00639195 0.225847 0.255678 58.0581 -87.8997 126.127 15.9297 145.039 0.000142589 0.267343 192.703 0.31013 0.0673174 0.00409892 0.000562476 0.00138541 0.986956 0.991714 -2.9923e-06 -85.6557 0.0930979 31165.8 311.987 0.983495 0.319146 0.739682 0.739678 9.99958 2.98718e-06 1.19486e-05 0.134941 0.983439 0.93122 -0.0132914 4.93481e-06 0.518902 -2.03594e-20 7.55901e-24 -2.03519e-20 0.00139662 0.997814 8.60344e-05 0.152754 2.85292 0.00139662 0.997815 0.79994 0.00106977 0.00188161 0.000860344 0.455354 0.0018816 0.445183 0.000131579 1.02 0.88892 0.534333 0.28777 1.71984e-07 3.08745e-09 2368.55 3145.33 -0.0588234 0.482218 0.277235 0.255183 -0.592991 -0.169582 0.485651 -0.265499 -0.220161 2.799 1 0 294.784 0 2.25373 2.797 0.000298941 0.871114 0.706224 0.310322 0.437287 2.25391 140.181 83.5694 18.7005 60.6971 0.00403981 0 -40 10
1.898 5.48918e-08 2.54017e-06 0.151678 0.151677 0.0120244 2.49508e-05 0.00115462 0.189597 0.000658881 0.190251 0.964329 101.351 0.233467 0.873357 4.64949 0.0665332 0.0438631 0.956137 0.0193532 0.00466489 0.0186074 0.00444402 0.00564677 0.00639256 0.225871 0.255702 58.0582 -87.8997 126.126 15.9296 145.039 0.000142592 0.267343 192.703 0.31013 0.0673173 0.00409893 0.000562476 0.00138541 0.986956 0.991714 -2.99231e-06 -85.6557 0.093098 31165.7 312 0.983495 0.319146 0.739695 0.73969 9.99958 2.98718e-06 1.19486e-05 0.134946 0.98344 0.931219 -0.0132914 4.93484e-06 0.518923 -2.03611e-20 7.55968e-24 -2.03535e-20 0.00139662 0.997814 8.60345e-05 0.152754 2.85292 0.00139662 0.997815 0.800009 0.00106978 0.00188161 0.000860345 0.455354 0.00188161 0.445188 0.000131582 1.02 0.888921 0.534333 0.287772 1.71984e-07 3.08747e-09 2368.53 3145.38 -0.0588285 0.482218 0.277235 0.255186 -0.59299 -0.169582 0.485635 -0.265497 -0.220147 2.8 1 0 294.779 0 2.25387 2.798 0.00029894 0.871143 0.706267 0.310286 0.437309 2.25404 140.188 83.5688 18.7005 60.6968 0.00403984 0 -40 10
1.899 5.49207e-08 2.54017e-06 0.151707 0.151707 0.0120244 2.49639e-05 0.00115462 0.189634 0.000658882 0.190288 0.964421 101.35 0.233456 0.873492 4.65018 0.0665441 0.0438696 0.95613 0.0193526 0.00466537 0.0186068 0.00444444 0.00564736 0.00639317 0.225895 0.255727 58.0583 -87.8997 126.126 15.9296 145.039 0.000142594 0.267343 192.703 0.310129 0.0673173 0.00409893 0.000562477 0.00138541 0.986956 0.991714 -2.99233e-06 -85.6557 0.0930981 31165.7 312.013 0.983495 0.319146 0.739707 0.739702 9.99958 2.98719e-06 1.19486e-05 0.134951 0.98344 0.931218 -0.0132914 4.93487e-06 0.518944 -2.03628e-20 7.56035e-24 -2.03552e-20 0.00139662 0.997814 8.60346e-05 0.152754 2.85292 0.00139662 0.997815 0.800078 0.0010698 0.00188161 0.000860346 0.455354 0.00188161 0.445192 0.000131584 1.02 0.888923 0.534333 0.287773 1.71984e-07 3.08749e-09 2368.51 3145.43 -0.0588336 0.482219 0.277235 0.255189 -0.592989 -0.169582 0.485618 -0.265495 -0.220133 2.801 1 0 294.775 0 2.254 2.799 0.000298939 0.871173 0.706309 0.310249 0.437331 2.25418 140.196 83.5682 18.7005 60.6965 0.00403986 0 -40 10
1.9 5.49495e-08 2.54017e-06 0.151737 0.151736 0.0120244 2.4977e-05 0.00115462 0.189671 0.000658882 0.190325 0.964513 101.349 0.233445 0.873626 4.65087 0.066555 0.0438761 0.956124 0.019352 0.00466586 0.0186062 0.00444486 0.00564796 0.00639379 0.225918 0.255751 58.0583 -87.8997 126.126 15.9296 145.039 0.000142596 0.267343 192.703 0.310129 0.0673172 0.00409893 0.000562478 0.00138541 0.986956 0.991714 -2.99234e-06 -85.6557 0.0930982 31165.7 312.026 0.983495 0.319146 0.739719 0.739715 9.99958 2.98719e-06 1.19487e-05 0.134956 0.98344 0.931217 -0.0132914 4.9349e-06 0.518965 -2.03644e-20 7.56102e-24 -2.03569e-20 0.00139663 0.997814 8.60347e-05 0.152755 2.85292 0.00139663 0.997815 0.800148 0.00106981 0.00188161 0.000860347 0.455354 0.00188161 0.445197 0.000131586 1.02 0.888924 0.534332 0.287775 1.71984e-07 3.08752e-09 2368.5 3145.48 -0.0588388 0.482219 0.277235 0.255193 -0.592989 -0.169583 0.485602 -0.265493 -0.220119 2.802 1 0 294.77 0 2.25414 2.8 0.000298937 0.871203 0.706352 0.310212 0.437353 2.25431 140.203 83.5676 18.7004 60.6962 0.00403988 0 -40 10
1.901 5.49783e-08 2.54018e-06 0.151766 0.151765 0.0120244 2.49901e-05 0.00115463 0.189707 0.000658883 0.190362 0.964605 101.348 0.233434 0.87376 4.65156 0.0665659 0.0438826 0.956117 0.0193514 0.00466634 0.0186056 0.00444527 0.00564855 0.0063944 0.225942 0.255776 58.0584 -87.8997 126.126 15.9295 145.039 0.000142599 0.267344 192.703 0.310129 0.0673172 0.00409894 0.000562478 0.00138542 0.986956 0.991714 -2.99236e-06 -85.6556 0.0930983 31165.7 312.039 0.983495 0.319146 0.739731 0.739727 9.99958 2.9872e-06 1.19487e-05 0.134961 0.98344 0.931216 -0.0132914 4.93493e-06 0.518986 -2.03661e-20 7.56169e-24 -2.03586e-20 0.00139663 0.997814 8.60347e-05 0.152755 2.85292 0.00139663 0.997815 0.800217 0.00106983 0.00188161 0.000860347 0.455353 0.00188161 0.445202 0.000131588 1.02 0.888925 0.534332 0.287776 1.71985e-07 3.08754e-09 2368.48 3145.53 -0.0588439 0.482219 0.277234 0.255196 -0.592988 -0.169583 0.485586 -0.265491 -0.220104 2.803 1 0 294.765 0 2.25427 2.801 0.000298936 0.871233 0.706394 0.310175 0.437375 2.25445 140.21 83.567 18.7004 60.6959 0.00403991 0 -40 10
1.902 5.50071e-08 2.54018e-06 0.151795 0.151795 0.0120244 2.50032e-05 0.00115463 0.189744 0.000658883 0.190398 0.964697 101.348 0.233423 0.873895 4.65225 0.0665768 0.0438891 0.956111 0.0193509 0.00466682 0.018605 0.00444569 0.00564914 0.00639501 0.225966 0.255801 58.0585 -87.8997 126.126 15.9295 145.039 0.000142601 0.267344 192.702 0.310128 0.0673171 0.00409894 0.000562479 0.00138542 0.986956 0.991714 -2.99237e-06 -85.6556 0.0930983 31165.6 312.052 0.983494 0.319146 0.739743 0.739739 9.99958 2.9872e-06 1.19487e-05 0.134966 0.98344 0.931215 -0.0132914 4.93496e-06 0.519007 -2.03678e-20 7.56236e-24 -2.03602e-20 0.00139663 0.997814 8.60348e-05 0.152755 2.85292 0.00139663 0.997815 0.800286 0.00106984 0.00188161 0.000860348 0.455353 0.00188161 0.445207 0.000131591 1.02 0.888926 0.534332 0.287778 1.71985e-07 3.08756e-09 2368.46 3145.58 -0.058849 0.482219 0.277234 0.255199 -0.592987 -0.169583 0.48557 -0.265489 -0.22009 2.804 1 0 294.761 0 2.25441 2.802 0.000298935 0.871262 0.706437 0.310139 0.437396 2.25458 140.218 83.5664 18.7004 60.6956 0.00403993 0 -40 10
1.903 5.5036e-08 2.54018e-06 0.151825 0.151824 0.0120244 2.50163e-05 0.00115463 0.189781 0.000658884 0.190435 0.964789 101.347 0.233412 0.874029 4.65294 0.0665878 0.0438957 0.956104 0.0193503 0.0046673 0.0186044 0.00444611 0.00564974 0.00639563 0.22599 0.255825 58.0585 -87.8997 126.125 15.9295 145.039 0.000142603 0.267344 192.702 0.310128 0.0673171 0.00409894 0.00056248 0.00138542 0.986956 0.991714 -2.99239e-06 -85.6556 0.0930984 31165.6 312.066 0.983494 0.319146 0.739756 0.739751 9.99958 2.98721e-06 1.19487e-05 0.13497 0.98344 0.931214 -0.0132914 4.93499e-06 0.519028 -2.03695e-20 7.56302e-24 -2.03619e-20 0.00139663 0.997814 8.60349e-05 0.152755 2.85293 0.00139663 0.997815 0.800355 0.00106986 0.00188161 0.000860349 0.455353 0.00188161 0.445212 0.000131593 1.02 0.888927 0.534331 0.287779 1.71985e-07 3.08759e-09 2368.45 3145.63 -0.0588541 0.482219 0.277234 0.255202 -0.592987 -0.169583 0.485553 -0.265487 -0.220076 2.805 1 0 294.756 0 2.25454 2.803 0.000298933 0.871292 0.706479 0.310102 0.437418 2.25472 140.225 83.5658 18.7003 60.6953 0.00403996 0 -40 10
1.904 5.50648e-08 2.54018e-06 0.151854 0.151853 0.0120243 2.50295e-05 0.00115463 0.189817 0.000658884 0.190472 0.964881 101.346 0.233401 0.874164 4.65363 0.0665987 0.0439022 0.956098 0.0193497 0.00466778 0.0186038 0.00444653 0.00565033 0.00639624 0.226013 0.25585 58.0586 -87.8997 126.125 15.9294 145.039 0.000142606 0.267344 192.702 0.310127 0.067317 0.00409894 0.00056248 0.00138542 0.986956 0.991714 -2.9924e-06 -85.6556 0.0930985 31165.6 312.079 0.983494 0.319146 0.739768 0.739763 9.99958 2.98721e-06 1.19487e-05 0.134975 0.983441 0.931213 -0.0132914 4.93502e-06 0.519049 -2.03712e-20 7.56369e-24 -2.03636e-20 0.00139663 0.997814 8.6035e-05 0.152755 2.85293 0.00139663 0.997815 0.800425 0.00106988 0.00188162 0.00086035 0.455353 0.00188162 0.445217 0.000131595 1.02 0.888928 0.534331 0.287781 1.71986e-07 3.08761e-09 2368.43 3145.69 -0.0588592 0.482219 0.277234 0.255206 -0.592986 -0.169583 0.485537 -0.265485 -0.220062 2.806 1 0 294.752 0 2.25468 2.804 0.000298932 0.871322 0.706522 0.310065 0.43744 2.25486 140.232 83.5652 18.7003 60.695 0.00403998 0 -40 10
1.905 5.50936e-08 2.54018e-06 0.151883 0.151883 0.0120243 2.50426e-05 0.00115463 0.189854 0.000658884 0.190508 0.964973 101.346 0.23339 0.874298 4.65432 0.0666096 0.0439087 0.956091 0.0193491 0.00466826 0.0186031 0.00444695 0.00565093 0.00639686 0.226037 0.255874 58.0586 -87.8997 126.125 15.9294 145.039 0.000142608 0.267344 192.702 0.310127 0.067317 0.00409895 0.000562481 0.00138542 0.986955 0.991714 -2.99242e-06 -85.6556 0.0930986 31165.6 312.092 0.983494 0.319146 0.73978 0.739776 9.99958 2.98722e-06 1.19488e-05 0.13498 0.983441 0.931212 -0.0132914 4.93505e-06 0.51907 -2.03728e-20 7.56436e-24 -2.03653e-20 0.00139663 0.997814 8.60351e-05 0.152755 2.85293 0.00139663 0.997815 0.800494 0.00106989 0.00188162 0.000860351 0.455352 0.00188162 0.445221 0.000131598 1.02 0.888929 0.534331 0.287782 1.71986e-07 3.08763e-09 2368.42 3145.74 -0.0588643 0.482219 0.277233 0.255209 -0.592985 -0.169583 0.485521 -0.265482 -0.220048 2.807 1 0 294.747 0 2.25481 2.805 0.000298931 0.871352 0.706564 0.310028 0.437462 2.25499 140.239 83.5646 18.7002 60.6947 0.00404001 0 -40 10
1.906 5.51225e-08 2.54019e-06 0.151912 0.151912 0.0120243 2.50557e-05 0.00115463 0.18989 0.000658885 0.190545 0.965065 101.345 0.233379 0.874432 4.65502 0.0666205 0.0439153 0.956085 0.0193485 0.00466875 0.0186025 0.00444736 0.00565152 0.00639747 0.226061 0.255899 58.0587 -87.8997 126.125 15.9294 145.039 0.000142611 0.267344 192.702 0.310126 0.0673169 0.00409895 0.000562482 0.00138543 0.986955 0.991714 -2.99243e-06 -85.6556 0.0930987 31165.6 312.105 0.983494 0.319146 0.739792 0.739788 9.99958 2.98722e-06 1.19488e-05 0.134985 0.983441 0.931211 -0.0132914 4.93508e-06 0.519091 -2.03745e-20 7.56503e-24 -2.03669e-20 0.00139663 0.997814 8.60351e-05 0.152755 2.85293 0.00139663 0.997815 0.800563 0.00106991 0.00188162 0.000860351 0.455352 0.00188162 0.445226 0.0001316 1.02 0.88893 0.53433 0.287784 1.71986e-07 3.08766e-09 2368.4 3145.79 -0.0588694 0.482219 0.277233 0.255212 -0.592985 -0.169583 0.485505 -0.26548 -0.220034 2.808 1 0 294.742 0 2.25495 2.806 0.000298929 0.871381 0.706606 0.309992 0.437484 2.25513 140.247 83.564 18.7002 60.6945 0.00404003 0 -40 10
1.907 5.51513e-08 2.54019e-06 0.151942 0.151941 0.0120243 2.50688e-05 0.00115463 0.189927 0.000658885 0.190581 0.965157 101.344 0.233369 0.874567 4.65571 0.0666315 0.0439218 0.956078 0.0193479 0.00466923 0.0186019 0.00444778 0.00565212 0.00639809 0.226085 0.255923 58.0588 -87.8997 126.124 15.9293 145.039 0.000142613 0.267345 192.702 0.310126 0.0673169 0.00409895 0.000562482 0.00138543 0.986955 0.991714 -2.99245e-06 -85.6556 0.0930988 31165.5 312.118 0.983494 0.319146 0.739804 0.7398 9.99958 2.98723e-06 1.19488e-05 0.13499 0.983441 0.93121 -0.0132914 4.93511e-06 0.519113 -2.03762e-20 7.56571e-24 -2.03686e-20 0.00139663 0.997814 8.60352e-05 0.152756 2.85293 0.00139663 0.997815 0.800632 0.00106992 0.00188162 0.000860352 0.455352 0.00188162 0.445231 0.000131602 1.02 0.888931 0.53433 0.287786 1.71986e-07 3.08768e-09 2368.38 3145.84 -0.0588745 0.482219 0.277233 0.255216 -0.592984 -0.169583 0.485488 -0.265478 -0.22002 2.809 1 0 294.738 0 2.25509 2.807 0.000298928 0.871411 0.706649 0.309955 0.437506 2.25526 140.254 83.5634 18.7002 60.6942 0.00404006 0 -40 10
1.908 5.51801e-08 2.54019e-06 0.151971 0.15197 0.0120243 2.50819e-05 0.00115463 0.189963 0.000658886 0.190618 0.96525 101.344 0.233358 0.874701 4.6564 0.0666424 0.0439283 0.956072 0.0193473 0.00466971 0.0186013 0.0044482 0.00565271 0.0063987 0.226108 0.255948 58.0588 -87.8997 126.124 15.9293 145.039 0.000142615 0.267345 192.701 0.310126 0.0673168 0.00409896 0.000562483 0.00138543 0.986955 0.991714 -2.99246e-06 -85.6556 0.0930989 31165.5 312.131 0.983494 0.319146 0.739817 0.739812 9.99958 2.98723e-06 1.19488e-05 0.134995 0.983441 0.931209 -0.0132914 4.93514e-06 0.519134 -2.03779e-20 7.56638e-24 -2.03703e-20 0.00139663 0.997814 8.60353e-05 0.152756 2.85293 0.00139663 0.997815 0.800701 0.00106994 0.00188162 0.000860353 0.455352 0.00188162 0.445236 0.000131605 1.02 0.888932 0.53433 0.287787 1.71987e-07 3.0877e-09 2368.37 3145.89 -0.0588797 0.482219 0.277232 0.255219 -0.592984 -0.169583 0.485472 -0.265476 -0.220005 2.81 1 0 294.733 0 2.25522 2.808 0.000298927 0.871441 0.706691 0.309919 0.437528 2.2554 140.261 83.5628 18.7001 60.6939 0.00404008 0 -40 10
1.909 5.52089e-08 2.54019e-06 0.152 0.151999 0.0120243 2.5095e-05 0.00115463 0.19 0.000658886 0.190654 0.965342 101.343 0.233347 0.874836 4.6571 0.0666533 0.0439349 0.956065 0.0193467 0.00467019 0.0186007 0.00444862 0.00565331 0.00639932 0.226132 0.255973 58.0589 -87.8997 126.124 15.9292 145.039 0.000142618 0.267345 192.701 0.310125 0.0673168 0.00409896 0.000562484 0.00138543 0.986955 0.991714 -2.99248e-06 -85.6556 0.093099 31165.5 312.144 0.983494 0.319146 0.739829 0.739824 9.99958 2.98724e-06 1.19488e-05 0.135 0.983441 0.931208 -0.0132914 4.93516e-06 0.519155 -2.03796e-20 7.56705e-24 -2.0372e-20 0.00139664 0.997814 8.60354e-05 0.152756 2.85293 0.00139664 0.997815 0.80077 0.00106995 0.00188162 0.000860354 0.455351 0.00188162 0.445241 0.000131607 1.02 0.888933 0.534329 0.287789 1.71987e-07 3.08772e-09 2368.35 3145.94 -0.0588848 0.482219 0.277232 0.255222 -0.592983 -0.169583 0.485456 -0.265474 -0.219991 2.811 1 0 294.729 0 2.25536 2.809 0.000298925 0.871471 0.706734 0.309882 0.437549 2.25553 140.269 83.5622 18.7001 60.6936 0.00404011 0 -40 10
1.91 5.52378e-08 2.54019e-06 0.152029 0.152029 0.0120243 2.51081e-05 0.00115463 0.190036 0.000658887 0.190691 0.965434 101.342 0.233336 0.87497 4.65779 0.0666642 0.0439414 0.956059 0.0193461 0.00467068 0.0186001 0.00444904 0.0056539 0.00639993 0.226156 0.255997 58.059 -87.8997 126.124 15.9292 145.039 0.00014262 0.267345 192.701 0.310125 0.0673167 0.00409896 0.000562484 0.00138544 0.986955 0.991714 -2.99249e-06 -85.6556 0.093099 31165.5 312.157 0.983494 0.319146 0.739841 0.739837 9.99958 2.98724e-06 1.19489e-05 0.135005 0.983442 0.931207 -0.0132914 4.93519e-06 0.519176 -2.03812e-20 7.56772e-24 -2.03737e-20 0.00139664 0.997814 8.60355e-05 0.152756 2.85293 0.00139664 0.997815 0.800839 0.00106997 0.00188163 0.000860355 0.455351 0.00188162 0.445246 0.000131609 1.02 0.888935 0.534329 0.28779 1.71987e-07 3.08775e-09 2368.33 3145.99 -0.0588899 0.482219 0.277232 0.255225 -0.592982 -0.169583 0.48544 -0.265472 -0.219977 2.812 1 0 294.724 0 2.25549 2.81 0.000298924 0.871501 0.706776 0.309846 0.437571 2.25567 140.276 83.5616 18.7001 60.6933 0.00404013 0 -40 10
1.911 5.52666e-08 2.5402e-06 0.152058 0.152058 0.0120242 2.51212e-05 0.00115463 0.190073 0.000658887 0.190727 0.965526 101.342 0.233325 0.875105 4.65849 0.0666752 0.043948 0.956052 0.0193455 0.00467116 0.0185995 0.00444946 0.0056545 0.00640055 0.22618 0.256022 58.059 -87.8997 126.124 15.9292 145.039 0.000142622 0.267345 192.701 0.310124 0.0673167 0.00409897 0.000562485 0.00138544 0.986955 0.991714 -2.99251e-06 -85.6555 0.0930991 31165.4 312.17 0.983494 0.319146 0.739853 0.739849 9.99958 2.98725e-06 1.19489e-05 0.13501 0.983442 0.931206 -0.0132914 4.93522e-06 0.519197 -2.03829e-20 7.56839e-24 -2.03754e-20 0.00139664 0.997814 8.60355e-05 0.152756 2.85293 0.00139664 0.997815 0.800908 0.00106999 0.00188163 0.000860355 0.455351 0.00188163 0.44525 0.000131611 1.02 0.888936 0.534329 0.287792 1.71987e-07 3.08777e-09 2368.32 3146.04 -0.058895 0.482219 0.277232 0.255229 -0.592982 -0.169583 0.485423 -0.26547 -0.219963 2.813 1 0 294.719 0 2.25563 2.811 0.000298923 0.871531 0.706819 0.309809 0.437593 2.2558 140.283 83.561 18.7 60.693 0.00404016 0 -40 10
1.912 5.52954e-08 2.5402e-06 0.152087 0.152087 0.0120242 2.51343e-05 0.00115464 0.190109 0.000658887 0.190763 0.965618 101.341 0.233314 0.875239 4.65918 0.0666861 0.0439545 0.956045 0.0193449 0.00467164 0.0185988 0.00444988 0.00565509 0.00640117 0.226204 0.256047 58.0591 -87.8997 126.123 15.9291 145.039 0.000142625 0.267346 192.701 0.310124 0.0673166 0.00409897 0.000562486 0.00138544 0.986955 0.991714 -2.99252e-06 -85.6555 0.0930992 31165.4 312.184 0.983494 0.319146 0.739865 0.739861 9.99958 2.98725e-06 1.19489e-05 0.135015 0.983442 0.931205 -0.0132914 4.93525e-06 0.519218 -2.03846e-20 7.56906e-24 -2.0377e-20 0.00139664 0.997814 8.60356e-05 0.152756 2.85293 0.00139664 0.997815 0.800977 0.00107 0.00188163 0.000860356 0.455351 0.00188163 0.445255 0.000131614 1.02 0.888937 0.534329 0.287793 1.71988e-07 3.08779e-09 2368.3 3146.09 -0.0589001 0.482219 0.277231 0.255232 -0.592981 -0.169583 0.485407 -0.265468 -0.219949 2.814 1 0 294.715 0 2.25576 2.812 0.000298921 0.87156 0.706861 0.309772 0.437615 2.25594 140.29 83.5604 18.7 60.6927 0.00404018 0 -40 10
1.913 5.53243e-08 2.5402e-06 0.152116 0.152116 0.0120242 2.51474e-05 0.00115464 0.190145 0.000658888 0.1908 0.96571 101.34 0.233303 0.875374 4.65988 0.066697 0.0439611 0.956039 0.0193443 0.00467213 0.0185982 0.0044503 0.00565569 0.00640178 0.226228 0.256071 58.0591 -87.8997 126.123 15.9291 145.039 0.000142627 0.267346 192.701 0.310123 0.0673166 0.00409897 0.000562486 0.00138544 0.986955 0.991714 -2.99254e-06 -85.6555 0.0930993 31165.4 312.197 0.983494 0.319146 0.739878 0.739873 9.99958 2.98726e-06 1.19489e-05 0.13502 0.983442 0.931204 -0.0132914 4.93528e-06 0.519239 -2.03863e-20 7.56973e-24 -2.03787e-20 0.00139664 0.997814 8.60357e-05 0.152757 2.85293 0.00139664 0.997815 0.801046 0.00107002 0.00188163 0.000860357 0.455351 0.00188163 0.44526 0.000131616 1.02 0.888938 0.534328 0.287795 1.71988e-07 3.08782e-09 2368.29 3146.15 -0.0589052 0.48222 0.277231 0.255235 -0.59298 -0.169583 0.485391 -0.265466 -0.219935 2.815 1 0 294.71 0 2.2559 2.813 0.00029892 0.87159 0.706904 0.309736 0.437637 2.25608 140.298 83.5598 18.7 60.6924 0.00404021 0 -40 10
1.914 5.53531e-08 2.5402e-06 0.152145 0.152145 0.0120242 2.51605e-05 0.00115464 0.190182 0.000658888 0.190836 0.965802 101.339 0.233292 0.875508 4.66057 0.066708 0.0439677 0.956032 0.0193437 0.00467261 0.0185976 0.00445072 0.00565629 0.0064024 0.226251 0.256096 58.0592 -87.8997 126.123 15.9291 145.039 0.000142629 0.267346 192.7 0.310123 0.0673165 0.00409897 0.000562487 0.00138544 0.986955 0.991714 -2.99255e-06 -85.6555 0.0930994 31165.4 312.21 0.983494 0.319146 0.73989 0.739885 9.99958 2.98726e-06 1.19489e-05 0.135025 0.983442 0.931203 -0.0132914 4.93531e-06 0.51926 -2.0388e-20 7.57041e-24 -2.03804e-20 0.00139664 0.997814 8.60358e-05 0.152757 2.85294 0.00139664 0.997815 0.801115 0.00107003 0.00188163 0.000860358 0.45535 0.00188163 0.445265 0.000131618 1.02 0.888939 0.534328 0.287796 1.71988e-07 3.08784e-09 2368.27 3146.2 -0.0589104 0.48222 0.277231 0.255239 -0.59298 -0.169583 0.485375 -0.265464 -0.21992 2.816 1 0 294.705 0 2.25604 2.814 0.000298919 0.87162 0.706946 0.3097 0.437659 2.25621 140.305 83.5592 18.6999 60.6921 0.00404023 0 -40 10
1.915 5.53819e-08 2.5402e-06 0.152174 0.152174 0.0120242 2.51736e-05 0.00115464 0.190218 0.000658889 0.190872 0.965895 101.339 0.233281 0.875643 4.66127 0.0667189 0.0439742 0.956026 0.0193431 0.00467309 0.018597 0.00445114 0.00565688 0.00640302 0.226275 0.256121 58.0593 -87.8997 126.123 15.929 145.039 0.000142632 0.267346 192.7 0.310123 0.0673165 0.00409898 0.000562488 0.00138545 0.986955 0.991714 -2.99257e-06 -85.6555 0.0930995 31165.4 312.223 0.983494 0.319146 0.739902 0.739898 9.99958 2.98727e-06 1.1949e-05 0.135029 0.983442 0.931202 -0.0132914 4.93534e-06 0.519281 -2.03897e-20 7.57108e-24 -2.03821e-20 0.00139664 0.997814 8.60359e-05 0.152757 2.85294 0.00139664 0.997815 0.801184 0.00107005 0.00188163 0.000860359 0.45535 0.00188163 0.44527 0.000131621 1.02 0.88894 0.534328 0.287798 1.71988e-07 3.08786e-09 2368.25 3146.25 -0.0589155 0.48222 0.27723 0.255242 -0.592979 -0.169583 0.485358 -0.265462 -0.219906 2.817 1 0 294.701 0 2.25617 2.815 0.000298917 0.87165 0.706989 0.309663 0.43768 2.25635 140.312 83.5586 18.6999 60.6918 0.00404026 0 -40 10
1.916 5.54107e-08 2.5402e-06 0.152203 0.152203 0.0120242 2.51867e-05 0.00115464 0.190254 0.000658889 0.190909 0.965987 101.338 0.23327 0.875777 4.66197 0.0667298 0.0439808 0.956019 0.0193425 0.00467358 0.0185964 0.00445156 0.00565748 0.00640363 0.226299 0.256145 58.0593 -87.8998 126.123 15.929 145.039 0.000142634 0.267346 192.7 0.310122 0.0673164 0.00409898 0.000562488 0.00138545 0.986955 0.991714 -2.99258e-06 -85.6555 0.0930996 31165.3 312.236 0.983494 0.319146 0.739914 0.73991 9.99958 2.98727e-06 1.1949e-05 0.135034 0.983443 0.931201 -0.0132914 4.93537e-06 0.519303 -2.03914e-20 7.57175e-24 -2.03838e-20 0.00139664 0.997814 8.60359e-05 0.152757 2.85294 0.00139664 0.997815 0.801253 0.00107007 0.00188163 0.000860359 0.45535 0.00188163 0.445274 0.000131623 1.02 0.888941 0.534327 0.287799 1.71989e-07 3.08788e-09 2368.24 3146.3 -0.0589206 0.48222 0.27723 0.255245 -0.592978 -0.169584 0.485342 -0.265459 -0.219892 2.818 1 0 294.696 0 2.25631 2.816 0.000298916 0.87168 0.707031 0.309627 0.437702 2.25648 140.32 83.558 18.6999 60.6916 0.00404028 0 -40 10
1.917 5.54396e-08 2.54021e-06 0.152232 0.152232 0.0120242 2.51998e-05 0.00115464 0.190291 0.00065889 0.190945 0.966079 101.337 0.233259 0.875912 4.66266 0.0667408 0.0439874 0.956013 0.0193419 0.00467406 0.0185957 0.00445198 0.00565808 0.00640425 0.226323 0.25617 58.0594 -87.8998 126.122 15.9289 145.039 0.000142636 0.267347 192.7 0.310122 0.0673163 0.00409898 0.000562489 0.00138545 0.986955 0.991714 -2.9926e-06 -85.6555 0.0930997 31165.3 312.249 0.983494 0.319146 0.739927 0.739922 9.99958 2.98728e-06 1.1949e-05 0.135039 0.983443 0.9312 -0.0132914 4.9354e-06 0.519324 -2.0393e-20 7.57242e-24 -2.03855e-20 0.00139664 0.997814 8.6036e-05 0.152757 2.85294 0.00139664 0.997815 0.801322 0.00107008 0.00188164 0.00086036 0.45535 0.00188163 0.445279 0.000131625 1.02 0.888942 0.534327 0.287801 1.71989e-07 3.08791e-09 2368.22 3146.35 -0.0589257 0.48222 0.27723 0.255248 -0.592978 -0.169584 0.485326 -0.265457 -0.219878 2.819 1 0 294.692 0 2.25644 2.817 0.000298915 0.87171 0.707074 0.30959 0.437724 2.25662 140.327 83.5574 18.6998 60.6913 0.00404031 0 -40 10
1.918 5.54684e-08 2.54021e-06 0.152261 0.152261 0.0120241 2.52129e-05 0.00115464 0.190327 0.00065889 0.190981 0.966171 101.337 0.233248 0.876046 4.66336 0.0667517 0.043994 0.956006 0.0193413 0.00467455 0.0185951 0.0044524 0.00565868 0.00640487 0.226347 0.256195 58.0595 -87.8998 126.122 15.9289 145.039 0.000142639 0.267347 192.7 0.310121 0.0673163 0.00409899 0.00056249 0.00138545 0.986955 0.991714 -2.99261e-06 -85.6555 0.0930997 31165.3 312.263 0.983494 0.319146 0.739939 0.739934 9.99958 2.98728e-06 1.1949e-05 0.135044 0.983443 0.931198 -0.0132914 4.93543e-06 0.519345 -2.03947e-20 7.5731e-24 -2.03872e-20 0.00139665 0.997814 8.60361e-05 0.152757 2.85294 0.00139665 0.997815 0.801391 0.0010701 0.00188164 0.000860361 0.455349 0.00188164 0.445284 0.000131628 1.02 0.888943 0.534327 0.287802 1.71989e-07 3.08793e-09 2368.2 3146.4 -0.0589308 0.48222 0.27723 0.255252 -0.592977 -0.169584 0.48531 -0.265455 -0.219864 2.82 1 0 294.687 0 2.25658 2.818 0.000298913 0.87174 0.707116 0.309554 0.437746 2.25675 140.334 83.5568 18.6998 60.691 0.00404033 0 -40 10
1.919 5.54972e-08 2.54021e-06 0.15229 0.15229 0.0120241 2.5226e-05 0.00115464 0.190363 0.000658891 0.191017 0.966263 101.336 0.233237 0.876181 4.66406 0.0667626 0.0440006 0.955999 0.0193407 0.00467503 0.0185945 0.00445282 0.00565927 0.00640549 0.226371 0.256219 58.0595 -87.8998 126.122 15.9289 145.039 0.000142641 0.267347 192.7 0.310121 0.0673162 0.00409899 0.00056249 0.00138545 0.986955 0.991714 -2.99263e-06 -85.6555 0.0930998 31165.3 312.276 0.983494 0.319146 0.739951 0.739947 9.99958 2.98729e-06 1.1949e-05 0.135049 0.983443 0.931197 -0.0132914 4.93546e-06 0.519366 -2.03964e-20 7.57377e-24 -2.03888e-20 0.00139665 0.997814 8.60362e-05 0.152757 2.85294 0.00139665 0.997815 0.80146 0.00107011 0.00188164 0.000860362 0.455349 0.00188164 0.445289 0.00013163 1.02 0.888944 0.534326 0.287804 1.7199e-07 3.08795e-09 2368.19 3146.45 -0.058936 0.48222 0.277229 0.255255 -0.592976 -0.169584 0.485293 -0.265453 -0.21985 2.821 1 0 294.682 0 2.25671 2.819 0.000298912 0.871769 0.707159 0.309518 0.437768 2.25689 140.341 83.5562 18.6998 60.6907 0.00404036 0 -40 10
1.92 5.5526e-08 2.54021e-06 0.152319 0.152319 0.0120241 2.52391e-05 0.00115464 0.190399 0.000658891 0.191053 0.966356 101.335 0.233226 0.876315 4.66476 0.0667736 0.0440072 0.955993 0.0193401 0.00467551 0.0185939 0.00445324 0.00565987 0.0064061 0.226395 0.256244 58.0596 -87.8998 126.122 15.9288 145.039 0.000142644 0.267347 192.699 0.31012 0.0673162 0.00409899 0.000562491 0.00138546 0.986955 0.991714 -2.99264e-06 -85.6555 0.0930999 31165.2 312.289 0.983494 0.319146 0.739963 0.739959 9.99958 2.98729e-06 1.19491e-05 0.135054 0.983443 0.931196 -0.0132914 4.93549e-06 0.519387 -2.03981e-20 7.57444e-24 -2.03905e-20 0.00139665 0.997814 8.60363e-05 0.152758 2.85294 0.00139665 0.997815 0.801529 0.00107013 0.00188164 0.000860363 0.455349 0.00188164 0.445294 0.000131632 1.02 0.888946 0.534326 0.287805 1.7199e-07 3.08798e-09 2368.17 3146.5 -0.0589411 0.48222 0.277229 0.255258 -0.592976 -0.169584 0.485277 -0.265451 -0.219835 2.822 1 0 294.678 0 2.25685 2.82 0.00029891 0.871799 0.707201 0.309481 0.43779 2.25702 140.349 83.5556 18.6997 60.6904 0.00404038 0 -40 10
1.921 5.55549e-08 2.54021e-06 0.152348 0.152348 0.0120241 2.52522e-05 0.00115464 0.190435 0.000658891 0.191089 0.966448 101.335 0.233215 0.87645 4.66546 0.0667845 0.0440138 0.955986 0.0193395 0.004676 0.0185933 0.00445366 0.00566047 0.00640672 0.226419 0.256269 58.0596 -87.8998 126.121 15.9288 145.039 0.000142646 0.267347 192.699 0.31012 0.0673161 0.004099 0.000562492 0.00138546 0.986955 0.991714 -2.99266e-06 -85.6555 0.0931 31165.2 312.302 0.983494 0.319146 0.739975 0.739971 9.99958 2.9873e-06 1.19491e-05 0.135059 0.983443 0.931195 -0.0132914 4.93552e-06 0.519408 -2.03998e-20 7.57512e-24 -2.03922e-20 0.00139665 0.997814 8.60364e-05 0.152758 2.85294 0.00139665 0.997815 0.801597 0.00107014 0.00188164 0.000860364 0.455349 0.00188164 0.445298 0.000131634 1.02 0.888947 0.534326 0.287807 1.7199e-07 3.088e-09 2368.16 3146.56 -0.0589462 0.48222 0.277229 0.255262 -0.592975 -0.169584 0.485261 -0.265449 -0.219821 2.823 1 0 294.673 0 2.25698 2.821 0.000298909 0.871829 0.707243 0.309445 0.437811 2.25716 140.356 83.555 18.6997 60.6901 0.00404041 0 -40 10
1.922 5.55837e-08 2.54022e-06 0.152377 0.152377 0.0120241 2.52653e-05 0.00115464 0.190471 0.000658892 0.191125 0.96654 101.334 0.233205 0.876584 4.66616 0.0667954 0.0440204 0.95598 0.0193389 0.00467648 0.0185927 0.00445408 0.00566107 0.00640734 0.226443 0.256294 58.0597 -87.8998 126.121 15.9288 145.039 0.000142648 0.267348 192.699 0.31012 0.0673161 0.004099 0.000562492 0.00138546 0.986955 0.991713 -2.99267e-06 -85.6554 0.0931001 31165.2 312.315 0.983494 0.319146 0.739988 0.739983 9.99958 2.9873e-06 1.19491e-05 0.135064 0.983443 0.931194 -0.0132914 4.93555e-06 0.51943 -2.04015e-20 7.57579e-24 -2.03939e-20 0.00139665 0.997814 8.60364e-05 0.152758 2.85294 0.00139665 0.997815 0.801666 0.00107016 0.00188164 0.000860364 0.455349 0.00188164 0.445303 0.000131637 1.02 0.888948 0.534325 0.287808 1.7199e-07 3.08802e-09 2368.14 3146.61 -0.0589513 0.48222 0.277228 0.255265 -0.592975 -0.169584 0.485245 -0.265447 -0.219807 2.824 1 0 294.669 0 2.25712 2.822 0.000298908 0.871859 0.707286 0.309409 0.437833 2.2573 140.363 83.5544 18.6997 60.6898 0.00404043 0 -40 10
1.923 5.56125e-08 2.54022e-06 0.152406 0.152405 0.0120241 2.52784e-05 0.00115464 0.190507 0.000658892 0.191162 0.966633 101.333 0.233194 0.876719 4.66686 0.0668064 0.044027 0.955973 0.0193383 0.00467697 0.018592 0.0044545 0.00566166 0.00640796 0.226467 0.256318 58.0598 -87.8998 126.121 15.9287 145.039 0.000142651 0.267348 192.699 0.310119 0.067316 0.004099 0.000562493 0.00138546 0.986955 0.991713 -2.99269e-06 -85.6554 0.0931002 31165.2 312.328 0.983494 0.319146 0.74 0.739995 9.99958 2.98731e-06 1.19491e-05 0.135069 0.983444 0.931193 -0.0132914 4.93558e-06 0.519451 -2.04032e-20 7.57647e-24 -2.03956e-20 0.00139665 0.997814 8.60365e-05 0.152758 2.85294 0.00139665 0.997815 0.801735 0.00107018 0.00188164 0.000860365 0.455348 0.00188164 0.445308 0.000131639 1.02 0.888949 0.534325 0.28781 1.71991e-07 3.08804e-09 2368.12 3146.66 -0.0589564 0.48222 0.277228 0.255268 -0.592974 -0.169584 0.485228 -0.265445 -0.219793 2.825 1 0 294.664 0 2.25725 2.823 0.000298906 0.871889 0.707328 0.309372 0.437855 2.25743 140.37 83.5538 18.6996 60.6895 0.00404046 0 -40 10
1.924 5.56414e-08 2.54022e-06 0.152435 0.152434 0.0120241 2.52915e-05 0.00115465 0.190543 0.000658893 0.191198 0.966725 101.332 0.233183 0.876854 4.66756 0.0668173 0.0440336 0.955966 0.0193377 0.00467746 0.0185914 0.00445493 0.00566226 0.00640858 0.226491 0.256343 58.0598 -87.8998 126.121 15.9287 145.039 0.000142653 0.267348 192.699 0.310119 0.067316 0.00409901 0.000562494 0.00138547 0.986955 0.991713 -2.9927e-06 -85.6554 0.0931003 31165.2 312.342 0.983494 0.319146 0.740012 0.740008 9.99958 2.98731e-06 1.19491e-05 0.135074 0.983444 0.931192 -0.0132914 4.93561e-06 0.519472 -2.04049e-20 7.57714e-24 -2.03973e-20 0.00139665 0.997814 8.60366e-05 0.152758 2.85295 0.00139665 0.997815 0.801804 0.00107019 0.00188165 0.000860366 0.455348 0.00188164 0.445313 0.000131641 1.02 0.88895 0.534325 0.287811 1.71991e-07 3.08807e-09 2368.11 3146.71 -0.0589616 0.48222 0.277228 0.255271 -0.592973 -0.169584 0.485212 -0.265443 -0.219779 2.826 1 0 294.659 0 2.25739 2.824 0.000298905 0.871919 0.707371 0.309336 0.437877 2.25757 140.378 83.5532 18.6996 60.6892 0.00404048 0 -40 10
1.925 5.56702e-08 2.54022e-06 0.152463 0.152463 0.012024 2.53046e-05 0.00115465 0.190579 0.000658893 0.191234 0.966817 101.332 0.233172 0.876988 4.66826 0.0668283 0.0440402 0.95596 0.0193371 0.00467794 0.0185908 0.00445535 0.00566286 0.0064092 0.226514 0.256368 58.0599 -87.8998 126.121 15.9286 145.039 0.000142655 0.267348 192.699 0.310118 0.0673159 0.00409901 0.000562494 0.00138547 0.986955 0.991713 -2.99272e-06 -85.6554 0.0931004 31165.1 312.355 0.983494 0.319146 0.740024 0.74002 9.99958 2.98732e-06 1.19492e-05 0.135079 0.983444 0.931191 -0.0132914 4.93564e-06 0.519493 -2.04066e-20 7.57782e-24 -2.0399e-20 0.00139665 0.997814 8.60367e-05 0.152758 2.85295 0.00139665 0.997815 0.801872 0.00107021 0.00188165 0.000860367 0.455348 0.00188165 0.445317 0.000131644 1.02 0.888951 0.534325 0.287813 1.71991e-07 3.08809e-09 2368.09 3146.76 -0.0589667 0.48222 0.277228 0.255275 -0.592973 -0.169584 0.485196 -0.265441 -0.219765 2.827 1 0 294.655 0 2.25753 2.825 0.000298904 0.871949 0.707413 0.3093 0.437899 2.2577 140.385 83.5526 18.6995 60.6889 0.00404051 0 -40 10
1.926 5.5699e-08 2.54022e-06 0.152492 0.152492 0.012024 2.53177e-05 0.00115465 0.190615 0.000658894 0.19127 0.966909 101.331 0.233161 0.877123 4.66896 0.0668392 0.0440468 0.955953 0.0193365 0.00467843 0.0185902 0.00445577 0.00566346 0.00640982 0.226538 0.256393 58.06 -87.8998 126.12 15.9286 145.039 0.000142658 0.267348 192.698 0.310118 0.0673159 0.00409901 0.000562495 0.00138547 0.986955 0.991713 -2.99273e-06 -85.6554 0.0931004 31165.1 312.368 0.983494 0.319146 0.740037 0.740032 9.99958 2.98732e-06 1.19492e-05 0.135084 0.983444 0.93119 -0.0132914 4.93567e-06 0.519514 -2.04083e-20 7.57849e-24 -2.04007e-20 0.00139666 0.997814 8.60368e-05 0.152759 2.85295 0.00139666 0.997815 0.801941 0.00107022 0.00188165 0.000860368 0.455348 0.00188165 0.445322 0.000131646 1.02 0.888952 0.534324 0.287814 1.71991e-07 3.08811e-09 2368.07 3146.81 -0.0589718 0.482221 0.277227 0.255278 -0.592972 -0.169584 0.48518 -0.265439 -0.21975 2.828 1 0 294.65 0 2.25766 2.826 0.000298902 0.871979 0.707456 0.309264 0.43792 2.25784 140.392 83.552 18.6995 60.6887 0.00404053 0 -40 10
1.927 5.57278e-08 2.54022e-06 0.152521 0.152521 0.012024 2.53308e-05 0.00115465 0.190651 0.000658894 0.191305 0.967002 101.33 0.23315 0.877257 4.66966 0.0668502 0.0440534 0.955947 0.0193359 0.00467891 0.0185896 0.00445619 0.00566406 0.00641044 0.226562 0.256418 58.06 -87.8998 126.12 15.9286 145.039 0.00014266 0.267349 192.698 0.310117 0.0673158 0.00409901 0.000562496 0.00138547 0.986955 0.991713 -2.99275e-06 -85.6554 0.0931005 31165.1 312.381 0.983494 0.319146 0.740049 0.740044 9.99958 2.98733e-06 1.19492e-05 0.135089 0.983444 0.931189 -0.0132914 4.9357e-06 0.519536 -2.041e-20 7.57917e-24 -2.04024e-20 0.00139666 0.997814 8.60368e-05 0.152759 2.85295 0.00139666 0.997815 0.80201 0.00107024 0.00188165 0.000860368 0.455347 0.00188165 0.445327 0.000131648 1.02 0.888953 0.534324 0.287816 1.71992e-07 3.08814e-09 2368.06 3146.86 -0.0589769 0.482221 0.277227 0.255281 -0.592971 -0.169584 0.485163 -0.265436 -0.219736 2.829 1 0 294.645 0 2.2578 2.827 0.000298901 0.872009 0.707498 0.309228 0.437942 2.25797 140.4 83.5514 18.6995 60.6884 0.00404056 0 -40 10
1.928 5.57567e-08 2.54023e-06 0.15255 0.152549 0.012024 2.53439e-05 0.00115465 0.190687 0.000658894 0.191341 0.967094 101.33 0.233139 0.877392 4.67036 0.0668611 0.04406 0.95594 0.0193353 0.0046794 0.0185889 0.00445661 0.00566466 0.00641106 0.226586 0.256442 58.0601 -87.8998 126.12 15.9285 145.039 0.000142662 0.267349 192.698 0.310117 0.0673158 0.00409902 0.000562496 0.00138547 0.986955 0.991713 -2.99276e-06 -85.6554 0.0931006 31165.1 312.395 0.983494 0.319146 0.740061 0.740057 9.99958 2.98733e-06 1.19492e-05 0.135094 0.983444 0.931188 -0.0132913 4.93573e-06 0.519557 -2.04117e-20 7.57984e-24 -2.04041e-20 0.00139666 0.997814 8.60369e-05 0.152759 2.85295 0.00139666 0.997815 0.802078 0.00107025 0.00188165 0.000860369 0.455347 0.00188165 0.445332 0.00013165 1.02 0.888954 0.534324 0.287817 1.71992e-07 3.08816e-09 2368.04 3146.92 -0.058982 0.482221 0.277227 0.255284 -0.592971 -0.169584 0.485147 -0.265434 -0.219722 2.83 1 0 294.641 0 2.25793 2.828 0.0002989 0.872039 0.707541 0.309192 0.437964 2.25811 140.407 83.5508 18.6994 60.6881 0.00404058 0 -40 10
1.929 5.57855e-08 2.54023e-06 0.152578 0.152578 0.012024 2.5357e-05 0.00115465 0.190723 0.000658895 0.191377 0.967186 101.329 0.233128 0.877527 4.67107 0.066872 0.0440667 0.955933 0.0193347 0.00467988 0.0185883 0.00445704 0.00566526 0.00641168 0.22661 0.256467 58.0601 -87.8998 126.12 15.9285 145.039 0.000142665 0.267349 192.698 0.310117 0.0673157 0.00409902 0.000562497 0.00138548 0.986955 0.991713 -2.99278e-06 -85.6554 0.0931007 31165 312.408 0.983494 0.319146 0.740073 0.740069 9.99958 2.98734e-06 1.19492e-05 0.135098 0.983445 0.931187 -0.0132913 4.93576e-06 0.519578 -2.04133e-20 7.58052e-24 -2.04058e-20 0.00139666 0.997814 8.6037e-05 0.152759 2.85295 0.00139666 0.997815 0.802147 0.00107027 0.00188165 0.00086037 0.455347 0.00188165 0.445337 0.000131653 1.02 0.888955 0.534323 0.287819 1.71992e-07 3.08818e-09 2368.03 3146.97 -0.0589872 0.482221 0.277227 0.255288 -0.59297 -0.169584 0.485131 -0.265432 -0.219708 2.831 1 0 294.636 0 2.25807 2.829 0.000298898 0.872069 0.707583 0.309155 0.437986 2.25824 140.414 83.5502 18.6994 60.6878 0.00404061 0 -40 10
1.93 5.58143e-08 2.54023e-06 0.152607 0.152607 0.012024 2.53701e-05 0.00115465 0.190759 0.000658895 0.191413 0.967279 101.328 0.233117 0.877661 4.67177 0.066883 0.0440733 0.955927 0.0193341 0.00468037 0.0185877 0.00445746 0.00566586 0.0064123 0.226634 0.256492 58.0602 -87.8998 126.119 15.9285 145.039 0.000142667 0.267349 192.698 0.310116 0.0673157 0.00409902 0.000562498 0.00138548 0.986955 0.991713 -2.99279e-06 -85.6554 0.0931008 31165 312.421 0.983494 0.319146 0.740086 0.740081 9.99958 2.98734e-06 1.19493e-05 0.135103 0.983445 0.931186 -0.0132913 4.93579e-06 0.519599 -2.0415e-20 7.58119e-24 -2.04075e-20 0.00139666 0.997814 8.60371e-05 0.152759 2.85295 0.00139666 0.997815 0.802215 0.00107029 0.00188166 0.000860371 0.455347 0.00188165 0.445341 0.000131655 1.02 0.888957 0.534323 0.28782 1.71993e-07 3.0882e-09 2368.01 3147.02 -0.0589923 0.482221 0.277226 0.255291 -0.592969 -0.169584 0.485115 -0.26543 -0.219694 2.832 1 0 294.632 0 2.2582 2.83 0.000298897 0.872099 0.707625 0.309119 0.438008 2.25838 140.421 83.5496 18.6994 60.6875 0.00404063 0 -40 10
1.931 5.58431e-08 2.54023e-06 0.152636 0.152635 0.012024 2.53832e-05 0.00115465 0.190795 0.000658896 0.191449 0.967371 101.328 0.233106 0.877796 4.67247 0.0668939 0.0440799 0.95592 0.0193335 0.00468086 0.0185871 0.00445788 0.00566646 0.00641292 0.226658 0.256517 58.0603 -87.8998 126.119 15.9284 145.039 0.000142669 0.267349 192.698 0.310116 0.0673156 0.00409903 0.000562498 0.00138548 0.986955 0.991713 -2.99281e-06 -85.6554 0.0931009 31165 312.434 0.983494 0.319146 0.740098 0.740093 9.99958 2.98735e-06 1.19493e-05 0.135108 0.983445 0.931185 -0.0132913 4.93582e-06 0.519621 -2.04167e-20 7.58187e-24 -2.04092e-20 0.00139666 0.997814 8.60372e-05 0.152759 2.85295 0.00139666 0.997815 0.802284 0.0010703 0.00188166 0.000860372 0.455347 0.00188166 0.445346 0.000131657 1.02 0.888958 0.534323 0.287822 1.71993e-07 3.08823e-09 2367.99 3147.07 -0.0589974 0.482221 0.277226 0.255294 -0.592969 -0.169584 0.485098 -0.265428 -0.21968 2.833 1 0 294.627 0 2.25834 2.831 0.000298896 0.872129 0.707668 0.309083 0.438029 2.25851 140.429 83.549 18.6993 60.6872 0.00404066 0 -40 10
1.932 5.5872e-08 2.54023e-06 0.152664 0.152664 0.012024 2.53963e-05 0.00115465 0.19083 0.000658896 0.191485 0.967464 101.327 0.233095 0.877931 4.67318 0.0669049 0.0440866 0.955913 0.0193329 0.00468134 0.0185865 0.0044583 0.00566706 0.00641354 0.226682 0.256542 58.0603 -87.8998 126.119 15.9284 145.039 0.000142672 0.267349 192.697 0.310115 0.0673156 0.00409903 0.000562499 0.00138548 0.986955 0.991713 -2.99282e-06 -85.6554 0.093101 31165 312.447 0.983494 0.319146 0.74011 0.740106 9.99958 2.98735e-06 1.19493e-05 0.135113 0.983445 0.931184 -0.0132913 4.93585e-06 0.519642 -2.04184e-20 7.58255e-24 -2.04109e-20 0.00139666 0.997814 8.60372e-05 0.152759 2.85295 0.00139666 0.997815 0.802352 0.00107032 0.00188166 0.000860372 0.455346 0.00188166 0.445351 0.00013166 1.02 0.888959 0.534322 0.287823 1.71993e-07 3.08825e-09 2367.98 3147.12 -0.0590025 0.482221 0.277226 0.255298 -0.592968 -0.169584 0.485082 -0.265426 -0.219665 2.834 1 0 294.622 0 2.25847 2.832 0.000298894 0.872159 0.70771 0.309047 0.438051 2.25865 140.436 83.5484 18.6993 60.6869 0.00404068 0 -40 10
1.933 5.59008e-08 2.54024e-06 0.152693 0.152693 0.0120239 2.54095e-05 0.00115465 0.190866 0.000658896 0.19152 0.967556 101.326 0.233084 0.878065 4.67388 0.0669158 0.0440932 0.955907 0.0193323 0.00468183 0.0185858 0.00445873 0.00566766 0.00641416 0.226706 0.256567 58.0604 -87.8998 126.119 15.9284 145.04 0.000142674 0.26735 192.697 0.310115 0.0673155 0.00409903 0.0005625 0.00138548 0.986955 0.991713 -2.99284e-06 -85.6553 0.0931011 31165 312.461 0.983494 0.319146 0.740122 0.740118 9.99958 2.98735e-06 1.19493e-05 0.135118 0.983445 0.931183 -0.0132913 4.93588e-06 0.519663 -2.04201e-20 7.58323e-24 -2.04126e-20 0.00139666 0.997814 8.60373e-05 0.15276 2.85295 0.00139666 0.997815 0.802421 0.00107033 0.00188166 0.000860373 0.455346 0.00188166 0.445356 0.000131662 1.02 0.88896 0.534322 0.287825 1.71993e-07 3.08827e-09 2367.96 3147.17 -0.0590077 0.482221 0.277225 0.255301 -0.592967 -0.169585 0.485066 -0.265424 -0.219651 2.835 1 0 294.618 0 2.25861 2.833 0.000298893 0.872189 0.707753 0.309011 0.438073 2.25878 140.443 83.5478 18.6993 60.6866 0.00404071 0 -40 10
1.934 5.59296e-08 2.54024e-06 0.152722 0.152721 0.0120239 2.54226e-05 0.00115465 0.190902 0.000658897 0.191556 0.967648 101.325 0.233073 0.8782 4.67459 0.0669268 0.0440999 0.9559 0.0193317 0.00468232 0.0185852 0.00445915 0.00566826 0.00641479 0.22673 0.256591 58.0604 -87.8998 126.119 15.9283 145.04 0.000142677 0.26735 192.697 0.310114 0.0673155 0.00409904 0.0005625 0.00138549 0.986955 0.991713 -2.99285e-06 -85.6553 0.0931011 31164.9 312.474 0.983494 0.319146 0.740135 0.74013 9.99958 2.98736e-06 1.19493e-05 0.135123 0.983445 0.931182 -0.0132913 4.9359e-06 0.519684 -2.04218e-20 7.5839e-24 -2.04143e-20 0.00139666 0.997814 8.60374e-05 0.15276 2.85295 0.00139666 0.997815 0.802489 0.00107035 0.00188166 0.000860374 0.455346 0.00188166 0.44536 0.000131664 1.02 0.888961 0.534322 0.287826 1.71994e-07 3.0883e-09 2367.94 3147.22 -0.0590128 0.482221 0.277225 0.255304 -0.592967 -0.169585 0.48505 -0.265422 -0.219637 2.836 1 0 294.613 0 2.25874 2.834 0.000298891 0.872219 0.707795 0.308975 0.438095 2.25892 140.45 83.5472 18.6992 60.6863 0.00404073 0 -40 10
1.935 5.59584e-08 2.54024e-06 0.15275 0.15275 0.0120239 2.54357e-05 0.00115465 0.190938 0.000658897 0.191592 0.967741 101.325 0.233062 0.878335 4.67529 0.0669377 0.0441065 0.955893 0.0193311 0.00468281 0.0185846 0.00445957 0.00566886 0.00641541 0.226754 0.256616 58.0605 -87.8998 126.118 15.9283 145.04 0.000142679 0.26735 192.697 0.310114 0.0673154 0.00409904 0.000562501 0.00138549 0.986955 0.991713 -2.99287e-06 -85.6553 0.0931012 31164.9 312.487 0.983494 0.319146 0.740147 0.740142 9.99958 2.98736e-06 1.19494e-05 0.135128 0.983445 0.931181 -0.0132913 4.93593e-06 0.519706 -2.04235e-20 7.58458e-24 -2.04159e-20 0.00139667 0.997814 8.60375e-05 0.15276 2.85296 0.00139667 0.997815 0.802558 0.00107036 0.00188166 0.000860375 0.455346 0.00188166 0.445365 0.000131666 1.02 0.888962 0.534321 0.287828 1.71994e-07 3.08832e-09 2367.93 3147.27 -0.0590179 0.482221 0.277225 0.255307 -0.592966 -0.169585 0.485033 -0.26542 -0.219623 2.837 1 0 294.609 0 2.25888 2.835 0.00029889 0.872249 0.707837 0.308939 0.438117 2.25906 140.458 83.5466 18.6992 60.686 0.00404076 0 -40 10
1.936 5.59873e-08 2.54024e-06 0.152779 0.152778 0.0120239 2.54488e-05 0.00115466 0.190973 0.000658898 0.191628 0.967833 101.324 0.233051 0.878469 4.676 0.0669487 0.0441132 0.955887 0.0193305 0.00468329 0.018584 0.00446 0.00566946 0.00641603 0.226779 0.256641 58.0606 -87.8998 126.118 15.9282 145.04 0.000142681 0.26735 192.697 0.310114 0.0673153 0.00409904 0.000562502 0.00138549 0.986955 0.991713 -2.99288e-06 -85.6553 0.0931013 31164.9 312.5 0.983494 0.319146 0.740159 0.740155 9.99958 2.98737e-06 1.19494e-05 0.135133 0.983446 0.93118 -0.0132913 4.93596e-06 0.519727 -2.04252e-20 7.58526e-24 -2.04176e-20 0.00139667 0.997814 8.60376e-05 0.15276 2.85296 0.00139667 0.997815 0.802626 0.00107038 0.00188166 0.000860376 0.455345 0.00188166 0.44537 0.000131669 1.02 0.888963 0.534321 0.287829 1.71994e-07 3.08834e-09 2367.91 3147.33 -0.059023 0.482221 0.277225 0.255311 -0.592966 -0.169585 0.485017 -0.265418 -0.219609 2.838 1 0 294.604 0 2.25901 2.836 0.000298889 0.872279 0.70788 0.308903 0.438138 2.25919 140.465 83.546 18.6992 60.6858 0.00404078 0 -40 10
1.937 5.60161e-08 2.54024e-06 0.152807 0.152807 0.0120239 2.54619e-05 0.00115466 0.191009 0.000658898 0.191663 0.967926 101.323 0.23304 0.878604 4.67671 0.0669596 0.0441199 0.95588 0.0193299 0.00468378 0.0185833 0.00446042 0.00567006 0.00641665 0.226803 0.256666 58.0606 -87.8998 126.118 15.9282 145.04 0.000142684 0.26735 192.697 0.310113 0.0673153 0.00409904 0.000562502 0.00138549 0.986955 0.991713 -2.9929e-06 -85.6553 0.0931014 31164.9 312.514 0.983494 0.319146 0.740171 0.740167 9.99958 2.98737e-06 1.19494e-05 0.135138 0.983446 0.931179 -0.0132913 4.93599e-06 0.519748 -2.04269e-20 7.58594e-24 -2.04193e-20 0.00139667 0.997814 8.60376e-05 0.15276 2.85296 0.00139667 0.997815 0.802695 0.0010704 0.00188167 0.000860376 0.455345 0.00188166 0.445375 0.000131671 1.02 0.888964 0.534321 0.287831 1.71994e-07 3.08836e-09 2367.9 3147.38 -0.0590281 0.482221 0.277224 0.255314 -0.592965 -0.169585 0.485001 -0.265416 -0.219595 2.839 1 0 294.599 0 2.25915 2.837 0.000298887 0.872309 0.707922 0.308867 0.43816 2.25933 140.472 83.5454 18.6991 60.6855 0.00404081 0 -40 10
1.938 5.60449e-08 2.54025e-06 0.152836 0.152835 0.0120239 2.5475e-05 0.00115466 0.191045 0.000658899 0.191699 0.968018 101.323 0.233029 0.878739 4.67741 0.0669706 0.0441265 0.955873 0.0193293 0.00468427 0.0185827 0.00446084 0.00567067 0.00641728 0.226827 0.256691 58.0607 -87.8998 126.118 15.9282 145.04 0.000142686 0.267351 192.697 0.310113 0.0673152 0.00409905 0.000562503 0.0013855 0.986955 0.991713 -2.99291e-06 -85.6553 0.0931015 31164.8 312.527 0.983494 0.319146 0.740183 0.740179 9.99958 2.98738e-06 1.19494e-05 0.135143 0.983446 0.931178 -0.0132913 4.93602e-06 0.51977 -2.04286e-20 7.58661e-24 -2.0421e-20 0.00139667 0.997814 8.60377e-05 0.15276 2.85296 0.00139667 0.997815 0.802763 0.00107041 0.00188167 0.000860377 0.455345 0.00188167 0.445379 0.000131673 1.02 0.888965 0.534321 0.287833 1.71995e-07 3.08839e-09 2367.88 3147.43 -0.0590333 0.482221 0.277224 0.255317 -0.592964 -0.169585 0.484984 -0.265413 -0.21958 2.84 1 0 294.595 0 2.25929 2.838 0.000298886 0.872339 0.707965 0.308831 0.438182 2.25946 140.48 83.5448 18.6991 60.6852 0.00404083 0 -40 10
1.939 5.60737e-08 2.54025e-06 0.152864 0.152864 0.0120239 2.54881e-05 0.00115466 0.19108 0.000658899 0.191734 0.968111 101.322 0.233018 0.878873 4.67812 0.0669816 0.0441332 0.955867 0.0193287 0.00468476 0.0185821 0.00446127 0.00567127 0.0064179 0.226851 0.256716 58.0608 -87.8998 126.117 15.9281 145.04 0.000142688 0.267351 192.696 0.310112 0.0673152 0.00409905 0.000562504 0.0013855 0.986955 0.991713 -2.99293e-06 -85.6553 0.0931016 31164.8 312.54 0.983494 0.319146 0.740196 0.740191 9.99958 2.98738e-06 1.19494e-05 0.135148 0.983446 0.931177 -0.0132913 4.93605e-06 0.519791 -2.04303e-20 7.58729e-24 -2.04228e-20 0.00139667 0.997814 8.60378e-05 0.152761 2.85296 0.00139667 0.997815 0.802831 0.00107043 0.00188167 0.000860378 0.455345 0.00188167 0.445384 0.000131675 1.02 0.888966 0.53432 0.287834 1.71995e-07 3.08841e-09 2367.86 3147.48 -0.0590384 0.482222 0.277224 0.255321 -0.592964 -0.169585 0.484968 -0.265411 -0.219566 2.841 1 0 294.59 0 2.25942 2.839 0.000298885 0.872369 0.708007 0.308795 0.438204 2.2596 140.487 83.5442 18.6991 60.6849 0.00404086 0 -40 10
1.94 5.61026e-08 2.54025e-06 0.152893 0.152892 0.0120238 2.55012e-05 0.00115466 0.191116 0.000658899 0.19177 0.968203 101.321 0.233007 0.879008 4.67883 0.0669925 0.0441399 0.95586 0.0193281 0.00468524 0.0185815 0.00446169 0.00567187 0.00641852 0.226875 0.256741 58.0608 -87.8998 126.117 15.9281 145.04 0.000142691 0.267351 192.696 0.310112 0.0673151 0.00409905 0.000562504 0.0013855 0.986955 0.991713 -2.99294e-06 -85.6553 0.0931017 31164.8 312.553 0.983494 0.319146 0.740208 0.740204 9.99958 2.98739e-06 1.19495e-05 0.135153 0.983446 0.931176 -0.0132913 4.93608e-06 0.519812 -2.0432e-20 7.58797e-24 -2.04245e-20 0.00139667 0.997814 8.60379e-05 0.152761 2.85296 0.00139667 0.997815 0.8029 0.00107044 0.00188167 0.000860379 0.455344 0.00188167 0.445389 0.000131678 1.02 0.888967 0.53432 0.287836 1.71995e-07 3.08843e-09 2367.85 3147.53 -0.0590435 0.482222 0.277223 0.255324 -0.592963 -0.169585 0.484952 -0.265409 -0.219552 2.842 1 0 294.585 0 2.25956 2.84 0.000298883 0.872399 0.708049 0.30876 0.438225 2.25973 140.494 83.5436 18.699 60.6846 0.00404088 0 -40 10
1.941 5.61314e-08 2.54025e-06 0.152921 0.152921 0.0120238 2.55143e-05 0.00115466 0.191151 0.0006589 0.191806 0.968296 101.32 0.232997 0.879143 4.67954 0.0670035 0.0441466 0.955853 0.0193275 0.00468573 0.0185809 0.00446212 0.00567247 0.00641914 0.226899 0.256766 58.0609 -87.8998 126.117 15.9281 145.04 0.000142693 0.267351 192.696 0.310111 0.0673151 0.00409906 0.000562505 0.0013855 0.986955 0.991713 -2.99296e-06 -85.6553 0.0931018 31164.8 312.567 0.983494 0.319146 0.74022 0.740216 9.99958 2.98739e-06 1.19495e-05 0.135158 0.983446 0.931175 -0.0132913 4.93611e-06 0.519834 -2.04337e-20 7.58865e-24 -2.04262e-20 0.00139667 0.997814 8.6038e-05 0.152761 2.85296 0.00139667 0.997815 0.802968 0.00107046 0.00188167 0.00086038 0.455344 0.00188167 0.445394 0.00013168 1.02 0.888969 0.53432 0.287837 1.71996e-07 3.08846e-09 2367.83 3147.58 -0.0590487 0.482222 0.277223 0.255327 -0.592962 -0.169585 0.484936 -0.265407 -0.219538 2.843 1 0 294.581 0 2.25969 2.841 0.000298882 0.872429 0.708092 0.308724 0.438247 2.25987 140.501 83.543 18.699 60.6843 0.00404091 0 -40 10
1.942 5.61602e-08 2.54025e-06 0.152949 0.152949 0.0120238 2.55274e-05 0.00115466 0.191187 0.0006589 0.191841 0.968388 101.32 0.232986 0.879278 4.68024 0.0670144 0.0441533 0.955847 0.0193269 0.00468622 0.0185802 0.00446254 0.00567308 0.00641977 0.226923 0.256791 58.0609 -87.8998 126.117 15.928 145.04 0.000142695 0.267351 192.696 0.310111 0.067315 0.00409906 0.000562506 0.0013855 0.986954 0.991713 -2.99297e-06 -85.6553 0.0931018 31164.7 312.58 0.983494 0.319146 0.740232 0.740228 9.99958 2.9874e-06 1.19495e-05 0.135163 0.983447 0.931173 -0.0132913 4.93614e-06 0.519855 -2.04354e-20 7.58933e-24 -2.04279e-20 0.00139667 0.997814 8.6038e-05 0.152761 2.85296 0.00139667 0.997815 0.803036 0.00107047 0.00188167 0.00086038 0.455344 0.00188167 0.445398 0.000131682 1.02 0.88897 0.534319 0.287839 1.71996e-07 3.08848e-09 2367.81 3147.63 -0.0590538 0.482222 0.277223 0.25533 -0.592962 -0.169585 0.484919 -0.265405 -0.219524 2.844 1 0 294.576 0 2.25983 2.842 0.00029888 0.872459 0.708134 0.308688 0.438269 2.26 140.509 83.5424 18.699 60.684 0.00404093 0 -40 10
1.943 5.61891e-08 2.54025e-06 0.152978 0.152977 0.0120238 2.55405e-05 0.00115466 0.191222 0.000658901 0.191877 0.968481 101.319 0.232975 0.879412 4.68095 0.0670254 0.0441599 0.95584 0.0193263 0.00468671 0.0185796 0.00446297 0.00567368 0.00642039 0.226947 0.256816 58.061 -87.8999 126.117 15.928 145.04 0.000142698 0.267352 192.696 0.310111 0.067315 0.00409906 0.000562506 0.00138551 0.986954 0.991713 -2.99299e-06 -85.6552 0.0931019 31164.7 312.593 0.983494 0.319146 0.740245 0.74024 9.99958 2.9874e-06 1.19495e-05 0.135168 0.983447 0.931172 -0.0132913 4.93617e-06 0.519876 -2.04372e-20 7.59001e-24 -2.04296e-20 0.00139667 0.997814 8.60381e-05 0.152761 2.85296 0.00139667 0.997815 0.803105 0.00107049 0.00188167 0.000860381 0.455344 0.00188167 0.445403 0.000131685 1.02 0.888971 0.534319 0.28784 1.71996e-07 3.0885e-09 2367.8 3147.69 -0.0590589 0.482222 0.277223 0.255334 -0.592961 -0.169585 0.484903 -0.265403 -0.219509 2.845 1 0 294.572 0 2.25996 2.843 0.000298879 0.872489 0.708177 0.308652 0.438291 2.26014 140.516 83.5418 18.6989 60.6837 0.00404096 0 -40 10
1.944 5.62179e-08 2.54026e-06 0.153006 0.153006 0.0120238 2.55536e-05 0.00115466 0.191258 0.000658901 0.191912 0.968573 101.318 0.232964 0.879547 4.68166 0.0670363 0.0441666 0.955833 0.0193257 0.0046872 0.018579 0.00446339 0.00567428 0.00642102 0.226971 0.256841 58.0611 -87.8999 126.116 15.9279 145.04 0.0001427 0.267352 192.696 0.31011 0.0673149 0.00409907 0.000562507 0.00138551 0.986954 0.991713 -2.993e-06 -85.6552 0.093102 31164.7 312.607 0.983494 0.319146 0.740257 0.740253 9.99958 2.98741e-06 1.19495e-05 0.135173 0.983447 0.931171 -0.0132913 4.9362e-06 0.519898 -2.04389e-20 7.59069e-24 -2.04313e-20 0.00139668 0.997814 8.60382e-05 0.152761 2.85296 0.00139668 0.997815 0.803173 0.0010705 0.00188168 0.000860382 0.455344 0.00188167 0.445408 0.000131687 1.02 0.888972 0.534319 0.287842 1.71996e-07 3.08852e-09 2367.78 3147.74 -0.059064 0.482222 0.277222 0.255337 -0.59296 -0.169585 0.484887 -0.265401 -0.219495 2.846 1 0 294.567 0 2.2601 2.844 0.000298878 0.872519 0.708219 0.308616 0.438313 2.26027 140.523 83.5412 18.6989 60.6834 0.00404098 0 -40 10
1.945 5.62467e-08 2.54026e-06 0.153035 0.153034 0.0120238 2.55667e-05 0.00115466 0.191293 0.000658902 0.191947 0.968666 101.318 0.232953 0.879682 4.68237 0.0670473 0.0441733 0.955827 0.0193251 0.00468769 0.0185784 0.00446381 0.00567488 0.00642164 0.226995 0.256866 58.0611 -87.8999 126.116 15.9279 145.04 0.000142703 0.267352 192.695 0.31011 0.0673149 0.00409907 0.000562508 0.00138551 0.986954 0.991713 -2.99302e-06 -85.6552 0.0931021 31164.7 312.62 0.983494 0.319146 0.740269 0.740265 9.99958 2.98741e-06 1.19495e-05 0.135178 0.983447 0.93117 -0.0132913 4.93623e-06 0.519919 -2.04406e-20 7.59137e-24 -2.0433e-20 0.00139668 0.997814 8.60383e-05 0.152761 2.85296 0.00139668 0.997815 0.803241 0.00107052 0.00188168 0.000860383 0.455343 0.00188168 0.445413 0.000131689 1.02 0.888973 0.534318 0.287843 1.71997e-07 3.08855e-09 2367.77 3147.79 -0.0590692 0.482222 0.277222 0.25534 -0.59296 -0.169585 0.484871 -0.265399 -0.219481 2.847 1 0 294.562 0 2.26023 2.845 0.000298876 0.872549 0.708261 0.30858 0.438334 2.26041 140.53 83.5406 18.6988 60.6831 0.00404101 0 -40 10
1.946 5.62755e-08 2.54026e-06 0.153063 0.153062 0.0120238 2.55798e-05 0.00115466 0.191329 0.000658902 0.191983 0.968758 101.317 0.232942 0.879817 4.68308 0.0670583 0.04418 0.95582 0.0193245 0.00468818 0.0185777 0.00446424 0.00567549 0.00642227 0.227019 0.256891 58.0612 -87.8999 126.116 15.9279 145.04 0.000142705 0.267352 192.695 0.310109 0.0673148 0.00409907 0.000562508 0.00138551 0.986954 0.991713 -2.99303e-06 -85.6552 0.0931022 31164.7 312.633 0.983494 0.319146 0.740281 0.740277 9.99958 2.98742e-06 1.19496e-05 0.135183 0.983447 0.931169 -0.0132913 4.93626e-06 0.519941 -2.04423e-20 7.59205e-24 -2.04347e-20 0.00139668 0.997814 8.60384e-05 0.152762 2.85297 0.00139668 0.997815 0.803309 0.00107054 0.00188168 0.000860384 0.455343 0.00188168 0.445417 0.000131691 1.02 0.888974 0.534318 0.287845 1.71997e-07 3.08857e-09 2367.75 3147.84 -0.0590743 0.482222 0.277222 0.255344 -0.592959 -0.169585 0.484854 -0.265397 -0.219467 2.848 1 0 294.558 0 2.26037 2.846 0.000298875 0.872579 0.708304 0.308545 0.438356 2.26054 140.538 83.54 18.6988 60.6828 0.00404103 0 -40 10
1.947 5.63044e-08 2.54026e-06 0.153091 0.153091 0.0120237 2.55929e-05 0.00115466 0.191364 0.000658902 0.192018 0.968851 101.316 0.232931 0.879952 4.68379 0.0670692 0.0441867 0.955813 0.0193239 0.00468867 0.0185771 0.00446467 0.00567609 0.00642289 0.227044 0.256916 58.0613 -87.8999 126.116 15.9278 145.04 0.000142707 0.267352 192.695 0.310109 0.0673148 0.00409907 0.000562509 0.00138552 0.986954 0.991713 -2.99305e-06 -85.6552 0.0931023 31164.6 312.647 0.983494 0.319146 0.740294 0.740289 9.99958 2.98742e-06 1.19496e-05 0.135188 0.983447 0.931168 -0.0132913 4.93629e-06 0.519962 -2.0444e-20 7.59273e-24 -2.04364e-20 0.00139668 0.997814 8.60384e-05 0.152762 2.85297 0.00139668 0.997815 0.803377 0.00107055 0.00188168 0.000860384 0.455343 0.00188168 0.445422 0.000131694 1.02 0.888975 0.534318 0.287846 1.71997e-07 3.08859e-09 2367.73 3147.89 -0.0590794 0.482222 0.277222 0.255347 -0.592958 -0.169585 0.484838 -0.265395 -0.219453 2.849 1 0 294.553 0 2.2605 2.847 0.000298874 0.872609 0.708346 0.308509 0.438378 2.26068 140.545 83.5393 18.6988 60.6826 0.00404106 0 -40 10
1.948 5.63332e-08 2.54026e-06 0.153119 0.153119 0.0120237 2.5606e-05 0.00115467 0.191399 0.000658903 0.192054 0.968943 101.315 0.23292 0.880086 4.68451 0.0670802 0.0441935 0.955807 0.0193233 0.00468915 0.0185765 0.00446509 0.00567669 0.00642352 0.227068 0.256941 58.0613 -87.8999 126.115 15.9278 145.04 0.00014271 0.267353 192.695 0.310108 0.0673147 0.00409908 0.00056251 0.00138552 0.986954 0.991713 -2.99306e-06 -85.6552 0.0931024 31164.6 312.66 0.983494 0.319146 0.740306 0.740302 9.99958 2.98743e-06 1.19496e-05 0.135193 0.983447 0.931167 -0.0132913 4.93632e-06 0.519983 -2.04457e-20 7.59341e-24 -2.04381e-20 0.00139668 0.997814 8.60385e-05 0.152762 2.85297 0.00139668 0.997815 0.803446 0.00107057 0.00188168 0.000860385 0.455343 0.00188168 0.445427 0.000131696 1.02 0.888976 0.534317 0.287848 1.71997e-07 3.08862e-09 2367.72 3147.94 -0.0590845 0.482222 0.277221 0.25535 -0.592958 -0.169585 0.484822 -0.265393 -0.219438 2.85 1 0 294.548 0 2.26064 2.848 0.000298872 0.872639 0.708388 0.308473 0.4384 2.26081 140.552 83.5387 18.6987 60.6823 0.00404108 0 -40 10
1.949 5.6362e-08 2.54027e-06 0.153148 0.153147 0.0120237 2.56191e-05 0.00115467 0.191435 0.000658903 0.192089 0.969036 101.315 0.232909 0.880221 4.68522 0.0670912 0.0442002 0.9558 0.0193227 0.00468964 0.0185759 0.00446552 0.0056773 0.00642414 0.227092 0.256966 58.0614 -87.8999 126.115 15.9278 145.04 0.000142712 0.267353 192.695 0.310108 0.0673147 0.00409908 0.00056251 0.00138552 0.986954 0.991713 -2.99308e-06 -85.6552 0.0931025 31164.6 312.673 0.983494 0.319146 0.740318 0.740314 9.99958 2.98743e-06 1.19496e-05 0.135198 0.983448 0.931166 -0.0132913 4.93635e-06 0.520005 -2.04474e-20 7.59409e-24 -2.04398e-20 0.00139668 0.997814 8.60386e-05 0.152762 2.85297 0.00139668 0.997815 0.803514 0.00107058 0.00188168 0.000860386 0.455342 0.00188168 0.445431 0.000131698 1.02 0.888977 0.534317 0.287849 1.71998e-07 3.08864e-09 2367.7 3147.99 -0.0590897 0.482222 0.277221 0.255354 -0.592957 -0.169586 0.484805 -0.26539 -0.219424 2.851 1 0 294.544 0 2.26077 2.849 0.000298871 0.872669 0.708431 0.308438 0.438421 2.26095 140.559 83.5381 18.6987 60.682 0.00404111 0 -40 10
1.95 5.63908e-08 2.54027e-06 0.153176 0.153175 0.0120237 2.56322e-05 0.00115467 0.19147 0.000658904 0.192124 0.969129 101.314 0.232898 0.880356 4.68593 0.0671021 0.0442069 0.955793 0.0193221 0.00469013 0.0185752 0.00446594 0.0056779 0.00642477 0.227116 0.256991 58.0614 -87.8999 126.115 15.9277 145.04 0.000142714 0.267353 192.695 0.310108 0.0673146 0.00409908 0.000562511 0.00138552 0.986954 0.991713 -2.99309e-06 -85.6552 0.0931025 31164.6 312.686 0.983494 0.319146 0.740331 0.740326 9.99958 2.98744e-06 1.19496e-05 0.135203 0.983448 0.931165 -0.0132913 4.93638e-06 0.520026 -2.04491e-20 7.59477e-24 -2.04415e-20 0.00139668 0.997814 8.60387e-05 0.152762 2.85297 0.00139668 0.997815 0.803582 0.0010706 0.00188168 0.000860387 0.455342 0.00188168 0.445436 0.0001317 1.02 0.888978 0.534317 0.287851 1.71998e-07 3.08866e-09 2367.68 3148.05 -0.0590948 0.482222 0.277221 0.255357 -0.592956 -0.169586 0.484789 -0.265388 -0.21941 2.852 1 0 294.539 0 2.26091 2.85 0.000298869 0.872699 0.708473 0.308402 0.438443 2.26108 140.567 83.5375 18.6987 60.6817 0.00404113 0 -40 10
1.951 5.64196e-08 2.54027e-06 0.153204 0.153204 0.0120237 2.56453e-05 0.00115467 0.191505 0.000658904 0.192159 0.969221 101.313 0.232887 0.880491 4.68664 0.0671131 0.0442136 0.955786 0.0193215 0.00469062 0.0185746 0.00446637 0.00567851 0.00642539 0.22714 0.257016 58.0615 -87.8999 126.115 15.9277 145.04 0.000142717 0.267353 192.694 0.310107 0.0673146 0.00409909 0.000562512 0.00138552 0.986954 0.991713 -2.99311e-06 -85.6552 0.0931026 31164.5 312.7 0.983493 0.319146 0.740343 0.740338 9.99958 2.98744e-06 1.19497e-05 0.135208 0.983448 0.931164 -0.0132913 4.93641e-06 0.520048 -2.04508e-20 7.59545e-24 -2.04432e-20 0.00139668 0.997814 8.60388e-05 0.152762 2.85297 0.00139668 0.997815 0.80365 0.00107061 0.00188169 0.000860388 0.455342 0.00188169 0.445441 0.000131703 1.02 0.88898 0.534317 0.287852 1.71998e-07 3.08869e-09 2367.67 3148.1 -0.0590999 0.482222 0.27722 0.25536 -0.592956 -0.169586 0.484773 -0.265386 -0.219396 2.853 1 0 294.535 0 2.26104 2.851 0.000298868 0.872729 0.708516 0.308366 0.438465 2.26122 140.574 83.5369 18.6986 60.6814 0.00404116 0 -40 10
1.952 5.64485e-08 2.54027e-06 0.153232 0.153232 0.0120237 2.56584e-05 0.00115467 0.19154 0.000658904 0.192195 0.969314 101.313 0.232876 0.880626 4.68736 0.0671241 0.0442203 0.95578 0.0193209 0.00469111 0.018574 0.00446679 0.00567911 0.00642602 0.227164 0.257041 58.0616 -87.8999 126.115 15.9276 145.04 0.000142719 0.267353 192.694 0.310107 0.0673145 0.00409909 0.000562512 0.00138553 0.986954 0.991713 -2.99312e-06 -85.6552 0.0931027 31164.5 312.713 0.983493 0.319146 0.740355 0.740351 9.99958 2.98745e-06 1.19497e-05 0.135213 0.983448 0.931163 -0.0132913 4.93644e-06 0.520069 -2.04525e-20 7.59613e-24 -2.04449e-20 0.00139668 0.997814 8.60388e-05 0.152763 2.85297 0.00139668 0.997815 0.803718 0.00107063 0.00188169 0.000860388 0.455342 0.00188169 0.445446 0.000131705 1.02 0.888981 0.534316 0.287854 1.71998e-07 3.08871e-09 2367.65 3148.15 -0.0591051 0.482222 0.27722 0.255363 -0.592955 -0.169586 0.484757 -0.265384 -0.219382 2.854 1 0 294.53 0 2.26118 2.852 0.000298867 0.872759 0.708558 0.308331 0.438487 2.26135 140.581 83.5363 18.6986 60.6811 0.00404118 0 -40 10
1.953 5.64773e-08 2.54027e-06 0.15326 0.15326 0.0120237 2.56715e-05 0.00115467 0.191575 0.000658905 0.19223 0.969406 101.312 0.232865 0.88076 4.68807 0.067135 0.0442271 0.955773 0.0193203 0.0046916 0.0185734 0.00446722 0.00567972 0.00642664 0.227189 0.257066 58.0616 -87.8999 126.114 15.9276 145.04 0.000142721 0.267353 192.694 0.310106 0.0673145 0.00409909 0.000562513 0.00138553 0.986954 0.991713 -2.99314e-06 -85.6552 0.0931028 31164.5 312.726 0.983493 0.319146 0.740367 0.740363 9.99958 2.98745e-06 1.19497e-05 0.135218 0.983448 0.931162 -0.0132913 4.93647e-06 0.520091 -2.04542e-20 7.59682e-24 -2.04466e-20 0.00139669 0.997814 8.60389e-05 0.152763 2.85297 0.00139669 0.997815 0.803786 0.00107065 0.00188169 0.000860389 0.455342 0.00188169 0.44545 0.000131707 1.02 0.888982 0.534316 0.287855 1.71999e-07 3.08873e-09 2367.64 3148.2 -0.0591102 0.482223 0.27722 0.255367 -0.592955 -0.169586 0.48474 -0.265382 -0.219368 2.855 1 0 294.525 0 2.26131 2.853 0.000298865 0.87279 0.7086 0.308295 0.438508 2.26149 140.588 83.5357 18.6986 60.6808 0.00404121 0 -40 10
1.954 5.65061e-08 2.54028e-06 0.153289 0.153288 0.0120236 2.56846e-05 0.00115467 0.191611 0.000658905 0.192265 0.969499 101.311 0.232854 0.880895 4.68878 0.067146 0.0442338 0.955766 0.0193197 0.00469209 0.0185727 0.00446765 0.00568032 0.00642727 0.227213 0.257091 58.0617 -87.8999 126.114 15.9276 145.04 0.000142724 0.267354 192.694 0.310106 0.0673144 0.0040991 0.000562514 0.00138553 0.986954 0.991713 -2.99315e-06 -85.6551 0.0931029 31164.5 312.74 0.983493 0.319146 0.74038 0.740375 9.99958 2.98746e-06 1.19497e-05 0.135223 0.983448 0.931161 -0.0132913 4.9365e-06 0.520112 -2.04559e-20 7.5975e-24 -2.04483e-20 0.00139669 0.997814 8.6039e-05 0.152763 2.85297 0.00139669 0.997815 0.803854 0.00107066 0.00188169 0.00086039 0.455341 0.00188169 0.445455 0.00013171 1.02 0.888983 0.534316 0.287857 1.71999e-07 3.08875e-09 2367.62 3148.25 -0.0591153 0.482223 0.27722 0.25537 -0.592954 -0.169586 0.484724 -0.26538 -0.219353 2.856 1 0 294.521 0 2.26145 2.854 0.000298864 0.87282 0.708643 0.30826 0.43853 2.26163 140.596 83.5351 18.6985 60.6805 0.00404123 0 -40 10
1.955 5.65349e-08 2.54028e-06 0.153317 0.153316 0.0120236 2.56977e-05 0.00115467 0.191646 0.000658906 0.1923 0.969592 101.311 0.232843 0.88103 4.6895 0.067157 0.0442405 0.955759 0.0193191 0.00469259 0.0185721 0.00446807 0.00568093 0.0064279 0.227237 0.257116 58.0618 -87.8999 126.114 15.9275 145.04 0.000142726 0.267354 192.694 0.310105 0.0673143 0.0040991 0.000562514 0.00138553 0.986954 0.991713 -2.99317e-06 -85.6551 0.093103 31164.5 312.753 0.983493 0.319146 0.740392 0.740387 9.99958 2.98746e-06 1.19497e-05 0.135228 0.983448 0.93116 -0.0132913 4.93653e-06 0.520133 -2.04577e-20 7.59818e-24 -2.04501e-20 0.00139669 0.997814 8.60391e-05 0.152763 2.85297 0.00139669 0.997815 0.803922 0.00107068 0.00188169 0.000860391 0.455341 0.00188169 0.44546 0.000131712 1.02 0.888984 0.534315 0.287858 1.71999e-07 3.08878e-09 2367.6 3148.3 -0.0591204 0.482223 0.277219 0.255373 -0.592953 -0.169586 0.484708 -0.265378 -0.219339 2.857 1 0 294.516 0 2.26158 2.855 0.000298863 0.87285 0.708685 0.308224 0.438552 2.26176 140.603 83.5345 18.6985 60.6802 0.00404126 0 -40 10
1.956 5.65638e-08 2.54028e-06 0.153345 0.153344 0.0120236 2.57108e-05 0.00115467 0.191681 0.000658906 0.192335 0.969684 101.31 0.232832 0.881165 4.69021 0.0671679 0.0442473 0.955753 0.0193185 0.00469308 0.0185715 0.0044685 0.00568153 0.00642852 0.227261 0.257141 58.0618 -87.8999 126.114 15.9275 145.04 0.000142728 0.267354 192.694 0.310105 0.0673143 0.0040991 0.000562515 0.00138553 0.986954 0.991713 -2.99318e-06 -85.6551 0.0931031 31164.4 312.766 0.983493 0.319146 0.740404 0.7404 9.99958 2.98747e-06 1.19498e-05 0.135233 0.983449 0.931159 -0.0132913 4.93656e-06 0.520155 -2.04594e-20 7.59886e-24 -2.04518e-20 0.00139669 0.997814 8.60392e-05 0.152763 2.85297 0.00139669 0.997815 0.80399 0.00107069 0.00188169 0.000860392 0.455341 0.00188169 0.445464 0.000131714 1.02 0.888985 0.534315 0.28786 1.72e-07 3.0888e-09 2367.59 3148.35 -0.0591256 0.482223 0.277219 0.255377 -0.592953 -0.169586 0.484691 -0.265376 -0.219325 2.858 1 0 294.512 0 2.26172 2.856 0.000298861 0.87288 0.708727 0.308188 0.438574 2.2619 140.61 83.5339 18.6985 60.6799 0.00404128 0 -40 10
1.957 5.65926e-08 2.54028e-06 0.153373 0.153372 0.0120236 2.57239e-05 0.00115467 0.191716 0.000658906 0.19237 0.969777 101.309 0.232821 0.8813 4.69093 0.0671789 0.044254 0.955746 0.0193179 0.00469357 0.0185708 0.00446893 0.00568214 0.00642915 0.227285 0.257166 58.0619 -87.8999 126.113 15.9275 145.04 0.000142731 0.267354 192.693 0.310105 0.0673142 0.00409911 0.000562516 0.00138554 0.986954 0.991713 -2.9932e-06 -85.6551 0.0931032 31164.4 312.78 0.983493 0.319146 0.740416 0.740412 9.99958 2.98747e-06 1.19498e-05 0.135238 0.983449 0.931158 -0.0132913 4.93659e-06 0.520176 -2.04611e-20 7.59954e-24 -2.04535e-20 0.00139669 0.997814 8.60393e-05 0.152763 2.85298 0.00139669 0.997815 0.804058 0.00107071 0.0018817 0.000860393 0.455341 0.00188169 0.445469 0.000131716 1.02 0.888986 0.534315 0.287861 1.72e-07 3.08882e-09 2367.57 3148.41 -0.0591307 0.482223 0.277219 0.25538 -0.592952 -0.169586 0.484675 -0.265374 -0.219311 2.859 1 0 294.507 0 2.26185 2.857 0.00029886 0.87291 0.70877 0.308153 0.438595 2.26203 140.617 83.5333 18.6984 60.6796 0.00404131 0 -40 10
1.958 5.66214e-08 2.54028e-06 0.153401 0.1534 0.0120236 2.5737e-05 0.00115467 0.191751 0.000658907 0.192405 0.96987 101.308 0.23281 0.881435 4.69164 0.0671899 0.0442608 0.955739 0.0193173 0.00469406 0.0185702 0.00446935 0.00568274 0.00642978 0.22731 0.257191 58.0619 -87.8999 126.113 15.9274 145.04 0.000142733 0.267354 192.693 0.310104 0.0673142 0.00409911 0.000562516 0.00138554 0.986954 0.991713 -2.99321e-06 -85.6551 0.0931032 31164.4 312.793 0.983493 0.319146 0.740429 0.740424 9.99958 2.98748e-06 1.19498e-05 0.135243 0.983449 0.931157 -0.0132913 4.93662e-06 0.520198 -2.04628e-20 7.60023e-24 -2.04552e-20 0.00139669 0.997814 8.60393e-05 0.152763 2.85298 0.00139669 0.997815 0.804126 0.00107072 0.0018817 0.000860393 0.45534 0.0018817 0.445474 0.000131719 1.02 0.888987 0.534314 0.287863 1.72e-07 3.08885e-09 2367.55 3148.46 -0.0591358 0.482223 0.277218 0.255383 -0.592951 -0.169586 0.484659 -0.265372 -0.219297 2.86 1 0 294.502 0 2.26199 2.858 0.000298858 0.87294 0.708812 0.308117 0.438617 2.26217 140.625 83.5327 18.6984 60.6794 0.00404133 0 -40 10
1.959 5.66502e-08 2.54029e-06 0.153429 0.153428 0.0120236 2.57501e-05 0.00115468 0.191786 0.000658907 0.19244 0.969962 101.308 0.232799 0.88157 4.69236 0.0672008 0.0442675 0.955732 0.0193167 0.00469455 0.0185696 0.00446978 0.00568335 0.00643041 0.227334 0.257216 58.062 -87.8999 126.113 15.9274 145.04 0.000142736 0.267355 192.693 0.310104 0.0673141 0.00409911 0.000562517 0.00138554 0.986954 0.991713 -2.99323e-06 -85.6551 0.0931033 31164.4 312.807 0.983493 0.319146 0.740441 0.740436 9.99958 2.98748e-06 1.19498e-05 0.135248 0.983449 0.931156 -0.0132913 4.93664e-06 0.520219 -2.04645e-20 7.60091e-24 -2.04569e-20 0.00139669 0.997814 8.60394e-05 0.152764 2.85298 0.00139669 0.997815 0.804193 0.00107074 0.0018817 0.000860394 0.45534 0.0018817 0.445478 0.000131721 1.02 0.888988 0.534314 0.287864 1.72e-07 3.08887e-09 2367.54 3148.51 -0.059141 0.482223 0.277218 0.255386 -0.592951 -0.169586 0.484643 -0.26537 -0.219282 2.861 1 0 294.498 0 2.26213 2.859 0.000298857 0.87297 0.708854 0.308082 0.438639 2.2623 140.632 83.5321 18.6984 60.6791 0.00404136 0 -40 10
1.96 5.66791e-08 2.54029e-06 0.153457 0.153456 0.0120236 2.57632e-05 0.00115468 0.191821 0.000658908 0.192475 0.970055 101.307 0.232788 0.881705 4.69308 0.0672118 0.0442743 0.955726 0.019316 0.00469504 0.018569 0.00447021 0.00568396 0.00643103 0.227358 0.257241 58.0621 -87.8999 126.113 15.9273 145.04 0.000142738 0.267355 192.693 0.310103 0.0673141 0.00409911 0.000562518 0.00138554 0.986954 0.991713 -2.99324e-06 -85.6551 0.0931034 31164.3 312.82 0.983493 0.319146 0.740453 0.740449 9.99958 2.98749e-06 1.19498e-05 0.135253 0.983449 0.931155 -0.0132913 4.93667e-06 0.520241 -2.04662e-20 7.60159e-24 -2.04586e-20 0.00139669 0.997814 8.60395e-05 0.152764 2.85298 0.00139669 0.997815 0.804261 0.00107076 0.0018817 0.000860395 0.45534 0.0018817 0.445483 0.000131723 1.02 0.888989 0.534314 0.287866 1.72001e-07 3.08889e-09 2367.52 3148.56 -0.0591461 0.482223 0.277218 0.25539 -0.59295 -0.169586 0.484626 -0.265367 -0.219268 2.862 1 0 294.493 0 2.26226 2.86 0.000298856 0.873001 0.708897 0.308047 0.438661 2.26244 140.639 83.5315 18.6983 60.6788 0.00404138 0 -40 10
1.961 5.67079e-08 2.54029e-06 0.153485 0.153484 0.0120235 2.57763e-05 0.00115468 0.191856 0.000658908 0.19251 0.970148 101.306 0.232777 0.881839 4.69379 0.0672228 0.0442811 0.955719 0.0193154 0.00469553 0.0185683 0.00447063 0.00568456 0.00643166 0.227382 0.257266 58.0621 -87.8999 126.113 15.9273 145.04 0.00014274 0.267355 192.693 0.310103 0.067314 0.00409912 0.000562518 0.00138555 0.986954 0.991713 -2.99326e-06 -85.6551 0.0931035 31164.3 312.833 0.983493 0.319146 0.740465 0.740461 9.99958 2.98749e-06 1.19499e-05 0.135258 0.983449 0.931154 -0.0132913 4.9367e-06 0.520262 -2.04679e-20 7.60228e-24 -2.04603e-20 0.0013967 0.997814 8.60396e-05 0.152764 2.85298 0.0013967 0.997815 0.804329 0.00107077 0.0018817 0.000860396 0.45534 0.0018817 0.445488 0.000131725 1.02 0.88899 0.534314 0.287867 1.72001e-07 3.08891e-09 2367.51 3148.61 -0.0591512 0.482223 0.277218 0.255393 -0.592949 -0.169586 0.48461 -0.265365 -0.219254 2.863 1 0 294.488 0 2.2624 2.861 0.000298854 0.873031 0.708939 0.308011 0.438682 2.26257 140.647 83.5309 18.6983 60.6785 0.00404141 0 -40 10
1.962 5.67367e-08 2.54029e-06 0.153513 0.153512 0.0120235 2.57894e-05 0.00115468 0.191891 0.000658909 0.192545 0.970241 101.305 0.232766 0.881974 4.69451 0.0672338 0.0442878 0.955712 0.0193148 0.00469602 0.0185677 0.00447106 0.00568517 0.00643229 0.227407 0.257292 58.0622 -87.8999 126.112 15.9273 145.04 0.000142743 0.267355 192.693 0.310102 0.067314 0.00409912 0.000562519 0.00138555 0.986954 0.991713 -2.99327e-06 -85.6551 0.0931036 31164.3 312.847 0.983493 0.319146 0.740478 0.740473 9.99958 2.9875e-06 1.19499e-05 0.135263 0.983449 0.931153 -0.0132913 4.93673e-06 0.520284 -2.04697e-20 7.60296e-24 -2.04621e-20 0.0013967 0.997814 8.60397e-05 0.152764 2.85298 0.0013967 0.997815 0.804397 0.00107079 0.0018817 0.000860397 0.45534 0.0018817 0.445493 0.000131728 1.02 0.888992 0.534313 0.287869 1.72001e-07 3.08894e-09 2367.49 3148.66 -0.0591564 0.482223 0.277217 0.255396 -0.592949 -0.169586 0.484594 -0.265363 -0.21924 2.864 1 0 294.484 0 2.26253 2.862 0.000298853 0.873061 0.708981 0.307976 0.438704 2.26271 140.654 83.5303 18.6983 60.6782 0.00404143 0 -40 10
1.963 5.67655e-08 2.54029e-06 0.153541 0.15354 0.0120235 2.58025e-05 0.00115468 0.191926 0.000658909 0.19258 0.970333 101.305 0.232755 0.882109 4.69523 0.0672447 0.0442946 0.955705 0.0193142 0.00469652 0.0185671 0.00447149 0.00568578 0.00643292 0.227431 0.257317 58.0623 -87.8999 126.112 15.9272 145.04 0.000142745 0.267355 192.692 0.310102 0.0673139 0.00409912 0.00056252 0.00138555 0.986954 0.991713 -2.99329e-06 -85.6551 0.0931037 31164.3 312.86 0.983493 0.319146 0.74049 0.740486 9.99958 2.9875e-06 1.19499e-05 0.135268 0.98345 0.931151 -0.0132913 4.93676e-06 0.520305 -2.04714e-20 7.60365e-24 -2.04638e-20 0.0013967 0.997814 8.60397e-05 0.152764 2.85298 0.0013967 0.997815 0.804465 0.0010708 0.0018817 0.000860397 0.455339 0.0018817 0.445497 0.00013173 1.02 0.888993 0.534313 0.28787 1.72001e-07 3.08896e-09 2367.47 3148.71 -0.0591615 0.482223 0.277217 0.2554 -0.592948 -0.169586 0.484577 -0.265361 -0.219226 2.865 1 0 294.479 0 2.26267 2.863 0.000298851 0.873091 0.709024 0.30794 0.438726 2.26284 140.661 83.5297 18.6982 60.6779 0.00404146 0 -40 10
1.964 5.67944e-08 2.54029e-06 0.153569 0.153568 0.0120235 2.58156e-05 0.00115468 0.191961 0.000658909 0.192615 0.970426 101.304 0.232744 0.882244 4.69595 0.0672557 0.0443014 0.955699 0.0193136 0.00469701 0.0185665 0.00447192 0.00568638 0.00643355 0.227455 0.257342 58.0623 -87.8999 126.112 15.9272 145.04 0.000142747 0.267356 192.692 0.310102 0.0673139 0.00409913 0.00056252 0.00138555 0.986954 0.991713 -2.9933e-06 -85.6551 0.0931038 31164.3 312.873 0.983493 0.319146 0.740502 0.740498 9.99958 2.98751e-06 1.19499e-05 0.135273 0.98345 0.93115 -0.0132913 4.93679e-06 0.520327 -2.04731e-20 7.60433e-24 -2.04655e-20 0.0013967 0.997814 8.60398e-05 0.152764 2.85298 0.0013967 0.997815 0.804533 0.00107082 0.00188171 0.000860398 0.455339 0.0018817 0.445502 0.000131732 1.02 0.888994 0.534313 0.287872 1.72002e-07 3.08898e-09 2367.46 3148.77 -0.0591666 0.482223 0.277217 0.255403 -0.592947 -0.169586 0.484561 -0.265359 -0.219211 2.866 1 0 294.475 0 2.2628 2.864 0.00029885 0.873121 0.709066 0.307905 0.438747 2.26298 140.668 83.5291 18.6982 60.6776 0.00404148 0 -40 10
1.965 5.68232e-08 2.5403e-06 0.153596 0.153596 0.0120235 2.58287e-05 0.00115468 0.191996 0.00065891 0.19265 0.970519 101.303 0.232733 0.882379 4.69667 0.0672667 0.0443082 0.955692 0.019313 0.0046975 0.0185658 0.00447235 0.00568699 0.00643418 0.22748 0.257367 58.0624 -87.8999 126.112 15.9272 145.04 0.00014275 0.267356 192.692 0.310101 0.0673138 0.00409913 0.000562521 0.00138555 0.986954 0.991713 -2.99332e-06 -85.655 0.0931038 31164.2 312.887 0.983493 0.319146 0.740515 0.74051 9.99958 2.98751e-06 1.19499e-05 0.135278 0.98345 0.931149 -0.0132913 4.93682e-06 0.520348 -2.04748e-20 7.60502e-24 -2.04672e-20 0.0013967 0.997814 8.60399e-05 0.152765 2.85298 0.0013967 0.997815 0.8046 0.00107083 0.00188171 0.000860399 0.455339 0.00188171 0.445507 0.000131734 1.02 0.888995 0.534312 0.287873 1.72002e-07 3.08901e-09 2367.44 3148.82 -0.0591717 0.482223 0.277217 0.255406 -0.592947 -0.169587 0.484545 -0.265357 -0.219197 2.867 1 0 294.47 0 2.26294 2.865 0.000298849 0.873151 0.709108 0.30787 0.438769 2.26311 140.676 83.5285 18.6981 60.6773 0.00404151 0 -40 10
1.966 5.6852e-08 2.5403e-06 0.153624 0.153624 0.0120235 2.58418e-05 0.00115468 0.19203 0.00065891 0.192685 0.970612 101.303 0.232722 0.882514 4.69739 0.0672777 0.044315 0.955685 0.0193124 0.00469799 0.0185652 0.00447277 0.0056876 0.00643481 0.227504 0.257392 58.0624 -87.8999 126.111 15.9271 145.04 0.000142752 0.267356 192.692 0.310101 0.0673138 0.00409913 0.000562522 0.00138556 0.986954 0.991713 -2.99333e-06 -85.655 0.0931039 31164.2 312.9 0.983493 0.319146 0.740527 0.740522 9.99958 2.98752e-06 1.195e-05 0.135283 0.98345 0.931148 -0.0132913 4.93685e-06 0.52037 -2.04765e-20 7.6057e-24 -2.04689e-20 0.0013967 0.997814 8.604e-05 0.152765 2.85298 0.0013967 0.997815 0.804668 0.00107085 0.00188171 0.0008604 0.455339 0.00188171 0.445511 0.000131737 1.02 0.888996 0.534312 0.287875 1.72002e-07 3.08903e-09 2367.42 3148.87 -0.0591769 0.482224 0.277216 0.255409 -0.592946 -0.169587 0.484529 -0.265355 -0.219183 2.868 1 0 294.465 0 2.26307 2.866 0.000298847 0.873182 0.709151 0.307834 0.438791 2.26325 140.683 83.5279 18.6981 60.677 0.00404153 0 -40 10
1.967 5.68808e-08 2.5403e-06 0.153652 0.153652 0.0120235 2.58549e-05 0.00115468 0.192065 0.000658911 0.192719 0.970704 101.302 0.232711 0.882649 4.69811 0.0672887 0.0443218 0.955678 0.0193118 0.00469849 0.0185646 0.0044732 0.00568821 0.00643543 0.227528 0.257417 58.0625 -87.8999 126.111 15.9271 145.04 0.000142755 0.267356 192.692 0.3101 0.0673137 0.00409914 0.000562523 0.00138556 0.986954 0.991713 -2.99335e-06 -85.655 0.093104 31164.2 312.914 0.983493 0.319146 0.740539 0.740535 9.99958 2.98752e-06 1.195e-05 0.135288 0.98345 0.931147 -0.0132913 4.93688e-06 0.520392 -2.04783e-20 7.60639e-24 -2.04706e-20 0.0013967 0.997814 8.60401e-05 0.152765 2.85298 0.0013967 0.997815 0.804736 0.00107086 0.00188171 0.000860401 0.455338 0.00188171 0.445516 0.000131739 1.02 0.888997 0.534312 0.287877 1.72003e-07 3.08905e-09 2367.41 3148.92 -0.059182 0.482224 0.277216 0.255413 -0.592946 -0.169587 0.484512 -0.265353 -0.219169 2.869 1 0 294.461 0 2.26321 2.867 0.000298846 0.873212 0.709193 0.307799 0.438813 2.26338 140.69 83.5273 18.6981 60.6767 0.00404156 0 -40 10
1.968 5.69096e-08 2.5403e-06 0.15368 0.15368 0.0120234 2.5868e-05 0.00115468 0.1921 0.000658911 0.192754 0.970797 101.301 0.2327 0.882784 4.69883 0.0672996 0.0443285 0.955671 0.0193112 0.00469898 0.0185639 0.00447363 0.00568881 0.00643606 0.227553 0.257443 58.0626 -87.8999 126.111 15.9271 145.04 0.000142757 0.267356 192.692 0.3101 0.0673137 0.00409914 0.000562523 0.00138556 0.986954 0.991713 -2.99336e-06 -85.655 0.0931041 31164.2 312.927 0.983493 0.319146 0.740551 0.740547 9.99958 2.98753e-06 1.195e-05 0.135293 0.98345 0.931146 -0.0132913 4.93691e-06 0.520413 -2.048e-20 7.60707e-24 -2.04724e-20 0.0013967 0.997814 8.60401e-05 0.152765 2.85299 0.0013967 0.997815 0.804803 0.00107088 0.00188171 0.000860401 0.455338 0.00188171 0.445521 0.000131741 1.02 0.888998 0.534311 0.287878 1.72003e-07 3.08907e-09 2367.39 3148.97 -0.0591871 0.482224 0.277216 0.255416 -0.592945 -0.169587 0.484496 -0.265351 -0.219155 2.87 1 0 294.456 0 2.26334 2.868 0.000298844 0.873242 0.709235 0.307764 0.438834 2.26352 140.697 83.5267 18.698 60.6764 0.00404158 0 -40 10
1.969 5.69385e-08 2.5403e-06 0.153708 0.153707 0.0120234 2.58811e-05 0.00115468 0.192135 0.000658911 0.192789 0.97089 101.3 0.232689 0.882919 4.69955 0.0673106 0.0443353 0.955665 0.0193106 0.00469947 0.0185633 0.00447406 0.00568942 0.00643669 0.227577 0.257468 58.0626 -87.8999 126.111 15.927 145.04 0.000142759 0.267357 192.691 0.3101 0.0673136 0.00409914 0.000562524 0.00138556 0.986954 0.991713 -2.99338e-06 -85.655 0.0931042 31164.1 312.94 0.983493 0.319146 0.740564 0.740559 9.99958 2.98753e-06 1.195e-05 0.135298 0.98345 0.931145 -0.0132913 4.93694e-06 0.520435 -2.04817e-20 7.60776e-24 -2.04741e-20 0.0013967 0.997814 8.60402e-05 0.152765 2.85299 0.0013967 0.997815 0.804871 0.0010709 0.00188171 0.000860402 0.455338 0.00188171 0.445525 0.000131743 1.02 0.888999 0.534311 0.28788 1.72003e-07 3.0891e-09 2367.38 3149.02 -0.0591923 0.482224 0.277215 0.255419 -0.592944 -0.169587 0.48448 -0.265349 -0.21914 2.871 1 0 294.451 0 2.26348 2.869 0.000298843 0.873272 0.709278 0.307728 0.438856 2.26365 140.705 83.5261 18.698 60.6762 0.00404161 0 -40 10
1.97 5.69673e-08 2.54031e-06 0.153736 0.153735 0.0120234 2.58942e-05 0.00115468 0.192169 0.000658912 0.192824 0.970983 101.3 0.232678 0.883054 4.70027 0.0673216 0.0443422 0.955658 0.01931 0.00469996 0.0185627 0.00447449 0.00569003 0.00643732 0.227601 0.257493 58.0627 -87.9 126.111 15.927 145.04 0.000142762 0.267357 192.691 0.310099 0.0673136 0.00409914 0.000562525 0.00138557 0.986954 0.991713 -2.99339e-06 -85.655 0.0931043 31164.1 312.954 0.983493 0.319146 0.740576 0.740571 9.99958 2.98754e-06 1.195e-05 0.135303 0.98345 0.931144 -0.0132913 4.93697e-06 0.520456 -2.04834e-20 7.60844e-24 -2.04758e-20 0.00139671 0.997814 8.60403e-05 0.152765 2.85299 0.00139671 0.997815 0.804939 0.00107091 0.00188171 0.000860403 0.455338 0.00188171 0.44553 0.000131746 1.02 0.889 0.534311 0.287881 1.72003e-07 3.08912e-09 2367.36 3149.07 -0.0591974 0.482224 0.277215 0.255423 -0.592944 -0.169587 0.484463 -0.265347 -0.219126 2.872 1 0 294.447 0 2.26361 2.87 0.000298842 0.873302 0.70932 0.307693 0.438878 2.26379 140.712 83.5255 18.698 60.6759 0.00404163 0 -40 10
1.971 5.69961e-08 2.54031e-06 0.153763 0.153763 0.0120234 2.59073e-05 0.00115469 0.192204 0.000658912 0.192858 0.971076 101.299 0.232667 0.883189 4.70099 0.0673326 0.044349 0.955651 0.0193094 0.00470046 0.018562 0.00447492 0.00569064 0.00643796 0.227626 0.257518 58.0627 -87.9 126.11 15.9269 145.04 0.000142764 0.267357 192.691 0.310099 0.0673135 0.00409915 0.000562525 0.00138557 0.986954 0.991713 -2.99341e-06 -85.655 0.0931044 31164.1 312.967 0.983493 0.319146 0.740588 0.740584 9.99958 2.98754e-06 1.19501e-05 0.135308 0.983451 0.931143 -0.0132913 4.937e-06 0.520478 -2.04851e-20 7.60913e-24 -2.04775e-20 0.00139671 0.997814 8.60404e-05 0.152765 2.85299 0.00139671 0.997815 0.805006 0.00107093 0.00188172 0.000860404 0.455337 0.00188171 0.445535 0.000131748 1.02 0.889001 0.53431 0.287883 1.72004e-07 3.08914e-09 2367.34 3149.13 -0.0592025 0.482224 0.277215 0.255426 -0.592943 -0.169587 0.484447 -0.265344 -0.219112 2.873 1 0 294.442 0 2.26375 2.871 0.00029884 0.873333 0.709362 0.307658 0.438899 2.26392 140.719 83.5249 18.6979 60.6756 0.00404166 0 -40 10
1.972 5.70249e-08 2.54031e-06 0.153791 0.153791 0.0120234 2.59204e-05 0.00115469 0.192239 0.000658913 0.192893 0.971169 101.298 0.232656 0.883324 4.70171 0.0673436 0.0443558 0.955644 0.0193088 0.00470095 0.0185614 0.00447535 0.00569125 0.00643859 0.22765 0.257543 58.0628 -87.9 126.11 15.9269 145.04 0.000142766 0.267357 192.691 0.310098 0.0673135 0.00409915 0.000562526 0.00138557 0.986954 0.991713 -2.99342e-06 -85.655 0.0931045 31164.1 312.981 0.983493 0.319146 0.7406 0.740596 9.99958 2.98755e-06 1.19501e-05 0.135313 0.983451 0.931142 -0.0132913 4.93703e-06 0.5205 -2.04869e-20 7.60982e-24 -2.04793e-20 0.00139671 0.997814 8.60405e-05 0.152766 2.85299 0.00139671 0.997815 0.805074 0.00107094 0.00188172 0.000860405 0.455337 0.00188172 0.445539 0.00013175 1.02 0.889003 0.53431 0.287884 1.72004e-07 3.08917e-09 2367.33 3149.18 -0.0592077 0.482224 0.277215 0.255429 -0.592942 -0.169587 0.484431 -0.265342 -0.219098 2.874 1 0 294.438 0 2.26388 2.872 0.000298839 0.873363 0.709404 0.307623 0.438921 2.26406 140.726 83.5243 18.6979 60.6753 0.00404168 0 -40 10
1.973 5.70538e-08 2.54031e-06 0.153819 0.153818 0.0120234 2.59335e-05 0.00115469 0.192273 0.000658913 0.192928 0.971261 101.298 0.232645 0.883459 4.70243 0.0673546 0.0443626 0.955637 0.0193081 0.00470145 0.0185608 0.00447578 0.00569186 0.00643922 0.227674 0.257569 58.0629 -87.9 126.11 15.9269 145.04 0.000142769 0.267357 192.691 0.310098 0.0673134 0.00409915 0.000562527 0.00138557 0.986954 0.991713 -2.99344e-06 -85.655 0.0931045 31164.1 312.994 0.983493 0.319146 0.740613 0.740608 9.99958 2.98755e-06 1.19501e-05 0.135318 0.983451 0.931141 -0.0132913 4.93706e-06 0.520521 -2.04886e-20 7.6105e-24 -2.0481e-20 0.00139671 0.997814 8.60405e-05 0.152766 2.85299 0.00139671 0.997815 0.805141 0.00107096 0.00188172 0.000860405 0.455337 0.00188172 0.445544 0.000131752 1.02 0.889004 0.53431 0.287886 1.72004e-07 3.08919e-09 2367.31 3149.23 -0.0592128 0.482224 0.277214 0.255432 -0.592942 -0.169587 0.484414 -0.26534 -0.219084 2.875 1 0 294.433 0 2.26402 2.873 0.000298837 0.873393 0.709447 0.307588 0.438943 2.26419 140.734 83.5237 18.6979 60.675 0.00404171 0 -40 10
1.974 5.70826e-08 2.54031e-06 0.153846 0.153846 0.0120234 2.59466e-05 0.00115469 0.192308 0.000658913 0.192962 0.971354 101.297 0.232634 0.883594 4.70316 0.0673655 0.0443694 0.955631 0.0193075 0.00470194 0.0185602 0.0044762 0.00569246 0.00643985 0.227699 0.257594 58.0629 -87.9 126.11 15.9268 145.04 0.000142771 0.267357 192.691 0.310097 0.0673133 0.00409916 0.000562527 0.00138557 0.986954 0.991713 -2.99345e-06 -85.655 0.0931046 31164 313.008 0.983493 0.319146 0.740625 0.740621 9.99958 2.98756e-06 1.19501e-05 0.135323 0.983451 0.93114 -0.0132913 4.93709e-06 0.520543 -2.04903e-20 7.61119e-24 -2.04827e-20 0.00139671 0.997814 8.60406e-05 0.152766 2.85299 0.00139671 0.997815 0.805209 0.00107097 0.00188172 0.000860406 0.455337 0.00188172 0.445549 0.000131755 1.02 0.889005 0.53431 0.287887 1.72004e-07 3.08921e-09 2367.29 3149.28 -0.0592179 0.482224 0.277214 0.255436 -0.592941 -0.169587 0.484398 -0.265338 -0.219069 2.876 1 0 294.428 0 2.26415 2.874 0.000298836 0.873423 0.709489 0.307552 0.438965 2.26433 140.741 83.5231 18.6978 60.6747 0.00404173 0 -40 10
1.975 5.71114e-08 2.54032e-06 0.153874 0.153874 0.0120234 2.59597e-05 0.00115469 0.192343 0.000658914 0.192997 0.971447 101.296 0.232623 0.883729 4.70388 0.0673765 0.0443762 0.955624 0.0193069 0.00470243 0.0185595 0.00447663 0.00569307 0.00644048 0.227723 0.257619 58.063 -87.9 126.109 15.9268 145.04 0.000142773 0.267358 192.69 0.310097 0.0673133 0.00409916 0.000562528 0.00138558 0.986954 0.991713 -2.99347e-06 -85.6549 0.0931047 31164 313.021 0.983493 0.319146 0.740637 0.740633 9.99958 2.98756e-06 1.19501e-05 0.135328 0.983451 0.931139 -0.0132913 4.93712e-06 0.520564 -2.0492e-20 7.61188e-24 -2.04844e-20 0.00139671 0.997814 8.60407e-05 0.152766 2.85299 0.00139671 0.997815 0.805276 0.00107099 0.00188172 0.000860407 0.455337 0.00188172 0.445553 0.000131757 1.02 0.889006 0.534309 0.287889 1.72005e-07 3.08923e-09 2367.28 3149.33 -0.0592231 0.482224 0.277214 0.255439 -0.59294 -0.169587 0.484382 -0.265336 -0.219055 2.877 1 0 294.424 0 2.26429 2.875 0.000298835 0.873454 0.709531 0.307517 0.438986 2.26446 140.748 83.5225 18.6978 60.6744 0.00404176 0 -40 10
1.976 5.71402e-08 2.54032e-06 0.153902 0.153901 0.0120233 2.59728e-05 0.00115469 0.192377 0.000658914 0.193031 0.97154 101.295 0.232612 0.883864 4.7046 0.0673875 0.0443831 0.955617 0.0193063 0.00470293 0.0185589 0.00447706 0.00569368 0.00644111 0.227747 0.257644 58.0631 -87.9 126.109 15.9268 145.04 0.000142776 0.267358 192.69 0.310097 0.0673132 0.00409916 0.000562529 0.00138558 0.986954 0.991713 -2.99348e-06 -85.6549 0.0931048 31164 313.034 0.983493 0.319146 0.74065 0.740645 9.99958 2.98757e-06 1.19502e-05 0.135333 0.983451 0.931138 -0.0132913 4.93715e-06 0.520586 -2.04938e-20 7.61256e-24 -2.04861e-20 0.00139671 0.997814 8.60408e-05 0.152766 2.85299 0.00139671 0.997815 0.805344 0.001071 0.00188172 0.000860408 0.455336 0.00188172 0.445558 0.000131759 1.02 0.889007 0.534309 0.28789 1.72005e-07 3.08926e-09 2367.26 3149.38 -0.0592282 0.482224 0.277213 0.255442 -0.59294 -0.169587 0.484366 -0.265334 -0.219041 2.878 1 0 294.419 0 2.26442 2.876 0.000298833 0.873484 0.709574 0.307482 0.439008 2.2646 140.755 83.5219 18.6978 60.6741 0.00404178 0 -40 10
1.977 5.7169e-08 2.54032e-06 0.153929 0.153929 0.0120233 2.59859e-05 0.00115469 0.192412 0.000658915 0.193066 0.971633 101.295 0.232601 0.883999 4.70533 0.0673985 0.0443899 0.95561 0.0193057 0.00470342 0.0185583 0.00447749 0.00569429 0.00644174 0.227772 0.25767 58.0631 -87.9 126.109 15.9267 145.04 0.000142778 0.267358 192.69 0.310096 0.0673132 0.00409917 0.000562529 0.00138558 0.986954 0.991713 -2.9935e-06 -85.6549 0.0931049 31164 313.048 0.983493 0.319146 0.740662 0.740657 9.99958 2.98757e-06 1.19502e-05 0.135338 0.983451 0.931137 -0.0132913 4.93718e-06 0.520608 -2.04955e-20 7.61325e-24 -2.04879e-20 0.00139671 0.997814 8.60409e-05 0.152766 2.85299 0.00139671 0.997815 0.805411 0.00107102 0.00188173 0.000860409 0.455336 0.00188172 0.445563 0.000131761 1.02 0.889008 0.534309 0.287892 1.72005e-07 3.08928e-09 2367.25 3149.43 -0.0592333 0.482224 0.277213 0.255446 -0.592939 -0.169587 0.484349 -0.265332 -0.219027 2.879 1 0 294.414 0 2.26456 2.877 0.000298832 0.873514 0.709616 0.307447 0.43903 2.26473 140.763 83.5213 18.6977 60.6738 0.00404181 0 -40 10
1.978 5.71979e-08 2.54032e-06 0.153957 0.153956 0.0120233 2.5999e-05 0.00115469 0.192446 0.000658915 0.1931 0.971726 101.294 0.232591 0.884134 4.70605 0.0674095 0.0443967 0.955603 0.0193051 0.00470392 0.0185576 0.00447792 0.0056949 0.00644237 0.227796 0.257695 58.0632 -87.9 126.109 15.9267 145.04 0.000142781 0.267358 192.69 0.310096 0.0673131 0.00409917 0.00056253 0.00138558 0.986954 0.991713 -2.99351e-06 -85.6549 0.093105 31163.9 313.061 0.983493 0.319146 0.740674 0.74067 9.99958 2.98758e-06 1.19502e-05 0.135343 0.983452 0.931136 -0.0132913 4.93721e-06 0.520629 -2.04972e-20 7.61394e-24 -2.04896e-20 0.00139671 0.997814 8.60409e-05 0.152767 2.85299 0.00139671 0.997815 0.805479 0.00107104 0.00188173 0.000860409 0.455336 0.00188173 0.445567 0.000131764 1.02 0.889009 0.534308 0.287893 1.72005e-07 3.0893e-09 2367.23 3149.49 -0.0592385 0.482224 0.277213 0.255449 -0.592938 -0.169587 0.484333 -0.26533 -0.219012 2.88 1 0 294.41 0 2.26469 2.878 0.00029883 0.873544 0.709658 0.307412 0.439051 2.26487 140.77 83.5207 18.6977 60.6735 0.00404183 0 -40 10
1.979 5.72267e-08 2.54032e-06 0.153984 0.153984 0.0120233 2.60121e-05 0.00115469 0.192481 0.000658915 0.193135 0.971819 101.293 0.23258 0.884269 4.70678 0.0674205 0.0444036 0.955596 0.0193045 0.00470441 0.018557 0.00447835 0.00569551 0.00644301 0.227821 0.25772 58.0632 -87.9 126.109 15.9266 145.04 0.000142783 0.267358 192.69 0.310095 0.0673131 0.00409917 0.000562531 0.00138558 0.986953 0.991713 -2.99353e-06 -85.6549 0.0931051 31163.9 313.075 0.983493 0.319146 0.740686 0.740682 9.99958 2.98758e-06 1.19502e-05 0.135348 0.983452 0.931135 -0.0132913 4.93724e-06 0.520651 -2.04989e-20 7.61463e-24 -2.04913e-20 0.00139672 0.997814 8.6041e-05 0.152767 2.853 0.00139672 0.997815 0.805546 0.00107105 0.00188173 0.00086041 0.455336 0.00188173 0.445572 0.000131766 1.02 0.88901 0.534308 0.287895 1.72006e-07 3.08933e-09 2367.21 3149.54 -0.0592436 0.482225 0.277213 0.255452 -0.592938 -0.169587 0.484317 -0.265328 -0.218998 2.881 1 0 294.405 0 2.26483 2.879 0.000298829 0.873575 0.7097 0.307377 0.439073 2.265 140.777 83.5201 18.6977 60.6732 0.00404186 0 -40 10
1.98 5.72555e-08 2.54033e-06 0.154012 0.154012 0.0120233 2.60252e-05 0.00115469 0.192515 0.000658916 0.193169 0.971912 101.292 0.232569 0.884404 4.7075 0.0674315 0.0444104 0.95559 0.0193039 0.00470491 0.0185564 0.00447878 0.00569612 0.00644364 0.227845 0.257746 58.0633 -87.9 126.108 15.9266 145.04 0.000142785 0.267359 192.69 0.310095 0.067313 0.00409918 0.000562531 0.00138559 0.986953 0.991713 -2.99354e-06 -85.6549 0.0931052 31163.9 313.088 0.983493 0.319146 0.740699 0.740694 9.99958 2.98759e-06 1.19502e-05 0.135353 0.983452 0.931134 -0.0132913 4.93727e-06 0.520673 -2.05007e-20 7.61532e-24 -2.04931e-20 0.00139672 0.997814 8.60411e-05 0.152767 2.853 0.00139672 0.997815 0.805613 0.00107107 0.00188173 0.000860411 0.455335 0.00188173 0.445577 0.000131768 1.02 0.889011 0.534308 0.287896 1.72006e-07 3.08935e-09 2367.2 3149.59 -0.0592487 0.482225 0.277212 0.255456 -0.592937 -0.169587 0.4843 -0.265326 -0.218984 2.882 1 0 294.401 0 2.26496 2.88 0.000298828 0.873605 0.709743 0.307342 0.439095 2.26514 140.784 83.5195 18.6976 60.673 0.00404188 0 -40 10
1.981 5.72843e-08 2.54033e-06 0.15404 0.154039 0.0120233 2.60383e-05 0.00115469 0.192549 0.000658916 0.193204 0.972005 101.292 0.232558 0.884539 4.70823 0.0674425 0.0444173 0.955583 0.0193033 0.0047054 0.0185557 0.00447922 0.00569673 0.00644427 0.227869 0.257771 58.0634 -87.9 126.108 15.9266 145.04 0.000142788 0.267359 192.689 0.310094 0.067313 0.00409918 0.000562532 0.00138559 0.986953 0.991713 -2.99356e-06 -85.6549 0.0931052 31163.9 313.102 0.983493 0.319146 0.740711 0.740707 9.99958 2.98759e-06 1.19503e-05 0.135358 0.983452 0.931133 -0.0132913 4.9373e-06 0.520694 -2.05024e-20 7.616e-24 -2.04948e-20 0.00139672 0.997814 8.60412e-05 0.152767 2.853 0.00139672 0.997815 0.805681 0.00107108 0.00188173 0.000860412 0.455335 0.00188173 0.445581 0.00013177 1.02 0.889012 0.534307 0.287898 1.72006e-07 3.08937e-09 2367.18 3149.64 -0.0592539 0.482225 0.277212 0.255459 -0.592936 -0.169588 0.484284 -0.265324 -0.21897 2.883 1 0 294.396 0 2.2651 2.881 0.000298826 0.873635 0.709785 0.307307 0.439116 2.26527 140.792 83.5189 18.6976 60.6727 0.00404191 0 -40 10
1.982 5.73132e-08 2.54033e-06 0.154067 0.154067 0.0120233 2.60514e-05 0.0011547 0.192584 0.000658917 0.193238 0.972098 101.291 0.232547 0.884674 4.70896 0.0674535 0.0444241 0.955576 0.0193027 0.0047059 0.0185551 0.00447965 0.00569735 0.0064449 0.227894 0.257796 58.0634 -87.9 126.108 15.9265 145.041 0.00014279 0.267359 192.689 0.310094 0.0673129 0.00409918 0.000562533 0.00138559 0.986953 0.991713 -2.99357e-06 -85.6549 0.0931053 31163.9 313.115 0.983493 0.319146 0.740723 0.740719 9.99958 2.9876e-06 1.19503e-05 0.135363 0.983452 0.931132 -0.0132913 4.93733e-06 0.520716 -2.05041e-20 7.61669e-24 -2.04965e-20 0.00139672 0.997814 8.60413e-05 0.152767 2.853 0.00139672 0.997815 0.805748 0.0010711 0.00188173 0.000860413 0.455335 0.00188173 0.445586 0.000131773 1.02 0.889014 0.534307 0.287899 1.72007e-07 3.08939e-09 2367.16 3149.69 -0.059259 0.482225 0.277212 0.255462 -0.592936 -0.169588 0.484268 -0.265322 -0.218956 2.884 1 0 294.391 0 2.26523 2.882 0.000298825 0.873665 0.709827 0.307272 0.439138 2.26541 140.799 83.5183 18.6976 60.6724 0.00404193 0 -40 10
1.983 5.7342e-08 2.54033e-06 0.154095 0.154094 0.0120232 2.60645e-05 0.0011547 0.192618 0.000658917 0.193272 0.972191 101.29 0.232536 0.884809 4.70968 0.0674645 0.044431 0.955569 0.019302 0.00470639 0.0185545 0.00448008 0.00569796 0.00644554 0.227918 0.257822 58.0635 -87.9 126.108 15.9265 145.041 0.000142792 0.267359 192.689 0.310094 0.0673129 0.00409918 0.000562533 0.00138559 0.986953 0.991713 -2.99359e-06 -85.6549 0.0931054 31163.8 313.129 0.983493 0.319146 0.740735 0.740731 9.99958 2.9876e-06 1.19503e-05 0.135368 0.983452 0.931131 -0.0132913 4.93736e-06 0.520738 -2.05059e-20 7.61738e-24 -2.04982e-20 0.00139672 0.997814 8.60413e-05 0.152767 2.853 0.00139672 0.997815 0.805815 0.00107111 0.00188173 0.000860413 0.455335 0.00188173 0.445591 0.000131775 1.02 0.889015 0.534307 0.287901 1.72007e-07 3.08942e-09 2367.15 3149.74 -0.0592641 0.482225 0.277212 0.255465 -0.592935 -0.169588 0.484251 -0.265319 -0.218941 2.885 1 0 294.387 0 2.26537 2.883 0.000298823 0.873696 0.70987 0.307237 0.43916 2.26554 140.806 83.5176 18.6975 60.6721 0.00404196 0 -40 10
1.984 5.73708e-08 2.54033e-06 0.154122 0.154122 0.0120232 2.60776e-05 0.0011547 0.192652 0.000658917 0.193307 0.972284 101.29 0.232525 0.884944 4.71041 0.0674755 0.0444378 0.955562 0.0193014 0.00470689 0.0185538 0.00448051 0.00569857 0.00644617 0.227943 0.257847 58.0636 -87.9 126.107 15.9265 145.041 0.000142795 0.267359 192.689 0.310093 0.0673128 0.00409919 0.000562534 0.0013856 0.986953 0.991712 -2.9936e-06 -85.6549 0.0931055 31163.8 313.142 0.983493 0.319146 0.740748 0.740743 9.99958 2.98761e-06 1.19503e-05 0.135373 0.983452 0.931129 -0.0132913 4.93738e-06 0.520759 -2.05076e-20 7.61807e-24 -2.05e-20 0.00139672 0.997814 8.60414e-05 0.152767 2.853 0.00139672 0.997814 0.805883 0.00107113 0.00188174 0.000860414 0.455335 0.00188173 0.445595 0.000131777 1.02 0.889016 0.534306 0.287902 1.72007e-07 3.08944e-09 2367.13 3149.79 -0.0592693 0.482225 0.277211 0.255469 -0.592935 -0.169588 0.484235 -0.265317 -0.218927 2.886 1 0 294.382 0 2.2655 2.884 0.000298822 0.873726 0.709912 0.307202 0.439181 2.26568 140.813 83.517 18.6975 60.6718 0.00404198 0 -40 10
1.985 5.73996e-08 2.54034e-06 0.154149 0.154149 0.0120232 2.60907e-05 0.0011547 0.192687 0.000658918 0.193341 0.972377 101.289 0.232514 0.885079 4.71114 0.0674864 0.0444447 0.955555 0.0193008 0.00470738 0.0185532 0.00448094 0.00569918 0.0064468 0.227967 0.257872 58.0636 -87.9 126.107 15.9264 145.041 0.000142797 0.26736 192.689 0.310093 0.0673128 0.00409919 0.000562535 0.0013856 0.986953 0.991712 -2.99362e-06 -85.6549 0.0931056 31163.8 313.156 0.983493 0.319146 0.74076 0.740756 9.99958 2.98761e-06 1.19503e-05 0.135378 0.983452 0.931128 -0.0132913 4.93741e-06 0.520781 -2.05093e-20 7.61876e-24 -2.05017e-20 0.00139672 0.997814 8.60415e-05 0.152768 2.853 0.00139672 0.997814 0.80595 0.00107114 0.00188174 0.000860415 0.455334 0.00188174 0.4456 0.000131779 1.02 0.889017 0.534306 0.287904 1.72007e-07 3.08946e-09 2367.12 3149.85 -0.0592744 0.482225 0.277211 0.255472 -0.592934 -0.169588 0.484219 -0.265315 -0.218913 2.887 1 0 294.377 0 2.26564 2.885 0.000298821 0.873756 0.709954 0.307167 0.439203 2.26581 140.821 83.5164 18.6974 60.6715 0.00404201 0 -40 10
1.986 5.74284e-08 2.54034e-06 0.154177 0.154176 0.0120232 2.61038e-05 0.0011547 0.192721 0.000658918 0.193375 0.97247 101.288 0.232503 0.885215 4.71187 0.0674974 0.0444516 0.955548 0.0193002 0.00470788 0.0185526 0.00448137 0.00569979 0.00644744 0.227992 0.257898 58.0637 -87.9 126.107 15.9264 145.041 0.000142799 0.26736 192.689 0.310092 0.0673127 0.00409919 0.000562535 0.0013856 0.986953 0.991712 -2.99363e-06 -85.6548 0.0931057 31163.8 313.169 0.983493 0.319146 0.740772 0.740768 9.99958 2.98762e-06 1.19504e-05 0.135383 0.983453 0.931127 -0.0132913 4.93744e-06 0.520803 -2.0511e-20 7.61945e-24 -2.05034e-20 0.00139672 0.997814 8.60416e-05 0.152768 2.853 0.00139672 0.997814 0.806017 0.00107116 0.00188174 0.000860416 0.455334 0.00188174 0.445604 0.000131782 1.02 0.889018 0.534306 0.287905 1.72008e-07 3.08949e-09 2367.1 3149.9 -0.0592796 0.482225 0.277211 0.255475 -0.592933 -0.169588 0.484203 -0.265313 -0.218899 2.888 1 0 294.373 0 2.26577 2.886 0.000298819 0.873787 0.709996 0.307132 0.439225 2.26595 140.828 83.5158 18.6974 60.6712 0.00404203 0 -40 10
1.987 5.74573e-08 2.54034e-06 0.154204 0.154204 0.0120232 2.61169e-05 0.0011547 0.192755 0.000658919 0.19341 0.972563 101.287 0.232492 0.88535 4.7126 0.0675084 0.0444585 0.955542 0.0192996 0.00470837 0.0185519 0.0044818 0.0057004 0.00644807 0.228016 0.257923 58.0637 -87.9 126.107 15.9264 145.041 0.000142802 0.26736 192.688 0.310092 0.0673127 0.0040992 0.000562536 0.0013856 0.986953 0.991712 -2.99365e-06 -85.6548 0.0931058 31163.7 313.183 0.983493 0.319146 0.740785 0.74078 9.99958 2.98762e-06 1.19504e-05 0.135388 0.983453 0.931126 -0.0132913 4.93747e-06 0.520824 -2.05128e-20 7.62014e-24 -2.05052e-20 0.00139672 0.997814 8.60417e-05 0.152768 2.853 0.00139672 0.997814 0.806084 0.00107118 0.00188174 0.000860417 0.455334 0.00188174 0.445609 0.000131784 1.02 0.889019 0.534306 0.287907 1.72008e-07 3.08951e-09 2367.08 3149.95 -0.0592847 0.482225 0.27721 0.255479 -0.592933 -0.169588 0.484186 -0.265311 -0.218885 2.889 1 0 294.368 0 2.26591 2.887 0.000298818 0.873817 0.710039 0.307097 0.439247 2.26608 140.835 83.5152 18.6974 60.6709 0.00404206 0 -40 10
1.988 5.74861e-08 2.54034e-06 0.154232 0.154231 0.0120232 2.613e-05 0.0011547 0.192789 0.000658919 0.193444 0.972656 101.287 0.232481 0.885485 4.71333 0.0675194 0.0444653 0.955535 0.019299 0.00470887 0.0185513 0.00448223 0.00570101 0.00644871 0.228041 0.257948 58.0638 -87.9 126.107 15.9263 145.041 0.000142804 0.26736 192.688 0.310091 0.0673126 0.0040992 0.000562537 0.0013856 0.986953 0.991712 -2.99366e-06 -85.6548 0.0931059 31163.7 313.196 0.983493 0.319146 0.740797 0.740792 9.99958 2.98763e-06 1.19504e-05 0.135393 0.983453 0.931125 -0.0132913 4.9375e-06 0.520846 -2.05145e-20 7.62083e-24 -2.05069e-20 0.00139673 0.997814 8.60417e-05 0.152768 2.853 0.00139673 0.997814 0.806152 0.00107119 0.00188174 0.000860417 0.455334 0.00188174 0.445614 0.000131786 1.02 0.88902 0.534305 0.287908 1.72008e-07 3.08953e-09 2367.07 3150 -0.0592898 0.482225 0.27721 0.255482 -0.592932 -0.169588 0.48417 -0.265309 -0.21887 2.89 1 0 294.364 0 2.26604 2.888 0.000298816 0.873847 0.710081 0.307062 0.439268 2.26622 140.842 83.5146 18.6973 60.6706 0.00404208 0 -40 10
1.989 5.75149e-08 2.54034e-06 0.154259 0.154259 0.0120232 2.61431e-05 0.0011547 0.192824 0.000658919 0.193478 0.972749 101.286 0.23247 0.88562 4.71405 0.0675304 0.0444722 0.955528 0.0192984 0.00470937 0.0185507 0.00448266 0.00570163 0.00644934 0.228065 0.257974 58.0639 -87.9 126.106 15.9263 145.041 0.000142807 0.26736 192.688 0.310091 0.0673126 0.0040992 0.000562537 0.00138561 0.986953 0.991712 -2.99368e-06 -85.6548 0.0931059 31163.7 313.21 0.983493 0.319146 0.740809 0.740805 9.99958 2.98763e-06 1.19504e-05 0.135398 0.983453 0.931124 -0.0132913 4.93753e-06 0.520868 -2.05162e-20 7.62152e-24 -2.05086e-20 0.00139673 0.997814 8.60418e-05 0.152768 2.853 0.00139673 0.997814 0.806219 0.00107121 0.00188174 0.000860418 0.455333 0.00188174 0.445618 0.000131788 1.02 0.889021 0.534305 0.28791 1.72008e-07 3.08955e-09 2367.05 3150.05 -0.059295 0.482225 0.27721 0.255485 -0.592931 -0.169588 0.484154 -0.265307 -0.218856 2.891 1 0 294.359 0 2.26618 2.889 0.000298815 0.873878 0.710123 0.307027 0.43929 2.26635 140.85 83.514 18.6973 60.6703 0.00404211 0 -40 10
1.99 5.75437e-08 2.54035e-06 0.154286 0.154286 0.0120231 2.61562e-05 0.0011547 0.192858 0.00065892 0.193512 0.972842 101.285 0.232459 0.885755 4.71478 0.0675414 0.0444791 0.955521 0.0192978 0.00470986 0.01855 0.0044831 0.00570224 0.00644998 0.22809 0.257999 58.0639 -87.9 126.106 15.9262 145.041 0.000142809 0.267361 192.688 0.310091 0.0673125 0.00409921 0.000562538 0.00138561 0.986953 0.991712 -2.99369e-06 -85.6548 0.093106 31163.7 313.223 0.983493 0.319146 0.740821 0.740817 9.99958 2.98764e-06 1.19504e-05 0.135403 0.983453 0.931123 -0.0132913 4.93756e-06 0.52089 -2.0518e-20 7.62221e-24 -2.05104e-20 0.00139673 0.997814 8.60419e-05 0.152768 2.85301 0.00139673 0.997814 0.806286 0.00107122 0.00188174 0.000860419 0.455333 0.00188174 0.445623 0.000131791 1.02 0.889022 0.534305 0.287911 1.72009e-07 3.08958e-09 2367.04 3150.1 -0.0593001 0.482225 0.27721 0.255489 -0.592931 -0.169588 0.484137 -0.265305 -0.218842 2.892 1 0 294.354 0 2.26631 2.89 0.000298814 0.873908 0.710165 0.306993 0.439312 2.26649 140.857 83.5134 18.6973 60.67 0.00404213 0 -40 10
1.991 5.75725e-08 2.54035e-06 0.154314 0.154313 0.0120231 2.61693e-05 0.0011547 0.192892 0.00065892 0.193546 0.972935 101.284 0.232448 0.88589 4.71552 0.0675524 0.044486 0.955514 0.0192971 0.00471036 0.0185494 0.00448353 0.00570285 0.00645061 0.228114 0.258024 58.064 -87.9 126.106 15.9262 145.041 0.000142811 0.267361 192.688 0.31009 0.0673125 0.00409921 0.000562539 0.00138561 0.986953 0.991712 -2.99371e-06 -85.6548 0.0931061 31163.6 313.237 0.983493 0.319146 0.740834 0.740829 9.99958 2.98764e-06 1.19505e-05 0.135408 0.983453 0.931122 -0.0132913 4.93759e-06 0.520911 -2.05197e-20 7.6229e-24 -2.05121e-20 0.00139673 0.997814 8.6042e-05 0.152769 2.85301 0.00139673 0.997814 0.806353 0.00107124 0.00188175 0.00086042 0.455333 0.00188174 0.445628 0.000131793 1.02 0.889023 0.534304 0.287913 1.72009e-07 3.0896e-09 2367.02 3150.16 -0.0593052 0.482225 0.277209 0.255492 -0.59293 -0.169588 0.484121 -0.265303 -0.218828 2.893 1 0 294.35 0 2.26645 2.891 0.000298812 0.873938 0.710208 0.306958 0.439333 2.26662 140.864 83.5128 18.6972 60.6698 0.00404216 0 -40 10
1.992 5.76014e-08 2.54035e-06 0.154341 0.15434 0.0120231 2.61824e-05 0.0011547 0.192926 0.000658921 0.19358 0.973028 101.284 0.232437 0.886025 4.71625 0.0675634 0.0444929 0.955507 0.0192965 0.00471086 0.0185488 0.00448396 0.00570346 0.00645125 0.228139 0.25805 58.0641 -87.9 126.106 15.9262 145.041 0.000142814 0.267361 192.688 0.31009 0.0673124 0.00409921 0.000562539 0.00138561 0.986953 0.991712 -2.99372e-06 -85.6548 0.0931062 31163.6 313.25 0.983493 0.319146 0.740846 0.740842 9.99958 2.98765e-06 1.19505e-05 0.135413 0.983453 0.931121 -0.0132913 4.93762e-06 0.520933 -2.05215e-20 7.62359e-24 -2.05138e-20 0.00139673 0.997814 8.60421e-05 0.152769 2.85301 0.00139673 0.997814 0.80642 0.00107125 0.00188175 0.000860421 0.455333 0.00188175 0.445632 0.000131795 1.02 0.889024 0.534304 0.287914 1.72009e-07 3.08962e-09 2367 3150.21 -0.0593104 0.482225 0.277209 0.255495 -0.592929 -0.169588 0.484105 -0.265301 -0.218814 2.894 1 0 294.345 0 2.26658 2.892 0.000298811 0.873969 0.71025 0.306923 0.439355 2.26675 140.871 83.5122 18.6972 60.6695 0.00404218 0 -40 10
1.993 5.76302e-08 2.54035e-06 0.154368 0.154368 0.0120231 2.61955e-05 0.00115471 0.19296 0.000658921 0.193614 0.973121 101.283 0.232426 0.88616 4.71698 0.0675744 0.0444998 0.9555 0.0192959 0.00471135 0.0185481 0.00448439 0.00570408 0.00645188 0.228163 0.258075 58.0641 -87.9 126.105 15.9261 145.041 0.000142816 0.267361 192.687 0.310089 0.0673124 0.00409921 0.00056254 0.00138561 0.986953 0.991712 -2.99374e-06 -85.6548 0.0931063 31163.6 313.264 0.983493 0.319146 0.740858 0.740854 9.99958 2.98765e-06 1.19505e-05 0.135418 0.983453 0.93112 -0.0132913 4.93765e-06 0.520955 -2.05232e-20 7.62429e-24 -2.05156e-20 0.00139673 0.997814 8.60422e-05 0.152769 2.85301 0.00139673 0.997814 0.806487 0.00107127 0.00188175 0.000860422 0.455333 0.00188175 0.445637 0.000131797 1.02 0.889026 0.534304 0.287916 1.7201e-07 3.08965e-09 2366.99 3150.26 -0.0593155 0.482226 0.277209 0.255498 -0.592929 -0.169588 0.484088 -0.265299 -0.218799 2.895 1 0 294.34 0 2.26671 2.893 0.000298809 0.873999 0.710292 0.306888 0.439377 2.26689 140.878 83.5116 18.6972 60.6692 0.00404221 0 -40 10
1.994 5.7659e-08 2.54035e-06 0.154395 0.154395 0.0120231 2.62086e-05 0.00115471 0.192994 0.000658921 0.193648 0.973214 101.282 0.232415 0.886296 4.71771 0.0675854 0.0445067 0.955493 0.0192953 0.00471185 0.0185475 0.00448483 0.00570469 0.00645252 0.228188 0.258101 58.0642 -87.9 126.105 15.9261 145.041 0.000142818 0.267361 192.687 0.310089 0.0673123 0.00409922 0.000562541 0.00138562 0.986953 0.991712 -2.99375e-06 -85.6548 0.0931064 31163.6 313.277 0.983493 0.319146 0.740871 0.740866 9.99958 2.98766e-06 1.19505e-05 0.135423 0.983454 0.931119 -0.0132913 4.93768e-06 0.520977 -2.05249e-20 7.62498e-24 -2.05173e-20 0.00139673 0.997814 8.60422e-05 0.152769 2.85301 0.00139673 0.997814 0.806554 0.00107128 0.00188175 0.000860422 0.455332 0.00188175 0.445641 0.0001318 1.02 0.889027 0.534303 0.287917 1.7201e-07 3.08967e-09 2366.97 3150.31 -0.0593206 0.482226 0.277208 0.255502 -0.592928 -0.169588 0.484072 -0.265296 -0.218785 2.896 1 0 294.336 0 2.26685 2.894 0.000298808 0.874029 0.710334 0.306853 0.439398 2.26702 140.886 83.511 18.6971 60.6689 0.00404223 0 -40 10
1.995 5.76878e-08 2.54036e-06 0.154423 0.154422 0.0120231 2.62217e-05 0.00115471 0.193028 0.000658922 0.193683 0.973307 101.282 0.232404 0.886431 4.71844 0.0675964 0.0445136 0.955486 0.0192947 0.00471235 0.0185468 0.00448526 0.0057053 0.00645315 0.228212 0.258126 58.0642 -87.9 126.105 15.9261 145.041 0.000142821 0.267361 192.687 0.310088 0.0673122 0.00409922 0.000562541 0.00138562 0.986953 0.991712 -2.99377e-06 -85.6548 0.0931065 31163.6 313.291 0.983493 0.319146 0.740883 0.740879 9.99958 2.98766e-06 1.19505e-05 0.135429 0.983454 0.931118 -0.0132913 4.93771e-06 0.520998 -2.05267e-20 7.62567e-24 -2.0519e-20 0.00139673 0.997814 8.60423e-05 0.152769 2.85301 0.00139673 0.997814 0.806621 0.0010713 0.00188175 0.000860423 0.455332 0.00188175 0.445646 0.000131802 1.02 0.889028 0.534303 0.287919 1.7201e-07 3.08969e-09 2366.95 3150.36 -0.0593258 0.482226 0.277208 0.255505 -0.592927 -0.169588 0.484056 -0.265294 -0.218771 2.897 1 0 294.331 0 2.26698 2.895 0.000298806 0.87406 0.710377 0.306819 0.43942 2.26716 140.893 83.5104 18.6971 60.6686 0.00404226 0 -40 10
1.996 5.77166e-08 2.54036e-06 0.15445 0.154449 0.0120231 2.62348e-05 0.00115471 0.193062 0.000658922 0.193717 0.9734 101.281 0.232393 0.886566 4.71917 0.0676075 0.0445205 0.955479 0.0192941 0.00471284 0.0185462 0.00448569 0.00570592 0.00645379 0.228237 0.258152 58.0643 -87.9 126.105 15.926 145.041 0.000142823 0.267362 192.687 0.310088 0.0673122 0.00409922 0.000562542 0.00138562 0.986953 0.991712 -2.99378e-06 -85.6548 0.0931066 31163.5 313.304 0.983493 0.319146 0.740895 0.740891 9.99958 2.98767e-06 1.19506e-05 0.135434 0.983454 0.931117 -0.0132913 4.93774e-06 0.52102 -2.05284e-20 7.62636e-24 -2.05208e-20 0.00139674 0.997814 8.60424e-05 0.152769 2.85301 0.00139674 0.997814 0.806688 0.00107132 0.00188175 0.000860424 0.455332 0.00188175 0.445651 0.000131804 1.02 0.889029 0.534303 0.28792 1.7201e-07 3.08971e-09 2366.94 3150.41 -0.0593309 0.482226 0.277208 0.255508 -0.592927 -0.169588 0.48404 -0.265292 -0.218757 2.898 1 0 294.327 0 2.26712 2.896 0.000298805 0.87409 0.710419 0.306784 0.439441 2.26729 140.9 83.5098 18.6971 60.6683 0.00404228 0 -40 10
1.997 5.77455e-08 2.54036e-06 0.154477 0.154477 0.012023 2.62479e-05 0.00115471 0.193096 0.000658923 0.19375 0.973493 101.28 0.232382 0.886701 4.71991 0.0676185 0.0445274 0.955473 0.0192935 0.00471334 0.0185456 0.00448612 0.00570653 0.00645443 0.228261 0.258177 58.0644 -87.9001 126.105 15.926 145.041 0.000142826 0.267362 192.687 0.310088 0.0673121 0.00409923 0.000562543 0.00138562 0.986953 0.991712 -2.9938e-06 -85.6547 0.0931066 31163.5 313.318 0.983493 0.319146 0.740908 0.740903 9.99958 2.98767e-06 1.19506e-05 0.135439 0.983454 0.931116 -0.0132913 4.93777e-06 0.521042 -2.05301e-20 7.62705e-24 -2.05225e-20 0.00139674 0.997814 8.60425e-05 0.152769 2.85301 0.00139674 0.997814 0.806755 0.00107133 0.00188175 0.000860425 0.455332 0.00188175 0.445655 0.000131806 1.02 0.88903 0.534302 0.287922 1.72011e-07 3.08974e-09 2366.92 3150.46 -0.0593361 0.482226 0.277208 0.255512 -0.592926 -0.169589 0.484023 -0.26529 -0.218742 2.899 1 0 294.322 0 2.26725 2.897 0.000298804 0.87412 0.710461 0.306749 0.439463 2.26743 140.907 83.5092 18.697 60.668 0.00404231 0 -40 10
1.998 5.77743e-08 2.54036e-06 0.154504 0.154504 0.012023 2.6261e-05 0.00115471 0.19313 0.000658923 0.193784 0.973586 101.279 0.232371 0.886836 4.72064 0.0676295 0.0445344 0.955466 0.0192929 0.00471384 0.0185449 0.00448656 0.00570715 0.00645506 0.228286 0.258202 58.0644 -87.9001 126.104 15.9259 145.041 0.000142828 0.267362 192.687 0.310087 0.0673121 0.00409923 0.000562543 0.00138563 0.986953 0.991712 -2.99381e-06 -85.6547 0.0931067 31163.5 313.331 0.983493 0.319146 0.74092 0.740915 9.99958 2.98768e-06 1.19506e-05 0.135444 0.983454 0.931115 -0.0132912 4.9378e-06 0.521064 -2.05319e-20 7.62775e-24 -2.05242e-20 0.00139674 0.997814 8.60426e-05 0.15277 2.85301 0.00139674 0.997814 0.806822 0.00107135 0.00188176 0.000860426 0.455331 0.00188176 0.44566 0.000131809 1.02 0.889031 0.534302 0.287923 1.72011e-07 3.08976e-09 2366.91 3150.52 -0.0593412 0.482226 0.277207 0.255515 -0.592925 -0.169589 0.484007 -0.265288 -0.218728 2.9 1 0 294.317 0 2.26739 2.898 0.000298802 0.874151 0.710503 0.306715 0.439485 2.26756 140.915 83.5086 18.697 60.6677 0.00404233 0 -40 10
1.999 5.78031e-08 2.54036e-06 0.154531 0.154531 0.012023 2.62741e-05 0.00115471 0.193164 0.000658923 0.193818 0.97368 101.279 0.23236 0.886971 4.72138 0.0676405 0.0445413 0.955459 0.0192922 0.00471434 0.0185443 0.00448699 0.00570776 0.0064557 0.22831 0.258228 58.0645 -87.9001 126.104 15.9259 145.041 0.00014283 0.267362 192.686 0.310087 0.067312 0.00409923 0.000562544 0.00138563 0.986953 0.991712 -2.99383e-06 -85.6547 0.0931068 31163.5 313.345 0.983493 0.319146 0.740932 0.740928 9.99958 2.98768e-06 1.19506e-05 0.135449 0.983454 0.931114 -0.0132912 4.93783e-06 0.521086 -2.05336e-20 7.62844e-24 -2.0526e-20 0.00139674 0.997814 8.60426e-05 0.15277 2.85301 0.00139674 0.997814 0.806889 0.00107136 0.00188176 0.000860426 0.455331 0.00188176 0.445664 0.000131811 1.02 0.889032 0.534302 0.287925 1.72011e-07 3.08978e-09 2366.89 3150.57 -0.0593463 0.482226 0.277207 0.255518 -0.592925 -0.169589 0.483991 -0.265286 -0.218714 2.901 1 0 294.313 0 2.26752 2.899 0.000298801 0.874181 0.710546 0.30668 0.439506 2.2677 140.922 83.508 18.697 60.6674 0.00404236 0 -40 10
2 5.78319e-08 2.54037e-06 0.154558 0.154558 0.012023 2.62872e-05 0.00115471 0.193198 0.000658924 0.193852 0.973773 101.278 0.232349 0.887107 4.72211 0.0676515 0.0445482 0.955452 0.0192916 0.00471483 0.0185437 0.00448742 0.00570837 0.00645634 0.228335 0.258253 58.0645 -87.9001 126.104 15.9259 145.041 0.000142833 0.267362 192.686 0.310086 0.067312 0.00409924 0.000562545 0.00138563 0.986953 0.991712 -2.99384e-06 -85.6547 0.0931069 31163.4 313.358 0.983493 0.319146 0.740944 0.74094 9.99958 2.98769e-06 1.19506e-05 0.135454 0.983454 0.931113 -0.0132912 4.93786e-06 0.521107 -2.05354e-20 7.62913e-24 -2.05277e-20 0.00139674 0.997814 8.60427e-05 0.15277 2.85301 0.00139674 0.997814 0.806956 0.00107138 0.00188176 0.000860427 0.455331 0.00188176 0.445669 0.000131813 1.02 0.889033 0.534302 0.287927 1.72011e-07 3.08981e-09 2366.87 3150.62 -0.0593515 0.482226 0.277207 0.255521 -0.592924 -0.169589 0.483974 -0.265284 -0.2187 2.902 1 0 294.308 0 2.26766 2.9 0.000298799 0.874212 0.710588 0.306645 0.439528 2.26783 140.929 83.5074 18.6969 60.6671 0.00404238 0 -40 10
2.001 5.78607e-08 2.54037e-06 0.154585 0.154585 0.012023 2.63003e-05 0.00115471 0.193232 0.000658924 0.193886 0.973866 101.277 0.232338 0.887242 4.72285 0.0676625 0.0445551 0.955445 0.019291 0.00471533 0.018543 0.00448786 0.00570899 0.00645697 0.22836 0.258279 58.0646 -87.9001 126.104 15.9258 145.041 0.000142835 0.267363 192.686 0.310086 0.0673119 0.00409924 0.000562545 0.00138563 0.986953 0.991712 -2.99386e-06 -85.6547 0.093107 31163.4 313.372 0.983492 0.319146 0.740957 0.740952 9.99958 2.98769e-06 1.19507e-05 0.135459 0.983454 0.931112 -0.0132912 4.93789e-06 0.521129 -2.05371e-20 7.62983e-24 -2.05295e-20 0.00139674 0.997814 8.60428e-05 0.15277 2.85302 0.00139674 0.997814 0.807023 0.00107139 0.00188176 0.000860428 0.455331 0.00188176 0.445674 0.000131815 1.02 0.889034 0.534301 0.287928 1.72012e-07 3.08983e-09 2366.86 3150.67 -0.0593566 0.482226 0.277207 0.255525 -0.592924 -0.169589 0.483958 -0.265282 -0.218686 2.903 1 0 294.303 0 2.26779 2.901 0.000298798 0.874242 0.71063 0.306611 0.43955 2.26797 140.936 83.5068 18.6969 60.6668 0.00404241 0 -40 10
2.002 5.78896e-08 2.54037e-06 0.154612 0.154612 0.012023 2.63134e-05 0.00115471 0.193266 0.000658924 0.19392 0.973959 101.276 0.232327 0.887377 4.72358 0.0676735 0.0445621 0.955438 0.0192904 0.00471583 0.0185424 0.00448829 0.0057096 0.00645761 0.228384 0.258304 58.0647 -87.9001 126.103 15.9258 145.041 0.000142837 0.267363 192.686 0.310085 0.0673119 0.00409924 0.000562546 0.00138563 0.986953 0.991712 -2.99387e-06 -85.6547 0.0931071 31163.4 313.385 0.983492 0.319146 0.740969 0.740965 9.99958 2.9877e-06 1.19507e-05 0.135464 0.983455 0.931111 -0.0132912 4.93792e-06 0.521151 -2.05388e-20 7.63052e-24 -2.05312e-20 0.00139674 0.997814 8.60429e-05 0.15277 2.85302 0.00139674 0.997814 0.80709 0.00107141 0.00188176 0.000860429 0.45533 0.00188176 0.445678 0.000131817 1.02 0.889035 0.534301 0.28793 1.72012e-07 3.08985e-09 2366.84 3150.72 -0.0593617 0.482226 0.277206 0.255528 -0.592923 -0.169589 0.483942 -0.26528 -0.218671 2.904 1 0 294.299 0 2.26793 2.902 0.000298797 0.874272 0.710672 0.306576 0.439571 2.2681 140.944 83.5062 18.6968 60.6665 0.00404243 0 -40 10
2.003 5.79184e-08 2.54037e-06 0.154639 0.154639 0.012023 2.63265e-05 0.00115471 0.193299 0.000658925 0.193954 0.974052 101.276 0.232315 0.887512 4.72432 0.0676845 0.044569 0.955431 0.0192898 0.00471633 0.0185418 0.00448873 0.00571022 0.00645825 0.228409 0.25833 58.0647 -87.9001 126.103 15.9258 145.041 0.00014284 0.267363 192.686 0.310085 0.0673118 0.00409924 0.000562547 0.00138564 0.986953 0.991712 -2.99389e-06 -85.6547 0.0931072 31163.4 313.399 0.983492 0.319146 0.740981 0.740977 9.99958 2.9877e-06 1.19507e-05 0.135469 0.983455 0.931109 -0.0132912 4.93795e-06 0.521173 -2.05406e-20 7.63121e-24 -2.05329e-20 0.00139674 0.997814 8.6043e-05 0.15277 2.85302 0.00139674 0.997814 0.807157 0.00107142 0.00188176 0.00086043 0.45533 0.00188176 0.445683 0.00013182 1.02 0.889037 0.534301 0.287931 1.72012e-07 3.08987e-09 2366.82 3150.77 -0.0593669 0.482226 0.277206 0.255531 -0.592922 -0.169589 0.483925 -0.265278 -0.218657 2.905 1 0 294.294 0 2.26806 2.903 0.000298795 0.874303 0.710714 0.306541 0.439593 2.26824 140.951 83.5056 18.6968 60.6663 0.00404246 0 -40 10
2.004 5.79472e-08 2.54037e-06 0.154667 0.154666 0.0120229 2.63396e-05 0.00115471 0.193333 0.000658925 0.193987 0.974145 101.275 0.232304 0.887647 4.72505 0.0676955 0.044576 0.955424 0.0192892 0.00471683 0.0185411 0.00448916 0.00571083 0.00645889 0.228433 0.258355 58.0648 -87.9001 126.103 15.9257 145.041 0.000142842 0.267363 192.686 0.310085 0.0673118 0.00409925 0.000562547 0.00138564 0.986953 0.991712 -2.9939e-06 -85.6547 0.0931073 31163.4 313.413 0.983492 0.319146 0.740994 0.740989 9.99958 2.98771e-06 1.19507e-05 0.135474 0.983455 0.931108 -0.0132912 4.93798e-06 0.521195 -2.05423e-20 7.63191e-24 -2.05347e-20 0.00139674 0.997814 8.6043e-05 0.152771 2.85302 0.00139674 0.997814 0.807223 0.00107144 0.00188177 0.00086043 0.45533 0.00188176 0.445687 0.000131822 1.02 0.889038 0.5343 0.287933 1.72012e-07 3.0899e-09 2366.81 3150.83 -0.059372 0.482226 0.277206 0.255535 -0.592922 -0.169589 0.483909 -0.265276 -0.218643 2.906 1 0 294.289 0 2.2682 2.904 0.000298794 0.874333 0.710757 0.306507 0.439615 2.26837 140.958 83.505 18.6968 60.666 0.00404248 0 -40 10
