time,L,R,Gs,b1ARtot,b1ARd,b1ARp,Gsagtptot,Gsagdp,Gsbg,Gsa_gtp,Fsk,AC,PDE,IBMX,cAMPtot,cAMP,PKACI,PKACII,PLBs,Inhib1ptot,Inhib1p,PP1,LCCap,LCCbp,m,h,j,v,w,x,y,z,rto,sto,ssto,rss,sss,Ca_nsr,Ca_jsr,Nai,Ki,Cai,Vm,trel
0 0.988 0.01079 3.829 0.01205 0 0.001154 0.02505 0.0006446 0.02569 0.02241 0 0.04706 0.0389 0 0.8453 0.2268 0.05868 0.008278 4.105 0.0526 6.3e-05 0.838 0.005103 0.005841 0.0014 0.99 0.99 0 0 0.13 0.96 0.92 0.0014 1 0.613 0.198 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
1.6828e-08 0.98801 5.5988e-05 3.8182 0.01205 2.2189e-13 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013999 0.99 0.99 1.5651e-09 3.131e-09 0.13 0.96 0.92 0.0014 1 0.613 0.198 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
3.3655e-08 0.98801 5.3039e-05 3.8182 0.01205 4.4384e-13 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013999 0.99 0.99 3.1294e-09 6.2613e-09 0.13 0.96 0.92 0.0014 1 0.613 0.19799 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
6.731e-08 0.98801 5.64e-05 3.8182 0.01205 8.8764e-13 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013998 0.99 0.99 6.2561e-09 1.252e-08 0.13 0.96 0.92 0.0014 1 0.613 0.19798 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
8.4138e-08 0.98801 5.2507e-05 3.8182 0.01205 1.1095e-12 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013997 0.99 0.99 7.8184e-09 1.5648e-08 0.13 0.96 0.92 0.0014 1 0.613 0.19798 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
1.1779e-07 0.98801 5.5256e-05 3.8182 0.01205 1.5533e-12 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013996 0.99 0.99 1.094e-08 2.1902e-08 0.13 0.96 0.92 0.0014 1 0.613 0.19797 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
1.851e-07 0.98801 5.5256e-05 3.8182 0.01205 2.4409e-12 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013995 0.99 0.99 1.7175e-08 3.44e-08 0.13 0.96 0.92 0.0014 1 0.613 0.19796 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
3.1972e-07 0.98801 5.5256e-05 3.8182 0.01205 4.2161e-12 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013991 0.99 0.99 2.9605e-08 5.9357e-08 0.13 0.96 0.92 0.0014 1 0.613 0.19793 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
5.8896e-07 0.98801 5.5256e-05 3.8182 0.01205 7.7669e-12 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013983 0.99 0.99 5.4311e-08 1.0912e-07 0.13 0.96 0.92 0.0014 1 0.613 0.19787 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
1.1274e-06 0.98801 5.5256e-05 3.8182 0.01205 1.4867e-11 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.001397 0.99 0.99 1.0309e-07 2.08e-07 0.13 0.96 0.92 0.0013999 1 0.613 0.19774 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
2.2044e-06 0.98801 5.5256e-05 3.8182 0.01205 2.9074e-11 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013946 0.99 0.99 1.9828e-07 4.0334e-07 0.13 0.96 0.92 0.0013999 1 0.613 0.1975 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
4.3583e-06 0.98801 5.5256e-05 3.8182 0.01205 5.7461e-11 0.001154 0.025051 0.0006446 0.025691 0.022414 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013912 0.99 0.99 3.791e-07 7.8408e-07 0.13 0.96 0.92 0.0013998 1 0.613 0.19701 0.43 1.92 1.92 16 145 0.000158 -85.6601 0.9
6.5123e-06 0.98801 5.5256e-05 3.8182 0.01205 8.5855e-11 0.001154 0.025051 0.0006446 0.025691 0.022414 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013889 0.98999 0.99 5.4823e-07 1.1523e-06 0.13001 0.96 0.92 0.0013997 1 0.613 0.19652 0.43 1.92 1.92 16 145 0.000158 -85.6601 0.90001
1.082e-05 0.98801 5.5256e-05 3.8182 0.01205 1.4262e-10 0.001154 0.025052 0.0006446 0.025692 0.022415 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013867 0.98999 0.99 8.5396e-07 1.8525e-06 0.13001 0.96 0.92 0.0013995 1 0.613 0.19555 0.43 1.92 1.92 16 145 0.000158 -85.6601 0.90001
1.5128e-05 0.98801 5.5256e-05 3.8182 0.01205 1.9941e-10 0.001154 0.025053 0.0006446 0.025693 0.022415 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013854 0.98999 0.99 1.1226e-06 2.508e-06 0.13002 0.96 0.92 0.0013994 1 0.613 0.19458 0.43 1.92 1.92 16 145 0.000158 -85.6602 0.90002
1.9436e-05 0.98801 5.5256e-05 3.8182 0.01205 2.5622e-10 0.001154 0.025053 0.0006446 0.025693 0.022416 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013847 0.98998 0.99 1.3574e-06 3.1211e-06 0.13002 0.96 0.92 0.0013992 1 0.613 0.19362 0.43 1.92 1.92 16 145 0.000158 -85.6603 0.90002
2.8051e-05 0.98801 5.5256e-05 3.8182 0.01205 3.6983e-10 0.001154 0.025055 0.0006446 0.025695 0.022417 0 0.047062 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013842 0.98997 0.99 1.7469e-06 4.2338e-06 0.13003 0.96 0.92 0.0013989 1 0.613 0.19171 0.43 1.92 1.92 16 145 0.000158 -85.6604 0.90003
3.6667e-05 0.98801 5.5256e-05 3.8182 0.01205 4.8344e-10 0.001154 0.025056 0.0006446 0.025696 0.022419 0 0.047062 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013842 0.98997 0.99 2.045e-06 5.2074e-06 0.13004 0.96 0.92 0.0013986 1 0.613 0.18981 0.43 1.92 1.92 16 145 0.000158 -85.6605 0.90004
5.3899e-05 0.98801 5.5256e-05 3.8182 0.01205 7.1067e-10 0.001154 0.025059 0.0006446 0.025699 0.022421 0 0.047062 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013842 0.98995 0.99001 2.4615e-06 6.8195e-06 0.13005 0.96 0.92 0.0013982 1 0.61301 0.18608 0.43 1.92 1.92 16 145 0.000158 -85.6607 0.90005
7.113e-05 0.98801 5.5256e-05 3.8182 0.01205 9.379e-10 0.001154 0.025062 0.0006446 0.025702 0.022424 0 0.047062 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013842 0.98993 0.99001 2.7016e-06 8.0526e-06 0.13007 0.96001 0.92 0.0013978 1 0.61301 0.18243 0.43 1.92 1.92 16 145 0.000158 -85.6609 0.90007
0.00010559 0.98801 5.5256e-05 3.8182 0.01205 1.3924e-09 0.001154 0.025068 0.0006446 0.025708 0.022429 0 0.047061 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013841 0.9899 0.99001 2.9471e-06 9.7751e-06 0.13009 0.96001 0.92 0.0013971 1 0.61301 0.17533 0.43 1.92 1.92 16 145 0.00015799 -85.6614 0.90011
0.00013661 0.98801 5.5256e-05 3.8182 0.01205 1.8014e-09 0.001154 0.025073 0.0006446 0.025713 0.022434 0 0.047061 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.001384 0.98987 0.99002 3.0034e-06 1.0681e-05 0.13012 0.96001 0.92001 0.0013967 1 0.61302 0.16919 0.43 1.9201 1.92 16 145 0.00015799 -85.6618 0.90014
0.00016763 0.98801 5.5256e-05 3.8182 0.01205 2.2104e-09 0.001154 0.025078 0.0006446 0.025718 0.022438 0 0.04706 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013839 0.98984 0.99002 3.0081e-06 1.1221e-05 0.13014 0.96001 0.92001 0.0013965 1 0.61302 0.16326 0.43 1.9201 1.92 16 145 0.00015799 -85.6621 0.90017
0.00019864 0.98801 5.5256e-05 3.8182 0.01205 2.6194e-09 0.001154 0.025084 0.0006446 0.025724 0.022443 0 0.04706 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013839 0.98982 0.99002 2.9997e-06 1.1535e-05 0.13016 0.96001 0.92001 0.0013963 1 0.61303 0.15753 0.43 1.9201 1.92 16 145 0.00015799 -85.6625 0.9002
0.00022966 0.98801 5.5256e-05 3.8182 0.01205 3.0284e-09 0.001154 0.025089 0.0006446 0.025729 0.022448 0 0.047059 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013838 0.98979 0.99003 2.9918e-06 1.1713e-05 0.13018 0.96002 0.92001 0.0013961 1 0.61303 0.15202 0.43 1.9201 1.92 16 145 0.00015799 -85.6628 0.90023
0.00029169 0.98801 5.5256e-05 3.8182 0.01205 3.8465e-09 0.001154 0.025099 0.0006446 0.025739 0.022457 0 0.047058 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013836 0.98973 0.99003 2.9792e-06 1.1829e-05 0.13021 0.96002 0.92001 0.0013959 0.99999 0.61304 0.14156 0.43 1.9201 1.92 16 145 0.00015798 -85.6634 0.90029
0.00035372 0.98801 5.5256e-05 3.8182 0.01205 4.6645e-09 0.001154 0.02511 0.0006446 0.02575 0.022467 0 0.047057 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013835 0.98968 0.99004 2.9785e-06 1.1858e-05 0.13024 0.96003 0.92002 0.0013958 0.99999 0.61305 0.13184 0.43 1.9201 1.92 16 145 0.00015798 -85.664 0.90035
0.00041576 0.98801 5.5256e-05 3.8182 0.01205 5.4826e-09 0.001154 0.02512 0.0006446 0.02576 0.022476 0 0.047056 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013834 0.98963 0.99005 2.982e-06 1.1899e-05 0.13027 0.96003 0.92002 0.0013957 0.99999 0.61306 0.12279 0.43001 1.9202 1.92 16 145 0.00015798 -85.6645 0.90042
0.00047779 0.98801 5.5256e-05 3.8182 0.01205 6.3006e-09 0.001154 0.025131 0.0006446 0.025771 0.022486 0 0.047055 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013833 0.98958 0.99006 2.9832e-06 1.1935e-05 0.13029 0.96004 0.92002 0.0013956 0.99999 0.61306 0.11437 0.43001 1.9202 1.92 16 145 0.00015797 -85.665 0.90048
0.00053982 0.98801 5.5256e-05 3.8182 0.01205 7.1186e-09 0.001154 0.025141 0.0006446 0.025781 0.022495 0 0.047054 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013832 0.98953 0.99006 2.9825e-06 1.1943e-05 0.13031 0.96004 0.92002 0.0013955 0.99999 0.61307 0.10654 0.43001 1.9202 1.92 16 145 0.00015797 -85.6655 0.90054
0.00062488 0.98801 5.5256e-05 3.8182 0.01205 8.2402e-09 0.001154 0.025155 0.0006446 0.025795 0.022508 0 0.047052 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.001383 0.98946 0.99007 2.9809e-06 1.1933e-05 0.13033 0.96005 0.92003 0.0013954 0.99999 0.61308 0.096677 0.43001 1.9203 1.92 16 145 0.00015796 -85.666 0.90062
0.00070993 0.98801 5.5256e-05 3.8182 0.01205 9.3618e-09 0.001154 0.02517 0.0006446 0.02581 0.022521 0 0.047051 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.9894 0.99008 2.9811e-06 1.1922e-05 0.13035 0.96005 0.92003 0.0013954 0.99999 0.6131 0.087744 0.43001 1.9203 1.9201 16 145 0.00015796 -85.6665 0.90071
0.00079498 0.98801 5.5256e-05 3.8182 0.01205 1.0483e-08 0.001154 0.025184 0.0006446 0.025824 0.022534 0 0.04705 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013828 0.98933 0.99009 2.9818e-06 1.1921e-05 0.13037 0.96006 0.92004 0.0013953 0.99999 0.61311 0.079653 0.43001 1.9203 1.9201 16 145 0.00015795 -85.667 0.90079
0.00088003 0.98801 5.5256e-05 3.8182 0.01205 1.1605e-08 0.001154 0.025199 0.0006446 0.025839 0.022547 0 0.047048 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013827 0.98927 0.9901 2.9812e-06 1.1925e-05 0.13038 0.96006 0.92004 0.0013952 0.99998 0.61312 0.072324 0.43001 1.9203 1.9201 16 145 0.00015795 -85.6674 0.90088
0.00096508 0.98801 5.5256e-05 3.8182 0.01205 1.2727e-08 0.001154 0.025213 0.0006446 0.025853 0.022559 0 0.047047 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013826 0.98921 0.99011 2.9805e-06 1.1925e-05 0.13039 0.96007 0.92004 0.0013952 0.99998 0.61313 0.065686 0.43001 1.9204 1.9201 16 145 0.00015794 -85.6678 0.90097
0.0010501 0.98801 5.5256e-05 3.8182 0.01205 1.3848e-08 0.001154 0.025227 0.0006446 0.025867 0.022572 0 0.047045 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013826 0.98915 0.99012 2.9806e-06 1.1924e-05 0.1304 0.96008 0.92005 0.0013952 0.99998 0.61314 0.059672 0.43001 1.9204 1.9201 16 145 0.00015794 -85.6681 0.90105
0.0011352 0.98801 5.5256e-05 3.8182 0.01205 1.497e-08 0.001154 0.025242 0.00064461 0.025882 0.022585 0 0.047044 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013825 0.98909 0.99013 2.9808e-06 1.1922e-05 0.13041 0.96008 0.92005 0.0013951 0.99998 0.61315 0.054226 0.43001 1.9204 1.9201 16 145 0.00015793 -85.6684 0.90114
0.0012202 0.98801 5.5256e-05 3.8182 0.01205 1.6091e-08 0.001154 0.025256 0.00064461 0.025896 0.022598 0 0.047042 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98904 0.99014 2.9805e-06 1.1921e-05 0.13041 0.96009 0.92006 0.0013951 0.99998 0.61316 0.049292 0.43001 1.9205 1.9202 16 145 0.00015793 -85.6686 0.90122
0.0013053 0.98801 5.5256e-05 3.8182 0.01205 1.7213e-08 0.001154 0.02527 0.00064461 0.02591 0.022611 0 0.047041 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98898 0.99015 2.9801e-06 1.1921e-05 0.13042 0.9601 0.92006 0.001395 0.99998 0.61318 0.044823 0.43002 1.9205 1.9202 16 145 0.00015792 -85.6688 0.90131
0.0013903 0.98801 5.5256e-05 3.8182 0.01205 1.8335e-08 0.001154 0.025285 0.00064461 0.025925 0.022624 0 0.047039 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013823 0.98893 0.99016 2.9801e-06 1.1921e-05 0.13042 0.9601 0.92006 0.001395 0.99997 0.61319 0.040776 0.43002 1.9205 1.9202 16 145 0.00015792 -85.669 0.90139
0.0014754 0.98801 5.5256e-05 3.8182 0.01205 1.9456e-08 0.001154 0.025299 0.00064461 0.025939 0.022637 0 0.047038 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013823 0.98888 0.99017 2.9802e-06 1.192e-05 0.13042 0.96011 0.92007 0.001395 0.99997 0.6132 0.03711 0.43002 1.9206 1.9202 16 145 0.00015791 -85.6692 0.90148
0.0015604 0.98801 5.5256e-05 3.8182 0.01205 2.0578e-08 0.001154 0.025313 0.00064461 0.025953 0.02265 0 0.047037 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98883 0.99017 2.98e-06 1.192e-05 0.13043 0.96011 0.92007 0.001395 0.99997 0.61321 0.033789 0.43002 1.9206 1.9202 16 145 0.00015791 -85.6694 0.90156
0.0016455 0.98801 5.5256e-05 3.8182 0.01205 2.1699e-08 0.001154 0.025328 0.00064461 0.025968 0.022663 0 0.047035 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98878 0.99018 2.9798e-06 1.192e-05 0.13043 0.96012 0.92008 0.001395 0.99997 0.61322 0.030781 0.43002 1.9206 1.9203 15.9999 145 0.0001579 -85.6695 0.90165
0.0018156 0.98801 5.5256e-05 3.8182 0.01205 2.3942e-08 0.001154 0.025356 0.00064461 0.025996 0.022689 0 0.047032 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98869 0.9902 2.9795e-06 1.1919e-05 0.13043 0.96013 0.92008 0.0013949 0.99997 0.61324 0.025589 0.43002 1.9207 1.9203 15.9999 145 0.00015789 -85.6697 0.90182
0.0019663 0.98801 5.5256e-05 3.8182 0.01205 2.5929e-08 0.001154 0.025382 0.00064461 0.026022 0.022711 0 0.04703 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98861 0.99022 2.9796e-06 1.1919e-05 0.13043 0.96014 0.92009 0.0013949 0.99996 0.61326 0.021774 0.43002 1.9207 1.9203 15.9999 145 0.00015788 -85.6698 0.90197
0.0021169 0.98801 5.5256e-05 3.8182 0.01205 2.7916e-08 0.001154 0.025407 0.00064461 0.026047 0.022734 0 0.047027 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98854 0.99023 2.9797e-06 1.1919e-05 0.13044 0.96016 0.9201 0.0013949 0.99996 0.61329 0.018574 0.43003 1.9208 1.9204 15.9999 145 0.00015787 -85.6699 0.90212
0.0022676 0.98801 5.5256e-05 3.8182 0.01205 2.9902e-08 0.001154 0.025432 0.00064461 0.026072 0.022757 0 0.047025 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98846 0.99025 2.9797e-06 1.1918e-05 0.13044 0.96017 0.9201 0.0013949 0.99996 0.61331 0.015889 0.43003 1.9208 1.9204 15.9999 145 0.00015786 -85.67 0.90227
0.0024182 0.98801 5.5256e-05 3.8182 0.01205 3.1889e-08 0.001154 0.025458 0.00064462 0.026098 0.02278 0 0.047022 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.9884 0.99026 2.9796e-06 1.1918e-05 0.13044 0.96018 0.92011 0.0013949 0.99996 0.61333 0.013636 0.43003 1.9209 1.9205 15.9999 145 0.00015786 -85.67 0.90242
0.0025689 0.98801 5.5256e-05 3.8182 0.01205 3.3876e-08 0.001154 0.025483 0.00064462 0.026123 0.022803 0 0.04702 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98833 0.99028 2.9796e-06 1.1918e-05 0.13044 0.96019 0.92012 0.0013949 0.99995 0.61335 0.011745 0.43003 1.9209 1.9205 15.9999 145.0001 0.00015785 -85.6701 0.90257
0.0027195 0.98801 5.5256e-05 3.8182 0.01205 3.5862e-08 0.001154 0.025509 0.00064462 0.026149 0.022826 0 0.047017 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98827 0.99029 2.9796e-06 1.1918e-05 0.13044 0.9602 0.92012 0.0013949 0.99995 0.61337 0.010158 0.43003 1.921 1.9206 15.9999 145.0001 0.00015784 -85.6701 0.90272
0.0028702 0.98801 5.5256e-05 3.8182 0.01205 3.7849e-08 0.001154 0.025534 0.00064462 0.026174 0.022848 0 0.047014 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98821 0.99031 2.9796e-06 1.1918e-05 0.13044 0.96021 0.92013 0.0013949 0.99995 0.61339 0.0088266 0.43004 1.9211 1.9206 15.9999 145.0001 0.00015783 -85.6701 0.90287
0.0030208 0.98801 5.5256e-05 3.8182 0.01205 3.9836e-08 0.001154 0.025559 0.00064462 0.026199 0.022871 0 0.047012 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98815 0.99032 2.9796e-06 1.1918e-05 0.13044 0.96022 0.92014 0.0013949 0.99994 0.61341 0.0077093 0.43004 1.9211 1.9206 15.9999 145.0001 0.00015782 -85.67 0.90302
0.0031715 0.98801 5.5256e-05 3.8182 0.01205 4.1822e-08 0.001154 0.025585 0.00064462 0.026225 0.022894 0 0.047009 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.9881 0.99034 2.9796e-06 1.1918e-05 0.13044 0.96023 0.92014 0.0013949 0.99994 0.61343 0.0067716 0.43004 1.9212 1.9207 15.9999 145.0001 0.00015781 -85.67 0.90317
0.0033221 0.98801 5.5256e-05 3.8182 0.01205 4.3809e-08 0.001154 0.02561 0.00064463 0.02625 0.022917 0 0.047007 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98805 0.99035 2.9796e-06 1.1918e-05 0.13044 0.96024 0.92015 0.0013949 0.99994 0.61345 0.0059847 0.43004 1.9212 1.9207 15.9999 145.0001 0.0001578 -85.67 0.90332
0.0034728 0.98801 5.5256e-05 3.8182 0.01205 4.5796e-08 0.001154 0.025635 0.00064463 0.026275 0.02294 0 0.047004 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.988 0.99036 2.9797e-06 1.1919e-05 0.13044 0.96025 0.92016 0.0013949 0.99994 0.61347 0.0053243 0.43004 1.9213 1.9208 15.9999 145.0001 0.00015779 -85.6699 0.90347
0.0036234 0.98801 5.5256e-05 3.8182 0.01205 4.7782e-08 0.001154 0.025661 0.00064463 0.026301 0.022963 0 0.047002 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98795 0.99038 2.9797e-06 1.1919e-05 0.13044 0.96027 0.92016 0.0013949 0.99993 0.61349 0.0047703 0.43004 1.9213 1.9208 15.9999 145.0001 0.00015778 -85.6699 0.90362
0.0037741 0.98801 5.5256e-05 3.8182 0.01205 4.9769e-08 0.001154 0.025686 0.00064463 0.026326 0.022985 0 0.046999 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98791 0.99039 2.9797e-06 1.1919e-05 0.13044 0.96028 0.92017 0.0013949 0.99993 0.61351 0.0043053 0.43005 1.9214 1.9209 15.9999 145.0001 0.00015778 -85.6698 0.90377
0.0039247 0.98801 5.5256e-05 3.8182 0.01205 5.1756e-08 0.001154 0.025711 0.00064463 0.026352 0.023008 0 0.046997 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98787 0.99041 2.9797e-06 1.1919e-05 0.13044 0.96029 0.92018 0.0013949 0.99993 0.61353 0.0039151 0.43005 1.9214 1.9209 15.9999 145.0001 0.00015777 -85.6698 0.90392
0.0040754 0.98801 5.5256e-05 3.8182 0.01205 5.3742e-08 0.001154 0.025737 0.00064464 0.026377 0.023031 0 0.046994 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98783 0.99042 2.9798e-06 1.1919e-05 0.13044 0.9603 0.92019 0.0013949 0.99993 0.61355 0.0035877 0.43005 1.9215 1.921 15.9999 145.0001 0.00015776 -85.6697 0.90408
0.004226 0.98801 5.5256e-05 3.8182 0.01205 5.5729e-08 0.001154 0.025762 0.00064464 0.026402 0.023054 0 0.046992 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98779 0.99043 2.9798e-06 1.1919e-05 0.13044 0.96031 0.92019 0.0013949 0.99992 0.61357 0.0033129 0.43005 1.9215 1.921 15.9999 145.0001 0.00015775 -85.6696 0.90423
0.0043767 0.98801 5.5256e-05 3.8182 0.01205 5.7715e-08 0.001154 0.025788 0.00064464 0.026428 0.023077 0 0.046989 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98775 0.99045 2.9798e-06 1.1919e-05 0.13044 0.96032 0.9202 0.0013949 0.99992 0.61359 0.0030824 0.43005 1.9216 1.9211 15.9999 145.0001 0.00015774 -85.6696 0.90438
0.0045273 0.98801 5.5256e-05 3.8182 0.01205 5.9702e-08 0.001154 0.025813 0.00064464 0.026453 0.023099 0 0.046987 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98772 0.99046 2.9799e-06 1.1919e-05 0.13044 0.96033 0.92021 0.0013949 0.99992 0.61361 0.0028889 0.43006 1.9216 1.9211 15.9999 145.0001 0.00015773 -85.6695 0.90453
0.004678 0.98801 5.5256e-05 3.8182 0.01205 6.1689e-08 0.001154 0.025838 0.00064465 0.026478 0.023122 0 0.046984 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013823 0.98768 0.99047 2.9799e-06 1.1919e-05 0.13044 0.96034 0.92021 0.0013949 0.99991 0.61363 0.0027265 0.43006 1.9217 1.9212 15.9999 145.0001 0.00015772 -85.6694 0.90468
0.0048286 0.98801 5.5256e-05 3.8182 0.01205 6.3675e-08 0.001154 0.025864 0.00064465 0.026504 0.023145 0 0.046982 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013821 0.98765 0.99049 2.9799e-06 1.192e-05 0.13044 0.96035 0.92022 0.0013949 0.99991 0.61365 0.0025903 0.43006 1.9217 1.9212 15.9998 145.0001 0.00015771 -85.6694 0.90483
0.0049793 0.98801 5.5256e-05 3.8182 0.01205 6.5662e-08 0.001154 0.025889 0.00064465 0.026529 0.023168 0 0.046979 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98762 0.9905 2.98e-06 1.192e-05 0.13044 0.96036 0.92023 0.001395 0.99991 0.61367 0.002476 0.43006 1.9218 1.9213 15.9998 145.0001 0.0001577 -85.6693 0.90498
0.0051299 0.98801 5.5256e-05 3.8182 0.01205 6.7649e-08 0.001154 0.025914 0.00064465 0.026554 0.023191 0 0.046976 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.001382 0.98759 0.99051 2.98e-06 1.192e-05 0.13044 0.96038 0.92023 0.001395 0.99991 0.61369 0.00238 0.43006 1.9218 1.9213 15.9998 145.0001 0.0001577 -85.6692 0.90513
0.0052806 0.98801 5.5256e-05 3.8182 0.01205 6.9635e-08 0.001154 0.02594 0.00064466 0.02658 0.023213 0 0.046974 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013822 0.98756 0.99052 2.98e-06 1.192e-05 0.13044 0.96039 0.92024 0.001395 0.9999 0.61371 0.0022996 0.43006 1.9219 1.9214 15.9998 145.0001 0.00015769 -85.6692 0.90528
0.0054312 0.98801 5.5256e-05 3.8182 0.01205 7.1622e-08 0.001154 0.025965 0.00064466 0.026605 0.023236 0 0.046971 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.001382 0.98754 0.99054 2.9801e-06 1.192e-05 0.13044 0.9604 0.92025 0.001395 0.9999 0.61373 0.002232 0.43007 1.9219 1.9214 15.9998 145.0001 0.00015768 -85.6691 0.90543
0.0055819 0.98801 5.5256e-05 3.8182 0.01205 7.3608e-08 0.001154 0.02599 0.00064466 0.02663 0.023259 0 0.046969 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013825 0.98751 0.99055 2.9801e-06 1.192e-05 0.13044 0.96041 0.92025 0.001395 0.9999 0.61375 0.0021753 0.43007 1.922 1.9215 15.9998 145.0001 0.00015767 -85.6691 0.90558
0.0057325 0.98801 5.5256e-05 3.8182 0.01205 7.5595e-08 0.001154 0.026015 0.00064467 0.026656 0.023282 0 0.046966 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.001382 0.98749 0.99056 2.9801e-06 1.192e-05 0.13044 0.96042 0.92026 0.001395 0.9999 0.61377 0.0021277 0.43007 1.922 1.9215 15.9998 145.0001 0.00015766 -85.669 0.90573
0.0058832 0.98801 5.5256e-05 3.8182 0.01205 7.7582e-08 0.001154 0.026041 0.00064467 0.026681 0.023305 0 0.046964 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013828 0.98747 0.99057 2.9802e-06 1.1921e-05 0.13044 0.96043 0.92027 0.001395 0.99989 0.61379 0.0020877 0.43007 1.9221 1.9216 15.9998 145.0001 0.00015765 -85.6689 0.90588
0.0060338 0.98801 5.5256e-05 3.8182 0.01205 7.9568e-08 0.001154 0.026066 0.00064467 0.026706 0.023327 0 0.046961 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98744 0.99058 2.9802e-06 1.1921e-05 0.13044 0.96044 0.92027 0.001395 0.99989 0.61381 0.002054 0.43007 1.9221 1.9216 15.9998 145.0001 0.00015764 -85.6689 0.90603
0.0061845 0.98801 5.5256e-05 3.8182 0.01205 8.1555e-08 0.001154 0.026091 0.00064468 0.026731 0.02335 0 0.046959 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98742 0.9906 2.9802e-06 1.1921e-05 0.13044 0.96045 0.92028 0.001395 0.99989 0.61383 0.0020257 0.43008 1.9222 1.9217 15.9998 145.0001 0.00015763 -85.6688 0.90618
0.0063351 0.98801 5.5256e-05 3.8182 0.01205 8.3542e-08 0.001154 0.026117 0.00064468 0.026757 0.023373 0 0.046956 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.9874 0.99061 2.9803e-06 1.1921e-05 0.13044 0.96046 0.92029 0.001395 0.99988 0.61385 0.0020019 0.43008 1.9222 1.9217 15.9998 145.0001 0.00015763 -85.6688 0.90634
0.0066364 0.98801 5.5256e-05 3.8182 0.01205 8.7515e-08 0.001154 0.026167 0.00064469 0.026807 0.023419 0 0.046951 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98737 0.99063 2.9803e-06 1.1921e-05 0.13044 0.96048 0.9203 0.001395 0.99988 0.61389 0.0019647 0.43008 1.9223 1.9218 15.9998 145.0001 0.00015761 -85.6686 0.90664
0.0069377 0.98801 5.5256e-05 3.8182 0.01205 9.1488e-08 0.001154 0.026218 0.00064469 0.026858 0.023464 0 0.046946 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013824 0.98733 0.99065 2.9804e-06 1.1921e-05 0.13044 0.96051 0.92031 0.001395 0.99987 0.61393 0.0019385 0.43008 1.9224 1.9219 15.9998 145.0001 0.00015759 -85.6685 0.90694
0.007239 0.98801 5.5256e-05 3.8182 0.01205 9.5461e-08 0.001154 0.026268 0.0006447 0.026909 0.02351 0 0.046941 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013825 0.9873 0.99067 2.9804e-06 1.1922e-05 0.13044 0.96053 0.92033 0.0013951 0.99987 0.61397 0.0019202 0.43009 1.9225 1.922 15.9998 145.0001 0.00015757 -85.6684 0.90724
0.0075403 0.98801 5.5256e-05 3.8182 0.01205 9.9435e-08 0.001154 0.026319 0.00064471 0.026959 0.023555 0 0.046936 0.0389 0 0.8453 0.22699 0.05879 0.0083355 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013825 0.98727 0.9907 2.9805e-06 1.1922e-05 0.13044 0.96055 0.92034 0.0013951 0.99986 0.61401 0.0019076 0.43009 1.9226 1.9221 15.9998 145.0002 0.00015755 -85.6683 0.90754
0.0081429 0.98801 5.5256e-05 3.8182 0.01205 1.0738e-07 0.001154 0.02642 0.00064472 0.02706 0.023646 0 0.046926 0.0389 0 0.8453 0.22699 0.058791 0.0083355 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013825 0.98722 0.99074 2.9806e-06 1.1922e-05 0.13044 0.96059 0.92037 0.0013951 0.99985 0.6141 0.0018938 0.4301 1.9228 1.9223 15.9997 145.0002 0.00015752 -85.6682 0.90814
0.0087456 0.98801 5.5256e-05 3.8182 0.01205 1.1533e-07 0.001154 0.026521 0.00064474 0.027161 0.023737 0 0.046916 0.0389 0 0.8453 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013826 0.98718 0.99078 2.9807e-06 1.1923e-05 0.13044 0.96064 0.92039 0.0013951 0.99984 0.61418 0.0018874 0.43011 1.923 1.9225 15.9997 145.0002 0.00015748 -85.668 0.90875
0.0093482 0.98801 5.5256e-05 3.8182 0.01205 1.2327e-07 0.001154 0.026622 0.00064475 0.027262 0.023828 0 0.046906 0.0389 0 0.84531 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013826 0.98715 0.99082 2.9808e-06 1.1923e-05 0.13044 0.96068 0.92042 0.0013951 0.99983 0.61426 0.0018834 0.43011 1.9232 1.9227 15.9997 145.0002 0.00015745 -85.6678 0.90935
0.0099508 0.98801 5.5255e-05 3.8182 0.01205 1.3122e-07 0.001154 0.026723 0.00064477 0.027363 0.023919 0 0.046896 0.0389 0 0.84531 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013826 0.98712 0.99085 2.9808e-06 1.1923e-05 0.13044 0.96072 0.92045 0.0013952 0.99982 0.61434 0.0018806 0.43012 1.9234 1.9229 15.9997 145.0002 0.00015741 -85.6677 0.90995
0.010951 0.98801 5.5255e-05 3.8182 0.01205 1.4441e-07 0.001154 0.026891 0.0006448 0.027531 0.02407 0 0.046879 0.0389 0 0.84531 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013827 0.98709 0.99091 2.9809e-06 1.1924e-05 0.13044 0.96079 0.92049 0.0013952 0.9998 0.61447 0.0018792 0.43013 1.9237 1.9233 15.9996 145.0002 0.00015736 -85.6675 0.91095
0.011951 0.98801 5.5255e-05 3.8182 0.01205 1.5759e-07 0.001154 0.027058 0.00064484 0.027698 0.02422 0 0.046862 0.0389 0 0.84531 0.227 0.058791 0.0083356 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013827 0.98706 0.99097 2.981e-06 1.1924e-05 0.13044 0.96086 0.92053 0.0013952 0.99979 0.61461 0.0018792 0.43015 1.9241 1.9236 15.9996 145.0002 0.0001573 -85.6673 0.91195
0.012951 0.98801 5.5255e-05 3.8182 0.01205 1.7078e-07 0.001154 0.027225 0.00064487 0.027865 0.024371 0 0.046846 0.0389 0 0.84531 0.227 0.058792 0.0083356 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013828 0.98704 0.99102 2.9811e-06 1.1924e-05 0.13044 0.96094 0.92058 0.0013952 0.99977 0.61474 0.0018795 0.43016 1.9244 1.9239 15.9996 145.0003 0.00015724 -85.6671 0.91295
0.013951 0.98801 5.5255e-05 3.8182 0.01205 1.8397e-07 0.001154 0.027392 0.00064491 0.028032 0.024521 0 0.046829 0.0389 0 0.84531 0.227 0.058792 0.0083356 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013828 0.98703 0.99106 2.9812e-06 1.1925e-05 0.13044 0.96101 0.92062 0.0013952 0.99975 0.61487 0.0018797 0.43017 1.9247 1.9242 15.9996 145.0003 0.00015718 -85.667 0.91395
0.014951 0.98801 5.5255e-05 3.8182 0.01205 1.9715e-07 0.001154 0.027559 0.00064495 0.028199 0.024671 0 0.046813 0.0389 0 0.84531 0.227 0.058792 0.0083357 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013828 0.98702 0.99111 2.9812e-06 1.1925e-05 0.13044 0.96108 0.92066 0.0013953 0.99974 0.61501 0.0018798 0.43018 1.9251 1.9246 15.9995 145.0003 0.00015713 -85.6669 0.91495
0.015951 0.98801 5.5255e-05 3.8182 0.01205 2.1034e-07 0.001154 0.027726 0.00064499 0.028366 0.024822 0 0.046796 0.0389 0 0.84532 0.227 0.058792 0.0083357 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013828 0.98701 0.99115 2.9813e-06 1.1925e-05 0.13044 0.96115 0.92071 0.0013953 0.99972 0.61514 0.0018798 0.43019 1.9254 1.9249 15.9995 145.0003 0.00015707 -85.6668 0.91595
0.016951 0.98801 5.5255e-05 3.8182 0.01205 2.2353e-07 0.001154 0.027892 0.00064504 0.028533 0.024972 0 0.04678 0.0389 0 0.84532 0.227 0.058793 0.0083358 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.987 0.99119 2.9813e-06 1.1925e-05 0.13044 0.96122 0.92075 0.0013953 0.9997 0.61528 0.0018798 0.43021 1.9257 1.9252 15.9995 145.0003 0.00015701 -85.6667 0.91695
0.017951 0.98801 5.5255e-05 3.8182 0.01205 2.3671e-07 0.001154 0.028059 0.00064508 0.028699 0.025122 0 0.046763 0.0389 0 0.84532 0.227 0.058793 0.0083358 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.987 0.99122 2.9814e-06 1.1925e-05 0.13044 0.96129 0.92079 0.0013953 0.99969 0.61541 0.0018798 0.43022 1.926 1.9256 15.9994 145.0004 0.00015696 -85.6667 0.91795
0.018951 0.98801 5.5255e-05 3.8182 0.01205 2.499e-07 0.001154 0.028225 0.00064513 0.028865 0.025272 0 0.046747 0.0389 0 0.84532 0.227 0.058794 0.0083358 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.987 0.99126 2.9814e-06 1.1925e-05 0.13044 0.96136 0.92083 0.0013953 0.99967 0.61554 0.0018799 0.43023 1.9264 1.9259 15.9994 145.0004 0.0001569 -85.6666 0.91895
0.019951 0.98801 5.5255e-05 3.8182 0.01205 2.6309e-07 0.001154 0.028391 0.00064518 0.029032 0.025421 0 0.04673 0.0389 0 0.84533 0.227 0.058794 0.0083359 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99129 2.9814e-06 1.1926e-05 0.13044 0.96143 0.92088 0.0013953 0.99965 0.61568 0.0018799 0.43024 1.9267 1.9262 15.9994 145.0004 0.00015685 -85.6666 0.91995
0.020951 0.98801 5.5255e-05 3.8182 0.01205 2.7627e-07 0.001154 0.028557 0.00064523 0.029198 0.025571 0 0.046714 0.0389 0 0.84533 0.22701 0.058794 0.0083359 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99132 2.9814e-06 1.1926e-05 0.13044 0.96149 0.92092 0.0013953 0.99964 0.61581 0.0018799 0.43025 1.927 1.9265 15.9993 145.0004 0.00015679 -85.6666 0.92095
0.021951 0.98801 5.5255e-05 3.8182 0.01205 2.8946e-07 0.001154 0.028723 0.00064528 0.029364 0.02572 0 0.046697 0.0389 0 0.84533 0.22701 0.058795 0.008336 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99134 2.9814e-06 1.1926e-05 0.13044 0.96156 0.92096 0.0013953 0.99962 0.61595 0.0018799 0.43027 1.9273 1.9269 15.9993 145.0005 0.00015673 -85.6666 0.92195
0.022951 0.98801 5.5255e-05 3.8182 0.01205 3.0264e-07 0.001154 0.028889 0.00064533 0.02953 0.02587 0 0.046681 0.0389 0 0.84533 0.22701 0.058795 0.0083361 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99137 2.9814e-06 1.1926e-05 0.13044 0.96163 0.921 0.0013953 0.9996 0.61608 0.0018799 0.43028 1.9277 1.9272 15.9993 145.0005 0.00015668 -85.6665 0.92295
0.023951 0.98801 5.5255e-05 3.8182 0.01205 3.1583e-07 0.001154 0.029055 0.00064538 0.029695 0.026019 0 0.046665 0.0389 0 0.84534 0.22701 0.058796 0.0083361 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99139 2.9814e-06 1.1926e-05 0.13044 0.9617 0.92104 0.0013953 0.99959 0.61621 0.0018799 0.43029 1.928 1.9275 15.9992 145.0005 0.00015662 -85.6665 0.92395
0.024951 0.98801 5.5255e-05 3.8182 0.01205 3.2902e-07 0.001154 0.02922 0.00064544 0.029861 0.026168 0 0.046648 0.0389 0 0.84534 0.22701 0.058796 0.0083362 4.105 0.0526 6.2734e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99142 2.9814e-06 1.1926e-05 0.13044 0.96177 0.92108 0.0013953 0.99957 0.61635 0.0018799 0.4303 1.9283 1.9278 15.9992 145.0005 0.00015657 -85.6665 0.92495
0.025951 0.98801 5.5254e-05 3.8182 0.01205 3.422e-07 0.001154 0.029386 0.00064549 0.030026 0.026317 0 0.046632 0.0389 0 0.84534 0.22701 0.058797 0.0083363 4.105 0.052601 6.2735e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99144 2.9814e-06 1.1926e-05 0.13044 0.96184 0.92112 0.0013953 0.99956 0.61648 0.0018799 0.43031 1.9286 1.9282 15.9992 145.0005 0.00015651 -85.6665 0.92595
0.026951 0.98801 5.5254e-05 3.8182 0.01205 3.5539e-07 0.001154 0.029551 0.00064555 0.030192 0.026466 0 0.046616 0.0389 0 0.84535 0.22701 0.058797 0.0083363 4.105 0.052601 6.2735e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99146 2.9814e-06 1.1926e-05 0.13044 0.9619 0.92116 0.0013953 0.99954 0.61661 0.0018799 0.43033 1.929 1.9285 15.9991 145.0006 0.00015646 -85.6665 0.92695
0.027951 0.98801 5.5254e-05 3.8182 0.01205 3.6857e-07 0.001154 0.029716 0.00064561 0.030357 0.026615 0 0.046599 0.0389 0 0.84535 0.22702 0.058798 0.0083364 4.105 0.052601 6.2735e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99147 2.9814e-06 1.1926e-05 0.13044 0.96197 0.92121 0.0013953 0.99953 0.61675 0.0018799 0.43034 1.9293 1.9288 15.9991 145.0006 0.0001564 -85.6665 0.92795
0.028951 0.98801 5.5254e-05 3.8182 0.01205 3.8176e-07 0.001154 0.029881 0.00064567 0.030522 0.026764 0 0.046583 0.0389 0 0.84535 0.22702 0.058798 0.0083365 4.105 0.052601 6.2735e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99149 2.9814e-06 1.1926e-05 0.13044 0.96204 0.92125 0.0013953 0.99951 0.61688 0.0018799 0.43035 1.9296 1.9291 15.9991 145.0006 0.00015635 -85.6666 0.92895
0.029951 0.98801 5.5254e-05 3.8182 0.01205 3.9495e-07 0.001154 0.030046 0.00064573 0.030687 0.026913 0 0.046567 0.0389 0 0.84536 0.22702 0.058799 0.0083365 4.105 0.052601 6.2735e-05 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99151 2.9814e-06 1.1926e-05 0.13044 0.96211 0.92129 0.0013953 0.9995 0.61701 0.0018799 0.43036 1.9299 1.9294 15.999 145.0006 0.00015629 -85.6666 0.92995
0.030951 0.98801 5.5254e-05 3.8182 0.01205 4.0813e-07 0.001154 0.030211 0.00064579 0.030852 0.027061 0 0.046551 0.0389 0 0.84536 0.22702 0.0588 0.0083366 4.105 0.052601 6.2735e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99152 2.9814e-06 1.1926e-05 0.13044 0.96217 0.92133 0.0013953 0.99948 0.61715 0.0018799 0.43038 1.9302 1.9298 15.999 145.0006 0.00015624 -85.6666 0.93095
0.031951 0.98801 5.5254e-05 3.8182 0.01205 4.2132e-07 0.001154 0.030375 0.00064585 0.031016 0.02721 0 0.046535 0.0389 0 0.84537 0.22702 0.0588 0.0083367 4.105 0.052601 6.2735e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99154 2.9814e-06 1.1926e-05 0.13044 0.96224 0.92137 0.0013953 0.99946 0.61728 0.0018799 0.43039 1.9306 1.9301 15.999 145.0007 0.00015619 -85.6666 0.93195
0.032951 0.98801 5.5254e-05 3.8182 0.01205 4.345e-07 0.001154 0.03054 0.00064591 0.031181 0.027358 0 0.046518 0.0389 0 0.84537 0.22702 0.058801 0.0083368 4.105 0.052601 6.2735e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99155 2.9814e-06 1.1925e-05 0.13044 0.96231 0.92141 0.0013953 0.99945 0.61741 0.0018799 0.4304 1.9309 1.9304 15.9989 145.0007 0.00015613 -85.6666 0.93295
0.033951 0.98801 5.5254e-05 3.8182 0.01205 4.4769e-07 0.001154 0.030704 0.00064597 0.031345 0.027506 0 0.046502 0.0389 0 0.84537 0.22703 0.058802 0.0083369 4.105 0.052601 6.2735e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99156 2.9814e-06 1.1925e-05 0.13044 0.96237 0.92145 0.0013953 0.99943 0.61755 0.0018799 0.43041 1.9312 1.9307 15.9989 145.0007 0.00015608 -85.6666 0.93395
0.034951 0.98801 5.5254e-05 3.8182 0.01205 4.6088e-07 0.001154 0.030868 0.00064604 0.03151 0.027654 0 0.046486 0.0389 0 0.84538 0.22703 0.058802 0.008337 4.105 0.052601 6.2736e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99157 2.9814e-06 1.1925e-05 0.13044 0.96244 0.92148 0.0013953 0.99942 0.61768 0.0018799 0.43042 1.9315 1.931 15.9989 145.0007 0.00015603 -85.6667 0.93495
0.035951 0.98801 5.5254e-05 3.8182 0.01205 4.7406e-07 0.001154 0.031032 0.0006461 0.031674 0.027802 0 0.04647 0.0389 0 0.84538 0.22703 0.058803 0.008337 4.105 0.052602 6.2736e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99158 2.9814e-06 1.1925e-05 0.13044 0.96251 0.92152 0.0013953 0.99941 0.61781 0.0018799 0.43044 1.9318 1.9314 15.9988 145.0007 0.00015597 -85.6667 0.93595
0.036951 0.98801 5.5254e-05 3.8182 0.01205 4.8725e-07 0.001154 0.031196 0.00064616 0.031838 0.02795 0 0.046454 0.0389 0 0.84539 0.22703 0.058804 0.0083371 4.105 0.052602 6.2736e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99159 2.9814e-06 1.1925e-05 0.13044 0.96257 0.92156 0.0013953 0.99939 0.61795 0.0018799 0.43045 1.9321 1.9317 15.9988 145.0008 0.00015592 -85.6667 0.93695
0.037951 0.98801 5.5254e-05 3.8182 0.012049 5.0043e-07 0.001154 0.03136 0.00064623 0.032002 0.028098 0 0.046438 0.0389 0 0.84539 0.22703 0.058805 0.0083372 4.105 0.052602 6.2736e-05 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.9916 2.9813e-06 1.1925e-05 0.13044 0.96264 0.9216 0.0013953 0.99938 0.61808 0.0018799 0.43046 1.9325 1.932 15.9988 145.0008 0.00015587 -85.6667 0.93795
0.038951 0.98801 5.5254e-05 3.8182 0.012049 5.1362e-07 0.001154 0.031524 0.00064629 0.032165 0.028246 0 0.046422 0.0389 0 0.8454 0.22704 0.058805 0.0083373 4.105 0.052602 6.2736e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99161 2.9813e-06 1.1925e-05 0.13044 0.9627 0.92164 0.0013953 0.99936 0.61821 0.0018798 0.43047 1.9328 1.9323 15.9987 145.0008 0.00015581 -85.6668 0.93895
0.039951 0.98801 5.5254e-05 3.8182 0.012049 5.268e-07 0.001154 0.031687 0.00064636 0.032329 0.028393 0 0.046406 0.0389 0 0.8454 0.22704 0.058806 0.0083374 4.105 0.052602 6.2737e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99162 2.9813e-06 1.1925e-05 0.13044 0.96277 0.92168 0.0013953 0.99935 0.61834 0.0018798 0.43048 1.9331 1.9326 15.9987 145.0008 0.00015576 -85.6668 0.93995
0.040951 0.98801 5.5254e-05 3.8182 0.012049 5.3999e-07 0.001154 0.031851 0.00064642 0.032493 0.028541 0 0.04639 0.0389 0 0.84541 0.22704 0.058807 0.0083375 4.105 0.052602 6.2737e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99163 2.9813e-06 1.1925e-05 0.13044 0.96283 0.92172 0.0013953 0.99933 0.61848 0.0018798 0.43049 1.9334 1.9329 15.9987 145.0008 0.00015571 -85.6668 0.94095
0.041951 0.98801 5.5254e-05 3.8182 0.012049 5.5317e-07 0.001154 0.032014 0.00064649 0.032656 0.028688 0 0.046374 0.0389 0 0.84541 0.22704 0.058808 0.0083376 4.105 0.052602 6.2737e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99163 2.9813e-06 1.1925e-05 0.13044 0.9629 0.92176 0.0013953 0.99932 0.61861 0.0018798 0.43051 1.9337 1.9333 15.9986 145.0009 0.00015566 -85.6668 0.94195
0.042951 0.98801 5.5253e-05 3.8182 0.012049 5.6636e-07 0.001154 0.032177 0.00064656 0.032819 0.028835 0 0.046358 0.0389 0 0.84542 0.22705 0.058809 0.0083378 4.105 0.052603 6.2737e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99164 2.9813e-06 1.1925e-05 0.13044 0.96296 0.92179 0.0013953 0.99931 0.61874 0.0018798 0.43052 1.934 1.9336 15.9986 145.0009 0.0001556 -85.6669 0.94295
0.043951 0.98801 5.5253e-05 3.8182 0.012049 5.7954e-07 0.001154 0.03234 0.00064662 0.032982 0.028982 0 0.046342 0.0389 0 0.84542 0.22705 0.05881 0.0083379 4.105 0.052603 6.2737e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99165 2.9813e-06 1.1925e-05 0.13044 0.96303 0.92183 0.0013953 0.99929 0.61888 0.0018798 0.43053 1.9343 1.9339 15.9986 145.0009 0.00015555 -85.6669 0.94395
0.044951 0.98801 5.5253e-05 3.8182 0.012049 5.9273e-07 0.001154 0.032503 0.00064669 0.033145 0.029129 0 0.046326 0.0389 0 0.84543 0.22705 0.05881 0.008338 4.1051 0.052603 6.2738e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99165 2.9812e-06 1.1925e-05 0.13044 0.96309 0.92187 0.0013952 0.99928 0.61901 0.0018798 0.43054 1.9347 1.9342 15.9985 145.0009 0.0001555 -85.6669 0.94495
0.045951 0.98801 5.5253e-05 3.8182 0.012049 6.0592e-07 0.001154 0.032666 0.00064676 0.033308 0.029276 0 0.04631 0.0389 0 0.84544 0.22705 0.058811 0.0083381 4.1051 0.052603 6.2738e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99166 2.9812e-06 1.1925e-05 0.13044 0.96315 0.92191 0.0013952 0.99926 0.61914 0.0018798 0.43055 1.935 1.9345 15.9985 145.0009 0.00015545 -85.667 0.94595
0.046951 0.98801 5.5253e-05 3.8182 0.012049 6.191e-07 0.001154 0.032829 0.00064682 0.033471 0.029423 0 0.046295 0.0389 0 0.84544 0.22706 0.058812 0.0083382 4.1051 0.052603 6.2738e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99166 2.9812e-06 1.1925e-05 0.13044 0.96322 0.92194 0.0013952 0.99925 0.61927 0.0018798 0.43057 1.9353 1.9348 15.9985 145.001 0.0001554 -85.667 0.94695
0.047951 0.98801 5.5253e-05 3.8182 0.012049 6.3229e-07 0.001154 0.032991 0.00064689 0.033633 0.02957 0 0.046279 0.0389 0 0.84545 0.22706 0.058813 0.0083383 4.1051 0.052604 6.2738e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99167 2.9812e-06 1.1925e-05 0.13044 0.96328 0.92198 0.0013952 0.99924 0.61941 0.0018798 0.43058 1.9356 1.9351 15.9984 145.001 0.00015535 -85.667 0.94795
0.048951 0.98801 5.5253e-05 3.8182 0.012049 6.4547e-07 0.001154 0.033153 0.00064696 0.033796 0.029717 0 0.046263 0.0389 0 0.84545 0.22706 0.058814 0.0083385 4.1051 0.052604 6.2739e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99167 2.9812e-06 1.1925e-05 0.13044 0.96334 0.92202 0.0013952 0.99922 0.61954 0.0018798 0.43059 1.9359 1.9354 15.9984 145.001 0.0001553 -85.667 0.94895
0.049951 0.98801 5.5253e-05 3.8182 0.012049 6.5866e-07 0.001154 0.033316 0.00064702 0.033958 0.029863 0 0.046247 0.0389 0 0.84546 0.22706 0.058815 0.0083386 4.1051 0.052604 6.2739e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99167 2.9812e-06 1.1925e-05 0.13044 0.96341 0.92206 0.0013952 0.99921 0.61967 0.0018798 0.4306 1.9362 1.9358 15.9984 145.001 0.00015525 -85.6671 0.94995
0.050951 0.98801 5.5253e-05 3.8182 0.012049 6.7184e-07 0.001154 0.033478 0.00064709 0.03412 0.030009 0 0.046232 0.0389 0 0.84547 0.22707 0.058816 0.0083387 4.1051 0.052604 6.2739e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99168 2.9812e-06 1.1925e-05 0.13044 0.96347 0.92209 0.0013952 0.9992 0.6198 0.0018798 0.43061 1.9365 1.9361 15.9983 145.001 0.0001552 -85.6671 0.95095
0.051951 0.98801 5.5253e-05 3.8182 0.012049 6.8503e-07 0.001154 0.03364 0.00064716 0.034282 0.030156 0 0.046216 0.0389 0 0.84547 0.22707 0.058817 0.0083388 4.1051 0.052605 6.274e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99168 2.9811e-06 1.1924e-05 0.13044 0.96353 0.92213 0.0013952 0.99918 0.61993 0.0018798 0.43063 1.9368 1.9364 15.9983 145.0011 0.00015514 -85.6671 0.95195
0.052951 0.98801 5.5253e-05 3.8182 0.012049 6.9821e-07 0.001154 0.033802 0.00064722 0.034444 0.030302 0 0.0462 0.0389 0 0.84548 0.22707 0.058818 0.008339 4.1051 0.052605 6.274e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99169 2.9811e-06 1.1924e-05 0.13044 0.9636 0.92217 0.0013952 0.99917 0.62007 0.0018798 0.43064 1.9371 1.9367 15.9983 145.0011 0.00015509 -85.6671 0.95295
0.053951 0.98801 5.5253e-05 3.8182 0.012049 7.114e-07 0.001154 0.033963 0.00064729 0.034606 0.030448 0 0.046184 0.0389 0 0.84549 0.22708 0.058819 0.0083391 4.1051 0.052605 6.274e-05 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99169 2.9811e-06 1.1924e-05 0.13044 0.96366 0.9222 0.0013952 0.99916 0.6202 0.0018798 0.43065 1.9374 1.937 15.9982 145.0011 0.00015504 -85.6672 0.95395
0.054951 0.98801 5.5253e-05 3.8182 0.012049 7.2458e-07 0.001154 0.034125 0.00064736 0.034768 0.030594 0 0.046169 0.0389 0 0.84549 0.22708 0.05882 0.0083393 4.1051 0.052605 6.2741e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99169 2.9811e-06 1.1924e-05 0.13044 0.96372 0.92224 0.0013952 0.99914 0.62033 0.0018798 0.43066 1.9378 1.9373 15.9982 145.0011 0.00015499 -85.6672 0.95495
0.055951 0.98801 5.5253e-05 3.8182 0.012049 7.3776e-07 0.001154 0.034287 0.00064742 0.034929 0.03074 0 0.046153 0.0389 0 0.8455 0.22708 0.058822 0.0083394 4.1051 0.052606 6.2741e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99169 2.9811e-06 1.1924e-05 0.13044 0.96378 0.92227 0.0013952 0.99913 0.62046 0.0018798 0.43067 1.9381 1.9376 15.9982 145.0011 0.00015494 -85.6672 0.95595
0.056951 0.98801 5.5253e-05 3.8182 0.012049 7.5095e-07 0.001154 0.034448 0.00064749 0.035091 0.030885 0 0.046138 0.0389 0 0.84551 0.22708 0.058823 0.0083395 4.1051 0.052606 6.2741e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.9811e-06 1.1924e-05 0.13044 0.96384 0.92231 0.0013952 0.99912 0.6206 0.0018798 0.43069 1.9384 1.9379 15.9981 145.0012 0.00015489 -85.6673 0.95695
0.057951 0.98801 5.5253e-05 3.8182 0.012049 7.6413e-07 0.001154 0.034609 0.00064755 0.035252 0.031031 0 0.046122 0.0389 0 0.84551 0.22709 0.058824 0.0083397 4.1051 0.052606 6.2742e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.9811e-06 1.1924e-05 0.13044 0.96391 0.92235 0.0013952 0.9991 0.62073 0.0018798 0.4307 1.9387 1.9382 15.9981 145.0012 0.00015485 -85.6673 0.95795
0.058951 0.98801 5.5252e-05 3.8182 0.012049 7.7732e-07 0.001154 0.03477 0.00064762 0.035413 0.031177 0 0.046106 0.0389 0 0.84552 0.22709 0.058825 0.0083398 4.1051 0.052607 6.2742e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.981e-06 1.1924e-05 0.13044 0.96397 0.92238 0.0013952 0.99909 0.62086 0.0018798 0.43071 1.939 1.9385 15.9981 145.0012 0.0001548 -85.6673 0.95895
0.059951 0.98801 5.5252e-05 3.8182 0.012049 7.905e-07 0.001154 0.034931 0.00064769 0.035574 0.031322 0 0.046091 0.0389 0 0.84553 0.22709 0.058826 0.00834 4.1051 0.052607 6.2743e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.981e-06 1.1924e-05 0.13044 0.96403 0.92242 0.0013952 0.99908 0.62099 0.0018798 0.43072 1.9393 1.9388 15.9981 145.0012 0.00015475 -85.6673 0.95995
0.060951 0.98801 5.5252e-05 3.8182 0.012049 8.0369e-07 0.001154 0.035092 0.00064775 0.035735 0.031467 0 0.046075 0.0389 0 0.84554 0.2271 0.058827 0.0083401 4.1051 0.052607 6.2743e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-06 1.1924e-05 0.13044 0.96409 0.92245 0.0013952 0.99907 0.62112 0.0018798 0.43073 1.9396 1.9391 15.998 145.0013 0.0001547 -85.6674 0.96095
0.061951 0.98801 5.5252e-05 3.8182 0.012049 8.1687e-07 0.001154 0.035253 0.00064782 0.035896 0.031612 0 0.04606 0.0389 0 0.84555 0.2271 0.058829 0.0083403 4.1051 0.052608 6.2743e-05 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-06 1.1924e-05 0.13044 0.96415 0.92249 0.0013952 0.99905 0.62126 0.0018798 0.43075 1.9399 1.9394 15.998 145.0013 0.00015465 -85.6674 0.96195
0.062951 0.98801 5.5252e-05 3.8182 0.012049 8.3006e-07 0.001154 0.035413 0.00064788 0.036057 0.031758 0 0.046044 0.0389 0 0.84555 0.2271 0.05883 0.0083405 4.1051 0.052608 6.2744e-05 0.83745 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-06 1.1924e-05 0.13044 0.96421 0.92252 0.0013952 0.99904 0.62139 0.0018797 0.43076 1.9402 1.9398 15.998 145.0013 0.0001546 -85.6674 0.96295
0.063951 0.98801 5.5252e-05 3.8182 0.012049 8.4324e-07 0.001154 0.035574 0.00064795 0.036217 0.031903 0 0.046029 0.0389 0 0.84556 0.22711 0.058831 0.0083406 4.1051 0.052608 6.2744e-05 0.83745 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-06 1.1924e-05 0.13044 0.96427 0.92256 0.0013952 0.99903 0.62152 0.0018797 0.43077 1.9405 1.9401 15.9979 145.0013 0.00015455 -85.6674 0.96395
0.064951 0.98801 5.5252e-05 3.8182 0.012049 8.5643e-07 0.001154 0.035734 0.00064801 0.036377 0.032047 0 0.046013 0.0389 0 0.84557 0.22711 0.058832 0.0083408 4.1051 0.052609 6.2745e-05 0.83745 0.0051032 0.0058411 0.0013827 0.98699 0.99171 2.981e-06 1.1924e-05 0.13044 0.96433 0.92259 0.0013952 0.99902 0.62165 0.0018797 0.43078 1.9408 1.9404 15.9979 145.0013 0.0001545 -85.6675 0.96495
0.065951 0.98801 5.5252e-05 3.8182 0.012049 8.6961e-07 0.001154 0.035894 0.00064807 0.036538 0.032192 0 0.045998 0.0389 0 0.84558 0.22712 0.058834 0.0083409 4.1051 0.052609 6.2745e-05 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99171 2.9809e-06 1.1924e-05 0.13044 0.96439 0.92263 0.0013952 0.99901 0.62178 0.0018797 0.43079 1.9411 1.9407 15.9979 145.0014 0.00015446 -85.6675 0.96595
0.066951 0.98801 5.5252e-05 3.8182 0.012049 8.8279e-07 0.001154 0.036054 0.00064814 0.036698 0.032337 0 0.045983 0.0389 0 0.84559 0.22712 0.058835 0.0083411 4.1051 0.052609 6.2746e-05 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-06 1.1924e-05 0.13044 0.96445 0.92266 0.0013952 0.99899 0.62191 0.0018797 0.4308 1.9414 1.941 15.9978 145.0014 0.00015441 -85.6675 0.96695
0.067951 0.98801 5.5252e-05 3.8182 0.012049 8.9598e-07 0.001154 0.036214 0.0006482 0.036858 0.032481 0 0.045967 0.0389 0 0.84559 0.22712 0.058836 0.0083413 4.1051 0.05261 6.2746e-05 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-06 1.1924e-05 0.13044 0.96451 0.92269 0.0013952 0.99898 0.62205 0.0018797 0.43082 1.9417 1.9413 15.9978 145.0014 0.00015436 -85.6675 0.96795
0.068951 0.98801 5.5252e-05 3.8182 0.012049 9.0916e-07 0.001154 0.036374 0.00064826 0.037018 0.032626 0 0.045952 0.0389 0 0.8456 0.22713 0.058838 0.0083415 4.1051 0.05261 6.2747e-05 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-06 1.1924e-05 0.13044 0.96457 0.92273 0.0013952 0.99897 0.62218 0.0018797 0.43083 1.942 1.9416 15.9978 145.0014 0.00015431 -85.6676 0.96895
0.069951 0.98801 5.5252e-05 3.8182 0.012049 9.2235e-07 0.001154 0.036534 0.00064833 0.037177 0.03277 0 0.045937 0.0389 0 0.84561 0.22713 0.058839 0.0083416 4.1051 0.052611 6.2747e-05 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-06 1.1923e-05 0.13044 0.96463 0.92276 0.0013952 0.99896 0.62231 0.0018797 0.43084 1.9423 1.9419 15.9977 145.0014 0.00015426 -85.6676 0.96995
0.070951 0.98801 5.5252e-05 3.8182 0.012049 9.3553e-07 0.001154 0.036693 0.00064839 0.037337 0.032914 0 0.045921 0.0389 0 0.84562 0.22713 0.058841 0.0083418 4.1051 0.052611 6.2748e-05 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-06 1.1923e-05 0.13044 0.96469 0.9228 0.0013952 0.99895 0.62244 0.0018797 0.43085 1.9426 1.9422 15.9977 145.0015 0.00015422 -85.6676 0.97095
0.071951 0.98801 5.5252e-05 3.8182 0.012049 9.4872e-07 0.001154 0.036853 0.00064845 0.037496 0.033059 0 0.045906 0.0389 0 0.84563 0.22714 0.058842 0.008342 4.1051 0.052611 6.2748e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9809e-06 1.1923e-05 0.13044 0.96475 0.92283 0.0013952 0.99894 0.62257 0.0018797 0.43086 1.9429 1.9425 15.9977 145.0015 0.00015417 -85.6676 0.97195
0.072951 0.98801 5.5252e-05 3.8182 0.012049 9.619e-07 0.001154 0.037012 0.00064851 0.037656 0.033203 0 0.045891 0.0389 0 0.84564 0.22714 0.058843 0.0083422 4.1051 0.052612 6.2749e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9809e-06 1.1923e-05 0.13044 0.96481 0.92286 0.0013952 0.99892 0.6227 0.0018797 0.43088 1.9432 1.9428 15.9976 145.0015 0.00015412 -85.6677 0.97295
0.073951 0.98801 5.5252e-05 3.8182 0.012049 9.7508e-07 0.001154 0.037171 0.00064857 0.037815 0.033347 0 0.045876 0.0389 0 0.84565 0.22715 0.058845 0.0083423 4.1051 0.052612 6.275e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-06 1.1923e-05 0.13044 0.96486 0.9229 0.0013952 0.99891 0.62283 0.0018797 0.43089 1.9435 1.9431 15.9976 145.0015 0.00015408 -85.6677 0.97395
0.074951 0.98801 5.5251e-05 3.8182 0.012049 9.8827e-07 0.001154 0.03733 0.00064863 0.037974 0.03349 0 0.04586 0.0389 0 0.84566 0.22715 0.058846 0.0083425 4.1051 0.052613 6.275e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-06 1.1923e-05 0.13044 0.96492 0.92293 0.0013952 0.9989 0.62297 0.0018797 0.4309 1.9438 1.9434 15.9976 145.0015 0.00015403 -85.6677 0.97495
0.075951 0.98801 5.5251e-05 3.8182 0.012049 1.0015e-06 0.001154 0.037489 0.00064869 0.038133 0.033634 0 0.045845 0.0389 0 0.84567 0.22715 0.058848 0.0083427 4.1051 0.052613 6.2751e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-06 1.1923e-05 0.13044 0.96498 0.92296 0.0013952 0.99889 0.6231 0.0018797 0.43091 1.9441 1.9437 15.9975 145.0016 0.00015398 -85.6677 0.97595
0.076951 0.98801 5.5251e-05 3.8182 0.012049 1.0146e-06 0.001154 0.037648 0.00064875 0.038292 0.033778 0 0.04583 0.0389 0 0.84568 0.22716 0.058849 0.0083429 4.1051 0.052614 6.2751e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-06 1.1923e-05 0.13044 0.96504 0.923 0.0013951 0.99888 0.62323 0.0018797 0.43092 1.9444 1.944 15.9975 145.0016 0.00015394 -85.6677 0.97695
0.077951 0.98801 5.5251e-05 3.8182 0.012049 1.0278e-06 0.001154 0.037806 0.00064881 0.038451 0.033921 0 0.045815 0.0389 0 0.84569 0.22716 0.058851 0.0083431 4.1051 0.052614 6.2752e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13044 0.9651 0.92303 0.0013951 0.99887 0.62336 0.0018797 0.43093 1.9447 1.9443 15.9975 145.0016 0.00015389 -85.6678 0.97795
0.078951 0.98801 5.5251e-05 3.8182 0.012049 1.041e-06 0.001154 0.037965 0.00064887 0.038609 0.034065 0 0.0458 0.0389 0 0.8457 0.22717 0.058853 0.0083433 4.1051 0.052615 6.2753e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13044 0.96515 0.92306 0.0013951 0.99886 0.62349 0.0018797 0.43095 1.945 1.9446 15.9974 145.0016 0.00015384 -85.6678 0.97895
0.079951 0.98801 5.5251e-05 3.8182 0.012049 1.0542e-06 0.001154 0.038123 0.00064893 0.038768 0.034208 0 0.045785 0.0389 0 0.84571 0.22717 0.058854 0.0083435 4.1051 0.052615 6.2753e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13044 0.96521 0.92309 0.0013951 0.99884 0.62362 0.0018797 0.43096 1.9453 1.9449 15.9974 145.0016 0.0001538 -85.6678 0.97995
0.080951 0.98801 5.5251e-05 3.8182 0.012049 1.0674e-06 0.001154 0.038282 0.00064899 0.038926 0.034351 0 0.045769 0.0389 0 0.84572 0.22718 0.058856 0.0083437 4.1051 0.052616 6.2754e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13044 0.96527 0.92313 0.0013951 0.99883 0.62375 0.0018797 0.43097 1.9456 1.9452 15.9974 145.0017 0.00015375 -85.6678 0.98095
0.081951 0.98801 5.5251e-05 3.8182 0.012049 1.0806e-06 0.001154 0.03844 0.00064904 0.039084 0.034494 0 0.045754 0.0389 0 0.84573 0.22718 0.058857 0.0083439 4.1051 0.052616 6.2755e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96533 0.92316 0.0013951 0.99882 0.62388 0.0018797 0.43098 1.9459 1.9455 15.9973 145.0017 0.0001537 -85.6679 0.98195
0.082951 0.98801 5.5251e-05 3.8182 0.012049 1.0937e-06 0.001154 0.038598 0.0006491 0.039242 0.034637 0 0.045739 0.0389 0 0.84574 0.22718 0.058859 0.0083441 4.1052 0.052617 6.2755e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96538 0.92319 0.0013951 0.99881 0.62401 0.0018797 0.43099 1.9462 1.9458 15.9973 145.0017 0.00015366 -85.6679 0.98295
0.083951 0.98801 5.5251e-05 3.8182 0.012049 1.1069e-06 0.001154 0.038756 0.00064916 0.0394 0.03478 0 0.045724 0.0389 0 0.84575 0.22719 0.058861 0.0083443 4.1052 0.052618 6.2756e-05 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96544 0.92322 0.0013951 0.9988 0.62414 0.0018797 0.431 1.9465 1.946 15.9973 145.0017 0.00015361 -85.6679 0.98395
0.084951 0.98801 5.5251e-05 3.8182 0.012049 1.1201e-06 0.001154 0.038913 0.00064921 0.039558 0.034923 0 0.045709 0.0389 0 0.84576 0.22719 0.058862 0.0083445 4.1052 0.052618 6.2757e-05 0.83744 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.9655 0.92326 0.0013951 0.99879 0.62428 0.0018797 0.43102 1.9468 1.9463 15.9972 145.0017 0.00015357 -85.6679 0.98495
0.085951 0.98801 5.5251e-05 3.8182 0.012049 1.1333e-06 0.001154 0.039071 0.00064927 0.039716 0.035065 0 0.045694 0.0389 0 0.84577 0.2272 0.058864 0.0083447 4.1052 0.052619 6.2758e-05 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96555 0.92329 0.0013951 0.99878 0.62441 0.0018797 0.43103 1.9471 1.9466 15.9972 145.0018 0.00015352 -85.6679 0.98595
0.086951 0.98801 5.5251e-05 3.8182 0.012049 1.1465e-06 0.001154 0.039229 0.00064932 0.039873 0.035208 0 0.045679 0.0389 0 0.84578 0.2272 0.058866 0.008345 4.1052 0.052619 6.2758e-05 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96561 0.92332 0.0013951 0.99877 0.62454 0.0018797 0.43104 1.9474 1.9469 15.9972 145.0018 0.00015348 -85.668 0.98695
0.087951 0.98801 5.5251e-05 3.8182 0.012049 1.1597e-06 0.001154 0.039386 0.00064938 0.040031 0.03535 0 0.045664 0.0389 0 0.84579 0.22721 0.058867 0.0083452 4.1052 0.05262 6.2759e-05 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96567 0.92335 0.0013951 0.99876 0.62467 0.0018797 0.43105 1.9477 1.9472 15.9971 145.0018 0.00015343 -85.668 0.98795
0.088951 0.98801 5.5251e-05 3.8182 0.012049 1.1728e-06 0.001154 0.039543 0.00064943 0.040188 0.035493 0 0.045649 0.0389 0 0.8458 0.22721 0.058869 0.0083454 4.1052 0.052621 6.276e-05 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96572 0.92338 0.0013951 0.99875 0.6248 0.0018797 0.43106 1.948 1.9475 15.9971 145.0018 0.00015339 -85.668 0.98895
0.089951 0.98801 5.5251e-05 3.8182 0.012049 1.186e-06 0.001154 0.0397 0.00064949 0.040345 0.035635 0 0.045635 0.0389 0 0.84581 0.22722 0.058871 0.0083456 4.1052 0.052621 6.2761e-05 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-06 1.1923e-05 0.13044 0.96578 0.92341 0.0013951 0.99874 0.62493 0.0018796 0.43107 1.9482 1.9478 15.997 145.0018 0.00015334 -85.668 0.98995
0.090951 0.98801 5.5251e-05 3.8182 0.012049 1.1992e-06 0.001154 0.039857 0.00064954 0.040502 0.035777 0 0.04562 0.0389 0 0.84582 0.22722 0.058873 0.0083458 4.1052 0.052622 6.2762e-05 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-06 1.1922e-05 0.13044 0.96583 0.92345 0.0013951 0.99873 0.62506 0.0018796 0.43109 1.9485 1.9481 15.997 145.0019 0.0001533 -85.668 0.99095
0.091951 0.98801 5.525e-05 3.8182 0.012049 1.2124e-06 0.001154 0.040014 0.00064959 0.040659 0.035919 0 0.045605 0.0389 0 0.84583 0.22723 0.058874 0.0083461 4.1052 0.052623 6.2762e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96589 0.92348 0.0013951 0.99872 0.62519 0.0018796 0.4311 1.9488 1.9484 15.997 145.0019 0.00015326 -85.6681 0.99195
0.092951 0.98801 5.525e-05 3.8182 0.012049 1.2256e-06 0.001154 0.040171 0.00064965 0.040816 0.036061 0 0.04559 0.0389 0 0.84584 0.22723 0.058876 0.0083463 4.1052 0.052623 6.2763e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96594 0.92351 0.0013951 0.99871 0.62532 0.0018796 0.43111 1.9491 1.9487 15.9969 145.0019 0.00015321 -85.6681 0.99295
0.093951 0.98801 5.525e-05 3.8182 0.012049 1.2388e-06 0.001154 0.040328 0.0006497 0.040973 0.036203 0 0.045575 0.0389 0 0.84586 0.22724 0.058878 0.0083465 4.1052 0.052624 6.2764e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.966 0.92354 0.0013951 0.9987 0.62545 0.0018796 0.43112 1.9494 1.949 15.9969 145.0019 0.00015317 -85.6681 0.99395
0.094951 0.98801 5.525e-05 3.8182 0.012049 1.2519e-06 0.001154 0.040484 0.00064975 0.041129 0.036345 0 0.04556 0.0389 0 0.84587 0.22724 0.05888 0.0083468 4.1052 0.052625 6.2765e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96605 0.92357 0.0013951 0.99869 0.62558 0.0018796 0.43113 1.9497 1.9493 15.9969 145.0019 0.00015312 -85.6681 0.99495
0.095951 0.98801 5.525e-05 3.8182 0.012049 1.2651e-06 0.001154 0.040641 0.0006498 0.041286 0.036486 0 0.045546 0.0389 0 0.84588 0.22725 0.058882 0.008347 4.1052 0.052625 6.2766e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96611 0.9236 0.0013951 0.99868 0.62571 0.0018796 0.43114 1.95 1.9496 15.9968 145.002 0.00015308 -85.6681 0.99595
0.096951 0.98801 5.525e-05 3.8182 0.012049 1.2783e-06 0.001154 0.040797 0.00064985 0.041442 0.036628 0 0.045531 0.0389 0 0.84589 0.22725 0.058884 0.0083472 4.1052 0.052626 6.2767e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96616 0.92363 0.0013951 0.99867 0.62584 0.0018796 0.43116 1.9503 1.9498 15.9968 145.002 0.00015304 -85.6682 0.99695
0.097951 0.98801 5.525e-05 3.8182 0.012049 1.2915e-06 0.001154 0.040953 0.0006499 0.041598 0.036769 0 0.045516 0.0389 0 0.8459 0.22726 0.058885 0.0083475 4.1052 0.052627 6.2768e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96622 0.92366 0.0013951 0.99866 0.62597 0.0018796 0.43117 1.9506 1.9501 15.9968 145.002 0.00015299 -85.6682 0.99795
0.098951 0.98801 5.525e-05 3.8182 0.012049 1.3047e-06 0.001154 0.041109 0.00064995 0.041754 0.03691 0 0.045501 0.0389 0 0.84592 0.22726 0.058887 0.0083477 4.1052 0.052627 6.2769e-05 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96627 0.92369 0.0013951 0.99865 0.6261 0.0018796 0.43118 1.9509 1.9504 15.9967 145.002 0.00015295 -85.6682 0.99895
0.099951 0.98801 5.525e-05 3.8182 0.012049 1.3179e-06 0.001154 0.041265 0.00065 0.04191 0.037051 0 0.045487 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96632 0.92372 0.0013951 0.99864 0.62623 0.0018796 0.43119 1.9511 1.9507 15.9967 145.0021 0.00015291 -85.6682 0.99995
0.099972 0.98801 5.525e-05 3.8182 0.012049 1.3181e-06 0.001154 0.041268 0.00065 0.041914 0.037054 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62623 0.0018796 0.43119 1.9511 1.9507 15.9967 145.0021 0.00015291 -85.6682 0.99997
0.09998 0.98801 5.525e-05 3.8182 0.012049 1.3182e-06 0.001154 0.041269 0.00065 0.041915 0.037056 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9511 1.9507 15.9967 145.0021 0.00015291 -85.6682 0.99998
0.099995 0.98801 5.525e-05 3.8182 0.012049 1.3184e-06 0.001154 0.041272 0.00065001 0.041917 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6682 0.99999
0.099997 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041272 0.00065001 0.041917 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6682 1
0.099998 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041272 0.00065001 0.041918 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6682 1
0.099998 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041272 0.00065001 0.041918 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6682 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041272 0.00065001 0.041918 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6682 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041272 0.00065001 0.041918 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6671 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041273 0.00065001 0.041918 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9806e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6641 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041273 0.00065001 0.041918 0.037059 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013828 0.98699 0.99173 2.9807e-06 1.1922e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.658 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041273 0.00065001 0.041918 0.037059 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013831 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6534 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3185e-06 0.001154 0.041273 0.00065001 0.041918 0.037059 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013838 0.98699 0.99173 2.9811e-06 1.1923e-05 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6443 1
0.1 0.98801 5.525e-05 3.8182 0.012049 1.3186e-06 0.001154 0.041273 0.00065001 0.041919 0.037059 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.001386 0.98699 0.99173 2.9823e-06 1.1926e-05 0.13044 0.96633 0.92372 0.0013952 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6261 1
0.10001 0.98801 5.525e-05 3.8182 0.012049 1.3186e-06 0.001154 0.041274 0.00065001 0.041919 0.03706 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013921 0.98699 0.99173 2.9863e-06 1.1934e-05 0.13044 0.96633 0.92372 0.0013956 0.99864 0.62624 0.0018797 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.5897 1
0.10001 0.98801 5.525e-05 3.8182 0.012049 1.3187e-06 0.001154 0.041274 0.00065001 0.04192 0.03706 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0013991 0.98699 0.99173 2.992e-06 1.1947e-05 0.13044 0.96633 0.92372 0.0013962 0.99864 0.62624 0.0018798 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.5534 1
0.10002 0.98801 5.525e-05 3.8182 0.012049 1.3187e-06 0.001154 0.041275 0.00065001 0.041921 0.037061 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.001415 0.98699 0.99173 3.0083e-06 1.1985e-05 0.13044 0.96633 0.92372 0.0013979 0.99864 0.62624 0.00188 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.4807 1
0.10003 0.98801 5.525e-05 3.8182 0.012049 1.3188e-06 0.001154 0.041277 0.00065001 0.041922 0.037062 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051033 0.0058413 0.0014317 0.98699 0.99173 3.0288e-06 1.2035e-05 0.13044 0.96633 0.92372 0.0014001 0.99864 0.62624 0.0018804 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.4081 1
0.10004 0.98801 5.525e-05 3.8182 0.012049 1.319e-06 0.001154 0.041279 0.00065001 0.041924 0.037064 0 0.045485 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.0014664 0.98698 0.99173 3.0818e-06 1.2174e-05 0.13044 0.96633 0.92372 0.0014064 0.99864 0.62624 0.0018814 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.2631 1
0.10006 0.98801 5.525e-05 3.8182 0.012049 1.3192e-06 0.001154 0.041281 0.00065001 0.041926 0.037066 0 0.045485 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.001502 0.98698 0.99173 3.1434e-06 1.2347e-05 0.13044 0.96633 0.92372 0.0014144 0.99864 0.62624 0.0018828 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.1185 1.0001
0.10007 0.98801 5.525e-05 3.8182 0.012049 1.3194e-06 0.001154 0.041283 0.00065001 0.041929 0.037068 0 0.045485 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.0015383 0.98697 0.99173 3.2116e-06 1.2548e-05 0.13044 0.96633 0.92372 0.0014237 0.99864 0.62625 0.0018845 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -84.9741 1.0001
0.1001 0.98801 5.525e-05 3.8182 0.012049 1.3198e-06 0.001154 0.041288 0.00065001 0.041933 0.037072 0 0.045484 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.0016135 0.98694 0.99173 3.3598e-06 1.3004e-05 0.13044 0.96633 0.92373 0.0014449 0.99864 0.62625 0.0018887 0.43119 1.9512 1.9508 15.9967 145.0021 0.0001529 -84.6859 1.0001
0.10013 0.98801 5.525e-05 3.8182 0.012049 1.3202e-06 0.001154 0.041292 0.00065001 0.041938 0.037076 0 0.045484 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.0016921 0.98692 0.99172 3.5234e-06 1.3537e-05 0.13044 0.96633 0.92373 0.0014697 0.99864 0.62625 0.001894 0.43119 1.9512 1.9508 15.9967 145.0021 0.0001529 -84.3986 1.0001
0.10016 0.98801 5.525e-05 3.8182 0.012049 1.3206e-06 0.001154 0.041297 0.00065001 0.041942 0.037081 0 0.045484 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.0017742 0.98688 0.99172 3.6996e-06 1.4137e-05 0.13044 0.96633 0.92373 0.0014976 0.99864 0.62626 0.0019005 0.43119 1.9512 1.9508 15.9967 145.0021 0.0001529 -84.1123 1.0002
0.10022 0.98801 5.525e-05 3.8182 0.012049 1.3213e-06 0.001154 0.041306 0.00065002 0.041951 0.037089 0 0.045483 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.0019493 0.98679 0.9917 4.0809e-06 1.5483e-05 0.13044 0.96634 0.92373 0.0015593 0.99864 0.62626 0.0019166 0.43119 1.9512 1.9508 15.9967 145.0021 0.0001529 -83.5427 1.0002
0.10027 0.98801 5.525e-05 3.8182 0.012049 1.3221e-06 0.001154 0.041315 0.00065002 0.041961 0.037097 0 0.045482 0.0389 0 0.84593 0.22727 0.05889 0.008348 4.1052 0.052628 6.277e-05 0.83743 0.0051034 0.0058413 0.00214 0.98667 0.99169 4.5011e-06 1.7009e-05 0.13044 0.96634 0.92373 0.0016275 0.99864 0.62627 0.0019365 0.43119 1.9512 1.9508 15.9967 145.0021 0.00015289 -82.9767 1.0003
0.10033 0.98801 5.525e-05 3.8182 0.012049 1.3229e-06 0.001154 0.041324 0.00065002 0.04197 0.037105 0 0.045481 0.0389 0 0.84593 0.22727 0.05889 0.0083481 4.1052 0.052629 6.277e-05 0.83743 0.0051034 0.0058413 0.0023474 0.98653 0.99166 4.9612e-06 1.8699e-05 0.13044 0.96634 0.92373 0.0017005 0.99863 0.62628 0.00196 0.43119 1.9512 1.9508 15.9967 145.0021 0.00015289 -82.4143 1.0003
0.10039 0.98801 5.525e-05 3.8182 0.012049 1.3236e-06 0.001154 0.041333 0.00065002 0.041979 0.037113 0 0.04548 0.0389 0 0.84593 0.22727 0.05889 0.0083481 4.1052 0.052629 6.277e-05 0.83743 0.0051034 0.0058413 0.002573 0.98637 0.99164 5.4643e-06 2.0552e-05 0.13044 0.96634 0.92373 0.0017773 0.99863 0.62629 0.0019866 0.43119 1.9513 1.9508 15.9967 145.0021 0.00015289 -81.8552 1.0004
0.10051 0.98801 5.525e-05 3.8182 0.012049 1.3252e-06 0.001154 0.041351 0.00065003 0.041997 0.03713 0 0.045478 0.0389 0 0.84594 0.22727 0.05889 0.0083481 4.1052 0.052629 6.277e-05 0.83743 0.0051034 0.0058413 0.0030852 0.98597 0.99157 6.6159e-06 2.4788e-05 0.13044 0.96634 0.92374 0.0019412 0.99863 0.6263 0.002048 0.43118 1.9513 1.9509 15.9967 145.0021 0.00015289 -80.7463 1.0005
0.10062 0.98801 5.525e-05 3.8182 0.012049 1.3267e-06 0.001154 0.04137 0.00065004 0.042015 0.037146 0 0.045477 0.0389 0 0.84594 0.22727 0.058891 0.0083481 4.1052 0.052629 6.277e-05 0.83743 0.0051034 0.0058413 0.0036893 0.98547 0.99147 7.9908e-06 2.9812e-05 0.13044 0.96634 0.92374 0.002117 0.99863 0.62631 0.0021188 0.43118 1.9513 1.9509 15.9967 145.0021 0.00015288 -79.6486 1.0006
0.10074 0.98801 5.525e-05 3.8182 0.012049 1.3283e-06 0.001154 0.041388 0.00065004 0.042033 0.037163 0 0.045475 0.0389 0 0.84594 0.22727 0.058891 0.0083482 4.1052 0.052629 6.277e-05 0.83743 0.0051034 0.0058413 0.0044004 0.98489 0.99136 9.6303e-06 3.576e-05 0.13044 0.96634 0.92374 0.0023046 0.99863 0.62632 0.0021973 0.43117 1.9514 1.9509 15.9967 145.0021 0.00015288 -78.5607 1.0007
0.10086 0.98801 5.525e-05 3.8182 0.012049 1.3298e-06 0.001154 0.041406 0.00065005 0.042051 0.037179 0 0.045473 0.0389 0 0.84594 0.22727 0.058891 0.0083482 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058413 0.0052366 0.98421 0.99121 1.1584e-05 4.2808e-05 0.13044 0.96634 0.92375 0.0025052 0.99862 0.62634 0.0022821 0.43116 1.9514 1.951 15.9967 145.002 0.00015288 -77.4815 1.0009
0.10097 0.98801 5.525e-05 3.8182 0.012049 1.3313e-06 0.001154 0.041424 0.00065005 0.04207 0.037196 0 0.045472 0.0389 0 0.84594 0.22727 0.058891 0.0083482 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058414 0.0062192 0.98344 0.99104 1.391e-05 5.1154e-05 0.13044 0.96633 0.92375 0.00272 0.99862 0.62635 0.0023727 0.43115 1.9514 1.951 15.9967 145.002 0.00015287 -76.4096 1.001
0.10109 0.98801 5.525e-05 3.8182 0.012049 1.3329e-06 0.001154 0.041442 0.00065006 0.042088 0.037212 0 0.04547 0.0389 0 0.84594 0.22728 0.058892 0.0083482 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058414 0.0073732 0.98257 0.99084 1.6679e-05 6.1024e-05 0.13044 0.96632 0.92375 0.0029496 0.99862 0.62636 0.0024683 0.43114 1.9515 1.951 15.9967 145.002 0.00015287 -75.3443 1.0011
0.10121 0.98801 5.525e-05 3.8182 0.012049 1.3344e-06 0.001154 0.04146 0.00065006 0.042106 0.037229 0 0.045468 0.0389 0 0.84594 0.22728 0.058892 0.0083483 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058414 0.0087252 0.98159 0.9906 1.9972e-05 7.267e-05 0.13044 0.96631 0.92376 0.003194 0.99861 0.62637 0.0025684 0.43113 1.9515 1.9511 15.9966 145.002 0.00015287 -74.2843 1.0012
0.10132 0.98801 5.525e-05 3.8182 0.012049 1.3359e-06 0.001154 0.041479 0.00065007 0.042124 0.037245 0 0.045466 0.0389 0 0.84595 0.22728 0.058892 0.0083483 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058414 0.010303 0.98051 0.99033 2.3879e-05 8.6383e-05 0.13044 0.96629 0.92376 0.0034534 0.99861 0.62638 0.0026725 0.43112 1.9515 1.9511 15.9966 145.002 0.00015287 -73.229 1.0013
0.10144 0.98801 5.525e-05 3.8182 0.012049 1.3375e-06 0.001154 0.041497 0.00065008 0.042142 0.037261 0 0.045465 0.0389 0 0.84595 0.22728 0.058892 0.0083483 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058414 0.012141 0.97931 0.99001 2.8508e-05 0.00010252 0.13044 0.96628 0.92377 0.0037288 0.9986 0.62639 0.00278 0.43111 1.9516 1.9511 15.9966 145.002 0.00015286 -72.1774 1.0014
0.10156 0.98801 5.525e-05 3.8182 0.012049 1.339e-06 0.001154 0.041515 0.00065008 0.04216 0.037278 0 0.045463 0.0389 0 0.84595 0.22728 0.058892 0.0083484 4.1052 0.052629 6.2771e-05 0.83743 0.0051034 0.0058414 0.014292 0.978 0.98964 3.4001e-05 0.0001215 0.13044 0.96625 0.92377 0.0040212 0.9986 0.62641 0.0028906 0.43109 1.9516 1.9512 15.9966 145.002 0.00015286 -71.1288 1.0016
0.10167 0.98801 5.525e-05 3.8182 0.012049 1.3406e-06 0.001154 0.041533 0.00065009 0.042178 0.037294 0 0.045461 0.0389 0 0.84595 0.22728 0.058893 0.0083484 4.1052 0.05263 6.2771e-05 0.83743 0.0051034 0.0058414 0.016799 0.97655 0.98922 4.0515e-05 0.00014382 0.13044 0.96622 0.92377 0.0043312 0.99859 0.62642 0.003004 0.43108 1.9516 1.9512 15.9966 145.002 0.00015286 -70.0824 1.0017
0.10179 0.98801 5.525e-05 3.8182 0.012049 1.3421e-06 0.001154 0.041551 0.00065009 0.042197 0.037311 0 0.04546 0.0389 0 0.84595 0.22728 0.058893 0.0083484 4.1052 0.05263 6.2771e-05 0.83743 0.0051034 0.0058414 0.01971 0.97497 0.98873 4.823e-05 0.00017002 0.13044 0.96619 0.92378 0.0046592 0.99858 0.62643 0.0031199 0.43106 1.9517 1.9512 15.9966 145.002 0.00015286 -69.0377 1.0018
0.10191 0.98801 5.525e-05 3.8182 0.012049 1.3436e-06 0.001154 0.041569 0.0006501 0.042215 0.037327 0 0.045458 0.0389 0 0.84595 0.22728 0.058893 0.0083485 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.023087 0.97324 0.98818 5.7357e-05 0.00020073 0.13044 0.96615 0.92378 0.0050054 0.99857 0.62644 0.0032381 0.43105 1.9517 1.9513 15.9966 145.002 0.00015286 -67.9939 1.0019
0.10202 0.98801 5.525e-05 3.8182 0.012049 1.3452e-06 0.001154 0.041587 0.0006501 0.042233 0.037344 0 0.045456 0.0389 0 0.84595 0.22728 0.058893 0.0083485 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.027 0.97135 0.98755 6.8148e-05 0.00023671 0.13044 0.9661 0.92378 0.0053706 0.99856 0.62645 0.0033583 0.43103 1.9517 1.9513 15.9966 145.002 0.00015286 -66.9504 1.002
0.10214 0.98801 5.525e-05 3.8182 0.012049 1.3467e-06 0.001154 0.041605 0.00065011 0.042251 0.03736 0 0.045455 0.0389 0 0.84596 0.22728 0.058894 0.0083485 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.031528 0.9693 0.98683 8.0905e-05 0.00027882 0.13044 0.96605 0.92379 0.0057551 0.99855 0.62646 0.0034804 0.43101 1.9518 1.9513 15.9966 145.002 0.00015286 -65.9065 1.0021
0.10226 0.98801 5.525e-05 3.8182 0.012049 1.3482e-06 0.001154 0.041624 0.00065012 0.042269 0.037376 0 0.045453 0.0389 0 0.84596 0.22728 0.058894 0.0083485 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.036757 0.96706 0.986 9.5982e-05 0.00032807 0.13044 0.96599 0.92379 0.0061595 0.99853 0.62647 0.0036041 0.43099 1.9518 1.9514 15.9966 145.002 0.00015286 -64.8613 1.0023
0.10237 0.98801 5.525e-05 3.8182 0.012049 1.3498e-06 0.001154 0.041642 0.00065012 0.042287 0.037393 0 0.045451 0.0389 0 0.84596 0.22728 0.058894 0.0083486 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.042786 0.96462 0.98507 0.0001138 0.00038567 0.13044 0.96592 0.92379 0.0065842 0.99851 0.62648 0.0037293 0.43097 1.9518 1.9514 15.9966 145.002 0.00015286 -63.8136 1.0024
0.10249 0.98801 5.525e-05 3.8182 0.012049 1.3513e-06 0.001154 0.04166 0.00065013 0.042305 0.037409 0 0.045449 0.0389 0 0.84596 0.22728 0.058894 0.0083486 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.049729 0.96196 0.98401 0.00013487 0.00045298 0.13044 0.96584 0.9238 0.0070297 0.99849 0.62649 0.0038559 0.43096 1.9519 1.9514 15.9965 145.002 0.00015286 -62.7619 1.0025
0.10261 0.98801 5.525e-05 3.8182 0.012049 1.3528e-06 0.001154 0.041678 0.00065013 0.042324 0.037426 0 0.045448 0.0389 0 0.84596 0.22728 0.058895 0.0083486 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.057712 0.95908 0.9828 0.00015978 0.00053164 0.13044 0.96574 0.9238 0.0074965 0.99846 0.6265 0.0039836 0.43094 1.9519 1.9515 15.9965 145.002 0.00015286 -61.7041 1.0026
0.10272 0.98801 5.525e-05 3.8182 0.012049 1.3544e-06 0.001154 0.041696 0.00065014 0.042342 0.037442 0 0.045446 0.0389 0 0.84596 0.22728 0.058895 0.0083487 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.066888 0.95593 0.98142 0.00018927 0.00062364 0.13044 0.96564 0.9238 0.0079853 0.99842 0.62651 0.0041125 0.43092 1.9519 1.9515 15.9965 145.002 0.00015286 -60.637 1.0027
0.10284 0.98801 5.525e-05 3.8182 0.012049 1.3559e-06 0.001154 0.041714 0.00065014 0.04236 0.037459 0 0.045444 0.0389 0 0.84596 0.22729 0.058895 0.0083487 4.1052 0.05263 6.2772e-05 0.83743 0.0051034 0.0058414 0.077443 0.95251 0.97986 0.00022428 0.00073138 0.13044 0.96553 0.92381 0.0084967 0.99837 0.62652 0.0042423 0.4309 1.952 1.9515 15.9965 145.002 0.00015287 -59.5558 1.0028
0.10295 0.98801 5.525e-05 3.8182 0.012049 1.3575e-06 0.001154 0.041732 0.00065015 0.042378 0.037475 0 0.045443 0.0389 0 0.84597 0.22729 0.058895 0.0083487 4.1052 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.089613 0.94878 0.97809 0.00026598 0.00085786 0.13044 0.9654 0.92381 0.0090318 0.99832 0.62653 0.0043731 0.43087 1.952 1.9516 15.9965 145.002 0.00015287 -58.4536 1.003
0.10307 0.98801 5.525e-05 3.8182 0.012049 1.359e-06 0.001154 0.04175 0.00065015 0.042396 0.037491 0 0.045441 0.0389 0 0.84597 0.22729 0.058896 0.0083487 4.1052 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.10371 0.9447 0.97607 0.00031593 0.0010069 0.13044 0.96526 0.92381 0.009592 0.99824 0.62654 0.0045048 0.43085 1.952 1.9516 15.9965 145.002 0.00015287 -57.3197 1.0031
0.10319 0.98801 5.525e-05 3.8182 0.012049 1.3605e-06 0.001154 0.041769 0.00065016 0.042414 0.037508 0 0.045439 0.0389 0 0.84597 0.22729 0.058896 0.0083488 4.1052 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.12017 0.94022 0.97377 0.00037629 0.0011838 0.13044 0.9651 0.92382 0.010179 0.99815 0.62654 0.0046374 0.43083 1.9521 1.9516 15.9965 145.002 0.00015287 -56.1377 1.0032
0.10329 0.98801 5.525e-05 3.8182 0.012049 1.3619e-06 0.001154 0.041785 0.00065017 0.04243 0.037523 0 0.045438 0.0389 0 0.84597 0.22729 0.058896 0.0083488 4.1052 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.13753 0.93579 0.97141 0.00044209 0.0013727 0.13044 0.96495 0.92382 0.010733 0.99804 0.62655 0.0047575 0.43081 1.9521 1.9517 15.9965 145.002 0.00015288 -55.0116 1.0033
0.10339 0.98801 5.525e-05 3.8182 0.012049 1.3632e-06 0.001154 0.0418 0.00065017 0.042445 0.037536 0 0.045436 0.0389 0 0.84597 0.22729 0.058896 0.0083488 4.1052 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.15582 0.93142 0.96901 0.00051347 0.0015734 0.13044 0.96479 0.92382 0.011255 0.99791 0.62656 0.0048664 0.4308 1.9521 1.9517 15.9965 145.002 0.00015288 -53.9225 1.0034
0.10346 0.98801 5.525e-05 3.8182 0.012049 1.3641e-06 0.001154 0.041811 0.00065017 0.042456 0.037546 0 0.045435 0.0389 0 0.84597 0.22729 0.058896 0.0083488 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.1721 0.92776 0.96696 0.00057858 0.0017527 0.13044 0.96467 0.92382 0.011674 0.99779 0.62656 0.0049506 0.43078 1.9521 1.9517 15.9965 145.002 0.00015288 -53.0148 1.0035
0.10353 0.98801 5.525e-05 3.8182 0.012049 1.3651e-06 0.001154 0.041822 0.00065018 0.042468 0.037556 0 0.045434 0.0389 0 0.84597 0.22729 0.058896 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.19087 0.92378 0.9647 0.00065529 0.0019595 0.13044 0.96453 0.92382 0.012109 0.99764 0.62656 0.0050354 0.43077 1.9522 1.9517 15.9965 145.002 0.00015288 -52.0209 1.0035
0.1036 0.98801 5.525e-05 3.8182 0.012049 1.3659e-06 0.001154 0.041832 0.00065018 0.042478 0.037565 0 0.045433 0.0389 0 0.84597 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.21053 0.91986 0.96244 0.00073731 0.0021758 0.13044 0.9644 0.92383 0.012518 0.99747 0.62656 0.0051122 0.43076 1.9522 1.9518 15.9965 145.002 0.00015289 -51.024 1.0036
0.10365 0.98801 5.525e-05 3.8182 0.012049 1.3666e-06 0.001154 0.041841 0.00065018 0.042486 0.037573 0 0.045432 0.0389 0 0.84597 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.22898 0.91637 0.96042 0.00081572 0.0023781 0.13044 0.96429 0.92383 0.012863 0.99731 0.62657 0.005175 0.43075 1.9522 1.9518 15.9966 145.002 0.00015289 -50.1174 1.0037
0.1037 0.98801 5.525e-05 3.8182 0.012049 1.3673e-06 0.001154 0.041849 0.00065019 0.042494 0.03758 0 0.045432 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.25032 0.91251 0.95821 0.00090817 0.0026115 0.13044 0.96417 0.92383 0.013222 0.9971 0.62657 0.0052384 0.43074 1.9522 1.9518 15.9966 145.002 0.00015289 -49.0914 1.0037
0.10375 0.98801 5.525e-05 3.8182 0.012049 1.368e-06 0.001154 0.041856 0.00065019 0.042502 0.037587 0 0.045431 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.27269 0.90862 0.95601 0.0010072 0.0028559 0.13044 0.96406 0.92383 0.013561 0.99688 0.62657 0.0052961 0.43073 1.9522 1.9518 15.9966 145.002 0.00015289 -48.0302 1.0038
0.10379 0.98801 5.525e-05 3.8182 0.012049 1.3685e-06 0.001154 0.041862 0.00065019 0.042508 0.037593 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.2935 0.90508 0.95407 0.0011016 0.0030838 0.13044 0.96397 0.92383 0.013845 0.99666 0.62657 0.0053431 0.43072 1.9522 1.9518 15.9967 145.002 0.0001529 -47.0479 1.0038
0.1038 0.98801 5.525e-05 3.8182 0.012049 1.3686e-06 0.001154 0.041864 0.00065019 0.042509 0.037594 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.2993 0.9041 0.95354 0.0011283 0.0031475 0.13044 0.96394 0.92383 0.01392 0.99659 0.62656 0.0053552 0.43072 1.9522 1.9518 15.9967 145.002 0.0001529 -46.7741 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3687e-06 0.001154 0.041865 0.00065019 0.04251 0.037595 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30314 0.90345 0.9532 0.0011461 0.0031897 0.13044 0.96393 0.92383 0.013968 0.99655 0.62656 0.005363 0.43072 1.9522 1.9518 15.9967 145.002 0.0001529 -46.593 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3687e-06 0.001154 0.041865 0.00065019 0.042511 0.037595 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.3057 0.90301 0.95297 0.001158 0.0032179 0.13044 0.96391 0.92383 0.014 0.99652 0.62656 0.0053681 0.43071 1.9522 1.9518 15.9967 145.002 0.0001529 -46.472 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042511 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30736 0.90273 0.95282 0.0011658 0.0032363 0.13044 0.96391 0.92383 0.014021 0.9965 0.62656 0.0053714 0.43071 1.9522 1.9518 15.9967 145.002 0.0001529 -46.3931 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042511 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30763 0.90269 0.9528 0.001167 0.0032392 0.13044 0.96391 0.92383 0.014024 0.9965 0.62656 0.005372 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3805 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30816 0.9026 0.95275 0.0011695 0.0032451 0.13044 0.9639 0.92383 0.014031 0.99649 0.62656 0.005373 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3552 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30826 0.90258 0.95274 0.0011699 0.0032461 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053732 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3508 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30827 0.90258 0.95274 0.00117 0.0032463 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053732 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3503 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30829 0.90257 0.95274 0.0011701 0.0032465 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053732 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3494 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30829 0.90257 0.95274 0.0011701 0.0032465 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053732 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3493 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30829 0.90257 0.95274 0.0011701 0.0032465 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053732 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3492 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30829 0.90257 0.95274 0.0011701 0.0032465 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053733 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3491 1.0038
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30829 0.90257 0.95274 0.0011701 0.0032466 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053733 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.349 1.0037
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.3083 0.90257 0.95274 0.0011701 0.0032466 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053733 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3488 1.0036
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30831 0.90257 0.95274 0.0011702 0.0032467 0.13044 0.9639 0.92383 0.014032 0.99649 0.62656 0.0053733 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3483 1.0035
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30833 0.90257 0.95273 0.0011703 0.003247 0.13044 0.9639 0.92383 0.014033 0.99649 0.62656 0.0053733 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3473 1.0031
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30837 0.90256 0.95273 0.0011705 0.0032474 0.13044 0.9639 0.92383 0.014033 0.99649 0.62656 0.0053734 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3453 1.0025
0.10381 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30846 0.90255 0.95272 0.0011709 0.0032483 0.13044 0.9639 0.92383 0.014034 0.99649 0.62656 0.0053736 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3413 1.0012
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30862 0.90252 0.95271 0.0011716 0.0032502 0.13044 0.9639 0.92383 0.014036 0.99649 0.62656 0.0053739 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3334 0.99853
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30879 0.90249 0.95269 0.0011724 0.003252 0.13044 0.9639 0.92383 0.014038 0.99649 0.62656 0.0053742 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3255 0.99591
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30896 0.90246 0.95268 0.0011732 0.0032539 0.13044 0.9639 0.92383 0.01404 0.99648 0.62656 0.0053746 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3175 0.99329
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.3093 0.9024 0.95265 0.0011748 0.0032576 0.13044 0.9639 0.92383 0.014044 0.99648 0.62656 0.0053752 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.3016 0.98806
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30963 0.90235 0.95262 0.0011764 0.0032613 0.13044 0.9639 0.92383 0.014049 0.99648 0.62656 0.0053759 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.2856 0.98286
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041866 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.30997 0.90229 0.95259 0.0011779 0.0032651 0.13044 0.9639 0.92383 0.014053 0.99647 0.62656 0.0053765 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.2697 0.97769
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3688e-06 0.001154 0.041867 0.00065019 0.042512 0.037596 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.31065 0.90217 0.95253 0.0011811 0.0032725 0.13044 0.96389 0.92383 0.014061 0.99647 0.62656 0.0053778 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.2376 0.96743
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3689e-06 0.001154 0.041867 0.00065019 0.042512 0.037597 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.31201 0.90194 0.95241 0.0011875 0.0032876 0.13044 0.96389 0.92383 0.014077 0.99645 0.62656 0.0053805 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.1731 0.94722
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3689e-06 0.001154 0.041867 0.00065019 0.042513 0.037597 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.31338 0.90171 0.95229 0.001194 0.0033028 0.13044 0.96388 0.92383 0.014094 0.99643 0.62656 0.0053831 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.108 0.92744
0.10382 0.98801 5.525e-05 3.8182 0.012049 1.3689e-06 0.001154 0.041868 0.00065019 0.042513 0.037597 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.31477 0.90147 0.95217 0.0012005 0.0033181 0.13044 0.96388 0.92383 0.014111 0.99642 0.62656 0.0053857 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -46.0423 0.90807
0.10383 0.98801 5.525e-05 3.8182 0.012049 1.3689e-06 0.001154 0.041868 0.00065019 0.042513 0.037598 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.31616 0.90123 0.95205 0.0012071 0.0033336 0.13044 0.96387 0.92383 0.014127 0.9964 0.62656 0.0053884 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -45.9761 0.8891
0.10383 0.98801 5.525e-05 3.8182 0.012049 1.369e-06 0.001154 0.041868 0.00065019 0.042514 0.037598 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.31899 0.90075 0.9518 0.0012205 0.0033649 0.13044 0.96386 0.92383 0.014161 0.99637 0.62656 0.0053936 0.43071 1.9523 1.9518 15.9967 145.002 0.0001529 -45.8418 0.85236
0.10384 0.98801 5.525e-05 3.8182 0.012049 1.3691e-06 0.001154 0.041869 0.00065019 0.042515 0.037599 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2773e-05 0.83743 0.0051034 0.0058414 0.32187 0.90026 0.95155 0.0012342 0.0033968 0.13044 0.96385 0.92383 0.014194 0.99634 0.62656 0.0053989 0.43071 1.9523 1.9518 15.9968 145.002 0.0001529 -45.7052 0.81713
0.10384 0.98801 5.525e-05 3.8182 0.012049 1.3691e-06 0.001154 0.04187 0.00065019 0.042515 0.037599 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.32479 0.89975 0.9513 0.0012481 0.0034293 0.13044 0.96384 0.92383 0.014228 0.9963 0.62656 0.0054042 0.43071 1.9523 1.9518 15.9968 145.002 0.0001529 -45.566 0.78336
0.10384 0.98801 5.525e-05 3.8182 0.012049 1.3692e-06 0.001154 0.041871 0.00065019 0.042516 0.0376 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.32857 0.8991 0.95098 0.0012662 0.0034714 0.13044 0.96382 0.92383 0.014271 0.99626 0.62656 0.0054109 0.43071 1.9523 1.9518 15.9968 145.002 0.0001529 -45.386 0.74257
0.10385 0.98801 5.525e-05 3.8182 0.012049 1.3693e-06 0.001154 0.041871 0.00065019 0.042517 0.037601 0 0.04543 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.33242 0.89843 0.95065 0.0012848 0.0035146 0.13044 0.96381 0.92383 0.014315 0.99621 0.62656 0.0054177 0.43071 1.9523 1.9518 15.9968 145.002 0.0001529 -45.2017 0.7039
0.10386 0.98801 5.525e-05 3.8182 0.012049 1.3693e-06 0.001154 0.041872 0.00065019 0.042518 0.037602 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.33637 0.89773 0.95032 0.001304 0.0035588 0.13044 0.96379 0.92383 0.014359 0.99617 0.62656 0.0054245 0.43071 1.9523 1.9518 15.9968 145.002 0.0001529 -45.0129 0.66724
0.10386 0.98801 5.525e-05 3.8182 0.012049 1.3694e-06 0.001154 0.041873 0.00065019 0.042519 0.037602 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.3404 0.89702 0.94998 0.0013237 0.0036041 0.13044 0.96378 0.92383 0.014403 0.99612 0.62656 0.0054313 0.4307 1.9523 1.9518 15.9968 145.002 0.0001529 -44.8195 0.63249
0.10387 0.98801 5.525e-05 3.8182 0.012049 1.3695e-06 0.001154 0.041874 0.00065019 0.04252 0.037603 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.34452 0.89629 0.94964 0.001344 0.0036507 0.13044 0.96376 0.92383 0.014447 0.99607 0.62656 0.0054381 0.4307 1.9523 1.9518 15.9968 145.002 0.0001529 -44.6212 0.59956
0.10387 0.98801 5.525e-05 3.8182 0.012049 1.3695e-06 0.001154 0.041875 0.00065019 0.04252 0.037604 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.0083489 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.34874 0.89553 0.94929 0.0013649 0.0036984 0.13044 0.96375 0.92383 0.014492 0.99602 0.62656 0.0054449 0.4307 1.9523 1.9518 15.9968 145.002 0.0001529 -44.4178 0.56833
0.10388 0.98801 5.525e-05 3.8182 0.012049 1.3697e-06 0.001154 0.041876 0.00065019 0.042522 0.037605 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.35747 0.89392 0.94858 0.0014086 0.0037979 0.13044 0.96372 0.92383 0.014583 0.99591 0.62656 0.0054587 0.4307 1.9523 1.9518 15.9968 145.002 0.0001529 -43.995 0.51068
0.10389 0.98801 5.525e-05 3.8182 0.012049 1.3698e-06 0.001154 0.041878 0.00065019 0.042523 0.037607 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.3654 0.89243 0.94794 0.0014489 0.0038891 0.13044 0.96369 0.92383 0.014664 0.99581 0.62656 0.0054707 0.4307 1.9523 1.9518 15.9969 145.002 0.0001529 -43.6084 0.46529
0.1039 0.98801 5.525e-05 3.8182 0.012049 1.3699e-06 0.001154 0.041879 0.00065019 0.042525 0.037608 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.37281 0.89099 0.94735 0.0014871 0.0039752 0.13044 0.96366 0.92383 0.014738 0.99572 0.62656 0.0054817 0.4307 1.9523 1.9519 15.9969 145.002 0.0001529 -43.2445 0.42789
0.10391 0.98801 5.525e-05 3.8182 0.012049 1.3701e-06 0.001154 0.041881 0.00065019 0.042527 0.03761 0 0.045429 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.38366 0.88879 0.9465 0.0015441 0.0041026 0.13044 0.96363 0.92383 0.014843 0.99558 0.62656 0.0054971 0.43069 1.9523 1.9519 15.9969 145.002 0.0001529 -42.708 0.38059
0.10392 0.98801 5.525e-05 3.8182 0.012049 1.3702e-06 0.001154 0.041883 0.0006502 0.042528 0.037611 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.3951 0.88635 0.94561 0.0016056 0.0042391 0.13044 0.96359 0.92383 0.014951 0.99543 0.62655 0.0055127 0.43069 1.9523 1.9519 15.997 145.002 0.0001529 -42.1365 0.33851
0.10394 0.98801 5.525e-05 3.8182 0.012049 1.3704e-06 0.001154 0.041885 0.0006502 0.04253 0.037613 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.40717 0.88358 0.94469 0.0016722 0.0043859 0.13044 0.96355 0.92383 0.015061 0.99527 0.62655 0.0055286 0.43069 1.9523 1.9519 15.997 145.002 0.0001529 -41.5265 0.30109
0.10395 0.98801 5.525e-05 3.8182 0.012049 1.3705e-06 0.001154 0.041886 0.0006502 0.042532 0.037615 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.4199 0.88041 0.94373 0.0017446 0.0045444 0.13044 0.96351 0.92383 0.015175 0.99509 0.62655 0.0055447 0.43069 1.9523 1.9519 15.997 145.002 0.0001529 -40.8741 0.2678
0.10396 0.98801 5.525e-05 3.8182 0.012049 1.3707e-06 0.001154 0.041888 0.0006502 0.042534 0.037616 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.43335 0.87671 0.94274 0.0018237 0.0047161 0.13044 0.96347 0.92383 0.015293 0.99491 0.62655 0.0055611 0.43069 1.9523 1.9519 15.9971 145.002 0.00015291 -40.1751 0.2382
0.10396 0.98801 5.525e-05 3.8182 0.012049 1.3707e-06 0.001154 0.041889 0.0006502 0.042534 0.037616 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.43531 0.87613 0.94259 0.0018354 0.0047415 0.13044 0.96347 0.92383 0.01531 0.99489 0.62655 0.0055635 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -40.0727 0.2343
0.10396 0.98801 5.525e-05 3.8182 0.012049 1.3707e-06 0.001154 0.041889 0.0006502 0.042535 0.037617 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.43926 0.87481 0.9423 0.0018593 0.0047932 0.13044 0.96346 0.92383 0.015344 0.99483 0.62655 0.0055682 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.8647 0.2267
0.10396 0.98801 5.525e-05 3.8182 0.012049 1.3708e-06 0.001154 0.041889 0.0006502 0.042535 0.037617 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.43999 0.87454 0.94225 0.0018637 0.0048027 0.13044 0.96345 0.92383 0.01535 0.99482 0.62655 0.005569 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.8264 0.22534
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3708e-06 0.001154 0.041889 0.0006502 0.042535 0.037617 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.44145 0.87399 0.94214 0.0018727 0.004822 0.13044 0.96345 0.92383 0.015362 0.9948 0.62655 0.0055708 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.7492 0.22265
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3708e-06 0.001154 0.04189 0.0006502 0.042535 0.037617 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.44292 0.87344 0.94203 0.0018817 0.0048414 0.13044 0.96345 0.92383 0.015375 0.99478 0.62655 0.0055725 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.6715 0.21999
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3708e-06 0.001154 0.04189 0.0006502 0.042535 0.037618 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.44439 0.87288 0.94193 0.0018908 0.004861 0.13044 0.96344 0.92383 0.015388 0.99476 0.62655 0.0055742 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.5933 0.21735
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3708e-06 0.001154 0.04189 0.0006502 0.042536 0.037618 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.44588 0.87232 0.94182 0.0019 0.0048808 0.13044 0.96344 0.92383 0.0154 0.99474 0.62655 0.005576 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.5144 0.21476
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3708e-06 0.001154 0.04189 0.0006502 0.042536 0.037618 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.44737 0.87176 0.94171 0.0019092 0.0049007 0.13044 0.96343 0.92383 0.015413 0.99472 0.62655 0.0055777 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.435 0.21219
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3709e-06 0.001154 0.04189 0.0006502 0.042536 0.037618 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.45039 0.87063 0.94149 0.0019281 0.0049412 0.13044 0.96342 0.92383 0.015438 0.99468 0.62654 0.0055812 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.2744 0.20714
0.10397 0.98801 5.525e-05 3.8182 0.012049 1.3709e-06 0.001154 0.041891 0.0006502 0.042536 0.037619 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.45344 0.86949 0.94126 0.0019473 0.0049825 0.13044 0.96342 0.92383 0.015464 0.99464 0.62654 0.0055847 0.43068 1.9523 1.9519 15.9971 145.002 0.00015291 -39.1114 0.20222
0.10398 0.98801 5.525e-05 3.8182 0.012049 1.371e-06 0.001154 0.041892 0.0006502 0.042537 0.037619 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.45963 0.86716 0.94081 0.001987 0.0050674 0.13044 0.9634 0.92383 0.015516 0.99455 0.62654 0.0055918 0.43068 1.9523 1.9519 15.9972 145.002 0.00015291 -38.7781 0.19272
0.10398 0.98801 5.525e-05 3.8182 0.012049 1.371e-06 0.001154 0.041892 0.0006502 0.042538 0.03762 0 0.045428 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.46597 0.86477 0.94035 0.0020283 0.0051556 0.13044 0.96338 0.92383 0.015569 0.99446 0.62654 0.005599 0.43068 1.9523 1.9519 15.9972 145.002 0.00015291 -38.4347 0.18366
0.10399 0.98801 5.525e-05 3.8182 0.012049 1.3711e-06 0.001154 0.041893 0.0006502 0.042539 0.037621 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.47245 0.86231 0.93988 0.0020715 0.0052475 0.13044 0.96336 0.92383 0.015623 0.99437 0.62654 0.0056062 0.43068 1.9523 1.9519 15.9972 145.002 0.00015291 -38.0809 0.17504
0.10399 0.98801 5.525e-05 3.8182 0.012049 1.3712e-06 0.001154 0.041894 0.0006502 0.042539 0.037621 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.47907 0.85979 0.93939 0.0021165 0.0053432 0.13044 0.96334 0.92383 0.015679 0.99428 0.62654 0.0056136 0.43068 1.9523 1.9519 15.9972 145.002 0.00015291 -37.7161 0.16681
0.104 0.98801 5.525e-05 3.8182 0.012049 1.3712e-06 0.001154 0.041895 0.0006502 0.04254 0.037622 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.48585 0.85719 0.9389 0.0021637 0.0054429 0.13044 0.96333 0.92383 0.015735 0.99418 0.62654 0.005621 0.43068 1.9523 1.9519 15.9973 145.002 0.00015291 -37.3401 0.15898
0.10401 0.98801 5.525e-05 3.8182 0.012049 1.3713e-06 0.001154 0.041896 0.0006502 0.042542 0.037623 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.49984 0.85177 0.93787 0.0022647 0.0056558 0.13044 0.96329 0.92383 0.015851 0.99399 0.62653 0.0056363 0.43068 1.9523 1.9519 15.9973 145.002 0.00015291 -36.5523 0.14439
0.10402 0.98801 5.525e-05 3.8182 0.012049 1.3715e-06 0.001154 0.041898 0.0006502 0.042543 0.037625 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.51443 0.84602 0.93679 0.0023758 0.0058888 0.13044 0.96325 0.92383 0.015972 0.99379 0.62653 0.0056521 0.43067 1.9523 1.9519 15.9974 145.002 0.00015291 -35.7141 0.13115
0.10403 0.98801 5.525e-05 3.8182 0.012049 1.3716e-06 0.001154 0.041899 0.0006502 0.042545 0.037626 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.52965 0.83988 0.93566 0.0024986 0.006145 0.13044 0.96321 0.92383 0.0161 0.99357 0.62653 0.0056685 0.43067 1.9523 1.9519 15.9974 145.002 0.00015291 -34.8219 0.11912
0.10404 0.98801 5.525e-05 3.8182 0.012049 1.3717e-06 0.001154 0.041901 0.0006502 0.042546 0.037627 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.54548 0.83333 0.93447 0.0026349 0.0064282 0.13044 0.96316 0.92384 0.016235 0.99336 0.62652 0.0056857 0.43067 1.9523 1.9519 15.9975 145.002 0.00015291 -33.8719 0.10819
0.10405 0.98801 5.525e-05 3.8182 0.012049 1.3719e-06 0.001154 0.041902 0.0006502 0.042548 0.037629 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.56194 0.82629 0.93321 0.0027872 0.0067428 0.13044 0.96312 0.92384 0.016378 0.99313 0.62652 0.0057038 0.43067 1.9523 1.9519 15.9976 145.002 0.00015291 -32.8607 0.098266
0.10406 0.98801 5.525e-05 3.8182 0.012049 1.372e-06 0.001154 0.041904 0.0006502 0.042549 0.03763 0 0.045426 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.579 0.81871 0.93189 0.0029581 0.0070945 0.13044 0.96307 0.92384 0.016532 0.9929 0.62651 0.0057229 0.43067 1.9523 1.9519 15.9976 145.002 0.00015291 -31.7846 0.089255
0.10407 0.98801 5.525e-05 3.8182 0.012049 1.3721e-06 0.001154 0.041905 0.0006502 0.042551 0.037631 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.59664 0.81053 0.93049 0.003151 0.0074898 0.13044 0.96302 0.92384 0.016699 0.99266 0.6265 0.0057433 0.43066 1.9523 1.9519 15.9977 145.002 0.00015291 -30.6407 0.08107
0.10408 0.98801 5.525e-05 3.8182 0.012049 1.3722e-06 0.001154 0.041907 0.0006502 0.042552 0.037633 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.61483 0.80165 0.92901 0.0033702 0.0079371 0.13044 0.96297 0.92384 0.01688 0.99241 0.6265 0.0057653 0.43066 1.9523 1.9519 15.9978 145.002 0.00015292 -29.426 0.073637
0.10409 0.98801 5.525e-05 3.8182 0.012049 1.3724e-06 0.001154 0.041908 0.0006502 0.042554 0.037634 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.63352 0.79201 0.92746 0.0036206 0.0084464 0.13044 0.96291 0.92384 0.017079 0.99217 0.62649 0.0057891 0.43066 1.9523 1.9519 15.9979 145.002 0.00015292 -28.1388 0.066886
0.1041 0.98801 5.525e-05 3.8182 0.012049 1.3725e-06 0.001154 0.04191 0.0006502 0.042555 0.037635 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.65265 0.78149 0.92582 0.0039087 0.0090304 0.13044 0.96285 0.92384 0.017299 0.99191 0.62648 0.0058153 0.43066 1.9523 1.9519 15.998 145.002 0.00015292 -26.7777 0.060755
0.1041 0.98801 5.525e-05 3.8182 0.012049 1.3726e-06 0.001154 0.041911 0.0006502 0.042557 0.037637 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052631 6.2774e-05 0.83743 0.0051034 0.0058414 0.67213 0.77001 0.9241 0.0042422 0.0097043 0.13044 0.96279 0.92384 0.017546 0.99166 0.62647 0.0058441 0.43066 1.9523 1.9519 15.9981 145.002 0.00015292 -25.3428 0.055187
0.10411 0.98801 5.525e-05 3.8182 0.012049 1.3727e-06 0.001154 0.041913 0.0006502 0.042558 0.037638 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.69188 0.75747 0.9223 0.0046308 0.010487 0.13044 0.96272 0.92384 0.017824 0.9914 0.62645 0.0058764 0.43065 1.9523 1.9519 15.9982 145.002 0.00015292 -23.8356 0.05013
0.10412 0.98801 5.525e-05 3.8182 0.012049 1.3729e-06 0.001154 0.041914 0.00065021 0.04256 0.03764 0 0.045426 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.71179 0.74375 0.92041 0.0050864 0.011403 0.13044 0.96264 0.92384 0.01814 0.99113 0.62644 0.0059126 0.43065 1.9523 1.9519 15.9983 145.002 0.00015292 -22.2591 0.045537
0.10413 0.98801 5.525e-05 3.8182 0.012049 1.373e-06 0.001154 0.041916 0.00065021 0.042561 0.037641 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.73173 0.72877 0.91844 0.0056237 0.012481 0.13044 0.96255 0.92384 0.018503 0.99087 0.62642 0.0059537 0.43065 1.9523 1.9519 15.9984 145.002 0.00015292 -20.6181 0.041366
0.10414 0.98801 5.525e-05 3.8182 0.012049 1.3731e-06 0.001154 0.041917 0.00065021 0.042563 0.037642 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.75156 0.71246 0.91639 0.0062607 0.013755 0.13044 0.96246 0.92384 0.018921 0.9906 0.62639 0.0060005 0.43065 1.9523 1.9519 15.9985 145.002 0.00015292 -18.9195 0.037578
0.10415 0.98801 5.525e-05 3.8182 0.012049 1.3732e-06 0.001154 0.041919 0.00065021 0.042564 0.037644 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.77114 0.69476 0.91427 0.0070194 0.01527 0.13044 0.96235 0.92384 0.019404 0.99034 0.62637 0.0060541 0.43065 1.9523 1.9519 15.9987 145.002 0.00015292 -17.1719 0.034137
0.10416 0.98801 5.525e-05 3.8182 0.012049 1.3734e-06 0.001154 0.04192 0.00065021 0.042566 0.037645 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.79032 0.67568 0.91209 0.0079264 0.017078 0.13044 0.96223 0.92384 0.019964 0.99007 0.62634 0.0061157 0.43064 1.9524 1.9519 15.9988 145.002 0.00015293 -15.3861 0.031013
0.10417 0.98801 5.525e-05 3.8182 0.012049 1.3735e-06 0.001154 0.041921 0.00065021 0.042567 0.037646 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.80897 0.65523 0.90985 0.0090134 0.019241 0.13044 0.9621 0.92384 0.020613 0.9898 0.6263 0.0061864 0.43064 1.9524 1.9519 15.9989 145.002 0.00015293 -13.574 0.028175
0.10418 0.98801 5.525e-05 3.8182 0.012049 1.3736e-06 0.001154 0.041923 0.00065021 0.042569 0.037648 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.82693 0.63351 0.90755 0.010318 0.021831 0.13044 0.96195 0.92384 0.021364 0.98953 0.62625 0.0062676 0.43064 1.9524 1.9519 15.9991 145.002 0.00015293 -11.7492 0.025598
0.10419 0.98801 5.525e-05 3.8182 0.012049 1.3738e-06 0.001154 0.041924 0.00065021 0.04257 0.037649 0 0.045425 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.84409 0.61066 0.90522 0.011884 0.024933 0.13044 0.96178 0.92384 0.022229 0.98926 0.6262 0.0063605 0.43064 1.9524 1.9519 15.9992 145.002 0.00015293 -9.9254 0.023257
0.1042 0.98801 5.525e-05 3.8182 0.012049 1.3739e-06 0.001154 0.041926 0.00065021 0.042572 0.03765 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.86033 0.58685 0.90284 0.01376 0.028643 0.13044 0.9616 0.92384 0.02322 0.98899 0.62613 0.0064662 0.43064 1.9524 1.9519 15.9993 145.002 0.00015293 -8.1167 0.021131
0.10421 0.98801 5.525e-05 3.8182 0.012049 1.374e-06 0.001154 0.041927 0.00065021 0.042573 0.037652 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.87556 0.56231 0.90044 0.016003 0.033065 0.13044 0.96139 0.92384 0.024349 0.98872 0.62606 0.0065859 0.43063 1.9524 1.9519 15.9994 145.002 0.00015293 -6.3366 0.0192
0.10422 0.98801 5.525e-05 3.8182 0.012049 1.3741e-06 0.001154 0.041929 0.00065021 0.042575 0.037653 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.88973 0.53727 0.89801 0.018672 0.038314 0.13044 0.96117 0.92384 0.025623 0.98845 0.62598 0.0067205 0.43063 1.9524 1.9519 15.9996 145.002 0.00015294 -4.5974 0.017447
0.10423 0.98801 5.525e-05 3.8182 0.012049 1.3743e-06 0.001154 0.04193 0.00065021 0.042576 0.037654 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.90279 0.51199 0.89557 0.021833 0.044509 0.13044 0.96092 0.92383 0.027052 0.98818 0.62588 0.0068707 0.43063 1.9524 1.9519 15.9997 145.002 0.00015294 -2.9102 0.015855
0.10424 0.98801 5.525e-05 3.8182 0.012049 1.3744e-06 0.001154 0.041932 0.00065021 0.042578 0.037656 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.91473 0.4867 0.89311 0.025552 0.051771 0.13044 0.96066 0.92383 0.028638 0.9879 0.62578 0.0070372 0.43063 1.9524 1.9519 15.9998 145.002 0.00015294 -1.2838 0.014408
0.10425 0.98801 5.525e-05 3.8182 0.012049 1.3745e-06 0.001154 0.041933 0.00065021 0.042579 0.037657 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.92452 0.46412 0.89089 0.029431 0.059316 0.13044 0.96041 0.92383 0.030204 0.98766 0.62567 0.0072011 0.43063 1.9524 1.9519 15.9999 145.002 0.00015294 0.12186 0.01322
0.10425 0.98801 5.525e-05 3.8182 0.012049 1.3745e-06 0.001154 0.041934 0.00065021 0.042579 0.037657 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.92613 0.46023 0.8905 0.03016 0.06073 0.13044 0.96036 0.92383 0.03049 0.98762 0.62565 0.007231 0.43063 1.9524 1.9519 15.9999 145.002 0.00015294 0.35996 0.013025
0.10425 0.98801 5.525e-05 3.8182 0.012049 1.3746e-06 0.001154 0.041934 0.00065021 0.04258 0.037658 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.92927 0.45248 0.88973 0.031668 0.063653 0.13044 0.96027 0.92383 0.031072 0.98753 0.62562 0.0072919 0.43063 1.9524 1.9519 15.9999 145.002 0.00015294 0.83076 0.012641
0.10426 0.98801 5.525e-05 3.8182 0.012049 1.3746e-06 0.001154 0.041934 0.00065021 0.04258 0.037658 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9323 0.44477 0.88895 0.033246 0.066706 0.13044 0.96018 0.92383 0.031671 0.98745 0.62558 0.0073545 0.43062 1.9524 1.9519 16 145.002 0.00015294 1.2942 0.01227
0.10426 0.98801 5.525e-05 3.8182 0.012049 1.3746e-06 0.001154 0.041935 0.00065021 0.042581 0.037658 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.93523 0.43712 0.88818 0.034896 0.069892 0.13044 0.96008 0.92383 0.032285 0.98736 0.62554 0.0074187 0.43062 1.9524 1.9519 16 145.002 0.00015295 1.7503 0.011909
0.10426 0.98801 5.525e-05 3.8182 0.012049 1.3747e-06 0.001154 0.041935 0.00065021 0.042581 0.037659 0 0.045424 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.93806 0.42953 0.8874 0.036619 0.073214 0.13044 0.95999 0.92383 0.032915 0.98728 0.6255 0.0074845 0.43062 1.9524 1.9519 16 145.002 0.00015295 2.1989 0.011559
0.10426 0.98801 5.525e-05 3.8182 0.012049 1.3747e-06 0.001154 0.041936 0.00065021 0.042581 0.037659 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.008349 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.94079 0.42199 0.88662 0.038418 0.076675 0.13044 0.95989 0.92383 0.033561 0.98719 0.62546 0.007552 0.43062 1.9524 1.9519 16.0001 145.002 0.00015295 2.6399 0.011219
0.10427 0.98801 5.525e-05 3.8182 0.012049 1.3748e-06 0.001154 0.041937 0.00065021 0.042582 0.03766 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.94595 0.40712 0.88507 0.042247 0.084021 0.13044 0.95969 0.92383 0.034899 0.98702 0.62537 0.0076918 0.43062 1.9524 1.9519 16.0001 145.002 0.00015295 3.4991 0.01057
0.10428 0.98801 5.525e-05 3.8182 0.012049 1.3749e-06 0.001154 0.041938 0.00065021 0.042583 0.037661 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.94996 0.39497 0.88378 0.045675 0.090574 0.13044 0.95952 0.92383 0.036059 0.98688 0.6253 0.0078131 0.43062 1.9524 1.9519 16.0002 145.002 0.00015295 4.1905 0.010059
0.10428 0.98801 5.525e-05 3.8182 0.012049 1.3749e-06 0.001154 0.041938 0.00065021 0.042584 0.037662 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.95371 0.38303 0.88249 0.049332 0.097536 0.13044 0.95935 0.92383 0.037262 0.98674 0.62523 0.0079388 0.43062 1.9524 1.9519 16.0002 145.002 0.00015295 4.8606 0.0095725
0.10429 0.98801 5.525e-05 3.8182 0.012049 1.375e-06 0.001154 0.041939 0.00065021 0.042585 0.037662 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.95722 0.37132 0.88119 0.053223 0.10491 0.13044 0.95918 0.92383 0.038507 0.9866 0.62515 0.0080689 0.43062 1.9524 1.9519 16.0003 145.002 0.00015296 5.5095 0.0091101
0.10429 0.98801 5.525e-05 3.8182 0.012049 1.3751e-06 0.001154 0.04194 0.00065021 0.042586 0.037663 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9605 0.35984 0.8799 0.057352 0.11271 0.13044 0.959 0.92383 0.039792 0.98646 0.62508 0.0082033 0.43062 1.9524 1.9518 16.0003 145.002 0.00015296 6.1373 0.0086702
0.1043 0.98801 5.525e-05 3.8182 0.012049 1.3751e-06 0.001154 0.041941 0.00065021 0.042586 0.037664 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.96356 0.34861 0.87861 0.061726 0.12093 0.13044 0.95882 0.92383 0.041117 0.98632 0.625 0.008342 0.43062 1.9524 1.9518 16.0004 145.002 0.00015296 6.7444 0.0082517
0.1043 0.98801 5.525e-05 3.8182 0.012049 1.3752e-06 0.001154 0.041941 0.00065021 0.042587 0.037664 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.96641 0.33763 0.87732 0.066346 0.12958 0.13044 0.95864 0.92383 0.042482 0.98618 0.62492 0.0084849 0.43062 1.9524 1.9517 16.0004 145.002 0.00015297 7.3309 0.0078537
0.10431 0.98801 5.525e-05 3.8182 0.012049 1.3753e-06 0.001154 0.041942 0.00065021 0.042588 0.037665 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.96905 0.3269 0.87602 0.071215 0.13864 0.13044 0.95845 0.92383 0.043885 0.98604 0.62484 0.0086319 0.43061 1.9524 1.9517 16.0004 145.002 0.00015297 7.8972 0.0074752
0.10431 0.98801 5.525e-05 3.8182 0.012049 1.3753e-06 0.001154 0.041943 0.00065021 0.042589 0.037666 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.97151 0.31644 0.87473 0.076336 0.14812 0.13044 0.95826 0.92383 0.045326 0.9859 0.62476 0.008783 0.43061 1.9524 1.9516 16.0005 145.002 0.00015297 8.4437 0.0071151
0.10432 0.98801 5.525e-05 3.8182 0.012049 1.3754e-06 0.001154 0.041944 0.00065021 0.042589 0.037667 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.97379 0.30623 0.87344 0.081709 0.15801 0.13044 0.95807 0.92382 0.046803 0.98575 0.62468 0.0089381 0.43061 1.9524 1.9515 16.0005 145.002 0.00015298 8.9709 0.0067726
0.10432 0.98801 5.525e-05 3.8182 0.012049 1.3755e-06 0.001154 0.041945 0.00065021 0.04259 0.037667 0 0.045423 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9759 0.29629 0.87215 0.087334 0.1683 0.13044 0.95788 0.92382 0.048316 0.98561 0.6246 0.0090971 0.43061 1.9524 1.9514 16.0005 145.002 0.00015299 9.4791 0.0064468
0.10433 0.98801 5.525e-05 3.8182 0.012049 1.3756e-06 0.001154 0.041946 0.00065021 0.042592 0.037669 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.97965 0.2772 0.86958 0.099333 0.19004 0.13044 0.95749 0.92382 0.051445 0.98533 0.62444 0.0094263 0.43061 1.9524 1.9511 16.0006 145.002 0.000153 10.4407 0.0058422
0.10434 0.98801 5.525e-05 3.8182 0.012049 1.3757e-06 0.001154 0.041948 0.00065022 0.042593 0.03767 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.98284 0.25914 0.867 0.11232 0.21324 0.13044 0.9571 0.92382 0.054704 0.98505 0.62427 0.0097702 0.43061 1.9524 1.9507 16.0007 145.002 0.00015303 11.3326 0.0052952
0.10435 0.98801 5.525e-05 3.8182 0.012049 1.3759e-06 0.001154 0.041949 0.00065022 0.042595 0.037671 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.98555 0.24211 0.86444 0.12625 0.23776 0.13044 0.9567 0.92382 0.058084 0.98477 0.6241 0.010128 0.43061 1.9524 1.9502 16.0007 145.002 0.00015305 12.159 0.0048002
0.10436 0.98801 5.525e-05 3.8182 0.012049 1.376e-06 0.001154 0.041951 0.00065022 0.042596 0.037673 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.98784 0.22607 0.86187 0.14109 0.26345 0.13044 0.9563 0.92381 0.061578 0.98449 0.62394 0.010499 0.4306 1.9524 1.9495 16.0008 145.002 0.00015309 12.9241 0.0043525
0.10437 0.98801 5.525e-05 3.8182 0.012049 1.3761e-06 0.001154 0.041952 0.00065022 0.042598 0.037674 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.98977 0.211 0.85932 0.15678 0.29013 0.13044 0.9559 0.92381 0.065178 0.98421 0.62376 0.010882 0.4306 1.9524 1.9487 16.0008 145.002 0.00015313 13.6321 0.0039474
0.10438 0.98801 5.525e-05 3.8182 0.012049 1.3763e-06 0.001154 0.041954 0.00065022 0.0426 0.037676 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99139 0.19684 0.85676 0.17326 0.31762 0.13044 0.95549 0.92381 0.068875 0.98392 0.62359 0.011277 0.4306 1.9524 1.9477 16.0009 145.002 0.00015319 14.2871 0.0035808
0.10439 0.98801 5.525e-05 3.8182 0.012049 1.3764e-06 0.001154 0.041955 0.00065022 0.042601 0.037677 0 0.045422 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99275 0.18356 0.85422 0.19046 0.34574 0.13044 0.95508 0.9238 0.072662 0.98364 0.62342 0.011682 0.4306 1.9524 1.9464 16.0009 145.002 0.00015325 14.893 0.0032492
0.1044 0.98801 5.525e-05 3.8182 0.012049 1.3765e-06 0.001154 0.041957 0.00065022 0.042603 0.037678 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99388 0.17113 0.85168 0.20829 0.37427 0.13044 0.95467 0.9238 0.076531 0.98336 0.62325 0.012098 0.43059 1.9524 1.9449 16.0009 145.002 0.00015333 15.4533 0.0029492
0.10441 0.98801 5.525e-05 3.8182 0.012049 1.3767e-06 0.001154 0.041959 0.00065022 0.042604 0.03768 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99483 0.15948 0.84915 0.22669 0.40303 0.13044 0.95426 0.92379 0.080476 0.98308 0.62308 0.012524 0.43059 1.9524 1.9432 16.001 145.002 0.00015342 15.9715 0.0026778
0.10442 0.98801 5.525e-05 3.8182 0.012049 1.3768e-06 0.001154 0.04196 0.00065022 0.042606 0.037681 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99561 0.14859 0.84662 0.24557 0.43184 0.13044 0.95384 0.92379 0.084489 0.9828 0.6229 0.012959 0.43059 1.9524 1.9412 16.001 145.002 0.00015352 16.4509 0.0024322
0.10443 0.98801 5.525e-05 3.8182 0.012049 1.3769e-06 0.001154 0.041962 0.00065022 0.042607 0.037683 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99627 0.13841 0.8441 0.26485 0.46052 0.13044 0.95343 0.92378 0.088565 0.98252 0.62273 0.013403 0.43059 1.9523 1.9389 16.001 145.002 0.00015364 16.8946 0.00221
0.10444 0.98801 5.525e-05 3.8182 0.012049 1.377e-06 0.001154 0.041963 0.00065022 0.042609 0.037684 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99681 0.1289 0.84159 0.28443 0.48891 0.13044 0.95301 0.92378 0.092696 0.98224 0.62256 0.013854 0.43059 1.9523 1.9363 16.0011 145.002 0.00015377 17.3051 0.002009
0.10445 0.98801 5.525e-05 3.8182 0.012049 1.3772e-06 0.001154 0.041965 0.00065022 0.04261 0.037686 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99726 0.12003 0.83908 0.30426 0.51685 0.13044 0.95259 0.92377 0.096878 0.98196 0.62238 0.014313 0.43058 1.9523 1.9333 16.0011 145.002 0.00015393 17.6852 0.0018272
0.10446 0.98801 5.525e-05 3.8182 0.012049 1.3773e-06 0.001154 0.041966 0.00065022 0.042612 0.037687 0 0.045421 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99763 0.11174 0.83658 0.32424 0.54422 0.13044 0.95218 0.92377 0.10111 0.98168 0.62221 0.014778 0.43058 1.9523 1.93 16.0011 145.002 0.0001541 18.0372 0.0016626
0.10447 0.98801 5.525e-05 3.8182 0.012049 1.3774e-06 0.001154 0.041968 0.00065022 0.042614 0.037688 0 0.04542 0.0389 0 0.84598 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99794 0.10401 0.83409 0.3443 0.5709 0.13044 0.95176 0.92376 0.10537 0.9814 0.62203 0.015251 0.43058 1.9522 1.9263 16.0011 145.002 0.00015429 18.3634 0.0015138
0.10448 0.98801 5.525e-05 3.8182 0.012049 1.3775e-06 0.001154 0.041969 0.00065022 0.042615 0.037689 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99814 0.098594 0.83224 0.35926 0.59026 0.13044 0.95145 0.92376 0.10857 0.98119 0.6219 0.015606 0.43058 1.9522 1.9233 16.0011 145.002 0.00015444 18.5908 0.0014582
0.10448 0.98801 5.525e-05 3.8182 0.012049 1.3776e-06 0.001154 0.04197 0.00065022 0.042616 0.03769 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99827 0.094646 0.83083 0.37066 0.60473 0.13044 0.95121 0.92375 0.11103 0.98103 0.6218 0.01588 0.43058 1.9522 1.9209 16.0011 145.002 0.00015457 18.756 0.0014553
0.10449 0.98801 5.525e-05 3.8182 0.012049 1.3777e-06 0.001154 0.041971 0.00065022 0.042616 0.037691 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99839 0.090853 0.82942 0.38205 0.61891 0.13044 0.95097 0.92375 0.11349 0.98087 0.6217 0.016155 0.43058 1.9521 1.9183 16.0011 145.002 0.0001547 18.9142 0.0014666
0.1045 0.98801 5.525e-05 3.8182 0.012049 1.3778e-06 0.001154 0.041972 0.00065022 0.042617 0.037692 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9985 0.087208 0.82801 0.39339 0.63278 0.13044 0.95073 0.92374 0.11597 0.98071 0.6216 0.016432 0.43058 1.9521 1.9157 16.0011 145.002 0.00015484 19.0659 0.0014767
0.1045 0.98801 5.525e-05 3.8182 0.012049 1.3778e-06 0.001154 0.041973 0.00065022 0.042618 0.037693 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99858 0.084051 0.82675 0.40357 0.64501 0.13044 0.95052 0.92374 0.1182 0.98056 0.62151 0.016683 0.43057 1.9521 1.9133 16.0012 145.002 0.00015497 19.197 0.0014819
0.10451 0.98801 5.525e-05 3.8182 0.012049 1.3779e-06 0.001154 0.041973 0.00065022 0.042619 0.037693 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99866 0.081005 0.82549 0.4137 0.65698 0.13044 0.9503 0.92373 0.12044 0.98042 0.62142 0.016935 0.43057 1.952 1.9108 16.0012 145.002 0.0001551 19.3233 0.0014857
0.10451 0.98801 5.525e-05 3.8182 0.012049 1.378e-06 0.001154 0.041974 0.00065022 0.04262 0.037694 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99873 0.078068 0.82423 0.42379 0.66869 0.13044 0.95009 0.92373 0.12269 0.98028 0.62133 0.017188 0.43057 1.952 1.9081 16.0012 145.002 0.00015524 19.445 0.00149
0.10452 0.98801 5.525e-05 3.8182 0.012049 1.378e-06 0.001154 0.041975 0.00065022 0.042621 0.037695 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9988 0.075236 0.82297 0.43382 0.68013 0.13044 0.94987 0.92372 0.12494 0.98013 0.62124 0.017442 0.43057 1.952 1.9054 16.0012 145.002 0.00015538 19.5622 0.0014951
0.10452 0.98801 5.525e-05 3.8182 0.012049 1.3781e-06 0.001154 0.041976 0.00065022 0.042621 0.037695 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99886 0.072504 0.82171 0.44379 0.69129 0.13044 0.94966 0.92372 0.12719 0.97999 0.62116 0.017698 0.43057 1.9519 1.9025 16.0012 145.002 0.00015554 19.6751 0.0015004
0.10453 0.98801 5.525e-05 3.8182 0.012049 1.3782e-06 0.001154 0.041976 0.00065022 0.042622 0.037696 0 0.04542 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99891 0.06987 0.82046 0.45368 0.70219 0.13044 0.94944 0.92371 0.12945 0.97985 0.62107 0.017955 0.43057 1.9519 1.8994 16.0012 145.002 0.0001557 19.7839 0.0015057
0.10454 0.98801 5.525e-05 3.8182 0.012049 1.3783e-06 0.001154 0.041978 0.00065022 0.042624 0.037698 0 0.045419 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99901 0.064882 0.81796 0.47326 0.72316 0.13044 0.94902 0.9237 0.13398 0.97956 0.62089 0.018471 0.43057 1.9518 1.8929 16.0012 145.002 0.00015605 19.99 0.0015163
0.10455 0.98801 5.525e-05 3.8182 0.012049 1.3784e-06 0.001154 0.04198 0.00065023 0.042625 0.037699 0 0.045419 0.0389 0 0.84599 0.22729 0.058898 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99908 0.060694 0.81571 0.49059 0.7411 0.13044 0.94863 0.92369 0.13807 0.9793 0.62072 0.01894 0.43057 1.9517 1.8863 16.0012 145.002 0.00015639 20.1632 0.0015257
0.10456 0.98801 5.525e-05 3.8182 0.012049 1.3785e-06 0.001154 0.041981 0.00065023 0.042627 0.0377 0 0.045419 0.0389 0 0.84599 0.22729 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99914 0.056773 0.81347 0.50764 0.75814 0.13044 0.94824 0.92368 0.14217 0.97904 0.62056 0.019411 0.43056 1.9516 1.879 16.0012 145.002 0.00015678 20.3258 0.0015349
0.10456 0.98801 5.525e-05 3.8182 0.012049 1.3787e-06 0.001154 0.041982 0.00065023 0.042628 0.037701 0 0.045419 0.0389 0 0.84599 0.22729 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99919 0.053102 0.81123 0.52436 0.77431 0.13044 0.94786 0.92367 0.14627 0.97879 0.6204 0.019885 0.43056 1.9515 1.8709 16.0012 145.002 0.00015722 20.4785 0.0015442
0.10457 0.98801 5.525e-05 3.8182 0.012049 1.3788e-06 0.001154 0.041984 0.00065023 0.042629 0.037703 0 0.045419 0.0389 0 0.84599 0.22729 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99923 0.049667 0.80901 0.54076 0.78961 0.13044 0.94747 0.92365 0.15037 0.97853 0.62024 0.020362 0.43056 1.9514 1.8617 16.0012 145.002 0.00015771 20.6221 0.0015534
0.10458 0.98801 5.525e-05 3.8182 0.012049 1.3789e-06 0.001154 0.041985 0.00065023 0.042631 0.037704 0 0.045419 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99927 0.046451 0.80678 0.5568 0.80406 0.13044 0.94708 0.92364 0.15448 0.97827 0.62008 0.020841 0.43056 1.9512 1.8514 16.0012 145.0019 0.00015827 20.7574 0.0015626
0.10459 0.98801 5.525e-05 3.8182 0.012049 1.379e-06 0.001154 0.041987 0.00065023 0.042632 0.037705 0 0.045419 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9993 0.043441 0.80457 0.57249 0.81769 0.13044 0.9467 0.92362 0.15859 0.97801 0.61992 0.021323 0.43056 1.9511 1.8398 16.0012 145.0019 0.0001589 20.885 0.0015718
0.1046 0.98801 5.525e-05 3.8182 0.012049 1.3792e-06 0.001154 0.041988 0.00065023 0.042634 0.037707 0 0.045419 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99933 0.040625 0.80235 0.5878 0.83052 0.13044 0.94631 0.9236 0.1627 0.97776 0.61976 0.021806 0.43055 1.9509 1.8267 16.0012 145.0019 0.00015962 21.0056 0.001581
0.10461 0.98801 5.525e-05 3.8182 0.012049 1.3793e-06 0.001154 0.04199 0.00065023 0.042635 0.037708 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99935 0.03799 0.80015 0.60273 0.84258 0.13044 0.94592 0.92359 0.16681 0.9775 0.61959 0.022292 0.43055 1.9507 1.812 16.0012 145.0019 0.00016043 21.1197 0.0015903
0.10462 0.98801 5.525e-05 3.8182 0.012049 1.3794e-06 0.001154 0.041991 0.00065023 0.042637 0.037709 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99937 0.035524 0.79795 0.61728 0.8539 0.13044 0.94554 0.92356 0.17092 0.97724 0.61943 0.02278 0.43055 1.9505 1.7955 16.0012 145.0019 0.00016134 21.2279 0.0015995
0.10463 0.98801 5.525e-05 3.8182 0.012049 1.3795e-06 0.001154 0.041992 0.00065023 0.042638 0.037711 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99939 0.033217 0.79576 0.63144 0.86452 0.13044 0.94515 0.92354 0.17502 0.97698 0.61927 0.02327 0.43055 1.9502 1.7772 16.0012 145.0019 0.00016237 21.3307 0.0016087
0.10464 0.98801 5.525e-05 3.8182 0.012049 1.3796e-06 0.001154 0.041994 0.00065023 0.042639 0.037712 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99941 0.031059 0.79357 0.64521 0.87445 0.13044 0.94477 0.92352 0.17912 0.97673 0.61911 0.023761 0.43055 1.95 1.757 16.0012 145.0019 0.00016352 21.4286 0.0016179
0.10465 0.98801 5.525e-05 3.8182 0.012049 1.3798e-06 0.001154 0.041995 0.00065023 0.042641 0.037713 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083491 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99942 0.029041 0.79139 0.65858 0.88374 0.13044 0.94438 0.92349 0.18321 0.97647 0.61895 0.024254 0.43054 1.9497 1.7349 16.0012 145.0019 0.00016479 21.5219 0.0016271
0.10466 0.98801 5.525e-05 3.8182 0.012049 1.3799e-06 0.001154 0.041997 0.00065023 0.042642 0.037714 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99943 0.027153 0.78921 0.67157 0.89241 0.13044 0.94399 0.92347 0.1873 0.97621 0.61879 0.024749 0.43054 1.9493 1.7112 16.0012 145.0019 0.00016618 21.6111 0.0016363
0.10467 0.98801 5.525e-05 3.8182 0.012049 1.38e-06 0.001154 0.041998 0.00065023 0.042644 0.037716 0 0.045418 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99945 0.025387 0.78704 0.68417 0.90051 0.13044 0.94361 0.92344 0.19137 0.97595 0.61863 0.025245 0.43054 1.9489 1.6859 16.0012 145.0019 0.00016768 21.6965 0.0016456
0.10467 0.98801 5.525e-05 3.8182 0.012049 1.3801e-06 0.001154 0.042 0.00065023 0.042645 0.037717 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99945 0.023735 0.78488 0.69638 0.90805 0.13044 0.94322 0.92341 0.19544 0.9757 0.61846 0.025742 0.43054 1.9485 1.6593 16.0012 145.0019 0.0001693 21.7785 0.0016548
0.10468 0.98801 5.525e-05 3.8182 0.012049 1.3803e-06 0.001154 0.042001 0.00065023 0.042647 0.037718 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99946 0.02219 0.78272 0.70821 0.91507 0.13044 0.94284 0.92338 0.19951 0.97544 0.6183 0.026241 0.43054 1.9481 1.6318 16.0012 145.0019 0.000171 21.8573 0.001664
0.10469 0.98801 5.525e-05 3.8182 0.012049 1.3804e-06 0.001154 0.042002 0.00065023 0.042648 0.03772 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99947 0.020745 0.78057 0.71966 0.92161 0.13044 0.94245 0.92334 0.20356 0.97518 0.61814 0.026741 0.43053 1.9476 1.6036 16.0012 145.0019 0.00017279 21.9334 0.0016732
0.1047 0.98801 5.525e-05 3.8182 0.012049 1.3805e-06 0.001154 0.042004 0.00065023 0.042649 0.037721 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99948 0.019394 0.77842 0.73074 0.92768 0.13044 0.94207 0.92331 0.2076 0.97493 0.61798 0.027243 0.43053 1.947 1.5752 16.0012 145.0019 0.00017464 22.0069 0.0016824
0.10471 0.98801 5.525e-05 3.8182 0.012049 1.3806e-06 0.001154 0.042005 0.00065023 0.042651 0.037722 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99948 0.01813 0.77628 0.74146 0.93332 0.13044 0.94168 0.92327 0.21164 0.97467 0.61782 0.027745 0.43053 1.9465 1.5466 16.0012 145.0019 0.00017654 22.078 0.0016917
0.10472 0.98801 5.525e-05 3.8182 0.012049 1.3807e-06 0.001154 0.042007 0.00065023 0.042652 0.037723 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99949 0.016948 0.77415 0.75182 0.93855 0.13044 0.9413 0.92323 0.21566 0.97441 0.61766 0.028249 0.43053 1.9458 1.5183 16.0012 145.0019 0.00017847 22.147 0.0017009
0.10473 0.98801 5.525e-05 3.8182 0.012049 1.3809e-06 0.001154 0.042008 0.00065023 0.042654 0.037725 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9995 0.015843 0.77202 0.76183 0.9434 0.13044 0.94091 0.92318 0.21967 0.97416 0.6175 0.028754 0.43053 1.9452 1.4903 16.0012 145.0019 0.00018043 22.2141 0.0017101
0.10474 0.98801 5.525e-05 3.8182 0.012049 1.381e-06 0.001154 0.04201 0.00065023 0.042655 0.037726 0 0.045417 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.9995 0.01481 0.7699 0.7715 0.94789 0.13044 0.94053 0.92314 0.22368 0.9739 0.61733 0.02926 0.43053 1.9445 1.463 16.0012 145.0019 0.0001824 22.2794 0.0017193
0.10475 0.98801 5.525e-05 3.8182 0.012049 1.3811e-06 0.001154 0.042011 0.00065023 0.042657 0.037727 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99951 0.013844 0.76778 0.78083 0.95205 0.13044 0.94014 0.92309 0.22767 0.97364 0.61717 0.029767 0.43052 1.9437 1.4363 16.0012 145.0019 0.00018437 22.3432 0.0017285
0.10476 0.98801 5.525e-05 3.8182 0.012049 1.3812e-06 0.001154 0.042012 0.00065024 0.042658 0.037729 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99951 0.012941 0.76567 0.78983 0.9559 0.13044 0.93976 0.92304 0.23165 0.97339 0.61701 0.030275 0.43052 1.9429 1.4104 16.0012 145.0019 0.00018634 22.4056 0.0017378
0.10477 0.98801 5.525e-05 3.8182 0.012049 1.3813e-06 0.001154 0.042014 0.00065024 0.042659 0.03773 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99951 0.012096 0.76356 0.79851 0.95946 0.13044 0.93937 0.92299 0.23561 0.97313 0.61685 0.030784 0.43052 1.9421 1.3853 16.0012 145.0018 0.0001883 22.4666 0.001747
0.10478 0.98801 5.525e-05 3.8182 0.012049 1.3815e-06 0.001154 0.042015 0.00065024 0.042661 0.037731 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99952 0.011306 0.76146 0.80688 0.96275 0.13044 0.93899 0.92293 0.23957 0.97288 0.61669 0.031294 0.43052 1.9412 1.361 16.0012 145.0018 0.00019024 22.5264 0.0017562
0.10479 0.98801 5.525e-05 3.8182 0.012049 1.3816e-06 0.001154 0.042017 0.00065024 0.042662 0.037733 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99952 0.010568 0.75937 0.81495 0.96578 0.13044 0.93861 0.92288 0.24351 0.97262 0.61653 0.031805 0.43052 1.9404 1.3376 16.0012 145.0018 0.00019217 22.5852 0.0017654
0.10479 0.98801 5.525e-05 3.8182 0.012049 1.3817e-06 0.001154 0.042018 0.00065024 0.042664 0.037734 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99953 0.0098779 0.75728 0.82272 0.96858 0.13044 0.93822 0.92282 0.24744 0.97236 0.61637 0.032317 0.43051 1.9394 1.3151 16.0012 145.0018 0.00019407 22.643 0.0017746
0.1048 0.98801 5.525e-05 3.8182 0.012049 1.3818e-06 0.001154 0.04202 0.00065024 0.042665 0.037735 0 0.045416 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2774e-05 0.83743 0.0051034 0.0058414 0.99953 0.0092326 0.7552 0.83021 0.97117 0.13044 0.93784 0.92276 0.25136 0.97211 0.61621 0.032829 0.43051 1.9385 1.2933 16.0012 145.0018 0.00019596 22.6998 0.0017839
0.10481 0.98801 5.525e-05 3.8182 0.012049 1.382e-06 0.001154 0.042021 0.00065024 0.042667 0.037736 0 0.045415 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99953 0.0086293 0.75312 0.83742 0.97355 0.13044 0.93746 0.92269 0.25527 0.97185 0.61605 0.033343 0.43051 1.9375 1.2724 16.0012 145.0018 0.00019782 22.7559 0.0017931
0.10482 0.98801 5.525e-05 3.8182 0.012049 1.3821e-06 0.001154 0.042022 0.00065024 0.042668 0.037738 0 0.045415 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99954 0.0080653 0.75105 0.84435 0.97574 0.13044 0.93707 0.92263 0.25916 0.97159 0.61588 0.033857 0.43051 1.9365 1.2523 16.0012 145.0018 0.00019966 22.8111 0.0018023
0.10483 0.98801 5.525e-05 3.8182 0.012049 1.3822e-06 0.001154 0.042024 0.00065024 0.04267 0.037739 0 0.045415 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99954 0.007538 0.74898 0.85103 0.97776 0.13044 0.93669 0.92256 0.26304 0.97134 0.61572 0.034373 0.43051 1.9354 1.2329 16.0012 145.0018 0.00020148 22.8656 0.0018115
0.10484 0.98801 5.525e-05 3.8182 0.012049 1.3823e-06 0.001154 0.042025 0.00065024 0.042671 0.03774 0 0.045415 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99954 0.0070451 0.74692 0.85745 0.97962 0.13044 0.93631 0.92249 0.26691 0.97108 0.61556 0.034889 0.4305 1.9343 1.2142 16.0012 145.0018 0.00020327 22.9194 0.0018207
0.10485 0.98801 5.525e-05 3.8182 0.012049 1.3824e-06 0.001154 0.042027 0.00065024 0.042672 0.037742 0 0.045415 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99955 0.0065843 0.74487 0.86362 0.98133 0.13044 0.93592 0.92241 0.27076 0.97083 0.6154 0.035406 0.4305 1.9332 1.1963 16.0012 145.0018 0.00020504 22.9726 0.0018299
0.10487 0.98801 5.525e-05 3.8182 0.012049 1.3827e-06 0.001154 0.04203 0.00065024 0.042675 0.037744 0 0.045415 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99955 0.0057509 0.74078 0.87525 0.98435 0.13044 0.93516 0.92226 0.27843 0.97032 0.61508 0.036442 0.4305 1.931 1.1623 16.0012 145.0018 0.00020852 23.0772 0.0018484
0.10489 0.98801 5.525e-05 3.8182 0.012049 1.3829e-06 0.001154 0.042032 0.00065024 0.042678 0.037747 0 0.045414 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99956 0.0050912 0.73711 0.88496 0.98666 0.13044 0.93447 0.92211 0.28528 0.96986 0.61479 0.037378 0.4305 1.9288 1.1338 16.0012 145.0018 0.00021157 23.1693 0.001865
0.1049 0.98801 5.525e-05 3.8182 0.012049 1.3831e-06 0.001154 0.042035 0.00065024 0.04268 0.037749 0 0.045414 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99956 0.004507 0.73347 0.89398 0.98864 0.13044 0.93378 0.92196 0.29209 0.9694 0.6145 0.038315 0.43049 1.9266 1.107 16.0012 145.0017 0.00021455 23.2597 0.0018816
0.10492 0.98801 5.525e-05 3.8182 0.012049 1.3833e-06 0.001154 0.042037 0.00065024 0.042683 0.037751 0 0.045414 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99956 0.0039897 0.72984 0.90236 0.99033 0.13044 0.93309 0.92179 0.29886 0.96894 0.61421 0.039256 0.43049 1.9244 1.0819 16.0012 145.0017 0.00021746 23.3483 0.0018982
0.10493 0.98801 5.525e-05 3.8182 0.012049 1.3836e-06 0.001154 0.04204 0.00065024 0.042686 0.037754 0 0.045414 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99957 0.0035316 0.72623 0.91013 0.99177 0.13044 0.93241 0.92163 0.30558 0.96848 0.61392 0.040198 0.43049 1.922 1.0583 16.0012 145.0017 0.00022032 23.4351 0.0019148
0.10495 0.98801 5.525e-05 3.8182 0.012049 1.3838e-06 0.001154 0.042042 0.00065024 0.042688 0.037756 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99957 0.0031259 0.72264 0.91734 0.993 0.13044 0.93172 0.92145 0.31225 0.96802 0.61363 0.041143 0.43048 1.9197 1.0361 16.0012 145.0017 0.00022311 23.5201 0.0019314
0.10497 0.98801 5.525e-05 3.8182 0.012049 1.384e-06 0.001154 0.042045 0.00065024 0.042691 0.037758 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0027668 0.71906 0.92401 0.99405 0.13044 0.93103 0.92127 0.31888 0.96756 0.61334 0.04209 0.43048 1.9172 1.0151 16.0012 145.0017 0.00022585 23.6033 0.001948
0.10498 0.98801 5.525e-05 3.8182 0.012049 1.3842e-06 0.001154 0.042048 0.00065025 0.042693 0.037761 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0024488 0.7155 0.93019 0.99494 0.13044 0.93035 0.92108 0.32546 0.9671 0.61305 0.043039 0.43048 1.9148 0.99531 16.0012 145.0017 0.00022853 23.6846 0.0019645
0.10499 0.98801 5.525e-05 3.8182 0.012049 1.3843e-06 0.001154 0.042049 0.00065025 0.042694 0.037761 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0023344 0.71412 0.93248 0.99525 0.13044 0.93008 0.921 0.32803 0.96692 0.61294 0.043412 0.43047 1.9138 0.98786 16.0012 145.0017 0.00022957 23.7158 0.001971
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.042049 0.00065025 0.042695 0.037762 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0022478 0.71302 0.93424 0.99548 0.13044 0.92987 0.92094 0.33005 0.96678 0.61285 0.043706 0.43047 1.913 0.98209 16.0012 145.0017 0.00023038 23.7403 0.0019762
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042695 0.037762 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0022312 0.71281 0.93458 0.99553 0.13044 0.92983 0.92093 0.33045 0.96675 0.61283 0.043764 0.43047 1.9128 0.98097 16.0012 145.0017 0.00023054 23.7451 0.0019772
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021984 0.71238 0.93525 0.99561 0.13044 0.92974 0.92091 0.33124 0.9667 0.6128 0.043879 0.43047 1.9125 0.97874 16.0012 145.0017 0.00023086 23.7546 0.0019792
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021913 0.71228 0.9354 0.99563 0.13044 0.92972 0.9209 0.33141 0.96668 0.61279 0.043905 0.43047 1.9125 0.97826 16.0012 145.0017 0.00023092 23.7567 0.0019796
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021882 0.71224 0.93547 0.99564 0.13044 0.92972 0.9209 0.33149 0.96668 0.61279 0.043916 0.43047 1.9124 0.97804 16.0012 145.0017 0.00023096 23.7576 0.0019798
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021818 0.71216 0.9356 0.99566 0.13044 0.9297 0.92089 0.33164 0.96667 0.61278 0.043938 0.43047 1.9124 0.97761 16.0012 145.0017 0.00023102 23.7578 0.0019802
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021807 0.71214 0.93562 0.99566 0.13044 0.9297 0.92089 0.33167 0.96667 0.61278 0.043942 0.43047 1.9124 0.97753 16.0012 145.0017 0.00023103 23.7574 0.0019803
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021784 0.71211 0.93567 0.99567 0.13044 0.92969 0.92089 0.33173 0.96666 0.61278 0.043951 0.43047 1.9123 0.97737 16.0012 145.0017 0.00023105 23.7565 0.0019804
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021761 0.71208 0.93572 0.99567 0.13044 0.92969 0.92089 0.33179 0.96666 0.61278 0.043959 0.43047 1.9123 0.97721 16.0012 145.0017 0.00023107 23.7557 0.0019806
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021738 0.71205 0.93576 0.99568 0.13044 0.92968 0.92089 0.33184 0.96665 0.61277 0.043967 0.43047 1.9123 0.97705 16.0012 145.0017 0.0002311 23.7549 0.0019807
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021715 0.71202 0.93581 0.99568 0.13044 0.92967 0.92089 0.3319 0.96665 0.61277 0.043975 0.43047 1.9123 0.9769 16.0012 145.0017 0.00023112 23.7542 0.0019809
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021692 0.71199 0.93586 0.99569 0.13044 0.92967 0.92088 0.33195 0.96665 0.61277 0.043984 0.43047 1.9123 0.97674 16.0012 145.0017 0.00023114 23.7534 0.001981
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021646 0.71193 0.93595 0.9957 0.13044 0.92966 0.92088 0.33207 0.96664 0.61276 0.044 0.43047 1.9122 0.97642 16.0012 145.0017 0.00023119 23.7519 0.0019813
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021555 0.71181 0.93614 0.99573 0.13044 0.92963 0.92087 0.33229 0.96662 0.61275 0.044033 0.43047 1.9121 0.97579 16.0012 145.0017 0.00023128 23.7489 0.0019819
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3844e-06 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021464 0.71168 0.93633 0.99575 0.13044 0.92961 0.92087 0.33252 0.96661 0.61274 0.044066 0.43047 1.912 0.97516 16.0012 145.0017 0.00023137 23.7458 0.0019825
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3845e-06 0.001154 0.042051 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021283 0.71144 0.93671 0.9958 0.13044 0.92956 0.92085 0.33297 0.96657 0.61272 0.044132 0.43047 1.9119 0.97391 16.0012 145.0017 0.00023155 23.7398 0.0019836
0.105 0.98801 5.525e-05 3.8182 0.012049 1.3845e-06 0.001154 0.042051 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0021105 0.7112 0.93708 0.99584 0.13044 0.92951 0.92084 0.33342 0.96654 0.6127 0.044198 0.43047 1.9117 0.97267 16.0012 145.0017 0.00023173 23.7337 0.0019848
0.10501 0.98801 5.525e-05 3.8182 0.012049 1.3845e-06 0.001154 0.042051 0.00065025 0.042697 0.037764 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0020927 0.71095 0.93745 0.99589 0.13044 0.92947 0.92083 0.33387 0.96651 0.61268 0.044264 0.43047 1.9115 0.97142 16.0012 145.0017 0.00023191 23.7276 0.0019859
0.10501 0.98801 5.525e-05 3.8182 0.012049 1.3845e-06 0.001154 0.042051 0.00065025 0.042697 0.037764 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0020577 0.71046 0.93818 0.99598 0.13044 0.92937 0.9208 0.33477 0.96645 0.61264 0.044396 0.43047 1.9112 0.96895 16.0012 145.0016 0.00023227 23.7154 0.0019882
0.10501 0.98801 5.525e-05 3.8182 0.012049 1.3846e-06 0.001154 0.042052 0.00065025 0.042697 0.037764 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0020231 0.70997 0.93891 0.99607 0.13044 0.92928 0.92077 0.33566 0.96638 0.6126 0.044527 0.43047 1.9108 0.9665 16.0012 145.0016 0.00023262 23.7033 0.0019905
0.10501 0.98801 5.525e-05 3.8182 0.012049 1.3846e-06 0.001154 0.042052 0.00065025 0.042698 0.037765 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0019891 0.70949 0.93962 0.99615 0.13044 0.92918 0.92074 0.33656 0.96632 0.61256 0.044659 0.43047 1.9104 0.96406 16.0012 145.0016 0.00023298 23.6911 0.0019928
0.10502 0.98801 5.525e-05 3.8182 0.012049 1.3846e-06 0.001154 0.042053 0.00065025 0.042698 0.037765 0 0.045412 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0019229 0.70851 0.94102 0.99632 0.13044 0.92899 0.92069 0.33834 0.96619 0.61248 0.044922 0.43047 1.9097 0.95924 16.0012 145.0016 0.00023369 23.6667 0.0019974
0.10503 0.98801 5.525e-05 3.8182 0.012049 1.3848e-06 0.001154 0.042054 0.00065025 0.0427 0.037766 0 0.045412 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0017968 0.70656 0.94372 0.99662 0.13044 0.92861 0.92057 0.34189 0.96594 0.61232 0.045447 0.43047 1.9083 0.94981 16.0012 145.0016 0.0002351 23.6178 0.0020066
0.10503 0.98801 5.525e-05 3.8182 0.012049 1.3849e-06 0.001154 0.042055 0.00065025 0.042701 0.037768 0 0.045412 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0016905 0.70482 0.94603 0.99687 0.13044 0.92827 0.92047 0.34506 0.96571 0.61218 0.045918 0.43046 1.907 0.94155 16.0011 145.0016 0.00023636 23.5737 0.0020149
0.10504 0.98801 5.525e-05 3.8182 0.012049 1.385e-06 0.001154 0.042057 0.00065025 0.042702 0.037769 0 0.045412 0.0389 0 0.84599 0.2273 0.058899 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0015904 0.70307 0.94823 0.9971 0.13044 0.92793 0.92036 0.34821 0.96548 0.61203 0.046388 0.43046 1.9057 0.93351 16.0011 145.0016 0.00023761 23.5295 0.0020232
0.10505 0.98801 5.525e-05 3.8182 0.012049 1.3851e-06 0.001154 0.042058 0.00065025 0.042704 0.03777 0 0.045412 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0014963 0.70134 0.95033 0.99731 0.13044 0.92759 0.92025 0.35133 0.96525 0.61189 0.046858 0.43046 1.9043 0.92568 16.0011 145.0016 0.00023884 23.4852 0.0020315
0.10506 0.98801 5.525e-05 3.8182 0.012049 1.3852e-06 0.001154 0.042059 0.00065025 0.042705 0.037771 0 0.045412 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99959 0.0014077 0.6996 0.95234 0.9975 0.13044 0.92725 0.92015 0.35443 0.96503 0.61175 0.047326 0.43046 1.903 0.91804 16.0011 145.0016 0.00024007 23.4407 0.0020398
0.10508 0.98801 5.525e-05 3.8182 0.012049 1.3854e-06 0.001154 0.042062 0.00065025 0.042708 0.037773 0 0.045412 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0012462 0.69615 0.95607 0.99783 0.13044 0.92657 0.91993 0.36057 0.96457 0.61146 0.048259 0.43046 1.9003 0.90335 16.0011 145.0016 0.00024249 23.3513 0.0020563
0.10509 0.98801 5.525e-05 3.8182 0.012049 1.3856e-06 0.001154 0.042064 0.00065025 0.04271 0.037776 0 0.045411 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.0011035 0.69271 0.95947 0.99811 0.13044 0.92589 0.9197 0.36663 0.96411 0.61117 0.049187 0.43045 1.8976 0.88937 16.0011 145.0016 0.00024487 23.2612 0.0020729
0.10511 0.98801 5.525e-05 3.8182 0.012049 1.3859e-06 0.001154 0.042067 0.00065025 0.042713 0.037778 0 0.045411 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99958 0.00097708 0.68929 0.96257 0.99834 0.13044 0.92521 0.91947 0.37259 0.96366 0.61088 0.050111 0.43045 1.8948 0.87606 16.0011 145.0015 0.00024721 23.1704 0.0020895
0.10513 0.98801 5.525e-05 3.8182 0.012049 1.3861e-06 0.001154 0.04207 0.00065025 0.042715 0.03778 0 0.045411 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99957 0.00086515 0.68589 0.9654 0.99854 0.13044 0.92453 0.91924 0.37848 0.9632 0.6106 0.051031 0.43045 1.8921 0.86338 16.0011 145.0015 0.00024951 23.0788 0.002106
0.10514 0.98801 5.525e-05 3.8182 0.012049 1.3863e-06 0.001154 0.042072 0.00065025 0.042718 0.037783 0 0.045411 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99957 0.00076602 0.6825 0.96798 0.9987 0.13044 0.92385 0.919 0.38428 0.96274 0.61031 0.051947 0.43044 1.8893 0.85129 16.0011 145.0015 0.00025177 22.9865 0.0021226
0.10517 0.98801 5.525e-05 3.8182 0.012049 1.3866e-06 0.001154 0.042076 0.00065025 0.042721 0.037786 0 0.04541 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99956 0.00064488 0.67773 0.97125 0.99889 0.13044 0.92289 0.91865 0.39235 0.9621 0.60991 0.053235 0.43044 1.8852 0.8351 16.0011 145.0015 0.00025492 22.8542 0.002146
0.10519 0.98801 5.525e-05 3.8182 0.012049 1.3869e-06 0.001154 0.042079 0.00065026 0.042725 0.037789 0 0.04541 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99956 0.00054296 0.673 0.97413 0.99903 0.13044 0.92193 0.9183 0.40026 0.96146 0.6095 0.054515 0.43043 1.8812 0.81993 16.0011 145.0015 0.00025801 22.7202 0.0021695
0.10521 0.98801 5.525e-05 3.8182 0.012049 1.3872e-06 0.001154 0.042083 0.00065026 0.042729 0.037793 0 0.04541 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99955 0.00045722 0.66831 0.97667 0.99915 0.13044 0.92097 0.91794 0.40801 0.96081 0.60909 0.055785 0.43043 1.8771 0.80569 16.0011 145.0014 0.00026102 22.5842 0.0021929
0.10524 0.98801 5.525e-05 3.8182 0.012049 1.3875e-06 0.001154 0.042087 0.00065026 0.042732 0.037796 0 0.045409 0.0389 0 0.84599 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99955 0.00038506 0.66364 0.97892 0.99923 0.13044 0.92001 0.91757 0.41561 0.96017 0.60869 0.057047 0.43042 1.873 0.7923 16.0011 145.0014 0.00026399 22.4464 0.0022164
0.10526 0.98801 5.525e-05 3.8182 0.012049 1.3878e-06 0.001154 0.04209 0.00065026 0.042736 0.037799 0 0.045409 0.0389 0 0.846 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99954 0.00032432 0.65901 0.98089 0.9993 0.13044 0.91906 0.91719 0.42305 0.95953 0.60829 0.0583 0.43042 1.8688 0.7797 16.0011 145.0014 0.00026689 22.3066 0.0022398
0.10528 0.98801 5.525e-05 3.8182 0.012049 1.3882e-06 0.001154 0.042094 0.00065026 0.04274 0.037803 0 0.045409 0.0389 0 0.846 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99953 0.00027319 0.65441 0.98264 0.99935 0.13044 0.91811 0.91681 0.43035 0.95888 0.60788 0.059544 0.43041 1.8646 0.76783 16.0011 145.0014 0.00026974 22.1648 0.0022633
0.10531 0.98801 5.525e-05 3.8182 0.012049 1.3885e-06 0.001154 0.042098 0.00065026 0.042743 0.037806 0 0.045408 0.0389 0 0.846 0.2273 0.0589 0.0083493 4.1053 0.052632 6.2775e-05 0.83743 0.0051034 0.0058414 0.99953 0.00023014 0.64985 0.98419 0.99939 0.13044 0.91715 0.91643 0.4375 0.95824 0.60748 0.06078 0.43041 1.8604 0.75663 16.001 145.0013 0.00027254 22.021 0.0022867
0.10535 0.98801 5.525e-05 3.8182 0.012049 1.3891e-06 0.001154 0.042105 0.00065026 0.042751 0.037812 0 0.045408 0.0389 0 0.846 0.2273 0.0589 0.0083493 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99951 0.00016329 0.64081 0.98678 0.99944 0.13044 0.91525 0.91563 0.45137 0.95696 0.60667 0.063223 0.4304 1.8519 0.73608 16.001 145.0013 0.00027799 21.7278 0.0023336
0.10539 0.98801 5.525e-05 3.8182 0.012049 1.3896e-06 0.001154 0.042111 0.00065026 0.042757 0.037818 0 0.045407 0.0389 0 0.846 0.2273 0.0589 0.0083493 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.9995 0.00012207 0.63325 0.98854 0.99947 0.13044 0.91364 0.91495 0.46269 0.95587 0.60599 0.065266 0.43039 1.8446 0.72036 16.001 145.0012 0.00028246 21.4735 0.0023733
0.10543 0.98801 5.525e-05 3.8182 0.012049 1.3901e-06 0.001154 0.042117 0.00065027 0.042763 0.037824 0 0.045406 0.0389 0 0.846 0.2273 0.0589 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99949 9.1334e-05 0.62578 0.98997 0.99947 0.13044 0.91204 0.91424 0.47362 0.95479 0.60531 0.067284 0.43038 1.8372 0.70604 16.001 145.0012 0.00028682 21.2141 0.0024131
0.10547 0.98801 5.525e-05 3.8182 0.012049 1.3906e-06 0.001154 0.042123 0.00065027 0.042769 0.037829 0 0.045406 0.0389 0 0.846 0.2273 0.0589 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99947 6.8422e-05 0.61839 0.99115 0.99947 0.13044 0.91044 0.91353 0.48418 0.9537 0.60463 0.069275 0.43038 1.8299 0.69297 16.001 145.0011 0.00029107 20.9502 0.0024529
0.10551 0.98801 5.525e-05 3.8182 0.012049 1.3912e-06 0.001154 0.04213 0.00065027 0.042775 0.037835 0 0.045405 0.0389 0 0.846 0.2273 0.0589 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99946 5.1287e-05 0.6111 0.99211 0.99947 0.13044 0.90884 0.9128 0.49437 0.95262 0.60395 0.07124 0.43037 1.8224 0.68101 16.001 145.0011 0.0002952 20.6821 0.0024926
0.10555 0.98801 5.525e-05 3.8182 0.012049 1.3917e-06 0.001154 0.042136 0.00065027 0.042781 0.03784 0 0.045405 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99944 3.8437e-05 0.60389 0.99289 0.99945 0.13044 0.90725 0.91206 0.50421 0.95154 0.60327 0.073179 0.43036 1.815 0.67007 16.0009 145.001 0.00029924 20.4102 0.0025324
0.10559 0.98801 5.525e-05 3.8182 0.012049 1.3922e-06 0.001154 0.042142 0.00065027 0.042788 0.037846 0 0.045404 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99942 2.8807e-05 0.59677 0.99354 0.99944 0.13044 0.90566 0.91131 0.51371 0.95046 0.6026 0.075092 0.43035 1.8076 0.66003 16.0009 145.001 0.00030318 20.135 0.0025721
0.10563 0.98801 5.525e-05 3.8182 0.012049 1.3927e-06 0.001154 0.042148 0.00065028 0.042794 0.037852 0 0.045404 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99941 2.1606e-05 0.58973 0.99406 0.99942 0.13044 0.90407 0.91055 0.52288 0.94938 0.60192 0.076978 0.43034 1.8001 0.65083 16.0009 145.0009 0.00030704 19.857 0.0026119
0.10567 0.98801 5.525e-05 3.8182 0.012049 1.3933e-06 0.001154 0.042154 0.00065028 0.0428 0.037857 0 0.045403 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99939 1.6221e-05 0.58278 0.99449 0.9994 0.13044 0.90249 0.90978 0.53174 0.9483 0.60125 0.078839 0.43033 1.7926 0.64238 16.0009 145.0008 0.00031081 19.5766 0.0026516
0.10571 0.98801 5.525e-05 3.8182 0.012049 1.3938e-06 0.001154 0.04216 0.00065028 0.042806 0.037863 0 0.045402 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99937 1.2179e-05 0.57591 0.99483 0.99937 0.13044 0.90092 0.909 0.54028 0.94723 0.60057 0.080674 0.43033 1.7851 0.63462 16.0009 145.0008 0.0003145 19.2943 0.0026914
0.10575 0.98801 5.525e-05 3.8182 0.012049 1.3943e-06 0.001154 0.042167 0.00065028 0.042812 0.037868 0 0.045402 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2775e-05 0.83743 0.0051034 0.0058414 0.99935 9.1419e-06 0.56912 0.9951 0.99935 0.13044 0.89934 0.90821 0.54852 0.94615 0.5999 0.082483 0.43032 1.7777 0.62749 16.0009 145.0007 0.00031811 19.0106 0.0027311
0.10579 0.98801 5.525e-05 3.8182 0.012049 1.3948e-06 0.001154 0.042173 0.00065028 0.042818 0.037874 0 0.045401 0.0389 0 0.846 0.2273 0.058901 0.0083494 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99933 6.8667e-06 0.56242 0.99532 0.99932 0.13044 0.89778 0.90741 0.55648 0.94508 0.59923 0.084267 0.43031 1.7702 0.62094 16.0009 145.0007 0.00032166 18.7259 0.0027709
0.10587 0.98801 5.525e-05 3.8182 0.012049 1.3959e-06 0.001154 0.042185 0.00065029 0.042831 0.037885 0 0.0454 0.0389 0 0.846 0.2273 0.058901 0.0083495 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99929 3.9024e-06 0.54925 0.99561 0.99926 0.13044 0.89466 0.90579 0.57157 0.94293 0.5979 0.08776 0.43029 1.7553 0.6094 16.0008 145.0006 0.00032854 18.1551 0.0028504
0.10595 0.98801 5.525e-05 3.8182 0.012049 1.3969e-06 0.001154 0.042197 0.00065029 0.042843 0.037896 0 0.045399 0.0389 0 0.846 0.2273 0.058901 0.0083495 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99925 2.2652e-06 0.53639 0.99575 0.99919 0.13044 0.89155 0.90413 0.58561 0.94079 0.59657 0.091155 0.43028 1.7404 0.5997 16.0008 145.0004 0.00033518 17.5851 0.0029299
0.10603 0.98801 5.525e-05 3.8182 0.012049 1.398e-06 0.001154 0.04221 0.00065029 0.042855 0.037907 0 0.045398 0.0389 0 0.84601 0.2273 0.058902 0.0083495 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.9992 1.3324e-06 0.52383 0.99578 0.99911 0.13044 0.88847 0.90245 0.5987 0.93866 0.59524 0.094454 0.43026 1.7257 0.59156 16.0008 145.0003 0.00034158 17.0187 0.0030094
0.10611 0.98801 5.525e-05 3.8182 0.012049 1.399e-06 0.001154 0.042222 0.0006503 0.042868 0.037919 0 0.045397 0.0389 0 0.84601 0.2273 0.058902 0.0083495 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99915 7.7133e-07 0.51158 0.99572 0.99903 0.13044 0.88541 0.90073 0.61088 0.93653 0.59393 0.097661 0.43024 1.711 0.58479 16.0007 145.0002 0.00034778 16.4585 0.0030889
0.10619 0.98801 5.525e-05 3.8182 0.012049 1.4001e-06 0.001154 0.042234 0.0006503 0.04288 0.03793 0 0.045395 0.0389 0 0.84601 0.2273 0.058902 0.0083495 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.9991 4.3628e-07 0.49962 0.99559 0.99893 0.13044 0.88237 0.89899 0.62223 0.9344 0.59261 0.10078 0.43023 1.6964 0.57921 16.0007 145.0001 0.00035379 15.9064 0.0031685
0.10627 0.98801 5.525e-05 3.8182 0.012049 1.4011e-06 0.001154 0.042247 0.00065031 0.042892 0.037941 0 0.045394 0.0389 0 0.84601 0.2273 0.058902 0.0083496 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99905 2.5175e-07 0.48794 0.99541 0.99884 0.13044 0.87935 0.89723 0.6328 0.93228 0.59131 0.10381 0.43021 1.682 0.57468 16.0007 144.9999 0.00035961 15.3644 0.003248
0.10635 0.98801 5.525e-05 3.8182 0.012049 1.4022e-06 0.001154 0.042259 0.00065031 0.042905 0.037952 0 0.045393 0.0389 0 0.84601 0.22731 0.058902 0.0083496 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99899 1.5327e-07 0.47654 0.99517 0.99873 0.13044 0.87636 0.89544 0.64265 0.93017 0.59001 0.10676 0.4302 1.6677 0.57106 16.0007 144.9998 0.00036526 14.8337 0.0033275
0.10643 0.98801 5.525e-05 3.8182 0.012049 1.4032e-06 0.001154 0.042271 0.00065031 0.042917 0.037963 0 0.045392 0.0389 0 0.84601 0.22731 0.058902 0.0083496 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99893 9.2783e-08 0.46541 0.99489 0.99862 0.13044 0.87338 0.89363 0.65182 0.92806 0.58872 0.10963 0.43018 1.6536 0.56827 16.0006 144.9997 0.00037076 14.3157 0.003407
0.10651 0.98801 5.525e-05 3.8182 0.012049 1.4043e-06 0.001154 0.042284 0.00065032 0.042929 0.037974 0 0.045391 0.0389 0 0.84601 0.22731 0.058902 0.0083496 4.1053 0.052633 6.2776e-05 0.83743 0.0051034 0.0058414 0.99887 5.1337e-08 0.45455 0.99458 0.9985 0.13044 0.87044 0.8918 0.66037 0.92595 0.58744 0.11242 0.43016 1.6396 0.56621 16.0006 144.9996 0.00037611 13.8111 0.0034865
0.10659 0.98801 5.525e-05 3.8182 0.012049 1.4053e-06 0.001154 0.042296 0.00065032 0.042942 0.037986 0 0.04539 0.0389 0 0.84601 0.22731 0.058903 0.0083497 4.1053 0.052634 6.2776e-05 0.83743 0.0051034 0.0058414 0.99881 2.7107e-08 0.44394 0.99423 0.99837 0.13044 0.86751 0.88995 0.66834 0.92385 0.58616 0.11514 0.43015 1.6258 0.56479 16.0006 144.9994 0.00038131 13.3207 0.003566
0.10667 0.98801 5.525e-05 3.8182 0.012049 1.4064e-06 0.001154 0.042308 0.00065032 0.042954 0.037997 0 0.045388 0.0389 0 0.84601 0.22731 0.058903 0.0083497 4.1053 0.052634 6.2776e-05 0.83743 0.0051034 0.0058414 0.99875 1.6627e-08 0.43359 0.99385 0.99824 0.13044 0.86462 0.88808 0.67576 0.92176 0.5849 0.1178 0.43013 1.6121 0.56397 16.0005 144.9993 0.00038639 12.8448 0.0036455
0.10682 0.98801 5.525e-05 3.8182 0.012049 1.4085e-06 0.001154 0.042333 0.00065033 0.042979 0.038019 0 0.045386 0.0389 0 0.84602 0.22731 0.058903 0.0083497 4.1053 0.052634 6.2777e-05 0.83743 0.0051034 0.0058414 0.99862 3.1677e-08 0.41362 0.99299 0.99794 0.13044 0.8589 0.88428 0.68913 0.91758 0.58239 0.12291 0.4301 1.5853 0.56386 16.0005 144.999 0.00039616 11.9375 0.0038045
0.10697 0.98801 5.525e-05 3.8182 0.012049 1.4104e-06 0.001154 0.042355 0.00065034 0.043001 0.038039 0 0.045384 0.0389 0 0.84602 0.22731 0.058903 0.0083498 4.1053 0.052634 6.2777e-05 0.83743 0.0051034 0.0058414 0.9985 3.6122e-08 0.39645 0.99214 0.99766 0.13044 0.85384 0.88082 0.69966 0.91384 0.58016 0.1273 0.43007 1.5618 0.56525 16.0004 144.9988 0.00040455 11.1717 0.0039477
0.10711 0.98801 5.525e-05 3.8182 0.012049 1.4122e-06 0.001154 0.042377 0.00065035 0.043023 0.038059 0 0.045382 0.0389 0 0.84602 0.22731 0.058904 0.0083498 4.1053 0.052634 6.2777e-05 0.83743 0.0051034 0.0058414 0.99838 1.7625e-08 0.38002 0.9912 0.99735 0.13044 0.84886 0.8773 0.70893 0.91011 0.57795 0.13151 0.43004 1.5389 0.56783 16.0004 144.9986 0.0004126 10.4528 0.0040908
0.10725 0.98801 5.525e-05 3.8182 0.012049 1.4141e-06 0.001154 0.042399 0.00065035 0.043045 0.038079 0 0.04538 0.0389 0 0.84602 0.22731 0.058904 0.0083498 4.1053 0.052634 6.2777e-05 0.83743 0.0051034 0.0058414 0.99825 -1.1718e-09 0.36427 0.99019 0.99703 0.13044 0.84397 0.87375 0.71709 0.90639 0.57578 0.13556 0.43001 1.5167 0.57141 16.0003 144.9984 0.00042031 9.7788 0.0042339
0.1074 0.98801 5.5249e-05 3.8182 0.012049 1.416e-06 0.001154 0.042422 0.00065036 0.043067 0.038099 0 0.045378 0.0389 0 0.84602 0.22731 0.058904 0.0083499 4.1053 0.052634 6.2777e-05 0.83743 0.0051034 0.0058414 0.99813 -3.3271e-09 0.3492 0.98912 0.99668 0.13044 0.83915 0.87016 0.72426 0.9027 0.57364 0.13946 0.42998 1.495 0.57586 16.0003 144.9981 0.00042772 9.1471 0.004377
0.10754 0.98801 5.5249e-05 3.8182 0.012049 1.4179e-06 0.001154 0.042444 0.00065036 0.04309 0.03812 0 0.045376 0.0389 0 0.84602 0.22731 0.058905 0.0083499 4.1053 0.052634 6.2777e-05 0.83743 0.0051034 0.0058414 0.998 2.9846e-09 0.33476 0.98799 0.99632 0.13044 0.83442 0.86653 0.73056 0.89902 0.57152 0.14322 0.42995 1.474 0.58104 16.0003 144.9979 0.00043484 8.5548 0.0045201
0.10768 0.98801 5.5249e-05 3.8182 0.012049 1.4198e-06 0.001154 0.042466 0.00065037 0.043112 0.03814 0 0.045374 0.0389 0 0.84603 0.22731 0.058905 0.0083499 4.1053 0.052634 6.2778e-05 0.83743 0.0051034 0.0058414 0.99787 4.1755e-09 0.32093 0.9868 0.99594 0.13044 0.82977 0.86288 0.73608 0.89535 0.56943 0.14685 0.42992 1.4536 0.58684 16.0002 144.9977 0.00044168 7.9991 0.0046633
0.10783 0.98801 5.5249e-05 3.8182 0.012049 1.4217e-06 0.001154 0.042488 0.00065038 0.043134 0.03816 0 0.045372 0.0389 0 0.84603 0.22731 0.058905 0.00835 4.1053 0.052635 6.2778e-05 0.83743 0.0051034 0.0058414 0.99775 -4.7849e-11 0.30769 0.98555 0.99554 0.13044 0.82519 0.8592 0.7409 0.8917 0.56737 0.15036 0.42989 1.4338 0.5932 16.0002 144.9974 0.00044826 7.4767 0.0048064
0.10797 0.98801 5.5249e-05 3.8182 0.012049 1.4236e-06 0.001154 0.04251 0.00065038 0.043156 0.03818 0 0.04537 0.0389 0 0.84603 0.22731 0.058906 0.00835 4.1053 0.052635 6.2778e-05 0.83743 0.0051034 0.0058414 0.99762 -2.2705e-09 0.295 0.98426 0.99513 0.13044 0.82068 0.8555 0.74509 0.88806 0.56534 0.15377 0.42986 1.4146 0.60001 16.0001 144.9972 0.00045458 6.9846 0.0049495
0.10811 0.98801 5.5249e-05 3.8182 0.012049 1.4254e-06 0.001154 0.042532 0.00065039 0.043178 0.0382 0 0.045367 0.0389 0 0.84603 0.22732 0.058906 0.0083501 4.1053 0.052635 6.2778e-05 0.83743 0.0051034 0.0058414 0.99749 -4.8461e-10 0.28285 0.98292 0.99471 0.13044 0.81625 0.85179 0.74872 0.88444 0.56334 0.15707 0.42983 1.3961 0.60723 16.0001 144.997 0.00046066 6.5202 0.0050926
0.10826 0.98801 5.5249e-05 3.8182 0.012049 1.4273e-06 0.001154 0.042555 0.0006504 0.0432 0.03822 0 0.045365 0.0389 0 0.84603 0.22732 0.058906 0.0083501 4.1053 0.052635 6.2778e-05 0.83743 0.0051034 0.0058414 0.99737 1.2542e-09 0.27121 0.98154 0.99428 0.13044 0.81189 0.84806 0.75184 0.88083 0.56137 0.16027 0.42981 1.3782 0.61478 16 144.9967 0.0004665 6.0806 0.0052357
0.1084 0.98801 5.5249e-05 3.8182 0.012049 1.4292e-06 0.001154 0.042577 0.0006504 0.043223 0.03824 0 0.045363 0.0389 0 0.84604 0.22732 0.058906 0.0083501 4.1053 0.052635 6.2778e-05 0.83743 0.0051034 0.0058414 0.99724 5.8673e-10 0.26006 0.98012 0.99383 0.13044 0.80759 0.84432 0.7545 0.87724 0.55942 0.16339 0.42978 1.3608 0.62262 16 144.9965 0.00047212 5.6634 0.0053789
0.10854 0.98801 5.5249e-05 3.8182 0.012049 1.4311e-06 0.001154 0.042599 0.00065041 0.043245 0.03826 0 0.045361 0.0389 0 0.84604 0.22732 0.058907 0.0083502 4.1053 0.052635 6.2778e-05 0.83743 0.0051034 0.0058414 0.99712 -6.2899e-10 0.24938 0.97866 0.99337 0.13044 0.80336 0.84057 0.75674 0.87366 0.55751 0.16642 0.42975 1.3441 0.6307 15.9999 144.9963 0.00047752 5.2664 0.005522
0.10869 0.98801 5.5249e-05 3.8182 0.012049 1.433e-06 0.001154 0.042621 0.00065042 0.043267 0.03828 0 0.045359 0.0389 0 0.84604 0.22732 0.058907 0.0083502 4.1053 0.052635 6.2779e-05 0.83743 0.0051034 0.0058414 0.997 -4.8718e-10 0.23914 0.97716 0.9929 0.13044 0.79919 0.83681 0.75861 0.8701 0.55561 0.16937 0.42972 1.328 0.63898 15.9999 144.9961 0.00048271 4.8873 0.0056651
0.10883 0.98801 5.5249e-05 3.8182 0.012049 1.4349e-06 0.001154 0.042643 0.00065042 0.043289 0.0383 0 0.045357 0.0389 0 0.84604 0.22732 0.058907 0.0083502 4.1053 0.052635 6.2779e-05 0.83743 0.0051034 0.0058414 0.99687 2.9922e-10 0.22934 0.97563 0.99243 0.13044 0.79509 0.83306 0.76013 0.86655 0.55375 0.17225 0.42969 1.3124 0.64742 15.9999 144.9958 0.0004877 4.5244 0.0058082
0.10897 0.98801 5.5249e-05 3.8182 0.012049 1.4368e-06 0.001154 0.042665 0.00065043 0.043311 0.03832 0 0.045355 0.0389 0 0.84604 0.22732 0.058908 0.0083503 4.1053 0.052636 6.2779e-05 0.83743 0.0051034 0.0058414 0.99675 3.6725e-10 0.21994 0.97407 0.99194 0.13044 0.79105 0.8293 0.76134 0.86302 0.55191 0.17506 0.42966 1.2974 0.65598 15.9998 144.9956 0.00049249 4.176 0.0059513
0.10911 0.98801 5.5249e-05 3.8182 0.012049 1.4387e-06 0.001154 0.042687 0.00065044 0.043333 0.03834 0 0.045353 0.0389 0 0.84605 0.22732 0.058908 0.0083503 4.1053 0.052636 6.2779e-05 0.83743 0.0051034 0.0058414 0.99663 -1.2377e-10 0.21094 0.97247 0.99144 0.13044 0.78707 0.82555 0.76225 0.8595 0.5501 0.1778 0.42963 1.2829 0.66464 15.9998 144.9954 0.0004971 3.8404 0.0060945
0.10926 0.98801 5.5249e-05 3.8182 0.012049 1.4405e-06 0.001154 0.04271 0.00065044 0.043355 0.03836 0 0.045351 0.0389 0 0.84605 0.22732 0.058908 0.0083504 4.1053 0.052636 6.2779e-05 0.83743 0.0051034 0.0058414 0.9965 -2.6054e-10 0.20231 0.97084 0.99093 0.13044 0.78314 0.82179 0.76291 0.85599 0.54831 0.18048 0.4296 1.269 0.67337 15.9997 144.9952 0.00050152 3.5164 0.0062376
0.10954 0.98801 5.5249e-05 3.8182 0.012049 1.4443e-06 0.001154 0.042754 0.00065046 0.0434 0.038401 0 0.045347 0.0389 0 0.84605 0.22732 0.058909 0.0083504 4.1053 0.052636 6.278e-05 0.83743 0.0051034 0.0058414 0.99625 4.7945e-10 0.18612 0.96748 0.98987 0.13044 0.77546 0.81432 0.7635 0.84903 0.5448 0.18565 0.42954 1.2428 0.69091 15.9996 144.9947 0.00050984 2.8979 0.0065238
0.10983 0.98801 5.5249e-05 3.8182 0.012049 1.4481e-06 0.001154 0.042798 0.00065047 0.043444 0.038441 0 0.045343 0.0389 0 0.84606 0.22733 0.058909 0.0083505 4.1053 0.052636 6.278e-05 0.83743 0.0051034 0.0058414 0.996 1.5934e-09 0.17125 0.96399 0.98877 0.13044 0.76799 0.80688 0.76326 0.84212 0.5414 0.19059 0.42948 1.2186 0.70843 15.9996 144.9943 0.00051751 2.3122 0.0068101
0.11012 0.98801 5.5249e-05 3.8182 0.012049 1.4519e-06 0.001154 0.042842 0.00065048 0.043488 0.038481 0 0.045338 0.0389 0 0.84606 0.22733 0.05891 0.0083506 4.1053 0.052637 6.278e-05 0.83743 0.0051034 0.0058414 0.99575 1.0515e-09 0.1576 0.96037 0.98763 0.13044 0.76073 0.7995 0.7623 0.83527 0.53809 0.19532 0.42942 1.1963 0.72577 15.9995 144.9939 0.00052458 1.7522 0.0070963
0.1104 0.98801 5.5249e-05 3.8182 0.012049 1.4556e-06 0.001154 0.042887 0.0006505 0.043533 0.038521 0 0.045334 0.0389 0 0.84606 0.22733 0.058911 0.0083507 4.1053 0.052637 6.2781e-05 0.83743 0.0051034 0.0058414 0.99549 -2.3476e-10 0.14505 0.9566 0.98643 0.13044 0.75367 0.79219 0.76072 0.82848 0.53488 0.19985 0.42937 1.1759 0.74278 15.9994 144.9935 0.00053108 1.2122 0.0073825
0.11066 0.98801 5.5249e-05 3.8182 0.012049 1.459e-06 0.001154 0.042926 0.00065051 0.043572 0.038557 0 0.04533 0.0389 0 0.84607 0.22733 0.058911 0.0083507 4.1053 0.052637 6.2781e-05 0.83743 0.0051034 0.0058414 0.99524 -3.2872e-10 0.13463 0.95308 0.9853 0.13044 0.74749 0.78568 0.75883 0.82241 0.53206 0.20377 0.42931 1.159 0.75773 15.9993 144.9931 0.00053648 0.73955 0.0076402
0.11092 0.98801 5.5249e-05 3.8182 0.012049 1.4624e-06 0.001154 0.042966 0.00065052 0.043612 0.038593 0 0.045327 0.0389 0 0.84607 0.22733 0.058912 0.0083508 4.1053 0.052637 6.2781e-05 0.83743 0.0051034 0.0058414 0.99499 2.3291e-10 0.12498 0.94943 0.98412 0.13044 0.74145 0.77924 0.75654 0.81639 0.52932 0.20755 0.42926 1.1434 0.77226 15.9993 144.9928 0.0005415 0.27644 0.0078978
0.11115 0.98801 5.5249e-05 3.8182 0.012049 1.4655e-06 0.001154 0.043002 0.00065053 0.043648 0.038625 0 0.045323 0.0389 0 0.84607 0.22733 0.058912 0.0083509 4.1053 0.052637 6.2781e-05 0.83743 0.0051034 0.0058414 0.99476 2.5153e-10 0.1169 0.94602 0.983 0.13044 0.73615 0.77352 0.75417 0.81101 0.52692 0.21082 0.42921 1.1304 0.78494 15.9992 144.9924 0.0005457 -0.13426 0.0081296
0.11138 0.98801 5.5249e-05 3.8182 0.012049 1.4685e-06 0.001154 0.043038 0.00065054 0.043684 0.038658 0 0.04532 0.0389 0 0.84608 0.22733 0.058913 0.0083509 4.1053 0.052638 6.2782e-05 0.83743 0.0051034 0.0058414 0.99452 -1.0925e-10 0.10935 0.94249 0.98184 0.13044 0.73097 0.76786 0.75154 0.80566 0.52457 0.21399 0.42917 1.1184 0.7972 15.9991 144.9921 0.00054962 -0.54086 0.0083615
0.11161 0.98801 5.5249e-05 3.8182 0.012049 1.4716e-06 0.001154 0.043074 0.00065055 0.04372 0.03869 0 0.045317 0.0389 0 0.84608 0.22734 0.058913 0.008351 4.1053 0.052638 6.2782e-05 0.83742 0.0051034 0.0058414 0.99427 -1.7727e-10 0.1023 0.93883 0.98062 0.13044 0.7259 0.76228 0.74866 0.80035 0.52229 0.21705 0.42912 1.1073 0.80901 15.9991 144.9918 0.00055329 -0.94482 0.0085933
0.11185 0.98801 5.5249e-05 3.8182 0.012049 1.4747e-06 0.001154 0.043109 0.00065056 0.043755 0.038723 0 0.045313 0.0389 0 0.84608 0.22734 0.058914 0.0083511 4.1053 0.052638 6.2782e-05 0.83742 0.0051034 0.0058414 0.99401 6.2439e-11 0.095719 0.93502 0.97935 0.13044 0.72095 0.75679 0.74555 0.79508 0.52006 0.22001 0.42907 1.0971 0.82037 15.999 144.9915 0.00055672 -1.3475 0.0088252
0.11208 0.98801 5.5249e-05 3.8182 0.012049 1.4777e-06 0.001154 0.043145 0.00065057 0.043791 0.038755 0 0.04531 0.0389 0 0.84609 0.22734 0.058914 0.0083511 4.1053 0.052638 6.2782e-05 0.83742 0.0051034 0.0058414 0.99373 1.2603e-10 0.08957 0.93107 0.978 0.13044 0.71611 0.75137 0.74223 0.78984 0.51789 0.22287 0.42902 1.0876 0.83124 15.9989 144.9912 0.00055992 -1.7502 0.009057
0.11231 0.98801 5.5249e-05 3.8182 0.012049 1.4808e-06 0.001154 0.043181 0.00065058 0.043827 0.038788 0 0.045307 0.0389 0 0.84609 0.22734 0.058915 0.0083512 4.1053 0.052639 6.2783e-05 0.83742 0.0051035 0.0058414 0.99345 -4.7358e-11 0.083826 0.92695 0.97659 0.13044 0.71139 0.74605 0.7387 0.78464 0.51578 0.22562 0.42898 1.079 0.84163 15.9989 144.9909 0.00056292 -2.154 0.0092889
0.11254 0.98801 5.5249e-05 3.8182 0.012049 1.4838e-06 0.001154 0.043217 0.00065059 0.043863 0.03882 0 0.045303 0.0389 0 0.84609 0.22734 0.058915 0.0083512 4.1053 0.052639 6.2783e-05 0.83742 0.0051035 0.0058414 0.99314 -1.0014e-10 0.078461 0.92266 0.9751 0.13044 0.70678 0.74081 0.73498 0.77947 0.51373 0.22829 0.42893 1.071 0.85152 15.9988 144.9906 0.00056573 -2.5602 0.0095207
0.11277 0.98801 5.5249e-05 3.8182 0.012049 1.4869e-06 0.001154 0.043252 0.0006506 0.043898 0.038852 0 0.0453 0.0389 0 0.8461 0.22734 0.058916 0.0083513 4.1053 0.052639 6.2783e-05 0.83742 0.0051035 0.0058414 0.99283 3.9147e-11 0.073449 0.91818 0.97352 0.13044 0.70228 0.73567 0.73108 0.77434 0.51173 0.23085 0.42888 1.0637 0.86093 15.9988 144.9903 0.00056836 -2.9698 0.0097526
0.113 0.98801 5.5249e-05 3.8182 0.012049 1.4899e-06 0.001154 0.043288 0.00065061 0.043934 0.038885 0 0.045297 0.0389 0 0.8461 0.22734 0.058916 0.0083514 4.1053 0.052639 6.2783e-05 0.83742 0.0051035 0.0058414 0.99249 8.6615e-11 0.068767 0.91349 0.97185 0.13044 0.69789 0.73063 0.72701 0.76924 0.5098 0.23333 0.42883 1.057 0.86984 15.9987 144.9901 0.00057082 -3.384 0.0099845
0.11324 0.98801 5.5249e-05 3.8182 0.012049 1.493e-06 0.001154 0.043324 0.00065062 0.04397 0.038917 0 0.045293 0.0389 0 0.8461 0.22735 0.058917 0.0083514 4.1053 0.052639 6.2784e-05 0.83742 0.0051035 0.0058415 0.99213 -3.3529e-11 0.064393 0.90859 0.97008 0.13044 0.6936 0.72569 0.72276 0.76418 0.50792 0.23571 0.42879 1.0509 0.87828 15.9986 144.9898 0.00057312 -3.8039 0.010216
0.11347 0.98801 5.5249e-05 3.8182 0.012049 1.496e-06 0.001154 0.04336 0.00065063 0.044006 0.03895 0 0.04529 0.0389 0 0.8461 0.22735 0.058917 0.0083515 4.1053 0.05264 6.2784e-05 0.83742 0.0051035 0.0058415 0.99175 -7.9735e-11 0.060307 0.90344 0.96819 0.13044 0.68943 0.72086 0.71834 0.75915 0.5061 0.238 0.42874 1.0453 0.88624 15.9986 144.9895 0.00057529 -4.2307 0.010448
0.11393 0.98801 5.5249e-05 3.8182 0.012048 1.5022e-06 0.001154 0.043431 0.00065065 0.044077 0.039014 0 0.045283 0.0389 0 0.84611 0.22735 0.058918 0.0083516 4.1053 0.05264 6.2785e-05 0.83742 0.0051035 0.0058415 0.9909 -1.3597e-10 0.052922 0.89236 0.96405 0.13044 0.68141 0.71151 0.70901 0.74919 0.50264 0.24231 0.42865 1.0357 0.9008 15.9985 144.989 0.00057922 -5.1097 0.010912
0.1144 0.98801 5.5249e-05 3.8182 0.012048 1.5083e-06 0.001154 0.043503 0.00065067 0.044149 0.039079 0 0.045277 0.0389 0 0.84612 0.22735 0.058919 0.0083518 4.1053 0.05264 6.2785e-05 0.83742 0.0051035 0.0058415 0.98992 -1.1989e-09 0.046477 0.88007 0.95931 0.13044 0.67383 0.70263 0.69903 0.73937 0.49942 0.24626 0.42855 1.0277 0.91364 15.9983 144.9885 0.00058268 -6.0312 0.011376
0.11486 0.98801 5.5249e-05 3.8182 0.012048 1.5144e-06 0.001154 0.043574 0.00065069 0.04422 0.039144 0 0.04527 0.0389 0 0.84612 0.22736 0.05892 0.0083519 4.1053 0.052641 6.2786e-05 0.83742 0.0051035 0.0058415 0.98877 -1.6291e-09 0.040851 0.86637 0.95385 0.13044 0.66669 0.69423 0.68838 0.72969 0.49645 0.24986 0.42846 1.0213 0.92491 15.9982 144.988 0.00058573 -7.0067 0.011839
0.11532 0.98801 5.5249e-05 3.8182 0.012048 1.5205e-06 0.001154 0.043645 0.00065071 0.044292 0.039209 0 0.045263 0.0389 0 0.84613 0.22736 0.058921 0.008352 4.1053 0.052641 6.2786e-05 0.83742 0.0051035 0.0058415 0.98739 1.0797e-09 0.035942 0.85098 0.9475 0.13044 0.65999 0.68634 0.67705 0.72014 0.49371 0.25311 0.42836 1.0161 0.93475 15.9981 144.9875 0.00058841 -8.0491 0.012303
0.11579 0.98801 5.5249e-05 3.8182 0.012048 1.5266e-06 0.001154 0.043717 0.00065073 0.044363 0.039273 0 0.045257 0.0389 0 0.84614 0.22736 0.058922 0.0083522 4.1053 0.052642 6.2787e-05 0.83742 0.0051035 0.0058415 0.98571 3.3579e-09 0.031658 0.8336 0.94006 0.13044 0.65374 0.67898 0.665 0.71072 0.49123 0.25601 0.42827 1.0119 0.94332 15.998 144.9871 0.00059076 -9.1737 0.012767
0.11625 0.98801 5.5249e-05 3.8182 0.012048 1.5327e-06 0.001154 0.043788 0.00065075 0.044434 0.039338 0 0.04525 0.0389 0 0.84614 0.22736 0.058923 0.0083523 4.1053 0.052642 6.2787e-05 0.83742 0.0051035 0.0058415 0.98363 -1.0427e-09 0.027924 0.81385 0.93126 0.13044 0.64795 0.67219 0.6522 0.70145 0.489 0.25855 0.42817 1.0087 0.95077 15.9979 144.9867 0.00059281 -10.3978 0.01323
0.11671 0.98801 5.5249e-05 3.8182 0.012048 1.5388e-06 0.001154 0.043859 0.00065077 0.044506 0.039403 0 0.045243 0.0389 0 0.84615 0.22737 0.058925 0.0083524 4.1053 0.052643 6.2788e-05 0.83742 0.0051035 0.0058415 0.98099 -7.3722e-09 0.024671 0.79125 0.92076 0.13044 0.64263 0.66598 0.63861 0.6923 0.48703 0.26073 0.42808 1.0062 0.95723 15.9978 144.9863 0.00059456 -11.7419 0.013694
0.11718 0.98801 5.5249e-05 3.8182 0.012048 1.5449e-06 0.001154 0.043931 0.00065079 0.044577 0.039467 0 0.045237 0.0389 0 0.84616 0.22737 0.058926 0.0083525 4.1053 0.052643 6.2788e-05 0.83742 0.0051035 0.0058415 0.97756 -5.3876e-09 0.021842 0.76525 0.90813 0.13044 0.63779 0.6604 0.62418 0.6833 0.4853 0.26256 0.42798 1.0043 0.96285 15.9977 144.9859 0.00059604 -13.2292 0.014158
0.1176 0.98801 5.5249e-05 3.8182 0.012048 1.5504e-06 0.001154 0.043995 0.00065081 0.044641 0.039525 0 0.045231 0.0389 0 0.84616 0.22737 0.058926 0.0083527 4.1053 0.052644 6.2789e-05 0.83742 0.0051035 0.0058415 0.97354 1.0512e-09 0.019616 0.73838 0.89446 0.13044 0.63384 0.65591 0.61045 0.67533 0.48396 0.26389 0.4279 1.0031 0.96729 15.9976 144.9856 0.00059714 -14.7111 0.014575
0.11793 0.98801 5.5249e-05 3.8182 0.012048 1.5549e-06 0.001154 0.044047 0.00065082 0.044693 0.039573 0 0.045226 0.0389 0 0.84617 0.22737 0.058927 0.0083528 4.1053 0.052644 6.2789e-05 0.83742 0.0051035 0.0058415 0.96936 1.5716e-09 0.018009 0.71374 0.8814 0.13044 0.63093 0.65266 0.59878 0.66895 0.48302 0.26476 0.42783 1.0024 0.97052 15.9975 144.9853 0.00059787 -16.0279 0.014914
0.11827 0.98801 5.5249e-05 3.8182 0.012048 1.5594e-06 0.001154 0.044099 0.00065084 0.044745 0.03962 0 0.045221 0.0389 0 0.84617 0.22738 0.058928 0.0083529 4.1053 0.052644 6.279e-05 0.83742 0.0051035 0.0058415 0.96408 -1.8857e-09 0.016567 0.6862 0.86622 0.13044 0.62827 0.64977 0.58663 0.66265 0.4822 0.26545 0.42776 1.0019 0.97348 15.9975 144.9851 0.00059845 -17.4572 0.015253
0.11861 0.98801 5.5249e-05 3.8182 0.012048 1.5638e-06 0.001154 0.044151 0.00065085 0.044797 0.039667 0 0.045216 0.0389 0 0.84618 0.22738 0.058929 0.008353 4.1053 0.052644 6.279e-05 0.83742 0.0051035 0.0058415 0.95733 -2.5606e-09 0.015275 0.6554 0.84853 0.13044 0.62587 0.64723 0.57401 0.65645 0.4815 0.26595 0.42769 1.0015 0.97621 15.9974 144.9848 0.00059887 -19.0075 0.015592
0.11895 0.98801 5.5249e-05 3.8182 0.012048 1.5683e-06 0.001154 0.044203 0.00065086 0.044849 0.039714 0 0.045211 0.0389 0 0.84618 0.22738 0.05893 0.0083531 4.1053 0.052645 6.2791e-05 0.83742 0.0051035 0.0058415 0.9486 1.1368e-09 0.014123 0.62098 0.82787 0.13044 0.62371 0.64504 0.56093 0.65036 0.4809 0.26628 0.42762 1.0013 0.97878 15.9973 144.9846 0.00059913 -20.6839 0.01593
0.11926 0.98801 5.5249e-05 3.8182 0.012048 1.5723e-06 0.001154 0.04425 0.00065088 0.044896 0.039757 0 0.045207 0.0389 0 0.84619 0.22738 0.05893 0.0083531 4.1054 0.052645 6.2791e-05 0.83742 0.0051035 0.0058415 0.93852 2.4602e-09 0.013198 0.58664 0.80632 0.13044 0.62196 0.64336 0.54877 0.64499 0.48045 0.26643 0.42756 1.0013 0.98098 15.9973 144.9844 0.00059923 -22.3011 0.016235
0.11956 0.98801 5.5249e-05 3.8182 0.012048 1.5764e-06 0.001154 0.044296 0.00065089 0.044943 0.039799 0 0.045202 0.0389 0 0.84619 0.22739 0.058931 0.0083532 4.1054 0.052645 6.2791e-05 0.83742 0.0051035 0.0058415 0.9257 -3.3563e-09 0.01237 0.54892 0.78155 0.13044 0.6204 0.64194 0.53624 0.63973 0.48008 0.26645 0.4275 1.0014 0.98306 15.9972 144.9843 0.0005992 -24.0163 0.01654
0.11987 0.98801 5.5249e-05 3.8182 0.012048 1.5804e-06 0.001154 0.044343 0.0006509 0.04499 0.039841 0 0.045198 0.0389 0 0.8462 0.22739 0.058932 0.0083533 4.1054 0.052646 6.2792e-05 0.83742 0.0051035 0.0058415 0.90942 -1.0688e-08 0.011635 0.50779 0.75317 0.13044 0.61899 0.64076 0.52334 0.63462 0.47976 0.26635 0.42744 1.0016 0.98499 15.9972 144.9841 0.00059906 -25.8186 0.016845
0.12014 0.98801 5.5249e-05 3.8182 0.012048 1.584e-06 0.001154 0.044385 0.00065091 0.045032 0.03988 0 0.045194 0.0389 0 0.8462 0.22739 0.058932 0.0083534 4.1054 0.052646 6.2792e-05 0.83742 0.0051035 0.0058415 0.89117 -9.4227e-09 0.011047 0.46794 0.72424 0.13044 0.61785 0.63988 0.51139 0.63016 0.47953 0.26617 0.42738 1.0018 0.98658 15.9972 144.984 0.00059886 -27.5009 0.01712
0.12039 0.98801 5.5249e-05 3.8182 0.012048 1.5872e-06 0.001154 0.044423 0.00065092 0.045069 0.039914 0 0.045191 0.0389 0 0.8462 0.22739 0.058933 0.0083535 4.1054 0.052646 6.2792e-05 0.83742 0.0051035 0.0058415 0.87136 -3.2446e-09 0.010572 0.43004 0.6953 0.13044 0.61692 0.63922 0.50032 0.6263 0.47936 0.26593 0.42733 1.002 0.9879 15.9971 144.9839 0.00059863 -29.0489 0.017366
0.12063 0.98801 5.5249e-05 3.8182 0.012048 1.5905e-06 0.001154 0.044461 0.00065093 0.045107 0.039948 0 0.045187 0.0389 0 0.84621 0.22739 0.058933 0.0083535 4.1054 0.052647 6.2793e-05 0.83742 0.0051035 0.0058415 0.84795 -3.5814e-10 0.010147 0.39054 0.66351 0.13044 0.61607 0.63867 0.48891 0.62259 0.47921 0.26563 0.42728 1.0023 0.98915 15.9971 144.9838 0.00059834 -30.6127 0.017613
0.12083 0.98801 5.5249e-05 3.8182 0.012048 1.5931e-06 0.001154 0.044491 0.00065094 0.045138 0.039976 0 0.045184 0.0389 0 0.84621 0.22739 0.058934 0.0083536 4.1054 0.052647 6.2793e-05 0.83742 0.0051035 0.0058415 0.82647 -2.2243e-09 0.0098396 0.35813 0.63603 0.13044 0.61544 0.63829 0.4795 0.61977 0.47911 0.26533 0.42724 1.0026 0.99008 15.9971 144.9837 0.00059809 -31.8644 0.017811
0.12103 0.98801 5.5249e-05 3.8182 0.012048 1.5957e-06 0.001154 0.044522 0.00065095 0.045168 0.040003 0 0.045181 0.0389 0 0.84621 0.22739 0.058934 0.0083537 4.1054 0.052647 6.2793e-05 0.83742 0.0051035 0.0058415 0.80255 -3.8772e-09 0.009559 0.32536 0.60681 0.13044 0.61484 0.63796 0.46981 0.61709 0.47903 0.265 0.4272 1.0029 0.99098 15.997 144.9836 0.00059782 -33.1061 0.018009
0.12123 0.98801 5.5249e-05 3.8182 0.012048 1.5983e-06 0.001154 0.044552 0.00065096 0.045198 0.040031 0 0.045179 0.0389 0 0.84622 0.2274 0.058935 0.0083537 4.1054 0.052647 6.2794e-05 0.83742 0.0051035 0.0058415 0.7763 -3.1299e-09 0.0093032 0.29262 0.57598 0.13044 0.61429 0.63766 0.4598 0.61457 0.47896 0.26462 0.42716 1.0032 0.99183 15.997 144.9835 0.00059753 -34.3295 0.018207
0.1214 0.98801 5.5249e-05 3.8182 0.012048 1.6007e-06 0.001154 0.044579 0.00065097 0.045226 0.040055 0 0.045176 0.0389 0 0.84622 0.2274 0.058935 0.0083538 4.1054 0.052647 6.2794e-05 0.83742 0.0051035 0.0058415 0.75082 -1.9727e-09 0.0090927 0.26355 0.54699 0.13044 0.61382 0.63742 0.4505 0.61245 0.4789 0.26424 0.42713 1.0035 0.99256 15.997 144.9835 0.00059725 -35.4088 0.018385
0.12158 0.98801 5.5249e-05 3.8182 0.012048 1.603e-06 0.001154 0.044606 0.00065097 0.045253 0.04008 0 0.045174 0.0389 0 0.84622 0.2274 0.058936 0.0083538 4.1054 0.052647 6.2794e-05 0.83742 0.0051035 0.0058415 0.72379 -1.7754e-09 0.0088993 0.23518 0.51703 0.13044 0.61337 0.63721 0.4409 0.6105 0.47886 0.26382 0.42709 1.0038 0.99326 15.997 144.9834 0.00059697 -36.4628 0.018562
0.12176 0.98801 5.5249e-05 3.8182 0.012048 1.6054e-06 0.001154 0.044634 0.00065098 0.04528 0.040105 0 0.045171 0.0389 0 0.84622 0.2274 0.058936 0.0083539 4.1054 0.052648 6.2794e-05 0.83742 0.0051035 0.0058415 0.69549 -2.0703e-09 0.0087215 0.20783 0.48628 0.13044 0.61295 0.637 0.43098 0.60871 0.47882 0.26336 0.42706 1.0041 0.99394 15.9969 144.9833 0.00059669 -37.4878 0.01874
0.12194 0.98801 5.5249e-05 3.8182 0.012048 1.6077e-06 0.001154 0.044661 0.00065099 0.045307 0.040129 0 0.045169 0.0389 0 0.84623 0.2274 0.058936 0.0083539 4.1054 0.052648 6.2794e-05 0.83741 0.0051035 0.0058415 0.66624 -2.0029e-09 0.0085579 0.18182 0.45499 0.13044 0.61254 0.63682 0.42073 0.60709 0.47879 0.26286 0.42702 1.0044 0.9946 15.9969 144.9833 0.0005964 -38.4815 0.018918
0.1221 0.98801 5.5249e-05 3.8182 0.012048 1.6098e-06 0.001154 0.044685 0.00065099 0.045332 0.040152 0 0.045166 0.0389 0 0.84623 0.2274 0.058937 0.008354 4.1054 0.052648 6.2795e-05 0.83741 0.0051035 0.0058415 0.63938 -1.6458e-09 0.0084218 0.15977 0.42658 0.13044 0.6122 0.63666 0.41121 0.60579 0.47876 0.26237 0.42699 1.0047 0.99518 15.9969 144.9832 0.00059613 -39.3477 0.019079
0.12226 0.98801 5.5249e-05 3.8182 0.012048 1.6119e-06 0.001154 0.04471 0.000651 0.045356 0.040174 0 0.045164 0.0389 0 0.84623 0.2274 0.058937 0.008354 4.1054 0.052648 6.2795e-05 0.83741 0.0051035 0.0058415 0.61225 2.6144e-05 0.0083012 0.13918 0.39815 0.13044 0.61187 0.63651 0.4014 0.60464 0.47874 0.26185 0.42696 1.005 0.99573 15.9969 144.9832 0.00059586 -40.1866 0.019239
0.12238 0.98801 5.5249e-05 3.8182 0.012048 1.6135e-06 0.001154 0.044729 0.000651 0.045375 0.040191 0 0.045162 0.0389 0 0.84623 0.2274 0.058938 0.0083541 4.1054 0.052648 6.2795e-05 0.83741 0.0051035 0.0058415 0.59164 6.9416e-05 0.0082218 0.12461 0.37668 0.13044 0.61163 0.63641 0.39378 0.60386 0.47873 0.26143 0.42693 1.0052 0.99615 15.9969 144.9831 0.00059566 -40.8047 0.01936
0.1225 0.98801 5.5249e-05 3.8182 0.012048 1.6151e-06 0.001154 0.044747 0.00065101 0.045394 0.040208 0 0.045161 0.0389 0 0.84623 0.2274 0.058938 0.0083541 4.1054 0.052648 6.2795e-05 0.83741 0.0051036 0.0058415 0.57112 0.00012234 0.0081512 0.111 0.35541 0.13044 0.6114 0.63631 0.386 0.60316 0.47872 0.26098 0.42691 1.0055 0.99655 15.9969 144.9831 0.00059545 -41.4069 0.019482
0.12262 0.98801 5.5249e-05 3.8182 0.012048 1.6167e-06 0.001154 0.044766 0.00065101 0.045412 0.040224 0 0.045159 0.0389 0 0.84624 0.2274 0.058938 0.0083541 4.1054 0.052649 6.2795e-05 0.83741 0.0051036 0.0058415 0.55078 0.00017911 0.0080882 0.098354 0.33441 0.13044 0.61117 0.63622 0.37806 0.60253 0.47871 0.26051 0.42689 1.0057 0.99695 15.9969 144.9831 0.00059524 -41.9935 0.019603
0.12274 0.98801 5.5249e-05 3.8182 0.012048 1.6183e-06 0.001154 0.044784 0.00065102 0.045431 0.040241 0 0.045157 0.0389 0 0.84624 0.22741 0.058938 0.0083542 4.1054 0.052649 6.2796e-05 0.83741 0.0051036 0.0058415 0.53071 0.00023786 0.0080324 0.086699 0.31377 0.13044 0.61095 0.63614 0.36996 0.60199 0.4787 0.26002 0.42686 1.0059 0.99734 15.9969 144.983 0.00059504 -42.5645 0.019725
0.12287 0.98801 5.5249e-05 3.8182 0.012048 1.6199e-06 0.001154 0.044803 0.00065102 0.045449 0.040258 0 0.045155 0.0389 0 0.84624 0.22741 0.058939 0.0083542 4.1054 0.052649 6.2796e-05 0.83741 0.0051036 0.0058415 0.51098 0.00029984 0.0079837 0.076028 0.29356 0.13044 0.61074 0.63607 0.36173 0.60151 0.4787 0.25951 0.42684 1.0062 0.99773 15.9968 144.983 0.00059483 -43.1202 0.019846
0.12299 0.98801 5.5249e-05 3.8182 0.012048 1.6215e-06 0.001154 0.044821 0.00065103 0.045468 0.040275 0 0.045154 0.0389 0 0.84624 0.22741 0.058939 0.0083542 4.1054 0.052649 6.2796e-05 0.83741 0.0051036 0.0058415 0.49166 0.00036659 0.0079422 0.066326 0.27388 0.13044 0.61054 0.636 0.35335 0.60109 0.4787 0.25897 0.42681 1.0064 0.99811 15.9968 144.983 0.00059462 -43.6609 0.019968
0.12311 0.98801 5.5249e-05 3.8182 0.012048 1.6231e-06 0.001154 0.04484 0.00065103 0.045486 0.040292 0 0.045152 0.0389 0 0.84624 0.22741 0.058939 0.0083543 4.1054 0.052649 6.2796e-05 0.83741 0.0051036 0.0058415 0.47281 0.00043918 0.0079081 0.057566 0.25477 0.13044 0.61035 0.63595 0.34485 0.60074 0.47869 0.2584 0.42679 1.0067 0.99848 15.9968 144.983 0.00059441 -44.1867 0.020089
0.12323 0.98801 5.5249e-05 3.8182 0.012048 1.6247e-06 0.001154 0.044859 0.00065104 0.045505 0.040309 0 0.04515 0.0389 0 0.84625 0.22741 0.05894 0.0083543 4.1054 0.052649 6.2796e-05 0.83741 0.0051036 0.0058415 0.45448 0.0005179 0.0078812 0.049713 0.23631 0.13044 0.61016 0.6359 0.33623 0.60045 0.47869 0.25781 0.42677 1.0069 0.99885 15.9968 144.9829 0.0005942 -44.698 0.020211
0.12335 0.98801 5.5249e-05 3.8182 0.012048 1.6263e-06 0.001154 0.044877 0.00065104 0.045524 0.040326 0 0.045148 0.0389 0 0.84625 0.22741 0.05894 0.0083543 4.1054 0.052649 6.2796e-05 0.83741 0.0051036 0.0058415 0.43671 0.00060272 0.0078617 0.04272 0.21855 0.13044 0.60998 0.63587 0.3275 0.6002 0.47869 0.25719 0.42674 1.0072 0.99921 15.9968 144.9829 0.00059399 -45.195 0.020332
0.12347 0.98801 5.5249e-05 3.8182 0.012048 1.6279e-06 0.001154 0.044896 0.00065105 0.045542 0.040342 0 0.045147 0.0389 0 0.84625 0.22741 0.05894 0.0083544 4.1054 0.052649 6.2797e-05 0.83741 0.0051036 0.0058415 0.41954 0.00069371 0.0078492 0.036539 0.20153 0.13044 0.6098 0.63585 0.31869 0.60001 0.4787 0.25655 0.42672 1.0075 0.99957 15.9968 144.9829 0.00059377 -45.678 0.020453
0.1236 0.98801 5.5248e-05 3.8182 0.012048 1.6295e-06 0.001154 0.044914 0.00065105 0.045561 0.040359 0 0.045145 0.0389 0 0.84625 0.22741 0.05894 0.0083544 4.1054 0.05265 6.2797e-05 0.83741 0.0051036 0.0058416 0.40298 0.0007912 0.0078437 0.031111 0.18529 0.13044 0.60963 0.63584 0.30979 0.59985 0.4787 0.25587 0.4267 1.0077 0.99993 15.9968 144.9829 0.00059356 -46.1474 0.020575
0.12372 0.98801 5.5248e-05 3.8182 0.012048 1.6311e-06 0.001154 0.044933 0.00065106 0.045579 0.040376 0 0.045143 0.0389 0 0.84625 0.22741 0.058941 0.0083545 4.1054 0.05265 6.2797e-05 0.83741 0.0051036 0.0058416 0.38705 0.00089564 0.0078453 0.026379 0.16987 0.13044 0.60947 0.63584 0.30082 0.59974 0.4787 0.25517 0.42667 1.008 1.0003 15.9968 144.9828 0.00059335 -46.6033 0.020696
0.12384 0.98801 5.5248e-05 3.8182 0.012048 1.6327e-06 0.001154 0.044952 0.00065106 0.045598 0.040393 0 0.045141 0.0389 0 0.84625 0.22741 0.058941 0.0083545 4.1054 0.05265 6.2797e-05 0.83741 0.0051036 0.0058416 0.37177 0.0010074 0.0078538 0.02228 0.15527 0.13044 0.60931 0.63586 0.29181 0.59966 0.47871 0.25445 0.42665 1.0082 1.0006 15.9968 144.9828 0.00059313 -47.0461 0.020818
0.12396 0.98801 5.5248e-05 3.8182 0.012048 1.6343e-06 0.001154 0.04497 0.00065107 0.045617 0.04041 0 0.04514 0.0389 0 0.84626 0.22741 0.058941 0.0083545 4.1054 0.05265 6.2797e-05 0.83741 0.0051036 0.0058416 0.35713 0.0011267 0.0078693 0.018754 0.14152 0.13044 0.60916 0.63588 0.28277 0.59961 0.47871 0.25369 0.42662 1.0085 1.001 15.9968 144.9828 0.00059292 -47.476 0.020939
0.12408 0.98801 5.5248e-05 3.8182 0.012048 1.6359e-06 0.001154 0.044989 0.00065107 0.045635 0.040427 0 0.045138 0.0389 0 0.84626 0.22741 0.058942 0.0083546 4.1054 0.05265 6.2797e-05 0.83741 0.0051036 0.0058416 0.34314 0.0012538 0.0078916 0.01574 0.12863 0.13044 0.60901 0.63592 0.27371 0.59959 0.47872 0.2529 0.4266 1.0088 1.0013 15.9968 144.9828 0.00059271 -47.8935 0.021061
0.1242 0.98801 5.5248e-05 3.8182 0.012048 1.6375e-06 0.001154 0.045007 0.00065108 0.045654 0.040444 0 0.045136 0.0389 0 0.84626 0.22742 0.058942 0.0083546 4.1054 0.05265 6.2797e-05 0.83741 0.0051036 0.0058416 0.32978 0.0013888 0.0079207 0.01318 0.11658 0.13044 0.60887 0.63597 0.26466 0.59959 0.47872 0.25209 0.42658 1.009 1.0016 15.9968 144.9828 0.00059249 -48.2987 0.021182
0.12432 0.98801 5.5248e-05 3.8182 0.012048 1.6391e-06 0.001154 0.045026 0.00065108 0.045672 0.04046 0 0.045135 0.0389 0 0.84626 0.22742 0.058942 0.0083546 4.1054 0.05265 6.2798e-05 0.83741 0.0051036 0.0058416 0.31705 0.0015321 0.0079565 0.011019 0.10536 0.13044 0.60874 0.63604 0.25563 0.59961 0.47873 0.25125 0.42655 1.0093 1.002 15.9968 144.9827 0.00059228 -48.6919 0.021304
0.12445 0.98801 5.5248e-05 3.8182 0.012048 1.6407e-06 0.001154 0.045044 0.00065109 0.045691 0.040477 0 0.045133 0.0389 0 0.84626 0.22742 0.058942 0.0083547 4.1054 0.05265 6.2798e-05 0.83741 0.0051036 0.0058416 0.30493 0.0016838 0.007999 0.0092063 0.094972 0.13044 0.60861 0.63611 0.24664 0.59965 0.47874 0.25038 0.42653 1.0096 1.0023 15.9967 144.9827 0.00059206 -49.0736 0.021425
0.12457 0.98801 5.5248e-05 3.8182 0.012048 1.6423e-06 0.001154 0.045063 0.00065109 0.045709 0.040494 0 0.045131 0.0389 0 0.84627 0.22742 0.058943 0.0083547 4.1054 0.052651 6.2798e-05 0.83741 0.0051036 0.0058416 0.2934 0.0018443 0.0080482 0.0076929 0.085382 0.13044 0.60849 0.6362 0.2377 0.5997 0.47875 0.24948 0.42651 1.0098 1.0026 15.9967 144.9827 0.00059184 -49.4439 0.021547
0.12469 0.98801 5.5248e-05 3.8182 0.012048 1.644e-06 0.001154 0.045081 0.0006511 0.045728 0.040511 0 0.045129 0.0389 0 0.84627 0.22742 0.058943 0.0083548 4.1054 0.052651 6.2798e-05 0.83741 0.0051036 0.0058416 0.28244 0.0020136 0.0081039 0.0064364 0.076566 0.13044 0.60837 0.63629 0.22884 0.59978 0.47876 0.24855 0.42648 1.0101 1.003 15.9967 144.9827 0.00059163 -49.8032 0.021668
0.12481 0.98801 5.5248e-05 3.8182 0.012048 1.6456e-06 0.001154 0.0451 0.0006511 0.045747 0.040528 0 0.045128 0.0389 0 0.84627 0.22742 0.058943 0.0083548 4.1054 0.052651 6.2798e-05 0.83741 0.0051036 0.0058416 0.27204 0.002192 0.0081662 0.0053985 0.068492 0.13044 0.60825 0.6364 0.22007 0.59986 0.47877 0.2476 0.42646 1.0104 1.0033 15.9967 144.9827 0.00059141 -50.1519 0.02179
0.12493 0.98801 5.5248e-05 3.8182 0.012048 1.6472e-06 0.001154 0.045119 0.00065111 0.045765 0.040545 0 0.045126 0.0389 0 0.84627 0.22742 0.058944 0.0083548 4.1054 0.052651 6.2798e-05 0.83741 0.0051036 0.0058416 0.26216 0.0023797 0.0082349 0.004545 0.061128 0.13044 0.60814 0.63651 0.21141 0.59995 0.47878 0.24662 0.42644 1.0107 1.0036 15.9967 144.9826 0.00059119 -50.4901 0.021911
0.12505 0.98801 5.5248e-05 3.8182 0.012048 1.6488e-06 0.001154 0.045137 0.00065111 0.045784 0.040561 0 0.045124 0.0389 0 0.84627 0.22742 0.058944 0.0083549 4.1054 0.052651 6.2799e-05 0.83741 0.0051036 0.0058416 0.25279 0.0025769 0.00831 0.0038455 0.054435 0.13044 0.60804 0.63664 0.20287 0.60005 0.47879 0.2456 0.42641 1.0109 1.0039 15.9967 144.9826 0.00059097 -50.8184 0.022033
0.12517 0.98801 5.5248e-05 3.8182 0.012048 1.6504e-06 0.001154 0.045156 0.00065112 0.045802 0.040578 0 0.045123 0.0389 0 0.84627 0.22742 0.058944 0.0083549 4.1054 0.052651 6.2799e-05 0.83741 0.0051036 0.0058416 0.24391 0.0027836 0.0083914 0.0032741 0.048375 0.13044 0.60794 0.63677 0.19448 0.60016 0.4788 0.24456 0.42639 1.0112 1.0042 15.9967 144.9826 0.00059075 -51.1369 0.022154
0.1253 0.98801 5.5248e-05 3.8182 0.012048 1.652e-06 0.001154 0.045174 0.00065112 0.045821 0.040595 0 0.045121 0.0389 0 0.84628 0.22742 0.058944 0.0083549 4.1054 0.052651 6.2799e-05 0.83741 0.0051036 0.0058416 0.23548 0.0030001 0.0084792 0.0028078 0.042909 0.13044 0.60784 0.63691 0.18624 0.60028 0.47881 0.2435 0.42637 1.0115 1.0046 15.9967 144.9826 0.00059054 -51.4461 0.022276
0.12542 0.98801 5.5248e-05 3.8182 0.012048 1.6536e-06 0.001154 0.045193 0.00065113 0.045839 0.040612 0 0.045119 0.0389 0 0.84628 0.22742 0.058945 0.008355 4.1054 0.052651 6.2799e-05 0.83741 0.0051036 0.0058416 0.22748 0.0032265 0.0085731 0.002428 0.037995 0.13044 0.60775 0.63705 0.17816 0.6004 0.47882 0.2424 0.42635 1.0118 1.0049 15.9967 144.9826 0.00059032 -51.7461 0.022397
0.12554 0.98801 5.5248e-05 3.8182 0.012048 1.6552e-06 0.001154 0.045211 0.00065113 0.045858 0.040629 0 0.045117 0.0389 0 0.84628 0.22742 0.058945 0.008355 4.1054 0.052652 6.2799e-05 0.83741 0.0051036 0.0058416 0.2199 0.0034629 0.0086733 0.0021186 0.033594 0.13044 0.60766 0.63721 0.17027 0.60053 0.47883 0.24128 0.42632 1.012 1.0052 15.9967 144.9826 0.0005901 -52.0375 0.022519
0.12566 0.98801 5.5248e-05 3.8182 0.012048 1.6568e-06 0.001154 0.04523 0.00065113 0.045876 0.040645 0 0.045116 0.0389 0 0.84628 0.22742 0.058945 0.008355 4.1054 0.052652 6.2799e-05 0.83741 0.0051036 0.0058416 0.21271 0.0037094 0.0087795 0.0018663 0.029664 0.13044 0.60758 0.63736 0.16257 0.60066 0.47884 0.24014 0.4263 1.0123 1.0055 15.9967 144.9826 0.00058988 -52.3204 0.02264
0.12578 0.98801 5.5248e-05 3.8182 0.012048 1.6584e-06 0.001154 0.045248 0.00065114 0.045895 0.040662 0 0.045114 0.0389 0 0.84628 0.22743 0.058946 0.0083551 4.1054 0.052652 6.28e-05 0.83741 0.0051036 0.0058416 0.20588 0.0039661 0.0088918 0.00166 0.026167 0.13044 0.6075 0.63753 0.15507 0.6008 0.47885 0.23896 0.42628 1.0126 1.0058 15.9967 144.9826 0.00058966 -52.5952 0.022762
0.1259 0.98801 5.5248e-05 3.8182 0.012048 1.66e-06 0.001154 0.045267 0.00065114 0.045913 0.040679 0 0.045112 0.0389 0 0.84629 0.22743 0.058946 0.0083551 4.1054 0.052652 6.28e-05 0.83741 0.0051036 0.0058416 0.1994 0.0042332 0.00901 0.001491 0.023065 0.13044 0.60743 0.63769 0.14778 0.60093 0.47887 0.23777 0.42625 1.0129 1.0061 15.9967 144.9825 0.00058944 -52.8623 0.022883
0.12602 0.98801 5.5248e-05 3.8182 0.012048 1.6616e-06 0.001154 0.045285 0.00065115 0.045932 0.040696 0 0.04511 0.0389 0 0.84629 0.22743 0.058946 0.0083552 4.1054 0.052652 6.28e-05 0.83741 0.0051036 0.0058416 0.19325 0.0045107 0.0091342 0.001352 0.020322 0.13044 0.60736 0.63787 0.14071 0.60107 0.47888 0.23654 0.42623 1.0132 1.0064 15.9967 144.9825 0.00058922 -53.1219 0.023005
0.12615 0.98801 5.5248e-05 3.8182 0.012048 1.6632e-06 0.001154 0.045304 0.00065115 0.045951 0.040713 0 0.045109 0.0389 0 0.84629 0.22743 0.058946 0.0083552 4.1054 0.052652 6.28e-05 0.83741 0.0051036 0.0058416 0.1874 0.0047987 0.0092643 0.0012367 0.017903 0.13044 0.60729 0.63804 0.13387 0.60122 0.47889 0.2353 0.42621 1.0134 1.0067 15.9967 144.9825 0.000589 -53.3743 0.023126
0.12627 0.98801 5.5248e-05 3.8182 0.012048 1.6648e-06 0.001154 0.045323 0.00065116 0.045969 0.04073 0 0.045107 0.0389 0 0.84629 0.22743 0.058947 0.0083552 4.1054 0.052652 6.28e-05 0.83741 0.0051036 0.0058416 0.18184 0.0050973 0.0094002 0.0011402 0.015776 0.13044 0.60722 0.63822 0.12725 0.60136 0.4789 0.23403 0.42619 1.0137 1.007 15.9967 144.9825 0.00058878 -53.62 0.023248
0.12639 0.98801 5.5248e-05 3.8182 0.012048 1.6664e-06 0.001154 0.045341 0.00065116 0.045988 0.040746 0 0.045105 0.0389 0 0.84629 0.22743 0.058947 0.0083553 4.1054 0.052653 6.28e-05 0.83741 0.0051036 0.0058416 0.17655 0.0054065 0.0095418 0.0010586 0.01391 0.13044 0.60716 0.6384 0.12087 0.60151 0.47892 0.23273 0.42616 1.014 1.0073 15.9967 144.9825 0.00058856 -53.859 0.023369
0.12651 0.98801 5.5248e-05 3.8182 0.012048 1.668e-06 0.001154 0.04536 0.00065117 0.046006 0.040763 0 0.045104 0.0389 0 0.84629 0.22743 0.058947 0.0083553 4.1054 0.052653 6.2801e-05 0.83741 0.0051036 0.0058416 0.17151 0.0057265 0.0096892 0.00098895 0.012277 0.13044 0.60711 0.63858 0.11472 0.60165 0.47893 0.23142 0.42614 1.0143 1.0076 15.9967 144.9825 0.00058833 -54.0919 0.02349
0.12663 0.98801 5.5248e-05 3.8182 0.012048 1.6696e-06 0.001154 0.045378 0.00065117 0.046025 0.04078 0 0.045102 0.0389 0 0.8463 0.22743 0.058948 0.0083553 4.1054 0.052653 6.2801e-05 0.83741 0.0051036 0.0058416 0.16671 0.0060572 0.0098422 0.00092873 0.010852 0.13044 0.60705 0.63877 0.10881 0.6018 0.47894 0.23008 0.42612 1.0146 1.0079 15.9967 144.9825 0.00058811 -54.3188 0.023612
0.12675 0.98801 5.5248e-05 3.8182 0.012048 1.6712e-06 0.001154 0.045397 0.00065118 0.046043 0.040797 0 0.0451 0.0389 0 0.8463 0.22743 0.058948 0.0083554 4.1054 0.052653 6.2801e-05 0.83741 0.0051036 0.0058416 0.16213 0.0063988 0.010001 0.00087622 0.0096097 0.13044 0.607 0.63895 0.10314 0.60195 0.47895 0.22872 0.4261 1.0148 1.0082 15.9967 144.9825 0.00058789 -54.5401 0.023733
0.12688 0.98801 5.5248e-05 3.8182 0.012048 1.6728e-06 0.001154 0.045415 0.00065118 0.046062 0.040814 0 0.045098 0.0389 0 0.8463 0.22743 0.058948 0.0083554 4.1054 0.052653 6.2801e-05 0.83741 0.0051036 0.0058416 0.15776 0.0067513 0.010165 0.00082995 0.0085292 0.13044 0.60695 0.63914 0.097711 0.6021 0.47897 0.22734 0.42607 1.0151 1.0085 15.9967 144.9825 0.00058767 -54.756 0.023855
0.127 0.98801 5.5248e-05 3.8182 0.012048 1.6744e-06 0.001154 0.045434 0.00065119 0.04608 0.04083 0 0.045097 0.0389 0 0.8463 0.22743 0.058949 0.0083555 4.1054 0.052653 6.2801e-05 0.83741 0.0051036 0.0058416 0.15359 0.0071147 0.010335 0.00078894 0.0075911 0.13044 0.60691 0.63933 0.092516 0.60225 0.47898 0.22593 0.42605 1.0154 1.0088 15.9967 144.9825 0.00058745 -54.9667 0.023976
0.12712 0.98801 5.5248e-05 3.8182 0.012048 1.676e-06 0.001154 0.045452 0.00065119 0.046099 0.040847 0 0.045095 0.0389 0 0.8463 0.22743 0.058949 0.0083555 4.1054 0.052653 6.2801e-05 0.83741 0.0051036 0.0058416 0.1496 0.0074892 0.01051 0.00075228 0.0067778 0.13044 0.60686 0.63952 0.087556 0.6024 0.479 0.22451 0.42603 1.0157 1.0091 15.9967 144.9825 0.00058723 -55.1727 0.024098
0.12724 0.98801 5.5248e-05 3.8182 0.012048 1.6776e-06 0.001154 0.045471 0.0006512 0.046117 0.040864 0 0.045093 0.0389 0 0.84631 0.22744 0.058949 0.0083555 4.1054 0.052653 6.2802e-05 0.83741 0.0051036 0.0058416 0.14578 0.0078747 0.010691 0.00071917 0.0060734 0.13044 0.60682 0.63972 0.082827 0.60255 0.47901 0.22307 0.42601 1.016 1.0094 15.9966 144.9825 0.000587 -55.374 0.024219
0.12736 0.98801 5.5248e-05 3.8182 0.012048 1.6792e-06 0.001154 0.045489 0.0006512 0.046136 0.040881 0 0.045092 0.0389 0 0.84631 0.22744 0.058949 0.0083556 4.1054 0.052654 6.2802e-05 0.83741 0.0051036 0.0058416 0.14211 0.0082714 0.010877 0.00068898 0.0054639 0.13044 0.60679 0.63991 0.078326 0.6027 0.47902 0.22161 0.42599 1.0163 1.0097 15.9966 144.9825 0.00058678 -55.5709 0.024341
0.12748 0.98801 5.5248e-05 3.8182 0.012048 1.6808e-06 0.001154 0.045508 0.00065121 0.046154 0.040898 0 0.04509 0.0389 0 0.84631 0.22744 0.05895 0.0083556 4.1054 0.052654 6.2802e-05 0.83741 0.0051036 0.0058416 0.1386 0.0086793 0.011068 0.00066132 0.0049368 0.13044 0.60675 0.6401 0.074047 0.60285 0.47904 0.22013 0.42596 1.0165 1.01 15.9966 144.9824 0.00058656 -55.7638 0.024462
0.1276 0.98801 5.5248e-05 3.8182 0.012048 1.6824e-06 0.001154 0.045526 0.00065121 0.046173 0.040914 0 0.045088 0.0389 0 0.84631 0.22744 0.05895 0.0083556 4.1054 0.052654 6.2802e-05 0.83741 0.0051036 0.0058416 0.13523 0.0090985 0.011265 0.00063577 0.0044808 0.13044 0.60672 0.64029 0.069987 0.603 0.47905 0.21864 0.42594 1.0168 1.0103 15.9966 144.9824 0.00058634 -55.9528 0.024584
0.12773 0.98801 5.5248e-05 3.8182 0.012048 1.684e-06 0.001154 0.045545 0.00065121 0.046191 0.040931 0 0.045086 0.0389 0 0.84631 0.22744 0.05895 0.0083557 4.1054 0.052654 6.2802e-05 0.83741 0.0051036 0.0058416 0.132 0.0095289 0.011467 0.00061206 0.0040862 0.13044 0.60669 0.64049 0.066139 0.60314 0.47906 0.21713 0.42592 1.0171 1.0106 15.9966 144.9824 0.00058611 -56.138 0.024705
0.12785 0.98801 5.5248e-05 3.8182 0.012048 1.6856e-06 0.001154 0.045563 0.00065122 0.04621 0.040948 0 0.045085 0.0389 0 0.84632 0.22744 0.058951 0.0083557 4.1054 0.052654 6.2802e-05 0.83741 0.0051036 0.0058416 0.12888 0.0099708 0.011674 0.00058993 0.0037442 0.13044 0.60667 0.64068 0.062498 0.60329 0.47908 0.2156 0.4259 1.0174 1.0109 15.9966 144.9824 0.00058589 -56.3199 0.024827
0.12797 0.98801 5.5248e-05 3.8182 0.012048 1.6872e-06 0.001154 0.045582 0.00065122 0.046228 0.040965 0 0.045083 0.0389 0 0.84632 0.22744 0.058951 0.0083558 4.1054 0.052654 6.2803e-05 0.83741 0.0051036 0.0058416 0.12589 0.010424 0.011887 0.00056921 0.0034474 0.13044 0.60664 0.64088 0.059057 0.60344 0.47909 0.21405 0.42588 1.0177 1.0112 15.9966 144.9824 0.00058567 -56.4984 0.024948
0.12809 0.98801 5.5248e-05 3.8182 0.012048 1.6888e-06 0.001154 0.0456 0.00065123 0.046247 0.040982 0 0.045081 0.0389 0 0.84632 0.22744 0.058951 0.0083558 4.1054 0.052654 6.2803e-05 0.83741 0.0051036 0.0058416 0.123 0.010889 0.012105 0.00054975 0.0031896 0.13044 0.60662 0.64107 0.055809 0.60359 0.47911 0.21249 0.42585 1.018 1.0115 15.9966 144.9824 0.00058544 -56.6739 0.02507
0.12821 0.98801 5.5248e-05 3.8182 0.012048 1.6904e-06 0.001154 0.045619 0.00065123 0.046265 0.040998 0 0.04508 0.0389 0 0.84632 0.22744 0.058952 0.0083558 4.1054 0.052655 6.2803e-05 0.83741 0.0051036 0.0058416 0.12021 0.011366 0.012328 0.00053142 0.002965 0.13044 0.6066 0.64127 0.052748 0.60374 0.47912 0.21092 0.42583 1.0182 1.0118 15.9966 144.9824 0.00058522 -56.8465 0.025191
0.12833 0.98801 5.5248e-05 3.8182 0.012048 1.692e-06 0.001154 0.045637 0.00065124 0.046284 0.041015 0 0.045078 0.0389 0 0.84632 0.22744 0.058952 0.0083559 4.1054 0.052655 6.2803e-05 0.83741 0.0051036 0.0058416 0.11752 0.011854 0.012556 0.00051411 0.002769 0.13044 0.60658 0.64146 0.049866 0.60388 0.47914 0.20933 0.42581 1.0185 1.0121 15.9966 144.9824 0.000585 -57.0164 0.025313
0.12845 0.98801 5.5248e-05 3.8182 0.012048 1.6936e-06 0.001154 0.045656 0.00065124 0.046303 0.041032 0 0.045076 0.0389 0 0.84632 0.22744 0.058952 0.0083559 4.1054 0.052655 6.2803e-05 0.83741 0.0051036 0.0058416 0.11493 0.012354 0.01279 0.00049771 0.0025971 0.13044 0.60657 0.64166 0.047156 0.60403 0.47915 0.20772 0.42579 1.0188 1.0124 15.9966 144.9824 0.00058477 -57.1837 0.025434
0.1287 0.98801 5.5248e-05 3.8182 0.012048 1.6968e-06 0.001154 0.045693 0.00065125 0.04634 0.041066 0 0.045073 0.0389 0 0.84633 0.22745 0.058953 0.008356 4.1054 0.052655 6.2804e-05 0.83741 0.0051036 0.0058416 0.10998 0.01339 0.013272 0.00046737 0.0023132 0.13044 0.60655 0.64205 0.042223 0.60432 0.47918 0.20447 0.42574 1.0194 1.013 15.9966 144.9824 0.00058432 -57.5112 0.025677
0.12892 0.98801 5.5248e-05 3.8182 0.012048 1.6997e-06 0.001154 0.045726 0.00065126 0.046373 0.041096 0 0.04507 0.0389 0 0.84633 0.22745 0.058953 0.008356 4.1054 0.052655 6.2804e-05 0.83741 0.0051036 0.0058416 0.1058 0.014364 0.013725 0.00044247 0.0021098 0.13044 0.60653 0.6424 0.038299 0.60458 0.4792 0.20151 0.42571 1.0199 1.0135 15.9966 144.9824 0.00058392 -57.7987 0.025896
0.12913 0.98801 5.5248e-05 3.8182 0.012048 1.7026e-06 0.001154 0.045759 0.00065127 0.046406 0.041126 0 0.045066 0.0389 0 0.84633 0.22745 0.058954 0.0083561 4.1054 0.052656 6.2804e-05 0.83741 0.0051036 0.0058416 0.10183 0.015377 0.014194 0.00041954 0.0019428 0.13044 0.60653 0.64275 0.03482 0.60484 0.47923 0.1985 0.42567 1.0204 1.014 15.9966 144.9824 0.00058352 -58.0801 0.026114
0.12935 0.98801 5.5248e-05 3.8182 0.012048 1.7054e-06 0.001154 0.045793 0.00065128 0.046439 0.041156 0 0.045063 0.0389 0 0.84634 0.22745 0.058954 0.0083562 4.1054 0.052656 6.2805e-05 0.83741 0.0051036 0.0058416 0.098074 0.016432 0.01468 0.00039834 0.0018032 0.13044 0.60653 0.6431 0.031744 0.60509 0.47926 0.19546 0.42563 1.0209 1.0146 15.9966 144.9824 0.00058311 -58.356 0.026333
0.12957 0.98801 5.5248e-05 3.8182 0.012048 1.7083e-06 0.001154 0.045826 0.00065129 0.046473 0.041186 0 0.04506 0.0389 0 0.84634 0.22745 0.058955 0.0083563 4.1054 0.052656 6.2805e-05 0.83741 0.0051036 0.0058416 0.094498 0.017528 0.015183 0.00037866 0.0016843 0.13044 0.60653 0.64345 0.029032 0.60535 0.47928 0.19239 0.42559 1.0214 1.0151 15.9966 144.9824 0.00058271 -58.6271 0.026552
0.12979 0.98801 5.5248e-05 3.8182 0.012048 1.7112e-06 0.001154 0.045859 0.00065129 0.046506 0.041217 0 0.045057 0.0389 0 0.84635 0.22745 0.058955 0.0083563 4.1054 0.052656 6.2805e-05 0.83741 0.0051036 0.0058416 0.091092 0.018666 0.015704 0.00036032 0.0015812 0.13044 0.60654 0.6438 0.026646 0.6056 0.47931 0.18928 0.42555 1.0219 1.0156 15.9966 144.9824 0.00058231 -58.8938 0.02677
0.13001 0.98801 5.5248e-05 3.8182 0.012048 1.7141e-06 0.001154 0.045893 0.0006513 0.046539 0.041247 0 0.045054 0.0389 0 0.84635 0.22745 0.058956 0.0083564 4.1054 0.052657 6.2806e-05 0.83741 0.0051036 0.0058416 0.08784 0.019848 0.016242 0.00034318 0.0014902 0.13044 0.60656 0.64415 0.024551 0.60585 0.47934 0.18615 0.42551 1.0225 1.0161 15.9966 144.9824 0.0005819 -59.1567 0.026989
0.13023 0.98801 5.5248e-05 3.8182 0.012048 1.717e-06 0.001154 0.045926 0.00065131 0.046573 0.041277 0 0.045051 0.0389 0 0.84635 0.22746 0.058956 0.0083565 4.1054 0.052657 6.2806e-05 0.83741 0.0051036 0.0058416 0.084732 0.021075 0.016797 0.00032712 0.0014088 0.13044 0.60658 0.6445 0.022715 0.6061 0.47936 0.18299 0.42548 1.023 1.0167 15.9966 144.9824 0.0005815 -59.4162 0.027208
0.13045 0.98801 5.5248e-05 3.8182 0.012048 1.7199e-06 0.001154 0.045959 0.00065132 0.046606 0.041307 0 0.045048 0.0389 0 0.84636 0.22746 0.058957 0.0083565 4.1054 0.052657 6.2806e-05 0.83741 0.0051036 0.0058416 0.081756 0.022346 0.01737 0.00031203 0.0013352 0.13044 0.60661 0.64485 0.021106 0.60635 0.47939 0.17981 0.42544 1.0235 1.0172 15.9966 144.9824 0.00058109 -59.6726 0.027426
0.13067 0.98801 5.5248e-05 3.8182 0.012048 1.7227e-06 0.001154 0.045992 0.00065133 0.046639 0.041337 0 0.045045 0.0389 0 0.84636 0.22746 0.058958 0.0083566 4.1054 0.052657 6.2806e-05 0.83741 0.0051036 0.0058416 0.078904 0.023665 0.017961 0.00029784 0.001268 0.13044 0.60665 0.6452 0.019697 0.60659 0.47942 0.1766 0.4254 1.024 1.0177 15.9966 144.9823 0.00058069 -59.9262 0.027645
0.13088 0.98801 5.5248e-05 3.8182 0.012048 1.7256e-06 0.001154 0.046026 0.00065133 0.046672 0.041367 0 0.045042 0.0389 0 0.84636 0.22746 0.058958 0.0083567 4.1054 0.052658 6.2807e-05 0.83741 0.0051036 0.0058416 0.076168 0.025031 0.018571 0.00028445 0.0012063 0.13044 0.60669 0.64554 0.018464 0.60683 0.47945 0.17338 0.42536 1.0245 1.0182 15.9966 144.9823 0.00058028 -60.1772 0.027864
0.1311 0.98801 5.5248e-05 3.8182 0.012048 1.7285e-06 0.001154 0.046059 0.00065134 0.046706 0.041398 0 0.045039 0.0389 0 0.84637 0.22746 0.058959 0.0083567 4.1054 0.052658 6.2807e-05 0.83741 0.0051036 0.0058416 0.07354 0.026447 0.019198 0.00027181 0.001149 0.13044 0.60673 0.64589 0.017383 0.60707 0.47947 0.17013 0.42533 1.025 1.0187 15.9966 144.9823 0.00057988 -60.4261 0.028082
0.13132 0.98801 5.5248e-05 3.8182 0.012048 1.7314e-06 0.001154 0.046092 0.00065135 0.046739 0.041428 0 0.045036 0.0389 0 0.84637 0.22746 0.058959 0.0083568 4.1054 0.052658 6.2807e-05 0.8374 0.0051036 0.0058416 0.071015 0.027913 0.019845 0.00025984 0.0010955 0.13044 0.60678 0.64624 0.016435 0.60731 0.4795 0.16688 0.42529 1.0255 1.0193 15.9966 144.9823 0.00057947 -60.6728 0.028301
0.13154 0.98801 5.5248e-05 3.8182 0.012048 1.7343e-06 0.001154 0.046125 0.00065136 0.046772 0.041458 0 0.045033 0.0389 0 0.84637 0.22747 0.05896 0.0083569 4.1054 0.052658 6.2808e-05 0.8374 0.0051036 0.0058416 0.068586 0.029431 0.02051 0.00024851 0.0010454 0.13044 0.60684 0.64658 0.015601 0.60755 0.47953 0.1636 0.42525 1.0261 1.0198 15.9966 144.9823 0.00057907 -60.9176 0.02852
0.13176 0.98801 5.5248e-05 3.8182 0.012048 1.7371e-06 0.001154 0.046158 0.00065137 0.046805 0.041488 0 0.04503 0.0389 0 0.84638 0.22747 0.05896 0.0083569 4.1054 0.052659 6.2808e-05 0.8374 0.0051037 0.0058416 0.066248 0.031002 0.021194 0.00023776 0.00099827 0.13044 0.60689 0.64693 0.014866 0.60778 0.47955 0.16032 0.42521 1.0266 1.0203 15.9966 144.9823 0.00057866 -61.1607 0.028738
0.13198 0.98801 5.5248e-05 3.8182 0.012048 1.74e-06 0.001154 0.046192 0.00065138 0.046838 0.041518 0 0.045026 0.0389 0 0.84638 0.22747 0.058961 0.008357 4.1054 0.052659 6.2808e-05 0.8374 0.0051037 0.0058416 0.063997 0.032627 0.021898 0.00022756 0.00095381 0.13044 0.60696 0.64727 0.014215 0.60801 0.47958 0.15703 0.42518 1.0271 1.0208 15.9966 144.9823 0.00057825 -61.4022 0.028957
0.1322 0.98801 5.5248e-05 3.8182 0.012048 1.7429e-06 0.001154 0.046225 0.00065138 0.046872 0.041548 0 0.045023 0.0389 0 0.84638 0.22747 0.058961 0.0083571 4.1055 0.052659 6.2809e-05 0.8374 0.0051037 0.0058416 0.06183 0.034309 0.022622 0.00021787 0.00091179 0.13044 0.60703 0.64762 0.013636 0.60824 0.47961 0.15373 0.42514 1.0276 1.0213 15.9966 144.9823 0.00057785 -61.6421 0.029176
0.13241 0.98801 5.5248e-05 3.8182 0.012048 1.7458e-06 0.001154 0.046258 0.00065139 0.046905 0.041578 0 0.04502 0.0389 0 0.84639 0.22747 0.058962 0.0083571 4.1055 0.052659 6.2809e-05 0.8374 0.0051037 0.0058416 0.059741 0.036049 0.023367 0.00020865 0.00087201 0.13044 0.6071 0.64796 0.013118 0.60847 0.47964 0.15043 0.4251 1.0281 1.0219 15.9966 144.9823 0.00057744 -61.8806 0.029394
0.13263 0.98801 5.5248e-05 3.8182 0.012048 1.7487e-06 0.001154 0.046291 0.0006514 0.046938 0.041608 0 0.045017 0.0389 0 0.84639 0.22747 0.058963 0.0083572 4.1055 0.05266 6.2809e-05 0.8374 0.0051037 0.0058416 0.057728 0.037848 0.024132 0.00019988 0.00083428 0.13044 0.60718 0.6483 0.012653 0.6087 0.47967 0.14712 0.42507 1.0286 1.0224 15.9966 144.9823 0.00057703 -62.1178 0.029613
0.13285 0.98801 5.5248e-05 3.8182 0.012048 1.7516e-06 0.001154 0.046324 0.00065141 0.046971 0.041639 0 0.045014 0.0389 0 0.84639 0.22747 0.058963 0.0083573 4.1055 0.05266 6.281e-05 0.8374 0.0051037 0.0058417 0.055788 0.039707 0.024917 0.00019153 0.00079846 0.13044 0.60726 0.64864 0.012232 0.60893 0.47969 0.14382 0.42503 1.0291 1.0229 15.9966 144.9823 0.00057663 -62.3536 0.029832
0.13307 0.98801 5.5248e-05 3.8182 0.012048 1.7544e-06 0.001154 0.046358 0.00065142 0.047004 0.041669 0 0.045011 0.0389 0 0.8464 0.22748 0.058964 0.0083574 4.1055 0.05266 6.281e-05 0.8374 0.0051037 0.0058417 0.053915 0.04163 0.025725 0.00018357 0.00076443 0.13044 0.60735 0.64899 0.011849 0.60915 0.47972 0.14052 0.425 1.0297 1.0234 15.9966 144.9823 0.00057622 -62.5882 0.03005
0.13329 0.98801 5.5248e-05 3.8182 0.012048 1.7573e-06 0.001154 0.046391 0.00065142 0.047038 0.041699 0 0.045008 0.0389 0 0.8464 0.22748 0.058964 0.0083574 4.1055 0.05266 6.281e-05 0.8374 0.0051037 0.0058417 0.052109 0.043616 0.026553 0.00017599 0.00073207 0.13044 0.60744 0.64933 0.011497 0.60937 0.47975 0.13722 0.42496 1.0302 1.0239 15.9966 144.9823 0.00057581 -62.8216 0.030269
0.13351 0.98801 5.5248e-05 3.8182 0.012048 1.7602e-06 0.001154 0.046424 0.00065143 0.047071 0.041729 0 0.045005 0.0389 0 0.8464 0.22748 0.058965 0.0083575 4.1055 0.052661 6.2811e-05 0.8374 0.0051037 0.0058417 0.05037 0.045669 0.027404 0.00016876 0.00070127 0.13044 0.60753 0.64967 0.011172 0.60959 0.47978 0.13392 0.42493 1.0307 1.0245 15.9966 144.9823 0.00057541 -63.0538 0.030488
0.13373 0.98801 5.5248e-05 3.8182 0.012048 1.7631e-06 0.001154 0.046457 0.00065144 0.047104 0.041759 0 0.045002 0.0389 0 0.84641 0.22748 0.058965 0.0083576 4.1055 0.052661 6.2811e-05 0.8374 0.0051037 0.0058417 0.048688 0.047789 0.028278 0.00016186 0.00067194 0.13044 0.60763 0.65001 0.010869 0.60981 0.4798 0.13064 0.42489 1.0312 1.025 15.9966 144.9823 0.000575 -63.285 0.030706
0.13395 0.98801 5.5248e-05 3.8182 0.012048 1.766e-06 0.001154 0.04649 0.00065145 0.047137 0.041789 0 0.044999 0.0389 0 0.84641 0.22748 0.058966 0.0083576 4.1055 0.052661 6.2811e-05 0.8374 0.0051037 0.0058417 0.047072 0.049979 0.029174 0.00015528 0.00064401 0.13044 0.60774 0.65035 0.010587 0.61003 0.47983 0.12737 0.42486 1.0317 1.0255 15.9966 144.9823 0.00057459 -63.5149 0.030925
0.13416 0.98801 5.5248e-05 3.8182 0.012048 1.7689e-06 0.001154 0.046523 0.00065146 0.04717 0.041819 0 0.044996 0.0389 0 0.84641 0.22748 0.058966 0.0083577 4.1055 0.052661 6.2812e-05 0.8374 0.0051037 0.0058417 0.045509 0.052241 0.030094 0.000149 0.00061741 0.13044 0.60784 0.65069 0.010322 0.61025 0.47986 0.12411 0.42482 1.0322 1.026 15.9966 144.9823 0.00057419 -63.7439 0.031144
0.13436 0.98801 5.5248e-05 3.8182 0.012048 1.7714e-06 0.001154 0.046553 0.00065146 0.0472 0.041846 0 0.044993 0.0389 0 0.84642 0.22748 0.058967 0.0083578 4.1055 0.052662 6.2812e-05 0.8374 0.0051037 0.0058417 0.044151 0.054334 0.03094 0.00014361 0.0005946 0.13044 0.60794 0.65099 0.010097 0.61044 0.47988 0.1212 0.42479 1.0327 1.0265 15.9966 144.9823 0.00057382 -63.9485 0.03134
0.13456 0.98801 5.5248e-05 3.8182 0.012048 1.774e-06 0.001154 0.046583 0.00065147 0.04723 0.041873 0 0.04499 0.0389 0 0.84642 0.22749 0.058967 0.0083578 4.1055 0.052662 6.2812e-05 0.8374 0.0051037 0.0058417 0.042838 0.056487 0.031805 0.00013843 0.00057273 0.13044 0.60804 0.65129 0.009882 0.61063 0.47991 0.1183 0.42476 1.0331 1.0269 15.9966 144.9822 0.00057345 -64.1523 0.031537
0.13475 0.98801 5.5248e-05 3.8182 0.012048 1.7766e-06 0.001154 0.046613 0.00065148 0.04726 0.0419 0 0.044988 0.0389 0 0.84642 0.22749 0.058968 0.0083579 4.1055 0.052662 6.2812e-05 0.8374 0.0051037 0.0058417 0.041565 0.058701 0.032691 0.00013347 0.00055177 0.13044 0.60815 0.6516 0.0096766 0.61083 0.47993 0.11541 0.42473 1.0336 1.0274 15.9966 144.9822 0.00057309 -64.3552 0.031733
0.13495 0.98801 5.5248e-05 3.8182 0.012048 1.7792e-06 0.001154 0.046642 0.00065148 0.047289 0.041927 0 0.044985 0.0389 0 0.84643 0.22749 0.058968 0.008358 4.1055 0.052662 6.2813e-05 0.8374 0.0051037 0.0058417 0.040333 0.060979 0.033596 0.0001287 0.00053169 0.13044 0.60826 0.6519 0.0094795 0.61102 0.47996 0.11254 0.4247 1.0341 1.0279 15.9967 144.9822 0.00057272 -64.5573 0.031929
0.13515 0.98801 5.5248e-05 3.8182 0.012048 1.7818e-06 0.001154 0.046672 0.00065149 0.047319 0.041954 0 0.044982 0.0389 0 0.84643 0.22749 0.058969 0.008358 4.1055 0.052663 6.2813e-05 0.8374 0.0051037 0.0058417 0.039139 0.06332 0.034522 0.00012412 0.00051242 0.13044 0.60837 0.6522 0.0092896 0.61121 0.47998 0.1097 0.42467 1.0345 1.0283 15.9967 144.9822 0.00057235 -64.7586 0.032126
0.13534 0.98801 5.5248e-05 3.8182 0.012048 1.7844e-06 0.001154 0.046702 0.0006515 0.047349 0.041981 0 0.044979 0.0389 0 0.84643 0.22749 0.058969 0.0083581 4.1055 0.052663 6.2813e-05 0.8374 0.0051037 0.0058417 0.037985 0.065727 0.035468 0.00011973 0.00049395 0.13044 0.60848 0.6525 0.0091066 0.6114 0.48001 0.10687 0.42464 1.035 1.0288 15.9967 144.9822 0.00057199 -64.959 0.032322
0.13554 0.98801 5.5248e-05 3.8182 0.012048 1.787e-06 0.001154 0.046732 0.0006515 0.047379 0.042008 0 0.044977 0.0389 0 0.84644 0.22749 0.05897 0.0083582 4.1055 0.052663 6.2814e-05 0.8374 0.0051037 0.0058417 0.036866 0.068201 0.036436 0.00011551 0.00047623 0.13044 0.60859 0.6528 0.0089297 0.61159 0.48004 0.10407 0.42461 1.0354 1.0293 15.9967 144.9822 0.00057162 -65.1586 0.032518
0.13573 0.98801 5.5248e-05 3.8182 0.012048 1.7896e-06 0.001154 0.046761 0.00065151 0.047408 0.042035 0 0.044974 0.0389 0 0.84644 0.22749 0.05897 0.0083582 4.1055 0.052663 6.2814e-05 0.8374 0.0051037 0.0058417 0.035782 0.070743 0.037425 0.00011145 0.00045923 0.13044 0.60871 0.6531 0.0087583 0.61177 0.48006 0.10128 0.42458 1.0359 1.0297 15.9967 144.9822 0.00057126 -65.3574 0.032715
0.13593 0.98801 5.5248e-05 3.8182 0.012048 1.7921e-06 0.001154 0.046791 0.00065152 0.047438 0.042062 0 0.044971 0.0389 0 0.84644 0.2275 0.058971 0.0083583 4.1055 0.052663 6.2814e-05 0.8374 0.0051037 0.0058417 0.034733 0.073354 0.038436 0.00010756 0.00044291 0.13044 0.60883 0.6534 0.0085921 0.61196 0.48009 0.098528 0.42455 1.0364 1.0302 15.9967 144.9822 0.00057089 -65.5553 0.032911
0.13613 0.98801 5.5248e-05 3.8182 0.012048 1.7947e-06 0.001154 0.046821 0.00065153 0.047468 0.042089 0 0.044968 0.0389 0 0.84645 0.2275 0.058971 0.0083583 4.1055 0.052664 6.2815e-05 0.8374 0.0051037 0.0058417 0.033716 0.076037 0.039469 0.00010382 0.00042724 0.13044 0.60896 0.6537 0.0084305 0.61215 0.48011 0.0958 0.42452 1.0368 1.0307 15.9967 144.9822 0.00057052 -65.7524 0.033108
0.13632 0.98801 5.5248e-05 3.8182 0.012048 1.7973e-06 0.001154 0.046851 0.00065153 0.047498 0.042116 0 0.044966 0.0389 0 0.84645 0.2275 0.058972 0.0083584 4.1055 0.052664 6.2815e-05 0.8374 0.0051037 0.0058417 0.032731 0.078792 0.040525 0.00010022 0.0004122 0.13044 0.60908 0.654 0.0082735 0.61233 0.48014 0.093099 0.42449 1.0373 1.0311 15.9967 144.9822 0.00057016 -65.9487 0.033304
0.13652 0.98801 5.5248e-05 3.8182 0.012048 1.7999e-06 0.001154 0.04688 0.00065154 0.047527 0.042143 0 0.044963 0.0389 0 0.84645 0.2275 0.058972 0.0083585 4.1055 0.052664 6.2815e-05 0.8374 0.0051037 0.0058417 0.031779 0.08162 0.041603 9.6765e-05 0.00039776 0.13044 0.60921 0.6543 0.0081206 0.61252 0.48016 0.090429 0.42446 1.0377 1.0316 15.9967 144.9822 0.00056979 -66.1441 0.0335
0.13681 0.98801 5.5248e-05 3.8182 0.012048 1.8037e-06 0.001154 0.046924 0.00065155 0.047571 0.042183 0 0.044959 0.0389 0 0.84646 0.2275 0.058973 0.0083586 4.1055 0.052665 6.2816e-05 0.8374 0.0051037 0.0058417 0.030429 0.085923 0.043234 9.1916e-05 0.00037752 0.13044 0.6094 0.65474 0.0079028 0.61279 0.4802 0.086553 0.42441 1.0384 1.0323 15.9967 144.9822 0.00056925 -66.4305 0.033789
0.1371 0.98801 5.5248e-05 3.8182 0.012048 1.8075e-06 0.001154 0.046968 0.00065156 0.047615 0.042223 0 0.044955 0.0389 0 0.84646 0.2275 0.058974 0.0083587 4.1055 0.052665 6.2816e-05 0.8374 0.0051037 0.0058417 0.029141 0.090394 0.044918 8.7341e-05 0.00035845 0.13044 0.6096 0.65518 0.0076931 0.61306 0.48024 0.08275 0.42437 1.0391 1.0329 15.9967 144.9822 0.00056871 -66.715 0.034079
0.13739 0.98801 5.5248e-05 3.8182 0.012048 1.8114e-06 0.001154 0.047012 0.00065157 0.047659 0.042262 0 0.044951 0.0389 0 0.84647 0.22751 0.058975 0.0083588 4.1055 0.052665 6.2817e-05 0.8374 0.0051037 0.0058417 0.027912 0.095036 0.046654 8.3023e-05 0.00034046 0.13044 0.6098 0.65561 0.007491 0.61333 0.48027 0.079024 0.42433 1.0398 1.0336 15.9967 144.9822 0.00056817 -66.9977 0.034368
0.13768 0.98801 5.5248e-05 3.8182 0.012048 1.8152e-06 0.001154 0.047055 0.00065158 0.047702 0.042302 0 0.044947 0.0389 0 0.84647 0.22751 0.058975 0.0083589 4.1055 0.052666 6.2817e-05 0.8374 0.0051037 0.0058417 0.026741 0.099853 0.048445 7.8945e-05 0.0003235 0.13044 0.61001 0.65605 0.0072961 0.6136 0.48031 0.075378 0.42429 1.0404 1.0343 15.9967 144.9822 0.00056763 -67.2785 0.034657
0.13797 0.98801 5.5248e-05 3.8182 0.012048 1.819e-06 0.001154 0.047099 0.00065159 0.047746 0.042342 0 0.044943 0.0389 0 0.84648 0.22751 0.058976 0.008359 4.1055 0.052666 6.2817e-05 0.8374 0.0051037 0.0058417 0.025623 0.10485 0.050292 7.5094e-05 0.0003075 0.13044 0.61022 0.65648 0.0071081 0.61387 0.48035 0.071818 0.42425 1.0411 1.035 15.9967 144.9822 0.00056709 -67.5575 0.034946
0.13854 0.98801 5.5248e-05 3.8182 0.012048 1.8266e-06 0.001154 0.047186 0.00065161 0.047833 0.042421 0 0.044935 0.0389 0 0.84649 0.22752 0.058978 0.0083591 4.1055 0.052667 6.2818e-05 0.8374 0.0051037 0.0058417 0.023539 0.1154 0.05416 6.8019e-05 0.00027815 0.13045 0.61066 0.65735 0.0067515 0.6144 0.48042 0.064965 0.42417 1.0425 1.0363 15.9968 144.9821 0.00056601 -68.1098 0.035525
0.13907 0.98801 5.5248e-05 3.8182 0.012048 1.8335e-06 0.001154 0.047265 0.00065163 0.047912 0.042492 0 0.044927 0.0389 0 0.84649 0.22752 0.058979 0.0083593 4.1055 0.052667 6.2819e-05 0.8374 0.0051037 0.0058417 0.021824 0.12555 0.057848 6.2298e-05 0.00025447 0.13045 0.61106 0.65812 0.006451 0.61488 0.48049 0.059121 0.42409 1.0437 1.0376 15.9968 144.9821 0.00056503 -68.6003 0.036045
0.13959 0.98801 5.5248e-05 3.8182 0.012048 1.8403e-06 0.001154 0.047344 0.00065165 0.047991 0.042564 0 0.04492 0.0389 0 0.8465 0.22752 0.05898 0.0083595 4.1055 0.052668 6.282e-05 0.83739 0.0051037 0.0058417 0.020248 0.13633 0.061741 5.7128e-05 0.00023309 0.13045 0.61148 0.6589 0.0061685 0.61536 0.48056 0.053599 0.42402 1.0449 1.0388 15.9968 144.9821 0.00056406 -69.0845 0.036566
0.14011 0.98801 5.5247e-05 3.8182 0.012048 1.8472e-06 0.001154 0.047422 0.00065167 0.048069 0.042635 0 0.044913 0.0389 0 0.84651 0.22753 0.058982 0.0083597 4.1055 0.052669 6.2821e-05 0.83739 0.0051038 0.0058417 0.018802 0.14778 0.065849 5.2449e-05 0.00021378 0.13045 0.61191 0.65967 0.0059028 0.61584 0.48063 0.048411 0.42395 1.0461 1.04 15.9968 144.9821 0.00056308 -69.5621 0.037087
0.14063 0.98801 5.5247e-05 3.8182 0.012048 1.8541e-06 0.001154 0.047501 0.00065168 0.048148 0.042706 0 0.044906 0.0389 0 0.84652 0.22753 0.058983 0.0083598 4.1055 0.052669 6.2822e-05 0.83739 0.0051038 0.0058417 0.017467 0.1599 0.070183 4.8214e-05 0.00019633 0.13045 0.61234 0.66043 0.0056527 0.61632 0.4807 0.043564 0.42389 1.0473 1.0412 15.9968 144.9821 0.00056211 -70.0329 0.037607
0.14115 0.98801 5.5247e-05 3.8182 0.012048 1.8609e-06 0.001154 0.047579 0.0006517 0.048226 0.042778 0 0.044898 0.0389 0 0.84653 0.22753 0.058985 0.00836 4.1055 0.05267 6.2822e-05 0.83739 0.0051038 0.0058418 0.016248 0.1727 0.074754 4.4375e-05 0.00018053 0.13045 0.61279 0.66119 0.0054173 0.61681 0.48077 0.039064 0.42382 1.0485 1.0425 15.9969 144.9821 0.00056114 -70.4969 0.038128
0.14159 0.98801 5.5247e-05 3.8182 0.012048 1.8668e-06 0.001154 0.047646 0.00065172 0.048293 0.042839 0 0.044892 0.0389 0 0.84654 0.22754 0.058986 0.0083602 4.1055 0.05267 6.2823e-05 0.83739 0.0051038 0.0058418 0.015283 0.18419 0.078855 4.138e-05 0.00016822 0.13045 0.61318 0.66184 0.005227 0.61722 0.48082 0.035495 0.42377 1.0496 1.0435 15.9969 144.982 0.00056031 -70.8875 0.038573
0.14198 0.98801 5.5247e-05 3.8182 0.012048 1.8718e-06 0.001154 0.047704 0.00065173 0.048351 0.042891 0 0.044887 0.0389 0 0.84654 0.22754 0.058987 0.0083603 4.1055 0.052671 6.2824e-05 0.83739 0.0051038 0.0058418 0.014502 0.19455 0.082558 3.8983e-05 0.00015837 0.13045 0.61353 0.6624 0.00507 0.61758 0.48088 0.032608 0.42372 1.0505 1.0444 15.9969 144.982 0.00055958 -71.2214 0.038958
0.14236 0.98801 5.5247e-05 3.8182 0.012048 1.8769e-06 0.001154 0.047762 0.00065174 0.04841 0.042944 0 0.044882 0.0389 0 0.84655 0.22754 0.058988 0.0083604 4.1055 0.052671 6.2824e-05 0.83739 0.0051038 0.0058418 0.013768 0.2053 0.086408 3.6752e-05 0.00014922 0.13045 0.61387 0.66296 0.0049197 0.61795 0.48093 0.029907 0.42367 1.0513 1.0453 15.9969 144.982 0.00055886 -71.5513 0.039343
0.14275 0.98801 5.5247e-05 3.8182 0.012048 1.882e-06 0.001154 0.04782 0.00065176 0.048468 0.042997 0 0.044876 0.0389 0 0.84656 0.22755 0.058989 0.0083606 4.1055 0.052672 6.2825e-05 0.83739 0.0051038 0.0058418 0.013078 0.21643 0.090408 3.4675e-05 0.0001407 0.13045 0.61422 0.66352 0.0047759 0.61831 0.48098 0.027389 0.42363 1.0522 1.0462 15.9969 144.982 0.00055815 -71.8769 0.039728
0.14313 0.98801 5.5247e-05 3.8182 0.012048 1.8871e-06 0.001154 0.047878 0.00065177 0.048525 0.043049 0 0.044871 0.0389 0 0.84656 0.22755 0.05899 0.0083607 4.1056 0.052672 6.2826e-05 0.83739 0.0051038 0.0058418 0.012431 0.22794 0.094564 3.2741e-05 0.00013278 0.13045 0.61458 0.66407 0.0046384 0.61868 0.48103 0.025049 0.42358 1.0531 1.0471 15.997 144.982 0.00055743 -72.1983 0.040113
0.14352 0.98801 5.5247e-05 3.8182 0.012048 1.8922e-06 0.001154 0.047936 0.00065178 0.048583 0.043102 0 0.044866 0.0389 0 0.84657 0.22755 0.058991 0.0083608 4.1056 0.052673 6.2826e-05 0.83739 0.0051038 0.0058418 0.011822 0.23983 0.09888 3.0941e-05 0.00012541 0.13045 0.61494 0.66462 0.0045068 0.61905 0.48108 0.022885 0.42354 1.054 1.048 15.997 144.982 0.00055671 -72.5153 0.040498
0.1439 0.98801 5.5247e-05 3.8182 0.012048 1.8972e-06 0.001154 0.047994 0.00065179 0.048641 0.043154 0 0.04486 0.0389 0 0.84658 0.22755 0.058992 0.008361 4.1056 0.052673 6.2827e-05 0.83739 0.0051038 0.0058418 0.011251 0.25209 0.10336 2.9262e-05 0.00011855 0.13045 0.6153 0.66518 0.0043809 0.61942 0.48113 0.020889 0.4235 1.0549 1.0489 15.997 144.982 0.00055599 -72.8278 0.040883
0.14429 0.98801 5.5247e-05 3.8182 0.012048 1.9023e-06 0.001154 0.048052 0.00065181 0.048699 0.043207 0 0.044855 0.0389 0 0.84658 0.22756 0.058993 0.0083611 4.1056 0.052674 6.2828e-05 0.83739 0.0051038 0.0058418 0.010713 0.26471 0.10801 2.7698e-05 0.00011216 0.13045 0.61567 0.66572 0.0042603 0.6198 0.48119 0.019055 0.42346 1.0558 1.0498 15.997 144.982 0.00055527 -73.1358 0.041268
0.14467 0.98801 5.5247e-05 3.8182 0.012048 1.9074e-06 0.001154 0.04811 0.00065182 0.048757 0.04326 0 0.04485 0.0389 0 0.84659 0.22756 0.058994 0.0083612 4.1056 0.052674 6.2828e-05 0.83739 0.0051038 0.0058418 0.010208 0.27769 0.11283 2.6238e-05 0.0001062 0.13045 0.61604 0.66627 0.004145 0.62018 0.48124 0.017376 0.42342 1.0567 1.0507 15.997 144.982 0.00055455 -73.4391 0.041653
0.14506 0.98801 5.5247e-05 3.8182 0.012048 1.9125e-06 0.001154 0.048168 0.00065183 0.048815 0.043312 0 0.044844 0.0389 0 0.8466 0.22756 0.058995 0.0083614 4.1056 0.052675 6.2829e-05 0.83739 0.0051038 0.0058418 0.009734 0.29102 0.11784 2.4877e-05 0.00010064 0.13045 0.61641 0.66682 0.0040346 0.62056 0.48129 0.015844 0.42338 1.0576 1.0516 15.9971 144.9819 0.00055383 -73.7377 0.042038
0.14544 0.98801 5.5247e-05 3.8182 0.012048 1.9175e-06 0.001154 0.048226 0.00065184 0.048873 0.043365 0 0.044839 0.0389 0 0.8466 0.22757 0.058996 0.0083615 4.1056 0.052675 6.283e-05 0.83739 0.0051038 0.0058418 0.0092881 0.30468 0.12302 2.3608e-05 9.5462e-05 0.13045 0.61678 0.66736 0.003929 0.62095 0.48134 0.014451 0.42334 1.0585 1.0525 15.9971 144.9819 0.00055311 -74.0313 0.042423
0.14583 0.98801 5.5247e-05 3.8182 0.012048 1.9226e-06 0.001154 0.048284 0.00065186 0.048931 0.043417 0 0.044834 0.0389 0 0.84661 0.22757 0.058997 0.0083616 4.1056 0.052676 6.283e-05 0.83739 0.0051038 0.0058418 0.0088691 0.31866 0.1284 2.2423e-05 9.0631e-05 0.13045 0.61716 0.6679 0.0038279 0.62134 0.4814 0.013188 0.4233 1.0594 1.0534 15.9971 144.9819 0.00055239 -74.3201 0.042808
0.14621 0.98801 5.5247e-05 3.8182 0.012048 1.9277e-06 0.001154 0.048341 0.00065187 0.048989 0.04347 0 0.044828 0.0389 0 0.84662 0.22757 0.058998 0.0083618 4.1056 0.052677 6.2831e-05 0.83739 0.0051038 0.0058418 0.0084749 0.33293 0.13396 2.1316e-05 8.6123e-05 0.13045 0.61754 0.66844 0.0037312 0.62173 0.48145 0.012049 0.42326 1.0603 1.0543 15.9971 144.9819 0.00055168 -74.6038 0.043193
0.1466 0.98801 5.5247e-05 3.8182 0.012048 1.9328e-06 0.001154 0.048399 0.00065188 0.049047 0.043522 0 0.044823 0.0389 0 0.84662 0.22758 0.058999 0.0083619 4.1056 0.052677 6.2831e-05 0.83739 0.0051038 0.0058418 0.008105 0.3475 0.13971 2.0283e-05 8.1916e-05 0.13045 0.61792 0.66898 0.0036387 0.62213 0.4815 0.011023 0.42322 1.0612 1.0552 15.9972 144.9819 0.00055096 -74.8824 0.043578
0.14698 0.98801 5.5247e-05 3.8182 0.012048 1.9378e-06 0.001154 0.048457 0.0006519 0.049104 0.043575 0 0.044818 0.0389 0 0.84663 0.22758 0.059001 0.008362 4.1056 0.052678 6.2832e-05 0.83739 0.0051038 0.0058418 0.0077559 0.36232 0.14566 1.9318e-05 7.7988e-05 0.13045 0.61831 0.66952 0.0035502 0.62254 0.48156 0.010102 0.42319 1.062 1.0561 15.9972 144.9819 0.00055024 -75.1559 0.043963
0.14737 0.98801 5.5247e-05 3.8182 0.012048 1.9429e-06 0.001154 0.048515 0.00065191 0.049162 0.043627 0 0.044812 0.0389 0 0.84664 0.22758 0.059002 0.0083622 4.1056 0.052678 6.2833e-05 0.83738 0.0051039 0.0058418 0.007431 0.37738 0.15181 1.8416e-05 7.432e-05 0.13045 0.6187 0.67006 0.0034656 0.62294 0.48161 0.0092787 0.42315 1.0629 1.057 15.9972 144.9819 0.00054952 -75.4241 0.044349
0.14775 0.98801 5.5247e-05 3.8182 0.012048 1.948e-06 0.001154 0.048573 0.00065192 0.04922 0.04368 0 0.044807 0.0389 0 0.84664 0.22758 0.059003 0.0083623 4.1056 0.052679 6.2833e-05 0.83738 0.0051039 0.0058418 0.0071211 0.39266 0.15815 1.7573e-05 7.0892e-05 0.13045 0.61908 0.67059 0.0033846 0.62336 0.48166 0.0085441 0.42312 1.0638 1.0579 15.9972 144.9819 0.00054881 -75.687 0.044734
0.14814 0.98801 5.5247e-05 3.8182 0.012048 1.9531e-06 0.001154 0.04863 0.00065193 0.049278 0.043732 0 0.044802 0.0389 0 0.84665 0.22759 0.059004 0.0083624 4.1056 0.052679 6.2834e-05 0.83738 0.0051039 0.0058418 0.0068324 0.40814 0.16469 1.6785e-05 6.7688e-05 0.13045 0.61948 0.67112 0.0033072 0.62377 0.48172 0.0078905 0.42309 1.0647 1.0588 15.9973 144.9819 0.00054809 -75.9446 0.045119
0.14849 0.98801 5.5247e-05 3.8182 0.012048 1.9576e-06 0.001154 0.048682 0.00065194 0.04933 0.043779 0 0.044797 0.0389 0 0.84666 0.22759 0.059005 0.0083626 4.1056 0.05268 6.2835e-05 0.83738 0.0051039 0.0058419 0.0065871 0.4222 0.17074 1.6119e-05 6.4983e-05 0.13045 0.61983 0.6716 0.0032404 0.62415 0.48177 0.0073654 0.42306 1.0655 1.0596 15.9973 144.9819 0.00054745 -76.1717 0.045465
0.14883 0.98801 5.5247e-05 3.8182 0.012048 1.9622e-06 0.001154 0.048734 0.00065195 0.049382 0.043826 0 0.044792 0.0389 0 0.84666 0.22759 0.059006 0.0083627 4.1056 0.05268 6.2835e-05 0.83738 0.0051039 0.0058419 0.0063538 0.43638 0.17695 1.5491e-05 6.2436e-05 0.13045 0.62018 0.67208 0.0031763 0.62454 0.48182 0.0068946 0.42303 1.0663 1.0604 15.9973 144.9818 0.00054681 -76.3945 0.045812
0.14918 0.98801 5.5247e-05 3.8182 0.012048 1.9668e-06 0.001154 0.048786 0.00065197 0.049433 0.043874 0 0.044788 0.0389 0 0.84667 0.2276 0.059007 0.0083628 4.1056 0.052681 6.2836e-05 0.83738 0.0051039 0.0058419 0.0061335 0.45065 0.18332 1.49e-05 6.0037e-05 0.13045 0.62054 0.67255 0.0031147 0.62493 0.48187 0.006473 0.423 1.0671 1.0612 15.9973 144.9818 0.00054616 -76.6129 0.046158
0.14952 0.98801 5.5247e-05 3.8182 0.012048 1.9713e-06 0.001154 0.048838 0.00065198 0.049485 0.043921 0 0.044783 0.0389 0 0.84667 0.2276 0.059008 0.0083629 4.1056 0.052681 6.2837e-05 0.83738 0.0051039 0.0058419 0.005923 0.46499 0.18984 1.4343e-05 5.7776e-05 0.13045 0.62089 0.67302 0.0030556 0.62532 0.48192 0.0060961 0.42298 1.0679 1.062 15.9974 144.9818 0.00054552 -76.8267 0.046505
0.14987 0.98801 5.5247e-05 3.8182 0.012048 1.9759e-06 0.001154 0.04889 0.00065199 0.049537 0.043968 0 0.044778 0.0389 0 0.84668 0.2276 0.059009 0.008363 4.1056 0.052681 6.2837e-05 0.83738 0.0051039 0.0058419 0.0057271 0.47938 0.19651 1.3818e-05 5.5646e-05 0.13045 0.62125 0.6735 0.0029988 0.62572 0.48197 0.0057594 0.42295 1.0687 1.0628 15.9974 144.9818 0.00054488 -77.0362 0.046851
0.15022 0.98801 5.5247e-05 3.8182 0.012048 1.9805e-06 0.001154 0.048942 0.000652 0.049589 0.044015 0 0.044773 0.0389 0 0.84669 0.2276 0.05901 0.0083632 4.1056 0.052682 6.2838e-05 0.83738 0.0051039 0.0058419 0.00554 0.4938 0.20333 1.3323e-05 5.3637e-05 0.13045 0.62161 0.67397 0.0029442 0.62612 0.48202 0.0054587 0.42292 1.0695 1.0636 15.9974 144.9818 0.00054424 -77.2411 0.047198
0.15056 0.98801 5.5247e-05 3.8182 0.012048 1.985e-06 0.001154 0.048994 0.00065201 0.049641 0.044062 0 0.044769 0.0389 0 0.84669 0.22761 0.059011 0.0083633 4.1056 0.052682 6.2838e-05 0.83738 0.0051039 0.0058419 0.0053628 0.50822 0.21029 1.2855e-05 5.1743e-05 0.13045 0.62197 0.67444 0.0028919 0.62653 0.48207 0.0051903 0.4229 1.0703 1.0644 15.9974 144.9818 0.0005436 -77.4416 0.047544
0.15091 0.98801 5.5247e-05 3.8182 0.012048 1.9896e-06 0.001154 0.049045 0.00065202 0.049693 0.044109 0 0.044764 0.0389 0 0.8467 0.22761 0.059012 0.0083634 4.1056 0.052683 6.2839e-05 0.83738 0.0051039 0.0058419 0.0051948 0.52261 0.2174 1.2414e-05 4.9956e-05 0.13045 0.62233 0.67491 0.0028416 0.62694 0.48212 0.0049508 0.42287 1.0711 1.0652 15.9975 144.9818 0.00054296 -77.6376 0.047891
0.15126 0.98801 5.5247e-05 3.8182 0.012048 1.9942e-06 0.001154 0.049097 0.00065203 0.049745 0.044156 0 0.044759 0.0389 0 0.84671 0.22761 0.059013 0.0083635 4.1056 0.052683 6.284e-05 0.83738 0.0051039 0.0058419 0.005035 0.53697 0.22464 1.1998e-05 4.827e-05 0.13045 0.62269 0.67537 0.0027933 0.62735 0.48217 0.004737 0.42285 1.0719 1.066 15.9975 144.9818 0.00054232 -77.8291 0.048238
0.15195 0.98801 5.5247e-05 3.8182 0.012048 2.0033e-06 0.001154 0.049201 0.00065205 0.049848 0.04425 0 0.04475 0.0389 0 0.84672 0.22762 0.059015 0.0083638 4.1056 0.052684 6.2841e-05 0.83738 0.0051039 0.0058419 0.0047411 0.56546 0.2395 1.1233e-05 4.5175e-05 0.13045 0.62342 0.6763 0.0027025 0.6282 0.48227 0.0043754 0.42281 1.0735 1.0676 15.9975 144.9818 0.00054104 -78.1989 0.048931
0.15257 0.98801 5.5247e-05 3.8182 0.012048 2.0115e-06 0.001154 0.049294 0.00065207 0.049942 0.044335 0 0.044741 0.0389 0 0.84673 0.22762 0.059016 0.008364 4.1056 0.052685 6.2842e-05 0.83738 0.0051039 0.0058419 0.0045019 0.59074 0.25329 1.0616e-05 4.2676e-05 0.13045 0.62407 0.67714 0.0026269 0.62898 0.48236 0.0041114 0.42277 1.0749 1.0691 15.9976 144.9818 0.00053989 -78.5166 0.049555
0.1532 0.98801 5.5247e-05 3.8182 0.012048 2.0197e-06 0.001154 0.049387 0.00065209 0.050035 0.04442 0 0.044732 0.0389 0 0.84674 0.22763 0.059018 0.0083642 4.1057 0.052686 6.2843e-05 0.83738 0.0051039 0.0058419 0.0042844 0.61554 0.26742 1.0057e-05 4.0417e-05 0.13045 0.62473 0.67796 0.0025567 0.62977 0.48245 0.0038934 0.42273 1.0763 1.0705 15.9976 144.9817 0.00053874 -78.8201 0.050178
0.15382 0.98801 5.5247e-05 3.8182 0.012048 2.028e-06 0.001154 0.04948 0.00065211 0.050128 0.044504 0 0.044724 0.0389 0 0.84675 0.22763 0.05902 0.0083645 4.1057 0.052687 6.2844e-05 0.83738 0.0051039 0.0058419 0.0040865 0.63974 0.28187 9.5519e-06 3.8374e-05 0.13045 0.62538 0.67879 0.0024915 0.63058 0.48254 0.0037117 0.42269 1.0778 1.0719 15.9977 144.9817 0.0005376 -79.1098 0.050802
0.15445 0.98801 5.5247e-05 3.8182 0.012048 2.0362e-06 0.001154 0.049573 0.00065213 0.050221 0.044589 0 0.044715 0.0389 0 0.84676 0.22764 0.059022 0.0083647 4.1057 0.052688 6.2845e-05 0.83737 0.005104 0.0058419 0.0039062 0.66325 0.29658 9.094e-06 3.6523e-05 0.13045 0.62604 0.67961 0.0024309 0.6314 0.48264 0.0035587 0.42266 1.0792 1.0734 15.9977 144.9817 0.00053646 -79.3858 0.051426
0.15507 0.98801 5.5247e-05 3.8182 0.012048 2.0444e-06 0.001154 0.049666 0.00065215 0.050314 0.044673 0 0.044707 0.0389 0 0.84678 0.22764 0.059023 0.0083649 4.1057 0.052689 6.2846e-05 0.83737 0.005104 0.0058419 0.0037418 0.68597 0.31151 8.6787e-06 3.4846e-05 0.13045 0.6267 0.68043 0.0023747 0.63224 0.48273 0.0034283 0.42263 1.0806 1.0748 15.9978 144.9817 0.00053532 -79.6485 0.05205
0.15569 0.98801 5.5247e-05 3.8182 0.012048 2.0526e-06 0.001154 0.049759 0.00065217 0.050407 0.044758 0 0.044698 0.0389 0 0.84679 0.22765 0.059025 0.0083652 4.1057 0.05269 6.2848e-05 0.83737 0.005104 0.005842 0.0035918 0.70782 0.32663 8.3015e-06 3.3323e-05 0.13045 0.62736 0.68124 0.0023225 0.63309 0.48283 0.0033159 0.4226 1.082 1.0762 15.9979 144.9817 0.00053418 -79.8981 0.052673
0.15632 0.98801 5.5246e-05 3.8182 0.012048 2.0609e-06 0.001154 0.049852 0.00065219 0.0505 0.044842 0 0.04469 0.0389 0 0.8468 0.22765 0.059027 0.0083654 4.1057 0.052691 6.2849e-05 0.83737 0.005104 0.005842 0.0034549 0.72873 0.34188 7.9587e-06 3.1939e-05 0.13045 0.62803 0.68205 0.002274 0.63396 0.48292 0.0032178 0.42257 1.0834 1.0777 15.9979 144.9817 0.00053305 -80.1352 0.053297
0.15694 0.98801 5.5246e-05 3.8182 0.012048 2.0691e-06 0.001154 0.049945 0.00065221 0.050593 0.044927 0 0.044682 0.0389 0 0.84681 0.22766 0.059029 0.0083656 4.1057 0.052692 6.285e-05 0.83737 0.005104 0.005842 0.0033298 0.74865 0.35723 7.6467e-06 3.068e-05 0.13045 0.62869 0.68285 0.0022289 0.63484 0.48302 0.0031315 0.42254 1.0849 1.0791 15.998 144.9817 0.00053192 -80.36 0.053921
0.15756 0.98801 5.5246e-05 3.8182 0.012048 2.0773e-06 0.001154 0.050038 0.00065222 0.050686 0.045011 0 0.044673 0.0389 0 0.84682 0.22766 0.059031 0.0083659 4.1057 0.052693 6.2851e-05 0.83737 0.005104 0.005842 0.0032154 0.76754 0.37263 7.3624e-06 2.9533e-05 0.13045 0.62935 0.68365 0.0021871 0.63573 0.48311 0.0030549 0.42252 1.0863 1.0805 15.998 144.9817 0.00053079 -80.5729 0.054545
0.15819 0.98801 5.5246e-05 3.8182 0.012048 2.0855e-06 0.001154 0.050131 0.00065224 0.050779 0.045095 0 0.044665 0.0389 0 0.84683 0.22767 0.059033 0.0083661 4.1057 0.052693 6.2852e-05 0.83737 0.005104 0.005842 0.0031106 0.78537 0.38805 7.1031e-06 2.8487e-05 0.13045 0.63002 0.68445 0.0021483 0.63664 0.48321 0.0029864 0.42249 1.0877 1.082 15.9981 144.9817 0.00052966 -80.7745 0.055169
0.15881 0.98801 5.5246e-05 3.8182 0.012048 2.0937e-06 0.001154 0.050224 0.00065226 0.050871 0.04518 0 0.044656 0.0389 0 0.84684 0.22767 0.059034 0.0083663 4.1057 0.052694 6.2853e-05 0.83737 0.005104 0.005842 0.0030146 0.80214 0.40344 6.8664e-06 2.7533e-05 0.13045 0.63068 0.68524 0.0021122 0.63756 0.48331 0.0029247 0.42247 1.0891 1.0834 15.9981 144.9817 0.00052854 -80.9651 0.055792
0.15981 0.98801 5.5246e-05 3.8182 0.012048 2.1069e-06 0.001154 0.050372 0.00065229 0.05102 0.045315 0 0.044643 0.0389 0 0.84686 0.22768 0.059037 0.0083667 4.1057 0.052696 6.2855e-05 0.83737 0.005104 0.005842 0.0028772 0.82679 0.428 6.5285e-06 2.6171e-05 0.13045 0.63174 0.68651 0.0020596 0.63906 0.48347 0.0028375 0.42243 1.0914 1.0857 15.9982 144.9817 0.00052674 -81.2489 0.056792
0.16081 0.98801 5.5246e-05 3.8182 0.012048 2.1201e-06 0.001154 0.050521 0.00065232 0.051168 0.04545 0 0.044629 0.0389 0 0.84688 0.22769 0.05904 0.0083671 4.1057 0.052697 6.2857e-05 0.83737 0.0051041 0.005842 0.002757 0.84876 0.45227 6.2349e-06 2.4988e-05 0.13045 0.63281 0.68776 0.0020128 0.6406 0.48362 0.002762 0.4224 1.0937 1.088 15.9983 144.9817 0.00052495 -81.5075 0.057792
0.16181 0.98801 5.5246e-05 3.8182 0.012048 2.1333e-06 0.001154 0.050669 0.00065235 0.051317 0.045585 0 0.044616 0.0389 0 0.8469 0.2277 0.059043 0.0083675 4.1058 0.052699 6.2859e-05 0.83736 0.0051041 0.0058421 0.0026531 0.86815 0.47617 5.9798e-06 2.396e-05 0.13045 0.63387 0.68901 0.0019712 0.64215 0.48378 0.0026962 0.42237 1.0959 1.0903 15.9984 144.9816 0.00052317 -81.7427 0.058792
0.16281 0.98801 5.5246e-05 3.8182 0.012048 2.1465e-06 0.001154 0.050817 0.00065238 0.051465 0.045719 0 0.044602 0.0389 0 0.84692 0.22771 0.059047 0.0083678 4.1058 0.0527 6.2861e-05 0.83736 0.0051041 0.0058421 0.0025602 0.88512 0.49957 5.7566e-06 2.3062e-05 0.13045 0.63493 0.69024 0.0019342 0.64374 0.48394 0.0026385 0.42235 1.0982 1.0925 15.9985 144.9816 0.0005214 -81.9565 0.059792
0.16381 0.98801 5.5246e-05 3.8182 0.012048 2.1596e-06 0.001154 0.050965 0.00065241 0.051613 0.045854 0 0.044589 0.0389 0 0.84694 0.22771 0.05905 0.0083682 4.1058 0.052702 6.2863e-05 0.83736 0.0051041 0.0058421 0.0024797 0.89985 0.52242 5.5615e-06 2.2277e-05 0.13045 0.63599 0.69147 0.0019012 0.64534 0.4841 0.0025877 0.42232 1.1004 1.0948 15.9986 144.9816 0.00051963 -82.1504 0.060792
0.16481 0.98801 5.5246e-05 3.8182 0.012048 2.1728e-06 0.001154 0.051113 0.00065243 0.051761 0.045988 0 0.044575 0.0389 0 0.84696 0.22772 0.059053 0.0083686 4.1058 0.052704 6.2865e-05 0.83736 0.0051041 0.0058421 0.0024081 0.91255 0.54464 5.3903e-06 2.1588e-05 0.13045 0.63705 0.69268 0.0018718 0.64697 0.48426 0.0025428 0.4223 1.1027 1.0971 15.9987 144.9816 0.00051788 -82.3263 0.061792
0.16581 0.98801 5.5246e-05 3.8182 0.012048 2.186e-06 0.001154 0.051261 0.00065246 0.051909 0.046123 0 0.044562 0.0389 0 0.84698 0.22773 0.059056 0.008369 4.1058 0.052705 6.2867e-05 0.83736 0.0051041 0.0058421 0.0023463 0.92343 0.56618 5.2399e-06 2.0982e-05 0.13045 0.63811 0.69389 0.0018456 0.64861 0.48443 0.0025031 0.42228 1.1049 1.0993 15.9987 144.9816 0.00051613 -82.4856 0.062792
0.16681 0.98801 5.5246e-05 3.8182 0.012048 2.1992e-06 0.001154 0.051409 0.00065249 0.052057 0.046257 0 0.044548 0.0389 0 0.847 0.22774 0.059059 0.0083694 4.1058 0.052707 6.2869e-05 0.83736 0.0051042 0.0058421 0.0022906 0.93269 0.58701 5.1072e-06 2.0449e-05 0.13045 0.63916 0.69509 0.0018221 0.65027 0.48459 0.0024679 0.42226 1.1072 1.1016 15.9988 144.9816 0.00051439 -82.6299 0.063792
0.16781 0.98801 5.5246e-05 3.8182 0.012048 2.2124e-06 0.001154 0.051557 0.00065252 0.052204 0.046391 0 0.044535 0.0389 0 0.84702 0.22775 0.059062 0.0083698 4.1058 0.052708 6.2871e-05 0.83735 0.0051042 0.0058422 0.0022421 0.94053 0.6071 4.99e-06 1.9978e-05 0.13045 0.64022 0.69628 0.0018012 0.65194 0.48475 0.0024365 0.42224 1.1094 1.1039 15.9989 144.9816 0.00051266 -82.7606 0.064792
0.16881 0.98801 5.5246e-05 3.8182 0.012048 2.2255e-06 0.001154 0.051704 0.00065254 0.052352 0.046526 0 0.044522 0.0389 0 0.84704 0.22776 0.059065 0.0083702 4.1058 0.05271 6.2873e-05 0.83735 0.0051042 0.0058422 0.0021975 0.94715 0.62643 4.8861e-06 1.956e-05 0.13045 0.64127 0.69746 0.0017824 0.65363 0.48492 0.0024086 0.42223 1.1116 1.1061 15.999 144.9816 0.00051094 -82.8789 0.065792
0.16981 0.98801 5.5246e-05 3.8182 0.012048 2.2387e-06 0.001154 0.051851 0.00065257 0.052499 0.04666 0 0.044508 0.0389 0 0.84706 0.22777 0.059068 0.0083706 4.1059 0.052712 6.2875e-05 0.83735 0.0051042 0.0058422 0.0021603 0.9527 0.64499 4.794e-06 1.919e-05 0.13045 0.64232 0.69863 0.0017656 0.65532 0.48508 0.0023837 0.42221 1.1139 1.1084 15.9991 144.9816 0.00050923 -82.9861 0.066792
0.17081 0.98801 5.5246e-05 3.8182 0.012048 2.2519e-06 0.001154 0.051999 0.0006526 0.052647 0.046794 0 0.044495 0.0389 0 0.84708 0.22778 0.059071 0.008371 4.1059 0.052713 6.2877e-05 0.83735 0.0051042 0.0058422 0.0021234 0.95736 0.66278 4.7118e-06 1.886e-05 0.13045 0.64337 0.6998 0.0017504 0.65702 0.48524 0.0023614 0.4222 1.1161 1.1106 15.9992 144.9816 0.00050752 -83.0833 0.067792
0.17171 0.98801 5.5246e-05 3.8182 0.012048 2.2638e-06 0.001154 0.052131 0.00065262 0.052779 0.046914 0 0.044483 0.0389 0 0.8471 0.22778 0.059074 0.0083713 4.1059 0.052715 6.2879e-05 0.83735 0.0051042 0.0058422 0.0020968 0.96089 0.67814 4.6456e-06 1.8593e-05 0.13045 0.64431 0.70084 0.0017382 0.65856 0.48539 0.0023434 0.42219 1.1181 1.1126 15.9993 144.9816 0.00050599 -83.1629 0.068692
0.17261 0.98801 5.5245e-05 3.8182 0.012048 2.2756e-06 0.001154 0.052264 0.00065265 0.052912 0.047034 0 0.044471 0.0389 0 0.84711 0.22779 0.059077 0.0083717 4.1059 0.052716 6.2881e-05 0.83735 0.0051043 0.0058422 0.0020705 0.96388 0.69288 4.5858e-06 1.8353e-05 0.13045 0.64525 0.70187 0.001727 0.66011 0.48554 0.002327 0.42218 1.1201 1.1147 15.9994 144.9816 0.00050448 -83.236 0.069592
0.17351 0.98801 5.5245e-05 3.8182 0.012048 2.2875e-06 0.001154 0.052396 0.00065267 0.053044 0.047155 0 0.044459 0.0389 0 0.84713 0.2278 0.05908 0.0083721 4.1059 0.052718 6.2883e-05 0.83735 0.0051043 0.0058423 0.0020503 0.96642 0.70703 4.5316e-06 1.8135e-05 0.13045 0.64618 0.7029 0.0017168 0.66165 0.48569 0.0023122 0.42217 1.1221 1.1167 15.9994 144.9816 0.00050296 -83.303 0.070492
0.17441 0.98801 5.5245e-05 3.8182 0.012048 2.2993e-06 0.001154 0.052528 0.00065269 0.053176 0.047275 0 0.044447 0.0389 0 0.84715 0.22781 0.059083 0.0083724 4.1059 0.052719 6.2885e-05 0.83734 0.0051043 0.0058423 0.0020261 0.96857 0.72058 4.4823e-06 1.7937e-05 0.13045 0.64712 0.70392 0.0017075 0.6632 0.48584 0.0022987 0.42216 1.1241 1.1187 15.9995 144.9816 0.00050146 -83.3645 0.071392
0.17522 0.98801 5.5245e-05 3.8182 0.012048 2.31e-06 0.001154 0.052647 0.00065271 0.053295 0.047383 0 0.044436 0.0389 0 0.84717 0.22781 0.059085 0.0083728 4.1059 0.052721 6.2887e-05 0.83734 0.0051043 0.0058423 0.0020108 0.97023 0.73229 4.4418e-06 1.7774e-05 0.13045 0.64795 0.70483 0.0016998 0.6646 0.48598 0.0022875 0.42215 1.1259 1.1205 15.9996 144.9816 0.00050011 -83.4156 0.072202
0.17595 0.98801 5.5245e-05 3.8182 0.012048 2.3196e-06 0.001154 0.052754 0.00065273 0.053402 0.04748 0 0.044427 0.0389 0 0.84718 0.22782 0.059088 0.0083731 4.1059 0.052722 6.2888e-05 0.83734 0.0051043 0.0058423 0.0019968 0.97152 0.74243 4.4081e-06 1.7639e-05 0.13045 0.64871 0.70564 0.0016933 0.66585 0.4861 0.0022783 0.42214 1.1275 1.1221 15.9996 144.9816 0.0004989 -83.4585 0.072931
0.17668 0.98801 5.5245e-05 3.8182 0.012048 2.3292e-06 0.001154 0.052861 0.00065275 0.053509 0.047577 0 0.044417 0.0389 0 0.8472 0.22783 0.05909 0.0083734 4.106 0.052723 6.289e-05 0.83734 0.0051043 0.0058423 0.0019837 0.97265 0.75221 4.3768e-06 1.7513e-05 0.13045 0.64946 0.70646 0.0016873 0.66711 0.48622 0.0022696 0.42214 1.1291 1.1237 15.9997 144.9817 0.0004977 -83.4986 0.07366
0.17741 0.98801 5.5245e-05 3.8182 0.012048 2.3388e-06 0.001154 0.052967 0.00065277 0.053616 0.047675 0 0.044407 0.0389 0 0.84721 0.22783 0.059093 0.0083737 4.106 0.052725 6.2892e-05 0.83734 0.0051044 0.0058423 0.0019711 0.97364 0.76164 4.3477e-06 1.7396e-05 0.13045 0.65021 0.70726 0.0016817 0.66837 0.48634 0.0022616 0.42213 1.1307 1.1253 15.9998 144.9817 0.0004965 -83.5362 0.074389
0.17814 0.98801 5.5245e-05 3.8182 0.012048 2.3485e-06 0.001154 0.053074 0.00065279 0.053722 0.047772 0 0.044398 0.0389 0 0.84723 0.22784 0.059095 0.008374 4.106 0.052726 6.2893e-05 0.83734 0.0051044 0.0058423 0.0019597 0.9745 0.77072 4.3205e-06 1.7287e-05 0.13045 0.65096 0.70807 0.0016765 0.66963 0.48646 0.0022541 0.42212 1.1323 1.127 15.9998 144.9817 0.0004953 -83.5715 0.075118
0.17887 0.98801 5.5245e-05 3.8182 0.012048 2.3581e-06 0.001154 0.053181 0.00065281 0.053829 0.047869 0 0.044388 0.0389 0 0.84724 0.22785 0.059097 0.0083743 4.106 0.052727 6.2895e-05 0.83734 0.0051044 0.0058424 0.0019488 0.97526 0.77947 4.2952e-06 1.7186e-05 0.13045 0.65171 0.70887 0.0016716 0.67088 0.48658 0.0022471 0.42212 1.1339 1.1286 15.9999 144.9817 0.00049411 -83.6047 0.075847
0.1796 0.98801 5.5245e-05 3.8182 0.012048 2.3677e-06 0.001154 0.053287 0.00065283 0.053936 0.047966 0 0.044378 0.0389 0 0.84726 0.22785 0.0591 0.0083746 4.106 0.052728 6.2897e-05 0.83733 0.0051044 0.0058424 0.0019389 0.97592 0.78789 4.2715e-06 1.7091e-05 0.13045 0.65245 0.70966 0.001667 0.67214 0.48671 0.0022406 0.42211 1.1355 1.1302 16 144.9817 0.00049293 -83.6358 0.076576
0.18033 0.98801 5.5245e-05 3.8182 0.012048 2.3773e-06 0.001154 0.053394 0.00065284 0.054042 0.048063 0 0.044369 0.0389 0 0.84727 0.22786 0.059102 0.0083749 4.106 0.05273 6.2898e-05 0.83733 0.0051044 0.0058424 0.0019294 0.97651 0.796 4.2493e-06 1.7001e-05 0.13045 0.6532 0.71046 0.0016627 0.67339 0.48683 0.0022345 0.42211 1.1371 1.1318 16 144.9817 0.00049175 -83.6652 0.077305
0.18105 0.98801 5.5245e-05 3.8182 0.012048 2.3869e-06 0.001154 0.0535 0.00065286 0.054149 0.04816 0 0.044359 0.0389 0 0.84729 0.22787 0.059105 0.0083752 4.106 0.052731 6.29e-05 0.83733 0.0051044 0.0058424 0.0019207 0.97702 0.80381 4.2285e-06 1.6918e-05 0.13045 0.65394 0.71124 0.0016587 0.67465 0.48695 0.0022287 0.4221 1.1387 1.1334 16.0001 144.9817 0.00049057 -83.6928 0.078034
0.18178 0.98801 5.5245e-05 3.8182 0.012048 2.3965e-06 0.001154 0.053607 0.00065288 0.054255 0.048256 0 0.04435 0.0389 0 0.8473 0.22787 0.059107 0.0083755 4.106 0.052732 6.2901e-05 0.83733 0.0051044 0.0058424 0.0019122 0.97748 0.81131 4.2089e-06 1.6839e-05 0.13045 0.65468 0.71203 0.0016548 0.6759 0.48707 0.0022233 0.4221 1.1403 1.135 16.0002 144.9817 0.0004894 -83.719 0.078763
0.18251 0.98801 5.5245e-05 3.8182 0.012048 2.4061e-06 0.001154 0.053713 0.0006529 0.054361 0.048353 0 0.04434 0.0389 0 0.84732 0.22788 0.05911 0.0083758 4.106 0.052734 6.2903e-05 0.83733 0.0051045 0.0058424 0.0019045 0.97788 0.81853 4.1905e-06 1.6766e-05 0.13045 0.65542 0.71281 0.0016512 0.67715 0.48719 0.0022183 0.42209 1.1419 1.1366 16.0002 144.9817 0.00048823 -83.7437 0.079492
0.18324 0.98801 5.5245e-05 3.8182 0.012048 2.4157e-06 0.001154 0.053819 0.00065292 0.054468 0.04845 0 0.04433 0.0389 0 0.84733 0.22789 0.059112 0.0083761 4.106 0.052735 6.2905e-05 0.83733 0.0051045 0.0058424 0.001897 0.97823 0.82547 4.1732e-06 1.6696e-05 0.13045 0.65616 0.71358 0.0016478 0.6784 0.48732 0.0022135 0.42209 1.1435 1.1382 16.0003 144.9817 0.00048707 -83.7671 0.080221
0.18397 0.98801 5.5245e-05 3.8182 0.012048 2.4253e-06 0.001154 0.053926 0.00065293 0.054574 0.048547 0 0.044321 0.0389 0 0.84735 0.22789 0.059114 0.0083764 4.1061 0.052736 6.2907e-05 0.83733 0.0051045 0.0058425 0.0018902 0.97855 0.83214 4.1568e-06 1.663e-05 0.13045 0.6569 0.71435 0.0016446 0.67965 0.48744 0.002209 0.42209 1.1451 1.1398 16.0003 144.9817 0.00048592 -83.7893 0.08095
0.1847 0.98801 5.5245e-05 3.8182 0.012048 2.4349e-06 0.001154 0.054032 0.00065295 0.05468 0.048643 0 0.044311 0.0389 0 0.84736 0.2279 0.059117 0.0083767 4.1061 0.052738 6.2908e-05 0.83733 0.0051045 0.0058425 0.0018835 0.97883 0.83856 4.1412e-06 1.6568e-05 0.13045 0.65763 0.71512 0.0016416 0.68089 0.48756 0.0022047 0.42208 1.1467 1.1414 16.0004 144.9817 0.00048476 -83.8103 0.081679
0.18543 0.98801 5.5245e-05 3.8182 0.012048 2.4445e-06 0.001154 0.054138 0.00065297 0.054786 0.04874 0 0.044302 0.0389 0 0.84738 0.22791 0.059119 0.0083771 4.1061 0.052739 6.291e-05 0.83732 0.0051045 0.0058425 0.0018773 0.97908 0.84472 4.1265e-06 1.6509e-05 0.13045 0.65837 0.71588 0.0016387 0.68213 0.48768 0.0022007 0.42208 1.1483 1.143 16.0005 144.9817 0.00048361 -83.8304 0.082408
0.18616 0.98801 5.5245e-05 3.8182 0.012048 2.4541e-06 0.001154 0.054244 0.00065299 0.054892 0.048836 0 0.044292 0.0389 0 0.8474 0.22792 0.059122 0.0083774 4.1061 0.05274 6.2912e-05 0.83732 0.0051045 0.0058425 0.0018712 0.9793 0.85064 4.1126e-06 1.6453e-05 0.13045 0.6591 0.71664 0.0016359 0.68337 0.48781 0.0021969 0.42207 1.1498 1.1446 16.0005 144.9817 0.00048247 -83.8495 0.083137
0.18689 0.98801 5.5245e-05 3.8182 0.012048 2.4637e-06 0.001154 0.05435 0.000653 0.054998 0.048933 0 0.044283 0.0389 0 0.84741 0.22792 0.059124 0.0083777 4.1061 0.052742 6.2913e-05 0.83732 0.0051046 0.0058425 0.0018657 0.9795 0.85633 4.0993e-06 1.6399e-05 0.13045 0.65983 0.7174 0.0016333 0.68461 0.48793 0.0021932 0.42207 1.1514 1.1462 16.0006 144.9817 0.00048133 -83.8678 0.083866
0.18762 0.98801 5.5245e-05 3.8182 0.012048 2.4734e-06 0.001154 0.054456 0.00065302 0.055104 0.049029 0 0.044273 0.0389 0 0.84743 0.22793 0.059127 0.008378 4.1061 0.052743 6.2915e-05 0.83732 0.0051046 0.0058425 0.0018602 0.97969 0.86179 4.0866e-06 1.6349e-05 0.13045 0.66056 0.71815 0.0016308 0.68584 0.48805 0.0021897 0.42207 1.153 1.1478 16.0007 144.9817 0.0004802 -83.8853 0.084595
0.18834 0.98801 5.5245e-05 3.8182 0.012048 2.483e-06 0.001154 0.054562 0.00065304 0.05521 0.049126 0 0.044264 0.0389 0 0.84744 0.22794 0.059129 0.0083783 4.1061 0.052744 6.2917e-05 0.83732 0.0051046 0.0058425 0.0018551 0.97985 0.86703 4.0745e-06 1.63e-05 0.13045 0.66129 0.7189 0.0016284 0.68707 0.48817 0.0021864 0.42207 1.1546 1.1494 16.0007 144.9817 0.00047907 -83.902 0.085324
0.18907 0.98801 5.5244e-05 3.8182 0.012048 2.4926e-06 0.001154 0.054668 0.00065306 0.055316 0.049222 0 0.044254 0.0389 0 0.84746 0.22794 0.059132 0.0083786 4.1061 0.052746 6.2919e-05 0.83732 0.0051046 0.0058426 0.00185 0.98 0.87207 4.0629e-06 1.6254e-05 0.13045 0.66201 0.71965 0.0016261 0.6883 0.4883 0.0021833 0.42206 1.1562 1.151 16.0008 144.9817 0.00047794 -83.918 0.086053
0.1898 0.98801 5.5244e-05 3.8182 0.012047 2.5022e-06 0.001154 0.054773 0.00065307 0.055422 0.049318 0 0.044245 0.0389 0 0.84748 0.22795 0.059134 0.008379 4.1062 0.052747 6.292e-05 0.83732 0.0051046 0.0058426 0.0018455 0.98014 0.87691 4.0518e-06 1.6209e-05 0.13045 0.66274 0.72039 0.0016239 0.68953 0.48842 0.0021802 0.42206 1.1577 1.1526 16.0008 144.9817 0.00047682 -83.9335 0.086782
0.19053 0.98801 5.5244e-05 3.8182 0.012047 2.5118e-06 0.001154 0.054879 0.00065309 0.055527 0.049414 0 0.044235 0.0389 0 0.84749 0.22796 0.059137 0.0083793 4.1062 0.052748 6.2922e-05 0.83731 0.0051046 0.0058426 0.0018407 0.98026 0.88155 4.0412e-06 1.6167e-05 0.13045 0.66346 0.72112 0.0016218 0.69075 0.48854 0.0021773 0.42206 1.1593 1.1542 16.0009 144.9817 0.0004757 -83.9483 0.087511
0.19126 0.98801 5.5244e-05 3.8182 0.012047 2.5214e-06 0.001154 0.054985 0.00065311 0.055633 0.04951 0 0.044226 0.0389 0 0.84751 0.22796 0.05914 0.0083796 4.1062 0.05275 6.2924e-05 0.83731 0.0051046 0.0058426 0.0018366 0.98038 0.886 4.0309e-06 1.6125e-05 0.13045 0.66418 0.72186 0.0016197 0.69197 0.48867 0.0021746 0.42205 1.1609 1.1558 16.001 144.9817 0.00047459 -83.9626 0.08824
0.19199 0.98801 5.5244e-05 3.8182 0.012047 2.531e-06 0.001154 0.05509 0.00065312 0.055739 0.049606 0 0.044216 0.0389 0 0.84752 0.22797 0.059142 0.0083799 4.1062 0.052751 6.2926e-05 0.83731 0.0051047 0.0058426 0.0018321 0.98048 0.89028 4.021e-06 1.6086e-05 0.13045 0.6649 0.72259 0.0016178 0.69319 0.48879 0.0021719 0.42205 1.1624 1.1573 16.001 144.9818 0.00047348 -83.9765 0.088969
0.19272 0.98801 5.5244e-05 3.8182 0.012047 2.5406e-06 0.001154 0.055196 0.00065314 0.055844 0.049703 0 0.044207 0.0389 0 0.84754 0.22798 0.059145 0.0083802 4.1062 0.052753 6.2927e-05 0.83731 0.0051047 0.0058426 0.0018283 0.98058 0.89438 4.0115e-06 1.6048e-05 0.13045 0.66562 0.72331 0.0016159 0.6944 0.48891 0.0021693 0.42205 1.164 1.1589 16.0011 144.9818 0.00047238 -83.9898 0.089698
0.19345 0.98801 5.5244e-05 3.8182 0.012047 2.5502e-06 0.001154 0.055301 0.00065316 0.05595 0.049799 0 0.044198 0.0389 0 0.84756 0.22799 0.059147 0.0083806 4.1062 0.052754 6.2929e-05 0.83731 0.0051047 0.0058427 0.0018241 0.98067 0.89832 4.0023e-06 1.6011e-05 0.13045 0.66633 0.72404 0.001614 0.69561 0.48903 0.0021668 0.42205 1.1656 1.1605 16.0011 144.9818 0.00047128 -84.0028 0.090427
0.19418 0.98801 5.5244e-05 3.8182 0.012047 2.5598e-06 0.001154 0.055406 0.00065317 0.056055 0.049894 0 0.044188 0.0389 0 0.84757 0.22799 0.05915 0.0083809 4.1062 0.052756 6.2931e-05 0.83731 0.0051047 0.0058427 0.0018207 0.98076 0.9021 3.9934e-06 1.5975e-05 0.13045 0.66705 0.72476 0.0016122 0.69682 0.48916 0.0021644 0.42205 1.1671 1.1621 16.0012 144.9818 0.00047019 -84.0153 0.091156
0.19491 0.98801 5.5244e-05 3.8182 0.012047 2.5694e-06 0.001154 0.055512 0.00065319 0.05616 0.04999 0 0.044179 0.0389 0 0.84759 0.228 0.059152 0.0083812 4.1062 0.052757 6.2933e-05 0.83731 0.0051047 0.0058427 0.0018166 0.98084 0.90572 3.9848e-06 1.5941e-05 0.13045 0.66776 0.72547 0.0016105 0.69802 0.48928 0.0021621 0.42204 1.1687 1.1636 16.0012 144.9818 0.0004691 -84.0275 0.091885
0.19563 0.98801 5.5244e-05 3.8182 0.012047 2.579e-06 0.001154 0.055617 0.00065321 0.056265 0.050086 0 0.044169 0.0389 0 0.84761 0.22801 0.059155 0.0083815 4.1062 0.052758 6.2935e-05 0.8373 0.0051047 0.0058427 0.0018135 0.98091 0.9092 3.9764e-06 1.5907e-05 0.13045 0.66847 0.72619 0.0016088 0.69922 0.4894 0.0021598 0.42204 1.1702 1.1652 16.0013 144.9818 0.00046801 -84.0394 0.092614
0.19636 0.98801 5.5244e-05 3.8182 0.012047 2.5886e-06 0.001154 0.055722 0.00065322 0.056371 0.050182 0 0.04416 0.0389 0 0.84762 0.22801 0.059158 0.0083819 4.1063 0.05276 6.2936e-05 0.8373 0.0051048 0.0058427 0.0018094 0.98098 0.91253 3.9683e-06 1.5875e-05 0.13045 0.66918 0.72689 0.0016072 0.70042 0.48953 0.0021576 0.42204 1.1718 1.1668 16.0014 144.9818 0.00046693 -84.051 0.093343
0.19709 0.98801 5.5244e-05 3.8182 0.012047 2.5983e-06 0.001154 0.055827 0.00065324 0.056476 0.050278 0 0.044151 0.0389 0 0.84764 0.22802 0.05916 0.0083822 4.1063 0.052761 6.2938e-05 0.8373 0.0051048 0.0058427 0.0018067 0.98105 0.91573 3.9604e-06 1.5843e-05 0.13045 0.66989 0.7276 0.0016056 0.70161 0.48965 0.0021555 0.42204 1.1733 1.1683 16.0014 144.9818 0.00046585 -84.0622 0.094072
0.19782 0.98801 5.5244e-05 3.8182 0.012047 2.6079e-06 0.001154 0.055932 0.00065326 0.056581 0.050373 0 0.044141 0.0389 0 0.84765 0.22803 0.059163 0.0083825 4.1063 0.052763 6.294e-05 0.8373 0.0051048 0.0058428 0.0018032 0.98111 0.9188 3.9527e-06 1.5812e-05 0.13045 0.6706 0.7283 0.0016041 0.7028 0.48977 0.0021534 0.42204 1.1749 1.1699 16.0015 144.9818 0.00046478 -84.0732 0.094801
0.19855 0.98801 5.5244e-05 3.8182 0.012047 2.6175e-06 0.001154 0.056037 0.00065327 0.056686 0.050469 0 0.044132 0.0389 0 0.84767 0.22804 0.059165 0.0083829 4.1063 0.052764 6.2942e-05 0.8373 0.0051048 0.0058428 0.0018001 0.98117 0.92175 3.9452e-06 1.5782e-05 0.13045 0.67131 0.729 0.0016026 0.70399 0.48989 0.0021514 0.42203 1.1764 1.1715 16.0015 144.9818 0.00046371 -84.084 0.09553
0.19928 0.98801 5.5244e-05 3.8182 0.012047 2.6271e-06 0.001154 0.056142 0.00065329 0.056791 0.050565 0 0.044122 0.0389 0 0.84769 0.22804 0.059168 0.0083832 4.1063 0.052766 6.2944e-05 0.8373 0.0051048 0.0058428 0.0017965 0.98123 0.92457 3.9378e-06 1.5753e-05 0.13045 0.67201 0.7297 0.0016011 0.70517 0.49002 0.0021494 0.42203 1.178 1.173 16.0016 144.9818 0.00046264 -84.0945 0.096259
0.20001 0.98801 5.5244e-05 3.8182 0.012047 2.6367e-06 0.001154 0.056247 0.0006533 0.056896 0.05066 0 0.044113 0.0389 0 0.8477 0.22805 0.059171 0.0083835 4.1063 0.052767 6.2946e-05 0.8373 0.0051048 0.0058428 0.0017938 0.98128 0.92728 3.9306e-06 1.5724e-05 0.13045 0.67271 0.73039 0.0015996 0.70635 0.49014 0.0021475 0.42203 1.1795 1.1746 16.0016 144.9818 0.00046158 -84.1048 0.096988
0.20074 0.98801 5.5244e-05 3.8182 0.012047 2.6463e-06 0.001154 0.056352 0.00065332 0.057001 0.050756 0 0.044104 0.0389 0 0.84772 0.22806 0.059173 0.0083839 4.1063 0.052769 6.2948e-05 0.83729 0.0051049 0.0058428 0.0017906 0.98134 0.92987 3.9236e-06 1.5696e-05 0.13045 0.67341 0.73108 0.0015982 0.70753 0.49026 0.0021456 0.42203 1.1811 1.1761 16.0017 144.9818 0.00046053 -84.1149 0.097717
0.20147 0.98801 5.5244e-05 3.8182 0.012047 2.6559e-06 0.001154 0.056457 0.00065333 0.057105 0.050851 0 0.044094 0.0389 0 0.84774 0.22807 0.059176 0.0083842 4.1064 0.05277 6.295e-05 0.83729 0.0051049 0.0058428 0.0017879 0.98139 0.93236 3.9167e-06 1.5668e-05 0.13045 0.67411 0.73176 0.0015968 0.7087 0.49039 0.0021437 0.42203 1.1826 1.1777 16.0018 144.9818 0.00045947 -84.1248 0.098446
0.2022 0.98801 5.5244e-05 3.8182 0.012047 2.6655e-06 0.001154 0.056561 0.00065335 0.05721 0.050946 0 0.044085 0.0389 0 0.84775 0.22807 0.059179 0.0083846 4.1064 0.052772 6.2951e-05 0.83729 0.0051049 0.0058429 0.0017846 0.98144 0.93475 3.91e-06 1.5641e-05 0.13045 0.67481 0.73245 0.0015955 0.70987 0.49051 0.0021419 0.42203 1.1841 1.1792 16.0018 144.9818 0.00045843 -84.1346 0.099175
0.20292 0.98801 5.5244e-05 3.8182 0.012047 2.6751e-06 0.001154 0.056666 0.00065337 0.057315 0.051042 0 0.044076 0.0389 0 0.84777 0.22808 0.059181 0.0083849 4.1064 0.052773 6.2953e-05 0.83729 0.0051049 0.0058429 0.0017821 0.98149 0.93703 3.9033e-06 1.5614e-05 0.13045 0.67551 0.73312 0.0015941 0.71104 0.49063 0.0021402 0.42203 1.1857 1.1808 16.0019 144.9818 0.00045738 -84.1442 0.099904
0.20365 0.98801 5.5244e-05 3.8182 0.012047 2.6847e-06 0.001154 0.05677 0.00065338 0.057419 0.051137 0 0.044066 0.0389 0 0.84779 0.22809 0.059184 0.0083852 4.1064 0.052775 6.2955e-05 0.83729 0.0051049 0.0058429 0.0017789 0.98153 0.93923 3.8968e-06 1.5588e-05 0.13046 0.6762 0.7338 0.0015928 0.7122 0.49076 0.0021384 0.42203 1.1872 1.1823 16.0019 144.9819 0.00045634 -84.1536 0.10063
0.20438 0.98801 5.5244e-05 3.8182 0.012047 2.6943e-06 0.001154 0.056875 0.0006534 0.057524 0.051232 0 0.044057 0.0389 0 0.84781 0.2281 0.059187 0.0083856 4.1064 0.052776 6.2957e-05 0.83729 0.005105 0.0058429 0.0017763 0.98158 0.94133 3.8904e-06 1.5563e-05 0.13046 0.67689 0.73447 0.0015915 0.71336 0.49088 0.0021367 0.42203 1.1887 1.1839 16.002 144.9819 0.00045531 -84.1629 0.10136
0.20511 0.98801 5.5243e-05 3.8182 0.012047 2.7039e-06 0.001154 0.056979 0.00065341 0.057628 0.051327 0 0.044048 0.0389 0 0.84782 0.2281 0.05919 0.0083859 4.1064 0.052778 6.2959e-05 0.83729 0.005105 0.0058429 0.0017735 0.98162 0.94335 3.8841e-06 1.5538e-05 0.13046 0.67759 0.73514 0.0015902 0.71451 0.491 0.002135 0.42203 1.1903 1.1854 16.002 144.9819 0.00045428 -84.172 0.10209
0.20584 0.98801 5.5243e-05 3.8182 0.012047 2.7135e-06 0.001154 0.057084 0.00065343 0.057733 0.051422 0 0.044039 0.0389 0 0.84784 0.22811 0.059192 0.0083863 4.1064 0.052779 6.2961e-05 0.83728 0.005105 0.0058429 0.0017712 0.98166 0.94528 3.878e-06 1.5513e-05 0.13046 0.67828 0.73581 0.001589 0.71566 0.49112 0.0021333 0.42202 1.1918 1.1869 16.0021 144.9819 0.00045325 -84.181 0.10282
0.20657 0.98801 5.5243e-05 3.8182 0.012047 2.7231e-06 0.001154 0.057188 0.00065344 0.057837 0.051517 0 0.044029 0.0389 0 0.84786 0.22812 0.059195 0.0083866 4.1064 0.052781 6.2963e-05 0.83728 0.005105 0.005843 0.0017683 0.9817 0.94713 3.8719e-06 1.5488e-05 0.13046 0.67897 0.73647 0.0015878 0.71681 0.49125 0.0021317 0.42202 1.1933 1.1885 16.0021 144.9819 0.00045222 -84.1899 0.10355
0.2073 0.98801 5.5243e-05 3.8182 0.012047 2.7328e-06 0.001154 0.057292 0.00065346 0.057941 0.051612 0 0.04402 0.0389 0 0.84787 0.22813 0.059198 0.0083869 4.1065 0.052782 6.2965e-05 0.83728 0.005105 0.005843 0.0017658 0.98174 0.94891 3.8658e-06 1.5464e-05 0.13046 0.67965 0.73713 0.0015865 0.71795 0.49137 0.0021301 0.42202 1.1948 1.19 16.0022 144.9819 0.0004512 -84.1987 0.10428
0.20803 0.98801 5.5243e-05 3.8182 0.012047 2.7424e-06 0.001154 0.057397 0.00065347 0.058045 0.051707 0 0.044011 0.0389 0 0.84789 0.22813 0.0592 0.0083873 4.1065 0.052784 6.2967e-05 0.83728 0.005105 0.005843 0.0017631 0.98178 0.95061 3.8599e-06 1.5441e-05 0.13046 0.68034 0.73779 0.0015853 0.71909 0.49149 0.0021285 0.42202 1.1964 1.1915 16.0023 144.9819 0.00045019 -84.2074 0.10501
0.20876 0.98801 5.5243e-05 3.8182 0.012047 2.752e-06 0.001154 0.057501 0.00065349 0.05815 0.051802 0 0.044002 0.0389 0 0.84791 0.22814 0.059203 0.0083876 4.1065 0.052785 6.2969e-05 0.83728 0.0051051 0.005843 0.0017609 0.98182 0.95224 3.8541e-06 1.5417e-05 0.13046 0.68102 0.73844 0.0015841 0.72023 0.49162 0.0021269 0.42202 1.1979 1.1931 16.0023 144.9819 0.00044918 -84.2159 0.10574
0.20949 0.98801 5.5243e-05 3.8182 0.012047 2.7616e-06 0.001154 0.057605 0.0006535 0.058254 0.051897 0 0.043992 0.0389 0 0.84793 0.22815 0.059206 0.008388 4.1065 0.052787 6.2971e-05 0.83728 0.0051051 0.005843 0.0017582 0.98186 0.95381 3.8483e-06 1.5394e-05 0.13046 0.6817 0.73909 0.001583 0.72136 0.49174 0.0021254 0.42202 1.1994 1.1946 16.0024 144.9819 0.00044817 -84.2244 0.10647
0.21021 0.98801 5.5243e-05 3.8182 0.012047 2.7712e-06 0.001154 0.057709 0.00065352 0.058358 0.051992 0 0.043983 0.0389 0 0.84794 0.22816 0.059209 0.0083883 4.1065 0.052789 6.2973e-05 0.83727 0.0051051 0.0058431 0.0017561 0.9819 0.9553 3.8426e-06 1.5371e-05 0.13046 0.68239 0.73974 0.0015818 0.72249 0.49186 0.0021239 0.42202 1.2009 1.1961 16.0024 144.9819 0.00044717 -84.2327 0.10719
0.21094 0.98801 5.5243e-05 3.8182 0.012047 2.7808e-06 0.001154 0.057813 0.00065353 0.058462 0.052087 0 0.043974 0.0389 0 0.84796 0.22816 0.059211 0.0083887 4.1065 0.05279 6.2975e-05 0.83727 0.0051051 0.0058431 0.0017535 0.98193 0.95674 3.837e-06 1.5349e-05 0.13046 0.68307 0.74039 0.0015807 0.72361 0.49199 0.0021224 0.42202 1.2024 1.1977 16.0025 144.9819 0.00044617 -84.241 0.10792
0.21167 0.98801 5.5243e-05 3.8182 0.012047 2.7904e-06 0.001154 0.057917 0.00065355 0.058566 0.052181 0 0.043965 0.0389 0 0.84798 0.22817 0.059214 0.008389 4.1065 0.052792 6.2977e-05 0.83727 0.0051051 0.0058431 0.0017512 0.98197 0.95812 3.8314e-06 1.5327e-05 0.13046 0.68374 0.74103 0.0015795 0.72473 0.49211 0.0021209 0.42202 1.2039 1.1992 16.0025 144.9819 0.00044517 -84.2492 0.10865
0.2124 0.98801 5.5243e-05 3.8182 0.012047 2.8e-06 0.001154 0.05802 0.00065356 0.058669 0.052276 0 0.043955 0.0389 0 0.848 0.22818 0.059217 0.0083894 4.1066 0.052793 6.2979e-05 0.83727 0.0051052 0.0058431 0.0017486 0.98201 0.95944 3.8259e-06 1.5305e-05 0.13046 0.68442 0.74167 0.0015784 0.72585 0.49223 0.0021194 0.42202 1.2054 1.2007 16.0026 144.9819 0.00044418 -84.2573 0.10938
0.21313 0.98801 5.5243e-05 3.8182 0.012047 2.8096e-06 0.001154 0.058124 0.00065358 0.058773 0.05237 0 0.043946 0.0389 0 0.84801 0.22819 0.05922 0.0083897 4.1066 0.052795 6.2981e-05 0.83727 0.0051052 0.0058431 0.0017465 0.98204 0.9607 3.8205e-06 1.5283e-05 0.13046 0.6851 0.7423 0.0015773 0.72697 0.49236 0.0021179 0.42202 1.2069 1.2022 16.0026 144.9819 0.00044319 -84.2654 0.11011
0.21386 0.98801 5.5243e-05 3.8182 0.012047 2.8192e-06 0.001154 0.058228 0.00065359 0.058877 0.052465 0 0.043937 0.0389 0 0.84803 0.2282 0.059223 0.0083901 4.1066 0.052797 6.2983e-05 0.83727 0.0051052 0.0058431 0.0017441 0.98207 0.96191 3.8151e-06 1.5261e-05 0.13046 0.68577 0.74293 0.0015762 0.72808 0.49248 0.0021165 0.42202 1.2084 1.2037 16.0027 144.9819 0.00044221 -84.2733 0.11084
0.21459 0.98801 5.5243e-05 3.8182 0.012047 2.8288e-06 0.001154 0.058332 0.00065361 0.058981 0.052559 0 0.043928 0.0389 0 0.84805 0.2282 0.059225 0.0083905 4.1066 0.052798 6.2985e-05 0.83726 0.0051052 0.0058432 0.001742 0.98211 0.96307 3.8098e-06 1.524e-05 0.13046 0.68644 0.74357 0.0015751 0.72918 0.4926 0.0021151 0.42202 1.2099 1.2052 16.0027 144.982 0.00044123 -84.2812 0.11157
0.21532 0.98801 5.5243e-05 3.8182 0.012047 2.8384e-06 0.001154 0.058435 0.00065362 0.059084 0.052654 0 0.043919 0.0389 0 0.84807 0.22821 0.059228 0.0083908 4.1066 0.0528 6.2987e-05 0.83726 0.0051052 0.0058432 0.0017394 0.98214 0.96419 3.8045e-06 1.5219e-05 0.13046 0.68711 0.74419 0.001574 0.73029 0.49272 0.0021137 0.42202 1.2114 1.2067 16.0028 144.982 0.00044025 -84.2891 0.1123
0.21605 0.98801 5.5243e-05 3.8182 0.012047 2.848e-06 0.001154 0.058539 0.00065363 0.059188 0.052748 0 0.04391 0.0389 0 0.84809 0.22822 0.059231 0.0083912 4.1066 0.052801 6.2989e-05 0.83726 0.0051053 0.0058432 0.0017375 0.98217 0.96525 3.7993e-06 1.5198e-05 0.13046 0.68778 0.74482 0.001573 0.73139 0.49285 0.0021122 0.42202 1.2129 1.2083 16.0028 144.982 0.00043928 -84.2968 0.11303
0.21678 0.98801 5.5243e-05 3.8182 0.012047 2.8576e-06 0.001154 0.058642 0.00065365 0.059291 0.052843 0 0.0439 0.0389 0 0.8481 0.22823 0.059234 0.0083915 4.1066 0.052803 6.2991e-05 0.83726 0.0051053 0.0058432 0.0017348 0.98221 0.96628 3.7941e-06 1.5177e-05 0.13046 0.68845 0.74544 0.0015719 0.73248 0.49297 0.0021109 0.42202 1.2144 1.2098 16.0029 144.982 0.00043831 -84.3045 0.11376
0.2175 0.98801 5.5243e-05 3.8182 0.012047 2.8672e-06 0.001154 0.058746 0.00065366 0.059395 0.052937 0 0.043891 0.0389 0 0.84812 0.22823 0.059237 0.0083919 4.1067 0.052805 6.2993e-05 0.83726 0.0051053 0.0058432 0.0017328 0.98224 0.96725 3.789e-06 1.5157e-05 0.13046 0.68911 0.74606 0.0015709 0.73357 0.49309 0.0021095 0.42202 1.2159 1.2113 16.0029 144.982 0.00043734 -84.3121 0.11448
0.21823 0.98801 5.5243e-05 3.8182 0.012047 2.8769e-06 0.001154 0.058849 0.00065368 0.059498 0.053031 0 0.043882 0.0389 0 0.84814 0.22824 0.05924 0.0083922 4.1067 0.052806 6.2996e-05 0.83726 0.0051053 0.0058433 0.0017305 0.98227 0.96819 3.7839e-06 1.5136e-05 0.13046 0.68978 0.74667 0.0015698 0.73466 0.49322 0.0021081 0.42202 1.2174 1.2128 16.003 144.982 0.00043638 -84.3197 0.11521
0.21923 0.98801 5.5243e-05 3.8182 0.012047 2.89e-06 0.001154 0.058991 0.0006537 0.05964 0.05316 0 0.04387 0.0389 0 0.84816 0.22825 0.059244 0.0083927 4.1067 0.052809 6.2998e-05 0.83725 0.0051053 0.0058433 0.0017276 0.98231 0.96942 3.777e-06 1.5109e-05 0.13046 0.69069 0.74751 0.0015684 0.73615 0.49339 0.0021063 0.42202 1.2195 1.2148 16.003 144.982 0.00043507 -84.33 0.11621
0.22023 0.98801 5.5243e-05 3.8182 0.012047 2.9032e-06 0.001154 0.059132 0.00065371 0.059781 0.053289 0 0.043857 0.0389 0 0.84819 0.22826 0.059248 0.0083932 4.1067 0.052811 6.3001e-05 0.83725 0.0051054 0.0058433 0.0017248 0.98236 0.97057 3.7702e-06 1.5082e-05 0.13046 0.6916 0.74835 0.001567 0.73763 0.49355 0.0021044 0.42202 1.2215 1.2169 16.0031 144.982 0.00043376 -84.3401 0.11721
0.22123 0.98801 5.5242e-05 3.8182 0.012047 2.9164e-06 0.001154 0.059274 0.00065373 0.059923 0.053418 0 0.043845 0.0389 0 0.84821 0.22828 0.059252 0.0083937 4.1067 0.052813 6.3004e-05 0.83725 0.0051054 0.0058433 0.0017219 0.9824 0.97166 3.7635e-06 1.5055e-05 0.13046 0.6925 0.74918 0.0015656 0.7391 0.49372 0.0021026 0.42203 1.2235 1.2189 16.0032 144.982 0.00043246 -84.3502 0.11821
0.22223 0.98801 5.5242e-05 3.8182 0.012047 2.9296e-06 0.001154 0.059415 0.00065375 0.060064 0.053547 0 0.043832 0.0389 0 0.84824 0.22829 0.059255 0.0083942 4.1068 0.052816 6.3007e-05 0.83725 0.0051054 0.0058434 0.0017191 0.98244 0.97269 3.7569e-06 1.5028e-05 0.13046 0.6934 0.75 0.0015643 0.74057 0.49389 0.0021008 0.42203 1.2256 1.221 16.0032 144.982 0.00043117 -84.3602 0.11921
0.22323 0.98801 5.5242e-05 3.8182 0.012047 2.9427e-06 0.001154 0.059556 0.00065377 0.060205 0.053676 0 0.04382 0.0389 0 0.84826 0.2283 0.059259 0.0083947 4.1068 0.052818 6.301e-05 0.83725 0.0051055 0.0058434 0.0017163 0.98248 0.97366 3.7503e-06 1.5002e-05 0.13046 0.6943 0.75082 0.0015629 0.74203 0.49406 0.0020991 0.42203 1.2276 1.223 16.0033 144.982 0.00042988 -84.3701 0.12021
0.22423 0.98801 5.5242e-05 3.8182 0.012047 2.9559e-06 0.001154 0.059697 0.00065379 0.060346 0.053805 0 0.043807 0.0389 0 0.84829 0.22831 0.059263 0.0083953 4.1068 0.05282 6.3013e-05 0.83724 0.0051055 0.0058434 0.0017136 0.98252 0.97457 3.7438e-06 1.4976e-05 0.13046 0.69519 0.75164 0.0015616 0.74348 0.49423 0.0020973 0.42203 1.2296 1.225 16.0034 144.9821 0.00042861 -84.3799 0.12121
0.22523 0.98801 5.5242e-05 3.8182 0.012047 2.9691e-06 0.001154 0.059838 0.00065381 0.060487 0.053933 0 0.043795 0.0389 0 0.84831 0.22832 0.059268 0.0083958 4.1068 0.052823 6.3016e-05 0.83724 0.0051055 0.0058435 0.0017106 0.98256 0.97543 3.7374e-06 1.495e-05 0.13046 0.69609 0.75245 0.0015602 0.74493 0.4944 0.0020956 0.42203 1.2316 1.2271 16.0034 144.9821 0.00042733 -84.3895 0.12221
0.22623 0.98801 5.5242e-05 3.8182 0.012047 2.9823e-06 0.001154 0.059979 0.00065383 0.060628 0.054062 0 0.043783 0.0389 0 0.84834 0.22833 0.059272 0.0083963 4.1069 0.052825 6.3019e-05 0.83724 0.0051056 0.0058435 0.0017083 0.9826 0.97624 3.7311e-06 1.4925e-05 0.13046 0.69698 0.75325 0.0015589 0.74637 0.49457 0.0020939 0.42203 1.2336 1.2291 16.0035 144.9821 0.00042607 -84.3992 0.12321
0.22723 0.98801 5.5242e-05 3.8182 0.012047 2.9954e-06 0.001154 0.06012 0.00065385 0.060769 0.05419 0 0.04377 0.0389 0 0.84837 0.22834 0.059276 0.0083968 4.1069 0.052827 6.3022e-05 0.83724 0.0051056 0.0058435 0.0017045 0.98264 0.97701 3.7248e-06 1.49e-05 0.13046 0.69787 0.75405 0.0015576 0.7478 0.49474 0.0020922 0.42203 1.2356 1.2311 16.0036 144.9821 0.00042481 -84.4087 0.12421
0.22823 0.98801 5.5242e-05 3.8182 0.012047 3.0086e-06 0.001154 0.060261 0.00065386 0.06091 0.054318 0 0.043758 0.0389 0 0.84839 0.22835 0.05928 0.0083973 4.1069 0.05283 6.3025e-05 0.83723 0.0051056 0.0058435 0.001702 0.98267 0.97773 3.7186e-06 1.4875e-05 0.13046 0.69875 0.75485 0.0015564 0.74923 0.49491 0.0020905 0.42204 1.2376 1.2331 16.0036 144.9821 0.00042356 -84.4181 0.12521
0.22923 0.98801 5.5242e-05 3.8182 0.012047 3.0218e-06 0.001154 0.060401 0.00065388 0.06105 0.054447 0 0.043746 0.0389 0 0.84842 0.22837 0.059284 0.0083978 4.1069 0.052832 6.3028e-05 0.83723 0.0051056 0.0058436 0.0016997 0.98271 0.97842 3.7124e-06 1.485e-05 0.13046 0.69963 0.75564 0.0015551 0.75065 0.49507 0.0020888 0.42204 1.2396 1.2352 16.0037 144.9821 0.00042231 -84.4275 0.12621
0.23023 0.98801 5.5242e-05 3.8182 0.012047 3.035e-06 0.001154 0.060541 0.0006539 0.061191 0.054575 0 0.043733 0.0389 0 0.84844 0.22838 0.059288 0.0083983 4.1069 0.052835 6.3031e-05 0.83723 0.0051057 0.0058436 0.0016972 0.98275 0.97906 3.7063e-06 1.4826e-05 0.13046 0.70051 0.75642 0.0015538 0.75206 0.49524 0.0020872 0.42204 1.2416 1.2372 16.0038 144.9821 0.00042107 -84.4367 0.12721
0.23123 0.98801 5.5242e-05 3.8182 0.012047 3.0482e-06 0.001154 0.060682 0.00065392 0.061331 0.054703 0 0.043721 0.0389 0 0.84847 0.22839 0.059292 0.0083988 4.107 0.052837 6.3034e-05 0.83723 0.0051057 0.0058436 0.0016949 0.98278 0.97967 3.7003e-06 1.4802e-05 0.13046 0.70139 0.7572 0.0015526 0.75346 0.49541 0.0020855 0.42204 1.2436 1.2392 16.0038 144.9821 0.00041984 -84.4459 0.12821
0.23223 0.98801 5.5242e-05 3.8182 0.012047 3.0613e-06 0.001154 0.060822 0.00065394 0.061471 0.054831 0 0.043709 0.0389 0 0.8485 0.2284 0.059296 0.0083994 4.107 0.052839 6.3037e-05 0.83722 0.0051057 0.0058437 0.0016923 0.98282 0.98024 3.6944e-06 1.4778e-05 0.13046 0.70226 0.75798 0.0015513 0.75486 0.49558 0.0020839 0.42204 1.2456 1.2412 16.0039 144.9821 0.00041862 -84.455 0.12921
0.23323 0.98801 5.5242e-05 3.8182 0.012047 3.0745e-06 0.001154 0.060962 0.00065395 0.061611 0.054958 0 0.043696 0.0389 0 0.84852 0.22841 0.0593 0.0083999 4.107 0.052842 6.304e-05 0.83722 0.0051058 0.0058437 0.00169 0.98286 0.98078 3.6885e-06 1.4755e-05 0.13046 0.70313 0.75875 0.0015501 0.75625 0.49575 0.0020823 0.42205 1.2476 1.2432 16.004 144.9822 0.0004174 -84.4641 0.13021
0.23423 0.98801 5.5242e-05 3.8182 0.012047 3.0877e-06 0.001154 0.061102 0.00065397 0.061751 0.055086 0 0.043684 0.0389 0 0.84855 0.22842 0.059304 0.0084004 4.107 0.052844 6.3044e-05 0.83722 0.0051058 0.0058437 0.0016867 0.98289 0.98129 3.6826e-06 1.4731e-05 0.13046 0.704 0.75952 0.0015489 0.75764 0.49592 0.0020807 0.42205 1.2496 1.2452 16.004 144.9822 0.00041618 -84.473 0.13121
0.23523 0.98801 5.5242e-05 3.8182 0.012047 3.1009e-06 0.001154 0.061242 0.00065399 0.061891 0.055214 0 0.043672 0.0389 0 0.84857 0.22843 0.059309 0.0084009 4.1071 0.052847 6.3047e-05 0.83722 0.0051058 0.0058438 0.0016856 0.98293 0.98177 3.6769e-06 1.4708e-05 0.13046 0.70487 0.76028 0.0015477 0.75902 0.49609 0.0020792 0.42205 1.2515 1.2472 16.0041 144.9822 0.00041498 -84.4819 0.13221
0.23623 0.98801 5.5242e-05 3.8182 0.012047 3.114e-06 0.001154 0.061382 0.00065401 0.062031 0.055341 0 0.04366 0.0389 0 0.8486 0.22845 0.059313 0.0084015 4.1071 0.052849 6.305e-05 0.83721 0.0051059 0.0058438 0.001683 0.98296 0.98223 3.6711e-06 1.4685e-05 0.13046 0.70573 0.76104 0.0015465 0.76039 0.49626 0.0020776 0.42205 1.2535 1.2492 16.0041 144.9822 0.00041378 -84.4907 0.13321
0.23723 0.98801 5.5242e-05 3.8182 0.012047 3.1272e-06 0.001154 0.061521 0.00065402 0.062171 0.055469 0 0.043647 0.0389 0 0.84863 0.22846 0.059317 0.008402 4.1071 0.052852 6.3053e-05 0.83721 0.0051059 0.0058438 0.0016796 0.983 0.98265 3.6654e-06 1.4662e-05 0.13046 0.70659 0.76179 0.0015453 0.76175 0.49642 0.0020761 0.42206 1.2555 1.2511 16.0042 144.9822 0.00041258 -84.4994 0.13421
0.23823 0.98801 5.5241e-05 3.8182 0.012047 3.1404e-06 0.001154 0.061661 0.00065404 0.06231 0.055596 0 0.043635 0.0389 0 0.84865 0.22847 0.059321 0.0084025 4.1071 0.052854 6.3056e-05 0.83721 0.0051059 0.0058439 0.0016782 0.98303 0.98306 3.6598e-06 1.464e-05 0.13046 0.70745 0.76254 0.0015441 0.76311 0.49659 0.0020745 0.42206 1.2574 1.2531 16.0043 144.9822 0.0004114 -84.5081 0.13521
0.23923 0.98801 5.5241e-05 3.8182 0.012047 3.1536e-06 0.001154 0.0618 0.00065406 0.06245 0.055723 0 0.043623 0.0389 0 0.84868 0.22848 0.059325 0.0084031 4.1072 0.052857 6.306e-05 0.83721 0.005106 0.0058439 0.0016745 0.98306 0.98344 3.6543e-06 1.4618e-05 0.13046 0.70831 0.76329 0.001543 0.76446 0.49676 0.002073 0.42206 1.2594 1.2551 16.0043 144.9822 0.00041021 -84.5167 0.13621
0.24023 0.98801 5.5241e-05 3.8182 0.012047 3.1668e-06 0.001154 0.06194 0.00065407 0.062589 0.05585 0 0.043611 0.0389 0 0.84871 0.22849 0.05933 0.0084036 4.1072 0.052859 6.3063e-05 0.8372 0.005106 0.0058439 0.0016729 0.9831 0.9838 3.6488e-06 1.4596e-05 0.13046 0.70916 0.76403 0.0015418 0.76581 0.49693 0.0020715 0.42206 1.2613 1.2571 16.0044 144.9822 0.00040904 -84.5252 0.13721
0.24123 0.98801 5.5241e-05 3.8182 0.012047 3.1799e-06 0.001154 0.062079 0.00065409 0.062728 0.055977 0 0.043599 0.0389 0 0.84873 0.2285 0.059334 0.0084041 4.1072 0.052862 6.3066e-05 0.8372 0.005106 0.0058439 0.0016709 0.98313 0.98414 3.6433e-06 1.4574e-05 0.13046 0.71001 0.76477 0.0015407 0.76715 0.4971 0.00207 0.42207 1.2633 1.259 16.0044 144.9822 0.00040787 -84.5337 0.13821
0.24223 0.98801 5.5241e-05 3.8182 0.012047 3.1931e-06 0.001154 0.062218 0.00065411 0.062867 0.056104 0 0.043587 0.0389 0 0.84876 0.22852 0.059338 0.0084047 4.1072 0.052865 6.3069e-05 0.8372 0.0051061 0.005844 0.0016676 0.98316 0.98446 3.6379e-06 1.4552e-05 0.13046 0.71086 0.7655 0.0015396 0.76848 0.49727 0.0020685 0.42207 1.2652 1.261 16.0045 144.9823 0.00040671 -84.5421 0.13921
0.24323 0.98801 5.5241e-05 3.8182 0.012047 3.2063e-06 0.001154 0.062357 0.00065412 0.063006 0.056231 0 0.043574 0.0389 0 0.84879 0.22853 0.059342 0.0084052 4.1073 0.052867 6.3072e-05 0.8372 0.0051061 0.005844 0.0016651 0.9832 0.98477 3.6325e-06 1.4531e-05 0.13046 0.7117 0.76623 0.0015384 0.76981 0.49744 0.0020671 0.42207 1.2672 1.2629 16.0046 144.9823 0.00040555 -84.5504 0.14021
0.24423 0.98801 5.5241e-05 3.8182 0.012047 3.2195e-06 0.001154 0.062496 0.00065414 0.063145 0.056358 0 0.043562 0.0389 0 0.84882 0.22854 0.059347 0.0084058 4.1073 0.05287 6.3076e-05 0.83719 0.0051061 0.005844 0.0016633 0.98323 0.98505 3.6272e-06 1.451e-05 0.13046 0.71255 0.76695 0.0015373 0.77112 0.49761 0.0020656 0.42208 1.2691 1.2649 16.0046 144.9823 0.0004044 -84.5586 0.14121
0.24523 0.98801 5.5241e-05 3.8182 0.012047 3.2326e-06 0.001154 0.062634 0.00065416 0.063284 0.056485 0 0.04355 0.0389 0 0.84884 0.22855 0.059351 0.0084063 4.1073 0.052872 6.3079e-05 0.83719 0.0051062 0.0058441 0.0016603 0.98326 0.98532 3.622e-06 1.4488e-05 0.13047 0.71339 0.76767 0.0015362 0.77244 0.49777 0.0020642 0.42208 1.2711 1.2668 16.0047 144.9823 0.00040325 -84.5668 0.14221
0.24623 0.98801 5.5241e-05 3.8182 0.012047 3.2458e-06 0.001154 0.062773 0.00065417 0.063423 0.056611 0 0.043538 0.0389 0 0.84887 0.22856 0.059355 0.0084069 4.1073 0.052875 6.3082e-05 0.83719 0.0051062 0.0058441 0.0016582 0.98329 0.98558 3.6168e-06 1.4468e-05 0.13047 0.71422 0.76838 0.0015351 0.77374 0.49794 0.0020627 0.42208 1.273 1.2688 16.0047 144.9823 0.00040211 -84.575 0.14321
0.24723 0.98801 5.5241e-05 3.8182 0.012047 3.259e-06 0.001154 0.062912 0.00065419 0.063561 0.056738 0 0.043526 0.0389 0 0.8489 0.22858 0.05936 0.0084074 4.1074 0.052878 6.3086e-05 0.83719 0.0051062 0.0058441 0.0016564 0.98332 0.98582 3.6116e-06 1.4447e-05 0.13047 0.71506 0.7691 0.0015341 0.77504 0.49811 0.0020613 0.42209 1.2749 1.2707 16.0048 144.9823 0.00040098 -84.583 0.14421
0.24823 0.98801 5.5241e-05 3.8182 0.012047 3.2722e-06 0.001154 0.06305 0.00065421 0.0637 0.056864 0 0.043514 0.0389 0 0.84892 0.22859 0.059364 0.008408 4.1074 0.05288 6.3089e-05 0.83718 0.0051063 0.0058442 0.001654 0.98335 0.98605 3.6065e-06 1.4427e-05 0.13047 0.71589 0.7698 0.001533 0.77633 0.49828 0.0020599 0.42209 1.2768 1.2726 16.0048 144.9823 0.00039985 -84.591 0.14521
0.24923 0.98801 5.5241e-05 3.8182 0.012047 3.2853e-06 0.001154 0.063188 0.00065422 0.063838 0.05699 0 0.043502 0.0389 0 0.84895 0.2286 0.059369 0.0084085 4.1074 0.052883 6.3092e-05 0.83718 0.0051063 0.0058442 0.0016519 0.98338 0.98626 3.6015e-06 1.4406e-05 0.13047 0.71672 0.77051 0.0015319 0.77762 0.49845 0.0020585 0.42209 1.2787 1.2746 16.0049 144.9823 0.00039873 -84.5989 0.14621
0.25023 0.98801 5.5241e-05 3.8182 0.012047 3.2985e-06 0.001154 0.063327 0.00065424 0.063976 0.057117 0 0.04349 0.0389 0 0.84898 0.22861 0.059373 0.0084091 4.1074 0.052886 6.3096e-05 0.83718 0.0051063 0.0058443 0.0016497 0.98341 0.98647 3.5964e-06 1.4386e-05 0.13047 0.71755 0.7712 0.0015309 0.7789 0.49862 0.0020572 0.4221 1.2806 1.2765 16.005 144.9824 0.00039761 -84.6068 0.14721
0.25123 0.98801 5.5241e-05 3.8182 0.012047 3.3117e-06 0.001154 0.063465 0.00065425 0.064114 0.057243 0 0.043478 0.0389 0 0.84901 0.22863 0.059377 0.0084096 4.1075 0.052888 6.3099e-05 0.83717 0.0051064 0.0058443 0.0016481 0.98344 0.98666 3.5915e-06 1.4366e-05 0.13047 0.71837 0.7719 0.0015298 0.78017 0.49879 0.0020558 0.4221 1.2826 1.2784 16.005 144.9824 0.0003965 -84.6146 0.14821
0.25223 0.98801 5.5241e-05 3.8182 0.012047 3.3249e-06 0.001154 0.063603 0.00065427 0.064252 0.057369 0 0.043466 0.0389 0 0.84904 0.22864 0.059382 0.0084102 4.1075 0.052891 6.3103e-05 0.83717 0.0051064 0.0058443 0.001645 0.98347 0.98684 3.5866e-06 1.4347e-05 0.13047 0.71919 0.77259 0.0015288 0.78144 0.49895 0.0020544 0.42211 1.2845 1.2803 16.0051 144.9824 0.0003954 -84.6224 0.14921
0.25323 0.98801 5.5241e-05 3.8182 0.012047 3.338e-06 0.001154 0.06374 0.00065428 0.06439 0.057495 0 0.043454 0.0389 0 0.84906 0.22865 0.059386 0.0084108 4.1075 0.052894 6.3106e-05 0.83717 0.0051064 0.0058444 0.001643 0.9835 0.98701 3.5817e-06 1.4327e-05 0.13047 0.72001 0.77328 0.0015278 0.7827 0.49912 0.0020531 0.42211 1.2864 1.2823 16.0051 144.9824 0.0003943 -84.63 0.15021
0.25423 0.98801 5.524e-05 3.8182 0.012047 3.3512e-06 0.001154 0.063878 0.0006543 0.064528 0.05762 0 0.043442 0.0389 0 0.84909 0.22866 0.059391 0.0084113 4.1076 0.052896 6.311e-05 0.83717 0.0051065 0.0058444 0.0016416 0.98353 0.98718 3.5769e-06 1.4308e-05 0.13047 0.72083 0.77396 0.0015267 0.78396 0.49929 0.0020518 0.42211 1.2882 1.2842 16.0052 144.9824 0.0003932 -84.6377 0.15121
0.25523 0.98802 5.524e-05 3.8182 0.012047 3.3644e-06 0.001154 0.064016 0.00065432 0.064666 0.057746 0 0.04343 0.0389 0 0.84912 0.22867 0.059395 0.0084119 4.1076 0.052899 6.3113e-05 0.83716 0.0051065 0.0058444 0.0016388 0.98356 0.98733 3.5721e-06 1.4289e-05 0.13047 0.72165 0.77464 0.0015257 0.7852 0.49946 0.0020504 0.42212 1.2901 1.2861 16.0052 144.9824 0.00039212 -84.6452 0.15221
0.25623 0.98802 5.524e-05 3.8182 0.012047 3.3776e-06 0.001154 0.064153 0.00065433 0.064803 0.057872 0 0.043418 0.0389 0 0.84915 0.22869 0.0594 0.0084124 4.1076 0.052902 6.3116e-05 0.83716 0.0051065 0.0058445 0.0016367 0.98359 0.98748 3.5673e-06 1.427e-05 0.13047 0.72246 0.77532 0.0015247 0.78645 0.49963 0.0020491 0.42212 1.292 1.288 16.0053 144.9824 0.00039103 -84.6527 0.15321
0.25723 0.98802 5.524e-05 3.8182 0.012047 3.3907e-06 0.001154 0.064291 0.00065435 0.064941 0.057997 0 0.043406 0.0389 0 0.84918 0.2287 0.059404 0.008413 4.1076 0.052905 6.312e-05 0.83716 0.0051066 0.0058445 0.0016353 0.98361 0.98762 3.5626e-06 1.4251e-05 0.13047 0.72327 0.77599 0.0015237 0.78768 0.4998 0.0020478 0.42213 1.2939 1.2899 16.0053 144.9824 0.00038996 -84.6602 0.15421
0.25823 0.98802 5.524e-05 3.8182 0.012047 3.4039e-06 0.001154 0.064428 0.00065436 0.065078 0.058123 0 0.043394 0.0389 0 0.84921 0.22871 0.059409 0.0084136 4.1077 0.052907 6.3123e-05 0.83716 0.0051066 0.0058445 0.0016328 0.98364 0.98775 3.558e-06 1.4232e-05 0.13047 0.72407 0.77666 0.0015227 0.78891 0.49997 0.0020465 0.42213 1.2958 1.2918 16.0054 144.9825 0.00038889 -84.6676 0.15521
0.25923 0.98802 5.524e-05 3.8182 0.012047 3.4171e-06 0.001154 0.064565 0.00065438 0.065215 0.058248 0 0.043383 0.0389 0 0.84923 0.22872 0.059413 0.0084142 4.1077 0.05291 6.3127e-05 0.83715 0.0051067 0.0058446 0.0016309 0.98367 0.98787 3.5534e-06 1.4214e-05 0.13047 0.72488 0.77732 0.0015218 0.79013 0.50013 0.0020453 0.42214 1.2977 1.2936 16.0054 144.9825 0.00038782 -84.6749 0.15621
0.26023 0.98802 5.524e-05 3.8182 0.012047 3.4303e-06 0.001154 0.064702 0.00065439 0.065352 0.058373 0 0.043371 0.0389 0 0.84926 0.22874 0.059418 0.0084147 4.1077 0.052913 6.3131e-05 0.83715 0.0051067 0.0058446 0.0016288 0.9837 0.98799 3.5488e-06 1.4196e-05 0.13047 0.72568 0.77798 0.0015208 0.79135 0.5003 0.002044 0.42214 1.2995 1.2955 16.0055 144.9825 0.00038676 -84.6822 0.15721
0.26123 0.98802 5.524e-05 3.8182 0.012047 3.4435e-06 0.001154 0.064839 0.00065441 0.065489 0.058498 0 0.043359 0.0389 0 0.84929 0.22875 0.059422 0.0084153 4.1077 0.052916 6.3134e-05 0.83715 0.0051067 0.0058446 0.0016281 0.98372 0.9881 3.5443e-06 1.4178e-05 0.13047 0.72648 0.77864 0.0015198 0.79256 0.50047 0.0020427 0.42215 1.3014 1.2974 16.0055 144.9825 0.00038571 -84.6894 0.15821
0.26223 0.98802 5.524e-05 3.8182 0.012047 3.4566e-06 0.001154 0.064976 0.00065442 0.065626 0.058623 0 0.043347 0.0389 0 0.84932 0.22876 0.059427 0.0084159 4.1078 0.052918 6.3138e-05 0.83714 0.0051068 0.0058447 0.0016261 0.98375 0.98821 3.5398e-06 1.416e-05 0.13047 0.72728 0.77929 0.0015189 0.79376 0.50064 0.0020415 0.42215 1.3032 1.2993 16.0056 144.9825 0.00038466 -84.6966 0.15921
0.26323 0.98802 5.524e-05 3.8182 0.012047 3.4698e-06 0.001154 0.065113 0.00065444 0.065763 0.058748 0 0.043335 0.0389 0 0.84935 0.22878 0.059431 0.0084165 4.1078 0.052921 6.3141e-05 0.83714 0.0051068 0.0058447 0.0016232 0.98378 0.98831 3.5353e-06 1.4142e-05 0.13047 0.72807 0.77994 0.0015179 0.79496 0.50081 0.0020403 0.42216 1.3051 1.3011 16.0056 144.9825 0.00038361 -84.7037 0.16021
0.26423 0.98802 5.524e-05 3.8182 0.012047 3.483e-06 0.001154 0.06525 0.00065445 0.065899 0.058873 0 0.043324 0.0389 0 0.84938 0.22879 0.059436 0.008417 4.1078 0.052924 6.3145e-05 0.83714 0.0051069 0.0058448 0.0016211 0.9838 0.9884 3.5309e-06 1.4124e-05 0.13047 0.72887 0.78059 0.001517 0.79615 0.50098 0.002039 0.42216 1.307 1.303 16.0057 144.9825 0.00038257 -84.7107 0.16121
0.26523 0.98802 5.524e-05 3.8182 0.012046 3.4962e-06 0.001154 0.065386 0.00065447 0.066036 0.058998 0 0.043312 0.0389 0 0.84941 0.2288 0.059441 0.0084176 4.1079 0.052927 6.3148e-05 0.83714 0.0051069 0.0058448 0.0016198 0.98383 0.98849 3.5265e-06 1.4107e-05 0.13047 0.72966 0.78123 0.0015161 0.79734 0.50114 0.0020378 0.42217 1.3088 1.3049 16.0057 144.9825 0.00038154 -84.7177 0.16221
0.26623 0.98802 5.524e-05 3.8182 0.012046 3.5093e-06 0.001154 0.065523 0.00065448 0.066172 0.059123 0 0.0433 0.0389 0 0.84944 0.22881 0.059445 0.0084182 4.1079 0.05293 6.3152e-05 0.83713 0.0051069 0.0058448 0.0016174 0.98386 0.98858 3.5222e-06 1.4089e-05 0.13047 0.73044 0.78187 0.0015152 0.79852 0.50131 0.0020366 0.42217 1.3106 1.3067 16.0058 144.9826 0.00038051 -84.7247 0.16321
0.26723 0.98802 5.524e-05 3.8182 0.012046 3.5225e-06 0.001154 0.065659 0.0006545 0.066309 0.059247 0 0.043288 0.0389 0 0.84947 0.22883 0.05945 0.0084188 4.1079 0.052933 6.3156e-05 0.83713 0.005107 0.0058449 0.0016156 0.98388 0.98866 3.5179e-06 1.4072e-05 0.13047 0.73123 0.78251 0.0015142 0.79969 0.50148 0.0020354 0.42218 1.3125 1.3086 16.0058 144.9826 0.00037949 -84.7315 0.16421
0.26823 0.98802 5.524e-05 3.8182 0.012046 3.5357e-06 0.001154 0.065795 0.00065451 0.066445 0.059372 0 0.043277 0.0389 0 0.8495 0.22884 0.059455 0.0084194 4.108 0.052936 6.3159e-05 0.83713 0.005107 0.0058449 0.0016142 0.98391 0.98874 3.5137e-06 1.4055e-05 0.13047 0.73201 0.78314 0.0015133 0.80086 0.50165 0.0020342 0.42218 1.3143 1.3104 16.0059 144.9826 0.00037847 -84.7384 0.16521
0.26923 0.98802 5.524e-05 3.8182 0.012046 3.5489e-06 0.001154 0.065931 0.00065452 0.066581 0.059496 0 0.043265 0.0389 0 0.84952 0.22885 0.059459 0.00842 4.108 0.052939 6.3163e-05 0.83712 0.005107 0.005845 0.0016121 0.98393 0.98881 3.5095e-06 1.4038e-05 0.13047 0.73279 0.78377 0.0015124 0.80202 0.50182 0.0020331 0.42219 1.3162 1.3123 16.0059 144.9826 0.00037746 -84.7452 0.16621
0.27023 0.98802 5.5239e-05 3.8182 0.012046 3.562e-06 0.001154 0.066067 0.00065454 0.066717 0.05962 0 0.043253 0.0389 0 0.84955 0.22887 0.059464 0.0084206 4.108 0.052941 6.3167e-05 0.83712 0.0051071 0.005845 0.0016103 0.98396 0.98888 3.5053e-06 1.4022e-05 0.13047 0.73357 0.7844 0.0015116 0.80317 0.50199 0.0020319 0.42219 1.318 1.3141 16.006 144.9826 0.00037645 -84.7519 0.16721
0.27123 0.98802 5.5239e-05 3.8182 0.012046 3.5752e-06 0.001154 0.066203 0.00065455 0.066853 0.059745 0 0.043241 0.0389 0 0.84958 0.22888 0.059469 0.0084212 4.108 0.052944 6.3171e-05 0.83712 0.0051071 0.005845 0.0016085 0.98398 0.98895 3.5011e-06 1.4005e-05 0.13047 0.73435 0.78502 0.0015107 0.80432 0.50215 0.0020308 0.4222 1.3198 1.316 16.006 144.9826 0.00037545 -84.7586 0.16821
0.27223 0.98802 5.5239e-05 3.8182 0.012046 3.5884e-06 0.001154 0.066339 0.00065457 0.066989 0.059869 0 0.04323 0.0389 0 0.84961 0.22889 0.059473 0.0084217 4.1081 0.052947 6.3174e-05 0.83712 0.0051072 0.0058451 0.0016074 0.98401 0.98901 3.497e-06 1.3989e-05 0.13047 0.73512 0.78564 0.0015098 0.80547 0.50232 0.0020296 0.4222 1.3216 1.3178 16.0061 144.9826 0.00037445 -84.7652 0.16921
0.27323 0.98802 5.5239e-05 3.8182 0.012046 3.6016e-06 0.001154 0.066475 0.00065458 0.067125 0.059993 0 0.043218 0.0389 0 0.84964 0.2289 0.059478 0.0084223 4.1081 0.05295 6.3178e-05 0.83711 0.0051072 0.0058451 0.0016044 0.98403 0.98907 3.493e-06 1.3972e-05 0.13047 0.73589 0.78626 0.0015089 0.8066 0.50249 0.0020285 0.42221 1.3234 1.3196 16.0061 144.9827 0.00037345 -84.7718 0.17021
0.27423 0.98802 5.5239e-05 3.8182 0.012046 3.6147e-06 0.001154 0.06661 0.0006546 0.06726 0.060117 0 0.043206 0.0389 0 0.84967 0.22892 0.059483 0.0084229 4.1081 0.052953 6.3182e-05 0.83711 0.0051073 0.0058451 0.0016026 0.98405 0.98913 3.4889e-06 1.3956e-05 0.13047 0.73666 0.78687 0.0015081 0.80773 0.50266 0.0020273 0.42221 1.3252 1.3214 16.0062 144.9827 0.00037247 -84.7783 0.17121
0.27523 0.98802 5.5239e-05 3.8182 0.012046 3.6279e-06 0.001154 0.066746 0.00065461 0.067396 0.06024 0 0.043195 0.0389 0 0.8497 0.22893 0.059488 0.0084235 4.1082 0.052956 6.3186e-05 0.83711 0.0051073 0.0058452 0.0016019 0.98408 0.98919 3.4849e-06 1.394e-05 0.13047 0.73742 0.78748 0.0015072 0.80886 0.50283 0.0020262 0.42222 1.327 1.3233 16.0062 144.9827 0.00037148 -84.7848 0.17221
0.27623 0.98802 5.5239e-05 3.8182 0.012046 3.6411e-06 0.001154 0.066881 0.00065462 0.067531 0.060364 0 0.043183 0.0389 0 0.84973 0.22894 0.059492 0.0084241 4.1082 0.052959 6.3189e-05 0.8371 0.0051073 0.0058452 0.0016006 0.9841 0.98924 3.481e-06 1.3924e-05 0.13047 0.73819 0.78808 0.0015064 0.80998 0.503 0.0020251 0.42223 1.3288 1.3251 16.0063 144.9827 0.00037051 -84.7912 0.17321
0.27723 0.98802 5.5239e-05 3.8182 0.012046 3.6543e-06 0.001154 0.067016 0.00065464 0.067666 0.060488 0 0.043172 0.0389 0 0.84976 0.22896 0.059497 0.0084248 4.1082 0.052962 6.3193e-05 0.8371 0.0051074 0.0058453 0.0015983 0.98412 0.98929 3.4771e-06 1.3909e-05 0.13048 0.73895 0.78869 0.0015055 0.81109 0.50316 0.002024 0.42223 1.3306 1.3269 16.0063 144.9827 0.00036953 -84.7976 0.17421
0.27823 0.98802 5.5239e-05 3.8182 0.012046 3.6674e-06 0.001154 0.067151 0.00065465 0.067801 0.060611 0 0.04316 0.0389 0 0.84979 0.22897 0.059502 0.0084254 4.1083 0.052965 6.3197e-05 0.8371 0.0051074 0.0058453 0.0015963 0.98415 0.98934 3.4732e-06 1.3893e-05 0.13048 0.73971 0.78929 0.0015047 0.8122 0.50333 0.0020229 0.42224 1.3324 1.3287 16.0064 144.9827 0.00036857 -84.8039 0.17521
0.27923 0.98802 5.5239e-05 3.8182 0.012046 3.6806e-06 0.001154 0.067286 0.00065466 0.067936 0.060735 0 0.043148 0.0389 0 0.84982 0.22898 0.059507 0.008426 4.1083 0.052968 6.3201e-05 0.83709 0.0051075 0.0058454 0.0015953 0.98417 0.98938 3.4693e-06 1.3878e-05 0.13048 0.74047 0.78988 0.0015039 0.8133 0.5035 0.0020219 0.42224 1.3342 1.3305 16.0064 144.9827 0.0003676 -84.8102 0.17621
0.28023 0.98802 5.5239e-05 3.8182 0.012046 3.6938e-06 0.001154 0.067421 0.00065468 0.068071 0.060858 0 0.043137 0.0389 0 0.84985 0.229 0.059512 0.0084266 4.1083 0.052971 6.3205e-05 0.83709 0.0051075 0.0058454 0.0015939 0.98419 0.98943 3.4655e-06 1.3862e-05 0.13048 0.74122 0.79048 0.001503 0.8144 0.50367 0.0020208 0.42225 1.336 1.3323 16.0065 144.9828 0.00036664 -84.8164 0.17721
0.28123 0.98802 5.5239e-05 3.8182 0.012046 3.707e-06 0.001154 0.067556 0.00065469 0.068206 0.060981 0 0.043125 0.0389 0 0.84989 0.22901 0.059516 0.0084272 4.1084 0.052974 6.3208e-05 0.83709 0.0051076 0.0058454 0.0015916 0.98421 0.98947 3.4617e-06 1.3847e-05 0.13048 0.74197 0.79107 0.0015022 0.81549 0.50384 0.0020197 0.42226 1.3378 1.3341 16.0065 144.9828 0.00036569 -84.8226 0.17821
0.28223 0.98802 5.5239e-05 3.8182 0.012046 3.7201e-06 0.001154 0.067691 0.00065471 0.068341 0.061105 0 0.043114 0.0389 0 0.84992 0.22902 0.059521 0.0084278 4.1084 0.052977 6.3212e-05 0.83709 0.0051076 0.0058455 0.0015897 0.98424 0.98951 3.4579e-06 1.3832e-05 0.13048 0.74272 0.79165 0.0015014 0.81657 0.504 0.0020187 0.42226 1.3396 1.3359 16.0065 144.9828 0.00036474 -84.8287 0.17921
0.28323 0.98802 5.5239e-05 3.8182 0.012046 3.7333e-06 0.001154 0.067825 0.00065472 0.068475 0.061228 0 0.043102 0.0389 0 0.84995 0.22904 0.059526 0.0084284 4.1084 0.05298 6.3216e-05 0.83708 0.0051076 0.0058455 0.0015887 0.98426 0.98955 3.4542e-06 1.3817e-05 0.13048 0.74347 0.79224 0.0015006 0.81765 0.50417 0.0020176 0.42227 1.3413 1.3376 16.0066 144.9828 0.0003638 -84.8348 0.18021
0.28423 0.98802 5.5239e-05 3.8182 0.012046 3.7465e-06 0.001154 0.06796 0.00065473 0.06861 0.061351 0 0.043091 0.0389 0 0.84998 0.22905 0.059531 0.008429 4.1085 0.052984 6.322e-05 0.83708 0.0051077 0.0058456 0.0015874 0.98428 0.98959 3.4505e-06 1.3802e-05 0.13048 0.74421 0.79282 0.0014998 0.81872 0.50434 0.0020166 0.42228 1.3431 1.3394 16.0066 144.9828 0.00036286 -84.8409 0.18121
0.28523 0.98802 5.5239e-05 3.8182 0.012046 3.7597e-06 0.001154 0.068094 0.00065475 0.068744 0.061474 0 0.043079 0.0389 0 0.85001 0.22907 0.059536 0.0084296 4.1085 0.052987 6.3224e-05 0.83708 0.0051077 0.0058456 0.0015852 0.9843 0.98962 3.4469e-06 1.3788e-05 0.13048 0.74496 0.7934 0.001499 0.81979 0.50451 0.0020156 0.42228 1.3449 1.3412 16.0067 144.9828 0.00036192 -84.8469 0.18221
0.28623 0.98802 5.5239e-05 3.8182 0.012046 3.7728e-06 0.001154 0.068228 0.00065476 0.068879 0.061596 0 0.043068 0.0389 0 0.85004 0.22908 0.059541 0.0084303 4.1085 0.05299 6.3228e-05 0.83707 0.0051078 0.0058457 0.0015845 0.98432 0.98966 3.4432e-06 1.3773e-05 0.13048 0.7457 0.79397 0.0014983 0.82085 0.50468 0.0020145 0.42229 1.3466 1.343 16.0067 144.9828 0.00036099 -84.8528 0.18321
0.28723 0.98802 5.5238e-05 3.8182 0.012046 3.786e-06 0.001154 0.068363 0.00065477 0.069013 0.061719 0 0.043056 0.0389 0 0.85007 0.22909 0.059546 0.0084309 4.1086 0.052993 6.3232e-05 0.83707 0.0051078 0.0058457 0.0015819 0.98435 0.98969 3.4396e-06 1.3759e-05 0.13048 0.74644 0.79454 0.0014975 0.8219 0.50484 0.0020135 0.4223 1.3484 1.3447 16.0068 144.9828 0.00036007 -84.8587 0.18421
0.28823 0.98802 5.5238e-05 3.8182 0.012046 3.7992e-06 0.001154 0.068497 0.00065478 0.069147 0.061842 0 0.043045 0.0389 0 0.8501 0.22911 0.059551 0.0084315 4.1086 0.052996 6.3236e-05 0.83707 0.0051079 0.0058457 0.0015811 0.98437 0.98972 3.4361e-06 1.3745e-05 0.13048 0.74717 0.79511 0.0014967 0.82295 0.50501 0.0020125 0.4223 1.3501 1.3465 16.0068 144.9829 0.00035915 -84.8646 0.18521
0.28923 0.98802 5.5238e-05 3.8182 0.012046 3.8124e-06 0.001154 0.068631 0.0006548 0.069281 0.061964 0 0.043034 0.0389 0 0.85013 0.22912 0.059556 0.0084321 4.1086 0.052999 6.324e-05 0.83706 0.0051079 0.0058458 0.0015788 0.98439 0.98975 3.4325e-06 1.373e-05 0.13048 0.74791 0.79568 0.001496 0.824 0.50518 0.0020115 0.42231 1.3519 1.3483 16.0068 144.9829 0.00035823 -84.8704 0.18621
0.29023 0.98802 5.5238e-05 3.8182 0.012046 3.8255e-06 0.001154 0.068764 0.00065481 0.069415 0.062087 0 0.043022 0.0389 0 0.85016 0.22913 0.059561 0.0084328 4.1087 0.053002 6.3244e-05 0.83706 0.005108 0.0058458 0.001578 0.98441 0.98978 3.429e-06 1.3716e-05 0.13048 0.74864 0.79624 0.0014952 0.82504 0.50535 0.0020105 0.42232 1.3536 1.35 16.0069 144.9829 0.00035732 -84.8762 0.18721
0.29123 0.98802 5.5238e-05 3.8182 0.012046 3.8387e-06 0.001154 0.068898 0.00065482 0.069548 0.062209 0 0.043011 0.0389 0 0.8502 0.22915 0.059566 0.0084334 4.1087 0.053005 6.3248e-05 0.83706 0.005108 0.0058459 0.0015768 0.98443 0.98981 3.4256e-06 1.3703e-05 0.13048 0.74937 0.7968 0.0014945 0.82607 0.50552 0.0020096 0.42232 1.3553 1.3518 16.0069 144.9829 0.00035641 -84.8819 0.18821
0.29223 0.98802 5.5238e-05 3.8182 0.012046 3.8519e-06 0.001154 0.069032 0.00065484 0.069682 0.062331 0 0.042999 0.0389 0 0.85023 0.22916 0.059571 0.008434 4.1087 0.053009 6.3252e-05 0.83705 0.005108 0.0058459 0.0015744 0.98445 0.98984 3.4221e-06 1.3689e-05 0.13048 0.75009 0.79736 0.0014937 0.8271 0.50568 0.0020086 0.42233 1.3571 1.3535 16.007 144.9829 0.00035551 -84.8876 0.18921
0.29323 0.98802 5.5238e-05 3.8182 0.012046 3.8651e-06 0.001154 0.069165 0.00065485 0.069816 0.062453 0 0.042988 0.0389 0 0.85026 0.22918 0.059576 0.0084347 4.1088 0.053012 6.3256e-05 0.83705 0.0051081 0.005846 0.0015725 0.98447 0.98986 3.4187e-06 1.3675e-05 0.13048 0.75082 0.79791 0.001493 0.82812 0.50585 0.0020076 0.42234 1.3588 1.3553 16.007 144.9829 0.00035461 -84.8932 0.19021
0.29423 0.98802 5.5238e-05 3.8182 0.012046 3.8782e-06 0.001154 0.069299 0.00065486 0.069949 0.062575 0 0.042977 0.0389 0 0.85029 0.22919 0.059581 0.0084353 4.1088 0.053015 6.326e-05 0.83705 0.0051081 0.005846 0.0015719 0.98449 0.98989 3.4153e-06 1.3662e-05 0.13048 0.75154 0.79846 0.0014922 0.82913 0.50602 0.0020067 0.42234 1.3605 1.357 16.007 144.983 0.00035372 -84.8988 0.19121
0.29523 0.98802 5.5238e-05 3.8182 0.012046 3.8914e-06 0.001154 0.069432 0.00065487 0.070082 0.062697 0 0.042965 0.0389 0 0.85032 0.2292 0.059586 0.0084359 4.1089 0.053018 6.3264e-05 0.83704 0.0051082 0.0058461 0.0015709 0.98451 0.98991 3.412e-06 1.3648e-05 0.13048 0.75226 0.79901 0.0014915 0.83014 0.50619 0.0020057 0.42235 1.3623 1.3587 16.0071 144.983 0.00035283 -84.9044 0.19221
0.29623 0.98802 5.5238e-05 3.8182 0.012046 3.9046e-06 0.001154 0.069565 0.00065489 0.070215 0.062819 0 0.042954 0.0389 0 0.85035 0.22922 0.059591 0.0084366 4.1089 0.053021 6.3268e-05 0.83704 0.0051082 0.0058461 0.0015686 0.98453 0.98994 3.4086e-06 1.3635e-05 0.13048 0.75298 0.79956 0.0014908 0.83115 0.50635 0.0020048 0.42236 1.364 1.3605 16.0071 144.983 0.00035194 -84.9099 0.19321
0.29723 0.98802 5.5238e-05 3.8182 0.012046 3.9178e-06 0.001154 0.069698 0.0006549 0.070349 0.062941 0 0.042943 0.0389 0 0.85039 0.22923 0.059596 0.0084372 4.1089 0.053025 6.3272e-05 0.83704 0.0051083 0.0058462 0.0015668 0.98455 0.98996 3.4053e-06 1.3622e-05 0.13048 0.7537 0.8001 0.0014901 0.83215 0.50652 0.0020038 0.42237 1.3657 1.3622 16.0072 144.983 0.00035106 -84.9153 0.19421
0.29823 0.98802 5.5238e-05 3.8182 0.012046 3.9309e-06 0.001154 0.069831 0.00065491 0.070482 0.063063 0 0.042932 0.0389 0 0.85042 0.22925 0.059601 0.0084378 4.109 0.053028 6.3277e-05 0.83704 0.0051083 0.0058462 0.0015662 0.98457 0.98998 3.4021e-06 1.3609e-05 0.13048 0.75441 0.80064 0.0014894 0.83314 0.50669 0.0020029 0.42237 1.3674 1.3639 16.0072 144.983 0.00035019 -84.9208 0.19521
0.29923 0.98802 5.5238e-05 3.8182 0.012046 3.9441e-06 0.001154 0.069964 0.00065492 0.070614 0.063184 0 0.04292 0.0389 0 0.85045 0.22926 0.059606 0.0084385 4.109 0.053031 6.3281e-05 0.83703 0.0051084 0.0058462 0.0015652 0.98459 0.99 3.3988e-06 1.3596e-05 0.13048 0.75512 0.80118 0.0014887 0.83413 0.50686 0.002002 0.42238 1.3691 1.3656 16.0072 144.983 0.00034931 -84.9262 0.19621
0.30023 0.98802 5.5238e-05 3.8182 0.012046 3.9573e-06 0.001154 0.070097 0.00065494 0.070747 0.063306 0 0.042909 0.0389 0 0.85048 0.22927 0.059611 0.0084391 4.109 0.053035 6.3285e-05 0.83703 0.0051084 0.0058463 0.0015629 0.9846 0.99003 3.3956e-06 1.3583e-05 0.13048 0.75583 0.80171 0.001488 0.83511 0.50702 0.0020011 0.42239 1.3708 1.3673 16.0073 144.983 0.00034845 -84.9315 0.19721
0.30123 0.98802 5.5238e-05 3.8182 0.012046 3.9705e-06 0.001154 0.07023 0.00065495 0.07088 0.063427 0 0.042898 0.0389 0 0.85051 0.22929 0.059616 0.0084398 4.1091 0.053038 6.3289e-05 0.83703 0.0051085 0.0058463 0.0015612 0.98462 0.99005 3.3924e-06 1.357e-05 0.13048 0.75654 0.80225 0.0014873 0.83609 0.50719 0.0020002 0.42239 1.3725 1.369 16.0073 144.9831 0.00034758 -84.9368 0.19821
0.30223 0.98802 5.5238e-05 3.8182 0.012046 3.9836e-06 0.001154 0.070362 0.00065496 0.071012 0.063549 0 0.042887 0.0389 0 0.85055 0.2293 0.059621 0.0084404 4.1091 0.053041 6.3293e-05 0.83702 0.0051085 0.0058464 0.0015607 0.98464 0.99007 3.3893e-06 1.3557e-05 0.13048 0.75724 0.80278 0.0014866 0.83706 0.50736 0.0019993 0.4224 1.3742 1.3707 16.0074 144.9831 0.00034672 -84.9421 0.19921
0.30323 0.98802 5.5237e-05 3.8182 0.012046 3.9968e-06 0.001154 0.070495 0.00065497 0.071145 0.06367 0 0.042875 0.0389 0 0.85058 0.22932 0.059627 0.0084411 4.1092 0.053044 6.3297e-05 0.83702 0.0051086 0.0058464 0.0015597 0.98466 0.99008 3.3861e-06 1.3545e-05 0.13049 0.75795 0.8033 0.0014859 0.83803 0.50753 0.0019984 0.42241 1.3759 1.3724 16.0074 144.9831 0.00034587 -84.9473 0.20021
0.30423 0.98802 5.5237e-05 3.8182 0.012046 4.01e-06 0.001154 0.070627 0.00065498 0.071277 0.063791 0 0.042864 0.0389 0 0.85061 0.22933 0.059632 0.0084417 4.1092 0.053048 6.3302e-05 0.83702 0.0051086 0.0058465 0.0015575 0.98468 0.9901 3.383e-06 1.3532e-05 0.13049 0.75865 0.80383 0.0014853 0.83899 0.50769 0.0019975 0.42242 1.3776 1.3741 16.0074 144.9831 0.00034502 -84.9525 0.20121
0.30523 0.98802 5.5237e-05 3.8182 0.012046 4.0231e-06 0.001154 0.070759 0.000655 0.071409 0.063912 0 0.042853 0.0389 0 0.85064 0.22935 0.059637 0.0084424 4.1092 0.053051 6.3306e-05 0.83701 0.0051087 0.0058465 0.0015558 0.9847 0.99012 3.3799e-06 1.352e-05 0.13049 0.75935 0.80435 0.0014846 0.83995 0.50786 0.0019966 0.42242 1.3792 1.3758 16.0075 144.9831 0.00034417 -84.9576 0.20221
0.30623 0.98802 5.5237e-05 3.8182 0.012046 4.0363e-06 0.001154 0.070891 0.00065501 0.071542 0.064033 0 0.042842 0.0389 0 0.85068 0.22936 0.059642 0.008443 4.1093 0.053054 6.331e-05 0.83701 0.0051087 0.0058466 0.0015553 0.98471 0.99014 3.3769e-06 1.3508e-05 0.13049 0.76004 0.80487 0.0014839 0.8409 0.50803 0.0019958 0.42243 1.3809 1.3775 16.0075 144.9831 0.00034333 -84.9627 0.20321
0.30723 0.98802 5.5237e-05 3.8182 0.012046 4.0495e-06 0.001154 0.071023 0.00065502 0.071674 0.064154 0 0.042831 0.0389 0 0.85071 0.22937 0.059647 0.0084437 4.1093 0.053058 6.3314e-05 0.83701 0.0051088 0.0058466 0.0015544 0.98473 0.99016 3.3739e-06 1.3496e-05 0.13049 0.76074 0.80538 0.0014833 0.84185 0.5082 0.0019949 0.42244 1.3826 1.3792 16.0075 144.9831 0.00034249 -84.9678 0.20421
0.30823 0.98802 5.5237e-05 3.8182 0.012046 4.0627e-06 0.001154 0.071155 0.00065503 0.071806 0.064275 0 0.042819 0.0389 0 0.85074 0.22939 0.059652 0.0084443 4.1093 0.053061 6.3319e-05 0.837 0.0051088 0.0058467 0.0015522 0.98475 0.99017 3.3709e-06 1.3484e-05 0.13049 0.76143 0.8059 0.0014826 0.84279 0.50836 0.0019941 0.42245 1.3842 1.3809 16.0076 144.9832 0.00034165 -84.9728 0.20521
0.30923 0.98802 5.5237e-05 3.8182 0.012046 4.0758e-06 0.001154 0.071287 0.00065504 0.071937 0.064395 0 0.042808 0.0389 0 0.85078 0.2294 0.059658 0.008445 4.1094 0.053065 6.3323e-05 0.837 0.0051089 0.0058467 0.0015505 0.98477 0.99019 3.3679e-06 1.3472e-05 0.13049 0.76212 0.80641 0.001482 0.84372 0.50853 0.0019932 0.42246 1.3859 1.3826 16.0076 144.9832 0.00034082 -84.9778 0.20621
0.31023 0.98802 5.5237e-05 3.8182 0.012046 4.089e-06 0.001154 0.071419 0.00065506 0.072069 0.064516 0 0.042797 0.0389 0 0.85081 0.22942 0.059663 0.0084457 4.1094 0.053068 6.3327e-05 0.837 0.0051089 0.0058468 0.0015502 0.98478 0.99021 3.3649e-06 1.346e-05 0.13049 0.76281 0.80692 0.0014813 0.84465 0.5087 0.0019924 0.42246 1.3876 1.3842 16.0076 144.9832 0.00034 -84.9828 0.20721
0.31123 0.98802 5.5237e-05 3.8182 0.012046 4.1022e-06 0.001154 0.07155 0.00065507 0.072201 0.064636 0 0.042786 0.0389 0 0.85084 0.22943 0.059668 0.0084463 4.1095 0.053071 6.3332e-05 0.83699 0.005109 0.0058468 0.0015482 0.9848 0.99022 3.362e-06 1.3448e-05 0.13049 0.76349 0.80743 0.0014807 0.84558 0.50887 0.0019915 0.42247 1.3892 1.3859 16.0077 144.9832 0.00033917 -84.9877 0.20821
0.31223 0.98802 5.5237e-05 3.8182 0.012046 4.1154e-06 0.001154 0.071682 0.00065508 0.072332 0.064757 0 0.042775 0.0389 0 0.85088 0.22945 0.059674 0.008447 4.1095 0.053075 6.3336e-05 0.83699 0.005109 0.0058469 0.0015477 0.98482 0.99024 3.3591e-06 1.3437e-05 0.13049 0.76418 0.80793 0.00148 0.8465 0.50903 0.0019907 0.42248 1.3909 1.3876 16.0077 144.9832 0.00033836 -84.9926 0.20921
0.31323 0.98802 5.5237e-05 3.8182 0.012046 4.1285e-06 0.001154 0.071813 0.00065509 0.072464 0.064877 0 0.042764 0.0389 0 0.85091 0.22946 0.059679 0.0084477 4.1095 0.053078 6.334e-05 0.83699 0.0051091 0.0058469 0.0015468 0.98484 0.99025 3.3562e-06 1.3425e-05 0.13049 0.76486 0.80843 0.0014794 0.84741 0.5092 0.0019899 0.42249 1.3925 1.3892 16.0078 144.9832 0.00033754 -84.9974 0.21021
0.31423 0.98802 5.5237e-05 3.8182 0.012046 4.1417e-06 0.001154 0.071944 0.0006551 0.072595 0.064997 0 0.042753 0.0389 0 0.85094 0.22948 0.059684 0.0084483 4.1096 0.053082 6.3345e-05 0.83698 0.0051091 0.005847 0.0015446 0.98485 0.99027 3.3534e-06 1.3414e-05 0.13049 0.76554 0.80893 0.0014788 0.84832 0.50937 0.0019891 0.4225 1.3942 1.3909 16.0078 144.9832 0.00033673 -85.0023 0.21121
0.31523 0.98802 5.5237e-05 3.8182 0.012046 4.1549e-06 0.001154 0.072076 0.00065511 0.072726 0.065117 0 0.042742 0.0389 0 0.85098 0.22949 0.059689 0.008449 4.1096 0.053085 6.3349e-05 0.83698 0.0051092 0.005847 0.001544 0.98487 0.99028 3.3505e-06 1.3402e-05 0.13049 0.76622 0.80943 0.0014782 0.84923 0.50953 0.0019883 0.4225 1.3958 1.3925 16.0078 144.9833 0.00033593 -85.007 0.21221
0.31623 0.98802 5.5237e-05 3.8182 0.012046 4.1681e-06 0.001154 0.072207 0.00065512 0.072857 0.065238 0 0.042731 0.0389 0 0.85101 0.22951 0.059695 0.0084497 4.1097 0.053089 6.3353e-05 0.83697 0.0051092 0.0058471 0.0015421 0.98489 0.9903 3.3477e-06 1.3391e-05 0.13049 0.76689 0.80992 0.0014776 0.85013 0.5097 0.0019875 0.42251 1.3974 1.3942 16.0079 144.9833 0.00033512 -85.0118 0.21321
0.31723 0.98802 5.5237e-05 3.8182 0.012046 4.1812e-06 0.001154 0.072338 0.00065514 0.072988 0.065357 0 0.04272 0.0389 0 0.85104 0.22952 0.0597 0.0084503 4.1097 0.053092 6.3358e-05 0.83697 0.0051093 0.0058471 0.0015405 0.9849 0.99031 3.3449e-06 1.338e-05 0.13049 0.76756 0.81041 0.001477 0.85102 0.50987 0.0019867 0.42252 1.3991 1.3958 16.0079 144.9833 0.00033432 -85.0165 0.21421
0.31823 0.98802 5.5237e-05 3.8182 0.012046 4.1944e-06 0.001154 0.072468 0.00065515 0.073119 0.065477 0 0.042709 0.0389 0 0.85108 0.22954 0.059705 0.008451 4.1097 0.053095 6.3362e-05 0.83697 0.0051093 0.0058472 0.0015403 0.98492 0.99032 3.3422e-06 1.3369e-05 0.13049 0.76824 0.8109 0.0014764 0.85191 0.51004 0.0019859 0.42253 1.4007 1.3974 16.0079 144.9833 0.00033353 -85.0211 0.21521
0.31923 0.98802 5.5236e-05 3.8182 0.012046 4.2076e-06 0.001154 0.072599 0.00065516 0.07325 0.065597 0 0.042698 0.0389 0 0.85111 0.22955 0.059711 0.0084517 4.1098 0.053099 6.3367e-05 0.83696 0.0051094 0.0058472 0.0015385 0.98493 0.99034 3.3394e-06 1.3358e-05 0.13049 0.7689 0.81139 0.0014758 0.8528 0.5102 0.0019851 0.42254 1.4023 1.3991 16.008 144.9833 0.00033274 -85.0258 0.21621
0.32023 0.98802 5.5236e-05 3.8182 0.012046 4.2208e-06 0.001154 0.07273 0.00065517 0.07338 0.065717 0 0.042687 0.0389 0 0.85114 0.22957 0.059716 0.0084524 4.1098 0.053102 6.3371e-05 0.83696 0.0051094 0.0058473 0.001538 0.98495 0.99035 3.3367e-06 1.3347e-05 0.13049 0.76957 0.81187 0.0014752 0.85368 0.51037 0.0019843 0.42255 1.4039 1.4007 16.008 144.9833 0.00033195 -85.0304 0.21721
0.32123 0.98802 5.5236e-05 3.8182 0.012046 4.2339e-06 0.001154 0.07286 0.00065518 0.073511 0.065836 0 0.042676 0.0389 0 0.85118 0.22958 0.059722 0.0084531 4.1099 0.053106 6.3376e-05 0.83696 0.0051095 0.0058473 0.0015361 0.98497 0.99036 3.334e-06 1.3336e-05 0.13049 0.77024 0.81235 0.0014746 0.85455 0.51054 0.0019836 0.42255 1.4055 1.4023 16.008 144.9834 0.00033117 -85.0349 0.21821
0.32223 0.98802 5.5236e-05 3.8182 0.012046 4.2471e-06 0.001154 0.072991 0.00065519 0.073641 0.065956 0 0.042665 0.0389 0 0.85121 0.2296 0.059727 0.0084537 4.1099 0.05311 6.338e-05 0.83695 0.0051096 0.0058474 0.0015357 0.98498 0.99037 3.3314e-06 1.3326e-05 0.13049 0.7709 0.81283 0.001474 0.85542 0.5107 0.0019828 0.42256 1.4071 1.4039 16.008 144.9834 0.00033039 -85.0394 0.21921
0.32323 0.98802 5.5236e-05 3.8182 0.012046 4.2603e-06 0.001154 0.073121 0.0006552 0.073772 0.066075 0 0.042654 0.0389 0 0.85125 0.22961 0.059732 0.0084544 4.11 0.053113 6.3385e-05 0.83695 0.0051096 0.0058475 0.0015338 0.985 0.99039 3.3287e-06 1.3315e-05 0.13049 0.77156 0.81331 0.0014734 0.85629 0.51087 0.001982 0.42257 1.4087 1.4056 16.0081 144.9834 0.00032961 -85.0439 0.22021
0.32423 0.98802 5.5236e-05 3.8182 0.012046 4.2734e-06 0.001154 0.073251 0.00065521 0.073902 0.066195 0 0.042643 0.0389 0 0.85128 0.22963 0.059738 0.0084551 4.11 0.053117 6.3389e-05 0.83695 0.0051097 0.0058475 0.0015334 0.98501 0.9904 3.3261e-06 1.3305e-05 0.13049 0.77222 0.81379 0.0014728 0.85715 0.51104 0.0019813 0.42258 1.4103 1.4072 16.0081 144.9834 0.00032884 -85.0484 0.22121
0.32523 0.98802 5.5236e-05 3.8182 0.012046 4.2866e-06 0.001154 0.073382 0.00065522 0.074032 0.066314 0 0.042632 0.0389 0 0.85132 0.22964 0.059743 0.0084558 4.11 0.05312 6.3394e-05 0.83694 0.0051097 0.0058476 0.0015315 0.98503 0.99041 3.3235e-06 1.3294e-05 0.13049 0.77288 0.81426 0.0014723 0.858 0.5112 0.0019805 0.42259 1.4119 1.4088 16.0081 144.9834 0.00032807 -85.0528 0.22221
0.32623 0.98802 5.5236e-05 3.8182 0.012046 4.2998e-06 0.001154 0.073512 0.00065524 0.074162 0.066433 0 0.042621 0.0389 0 0.85135 0.22966 0.059749 0.0084565 4.1101 0.053124 6.3398e-05 0.83694 0.0051098 0.0058476 0.0015312 0.98504 0.99042 3.3209e-06 1.3284e-05 0.1305 0.77353 0.81473 0.0014717 0.85885 0.51137 0.0019798 0.4226 1.4135 1.4104 16.0082 144.9834 0.00032731 -85.0572 0.22321
0.32723 0.98802 5.5236e-05 3.8182 0.012046 4.313e-06 0.001154 0.073642 0.00065525 0.074292 0.066552 0 0.04261 0.0389 0 0.85138 0.22967 0.059754 0.0084572 4.1101 0.053127 6.3403e-05 0.83694 0.0051098 0.0058477 0.0015293 0.98506 0.99043 3.3183e-06 1.3274e-05 0.1305 0.77418 0.8152 0.0014711 0.8597 0.51154 0.0019791 0.42261 1.4151 1.412 16.0082 144.9835 0.00032655 -85.0616 0.22421
0.32823 0.98802 5.5236e-05 3.8182 0.012046 4.3261e-06 0.001154 0.073771 0.00065526 0.074422 0.066671 0 0.0426 0.0389 0 0.85142 0.22969 0.05976 0.0084579 4.1102 0.053131 6.3407e-05 0.83693 0.0051099 0.0058477 0.001529 0.98507 0.99045 3.3158e-06 1.3263e-05 0.1305 0.77483 0.81566 0.0014706 0.86054 0.5117 0.0019783 0.42262 1.4167 1.4136 16.0082 144.9835 0.00032579 -85.0659 0.22521
0.32923 0.98802 5.5236e-05 3.8182 0.012046 4.3393e-06 0.001154 0.073901 0.00065527 0.074552 0.06679 0 0.042589 0.0389 0 0.85145 0.2297 0.059765 0.0084586 4.1102 0.053135 6.3412e-05 0.83693 0.0051099 0.0058478 0.0015271 0.98509 0.99046 3.3133e-06 1.3253e-05 0.1305 0.77548 0.81613 0.00147 0.86138 0.51187 0.0019776 0.42262 1.4183 1.4152 16.0083 144.9835 0.00032503 -85.0702 0.22621
0.33023 0.98802 5.5236e-05 3.8182 0.012046 4.3525e-06 0.001154 0.074031 0.00065528 0.074681 0.066909 0 0.042578 0.0389 0 0.85149 0.22972 0.059771 0.0084593 4.1103 0.053138 6.3416e-05 0.83693 0.00511 0.0058478 0.0015268 0.9851 0.99047 3.3108e-06 1.3243e-05 0.1305 0.77613 0.81659 0.0014695 0.86221 0.51204 0.0019769 0.42263 1.4199 1.4168 16.0083 144.9835 0.00032428 -85.0745 0.22721
0.33123 0.98802 5.5236e-05 3.8182 0.012046 4.3657e-06 0.001154 0.07416 0.00065529 0.074811 0.067027 0 0.042567 0.0389 0 0.85152 0.22973 0.059776 0.0084599 4.1103 0.053142 6.3421e-05 0.83692 0.0051101 0.0058479 0.0015249 0.98512 0.99048 3.3083e-06 1.3233e-05 0.1305 0.77677 0.81705 0.0014689 0.86304 0.5122 0.0019762 0.42264 1.4214 1.4183 16.0083 144.9835 0.00032354 -85.0787 0.22821
0.33223 0.98802 5.5236e-05 3.8182 0.012046 4.3788e-06 0.001154 0.07429 0.0006553 0.07494 0.067146 0 0.042556 0.0389 0 0.85156 0.22975 0.059782 0.0084606 4.1104 0.053145 6.3426e-05 0.83692 0.0051101 0.005848 0.0015247 0.98513 0.99049 3.3058e-06 1.3224e-05 0.1305 0.77742 0.8175 0.0014684 0.86386 0.51237 0.0019755 0.42265 1.423 1.4199 16.0083 144.9835 0.00032279 -85.0829 0.22921
0.33323 0.98802 5.5236e-05 3.8182 0.012046 4.392e-06 0.001154 0.074419 0.00065531 0.07507 0.067264 0 0.042546 0.0389 0 0.85159 0.22976 0.059787 0.0084613 4.1104 0.053149 6.343e-05 0.83691 0.0051102 0.005848 0.0015227 0.98514 0.9905 3.3034e-06 1.3214e-05 0.1305 0.77806 0.81796 0.0014679 0.86467 0.51254 0.0019748 0.42266 1.4246 1.4215 16.0084 144.9835 0.00032205 -85.0871 0.23021
0.33423 0.98802 5.5236e-05 3.8182 0.012046 4.4052e-06 0.001154 0.074548 0.00065532 0.075199 0.067383 0 0.042535 0.0389 0 0.85163 0.22978 0.059793 0.008462 4.1104 0.053153 6.3435e-05 0.83691 0.0051102 0.0058481 0.0015226 0.98516 0.99051 3.301e-06 1.3204e-05 0.1305 0.7787 0.81841 0.0014673 0.86549 0.5127 0.0019741 0.42267 1.4261 1.4231 16.0084 144.9836 0.00032132 -85.0912 0.23121
0.33523 0.98802 5.5235e-05 3.8182 0.012046 4.4183e-06 0.001154 0.074677 0.00065533 0.075328 0.067501 0 0.042524 0.0389 0 0.85166 0.22979 0.059798 0.0084628 4.1105 0.053157 6.344e-05 0.83691 0.0051103 0.0058481 0.0015206 0.98517 0.99052 3.2986e-06 1.3195e-05 0.1305 0.77933 0.81886 0.0014668 0.8663 0.51287 0.0019734 0.42268 1.4277 1.4246 16.0084 144.9836 0.00032059 -85.0953 0.23221
0.33623 0.98802 5.5235e-05 3.8182 0.012046 4.4315e-06 0.001154 0.074806 0.00065534 0.075457 0.067619 0 0.042513 0.0389 0 0.8517 0.22981 0.059804 0.0084635 4.1105 0.05316 6.3444e-05 0.8369 0.0051104 0.0058482 0.0015206 0.98519 0.99053 3.2962e-06 1.3185e-05 0.1305 0.77997 0.81931 0.0014663 0.8671 0.51304 0.0019727 0.42269 1.4292 1.4262 16.0085 144.9836 0.00031986 -85.0994 0.23321
0.33723 0.98802 5.5235e-05 3.8182 0.012046 4.4447e-06 0.001154 0.074935 0.00065535 0.075586 0.067738 0 0.042502 0.0389 0 0.85173 0.22983 0.05981 0.0084642 4.1106 0.053164 6.3449e-05 0.8369 0.0051104 0.0058482 0.0015185 0.9852 0.99054 3.2938e-06 1.3176e-05 0.1305 0.7806 0.81976 0.0014658 0.8679 0.5132 0.001972 0.4227 1.4308 1.4278 16.0085 144.9836 0.00031913 -85.1034 0.23421
0.33823 0.98802 5.5235e-05 3.8182 0.012046 4.4579e-06 0.001154 0.075064 0.00065536 0.075715 0.067856 0 0.042492 0.0389 0 0.85177 0.22984 0.059815 0.0084649 4.1106 0.053168 6.3454e-05 0.8369 0.0051105 0.0058483 0.0015186 0.98521 0.99055 3.2915e-06 1.3166e-05 0.1305 0.78123 0.8202 0.0014652 0.86869 0.51337 0.0019714 0.42271 1.4323 1.4293 16.0085 144.9836 0.00031841 -85.1075 0.23521
0.33923 0.98802 5.5235e-05 3.8182 0.012046 4.471e-06 0.001154 0.075193 0.00065537 0.075843 0.067974 0 0.042481 0.0389 0 0.85181 0.22986 0.059821 0.0084656 4.1107 0.053171 6.3458e-05 0.83689 0.0051105 0.0058484 0.0015165 0.98523 0.99056 3.2892e-06 1.3157e-05 0.1305 0.78186 0.82064 0.0014647 0.86948 0.51354 0.0019707 0.42272 1.4339 1.4309 16.0085 144.9836 0.00031769 -85.1115 0.23621
0.34023 0.98802 5.5235e-05 3.8182 0.012046 4.4842e-06 0.001154 0.075321 0.00065538 0.075972 0.068091 0 0.04247 0.0389 0 0.85184 0.22987 0.059827 0.0084663 4.1107 0.053175 6.3463e-05 0.83689 0.0051106 0.0058484 0.0015166 0.98524 0.99057 3.2869e-06 1.3148e-05 0.1305 0.78249 0.82108 0.0014642 0.87027 0.5137 0.00197 0.42272 1.4354 1.4324 16.0086 144.9837 0.00031698 -85.1154 0.23721
0.34123 0.98802 5.5235e-05 3.8182 0.012045 4.4974e-06 0.001154 0.07545 0.00065539 0.0761 0.068209 0 0.04246 0.0389 0 0.85188 0.22989 0.059832 0.008467 4.1108 0.053179 6.3468e-05 0.83688 0.0051107 0.0058485 0.001515 0.98525 0.99058 3.2846e-06 1.3139e-05 0.1305 0.78311 0.82152 0.0014637 0.87105 0.51387 0.0019694 0.42273 1.4369 1.4339 16.0086 144.9837 0.00031626 -85.1193 0.23821
0.34223 0.98802 5.5235e-05 3.8182 0.012045 4.5106e-06 0.001154 0.075578 0.0006554 0.076229 0.068327 0 0.042449 0.0389 0 0.85191 0.2299 0.059838 0.0084677 4.1108 0.053183 6.3473e-05 0.83688 0.0051107 0.0058485 0.0015141 0.98527 0.99059 3.2823e-06 1.313e-05 0.1305 0.78374 0.82195 0.0014632 0.87182 0.51404 0.0019687 0.42274 1.4385 1.4355 16.0086 144.9837 0.00031556 -85.1232 0.23921
0.34323 0.98802 5.5235e-05 3.8182 0.012045 4.5237e-06 0.001154 0.075706 0.00065541 0.076357 0.068444 0 0.042438 0.0389 0 0.85195 0.22992 0.059844 0.0084684 4.1109 0.053186 6.3478e-05 0.83688 0.0051108 0.0058486 0.0015131 0.98528 0.9906 3.2801e-06 1.3121e-05 0.1305 0.78436 0.82239 0.0014627 0.87259 0.5142 0.0019681 0.42275 1.44 1.437 16.0087 144.9837 0.00031485 -85.1271 0.24021
0.34423 0.98802 5.5235e-05 3.8182 0.012045 4.5369e-06 0.001154 0.075834 0.00065542 0.076485 0.068562 0 0.042428 0.0389 0 0.85198 0.22994 0.059849 0.0084692 4.1109 0.05319 6.3482e-05 0.83687 0.0051108 0.0058486 0.0015121 0.98529 0.99061 3.2779e-06 1.3112e-05 0.1305 0.78497 0.82282 0.0014622 0.87336 0.51437 0.0019674 0.42276 1.4415 1.4385 16.0087 144.9837 0.00031415 -85.1309 0.24121
0.34523 0.98802 5.5235e-05 3.8182 0.012045 4.5501e-06 0.001154 0.075962 0.00065543 0.076613 0.068679 0 0.042417 0.0389 0 0.85202 0.22995 0.059855 0.0084699 4.111 0.053194 6.3487e-05 0.83687 0.0051109 0.0058487 0.0015112 0.98531 0.99062 3.2757e-06 1.3103e-05 0.1305 0.78559 0.82325 0.0014618 0.87412 0.51453 0.0019668 0.42277 1.443 1.4401 16.0087 144.9837 0.00031345 -85.1347 0.24221
0.34623 0.98802 5.5235e-05 3.8182 0.012045 4.5632e-06 0.001154 0.07609 0.00065544 0.076741 0.068797 0 0.042406 0.0389 0 0.85206 0.22997 0.059861 0.0084706 4.111 0.053198 6.3492e-05 0.83687 0.005111 0.0058488 0.0015102 0.98532 0.99063 3.2735e-06 1.3094e-05 0.13051 0.78621 0.82368 0.0014613 0.87488 0.5147 0.0019662 0.42278 1.4445 1.4416 16.0087 144.9838 0.00031276 -85.1385 0.24321
0.34723 0.98802 5.5235e-05 3.8182 0.012045 4.5764e-06 0.001154 0.076218 0.00065545 0.076869 0.068914 0 0.042396 0.0389 0 0.85209 0.22998 0.059866 0.0084713 4.1111 0.053202 6.3497e-05 0.83686 0.005111 0.0058488 0.0015093 0.98533 0.99063 3.2713e-06 1.3085e-05 0.13051 0.78682 0.8241 0.0014608 0.87563 0.51487 0.0019655 0.42279 1.446 1.4431 16.0088 144.9838 0.00031207 -85.1423 0.24421
0.34823 0.98802 5.5235e-05 3.8182 0.012045 4.5896e-06 0.001154 0.076346 0.00065546 0.076997 0.069031 0 0.042385 0.0389 0 0.85213 0.23 0.059872 0.008472 4.1111 0.053205 6.3502e-05 0.83686 0.0051111 0.0058489 0.0015083 0.98534 0.99064 3.2691e-06 1.3077e-05 0.13051 0.78743 0.82453 0.0014603 0.87638 0.51503 0.0019649 0.4228 1.4475 1.4446 16.0088 144.9838 0.00031138 -85.146 0.24521
0.34923 0.98802 5.5235e-05 3.8182 0.012045 4.6028e-06 0.001154 0.076473 0.00065547 0.077124 0.069148 0 0.042375 0.0389 0 0.85216 0.23002 0.059878 0.0084728 4.1111 0.053209 6.3507e-05 0.83685 0.0051111 0.005849 0.0015074 0.98536 0.99065 3.267e-06 1.3068e-05 0.13051 0.78804 0.82495 0.0014598 0.87713 0.5152 0.0019643 0.42281 1.449 1.4461 16.0088 144.9838 0.00031069 -85.1497 0.24621
0.35023 0.98802 5.5235e-05 3.8182 0.012045 4.6159e-06 0.001154 0.076601 0.00065548 0.077252 0.069265 0 0.042364 0.0389 0 0.8522 0.23003 0.059884 0.0084735 4.1112 0.053213 6.3511e-05 0.83685 0.0051112 0.005849 0.0015065 0.98537 0.99066 3.2649e-06 1.306e-05 0.13051 0.78865 0.82537 0.0014594 0.87787 0.51536 0.0019637 0.42282 1.4505 1.4476 16.0088 144.9838 0.00031001 -85.1534 0.24721
0.35123 0.98802 5.5234e-05 3.8182 0.012045 4.6291e-06 0.001154 0.076728 0.00065549 0.077379 0.069382 0 0.042354 0.0389 0 0.85224 0.23005 0.05989 0.0084742 4.1112 0.053217 6.3516e-05 0.83685 0.0051113 0.0058491 0.0015055 0.98538 0.99067 3.2628e-06 1.3051e-05 0.13051 0.78926 0.82579 0.0014589 0.8786 0.51553 0.0019631 0.42283 1.452 1.4491 16.0089 144.9838 0.00030933 -85.157 0.24821
0.35223 0.98802 5.5234e-05 3.8182 0.012045 4.6423e-06 0.001154 0.076856 0.0006555 0.077507 0.069499 0 0.042343 0.0389 0 0.85227 0.23006 0.059895 0.008475 4.1113 0.053221 6.3521e-05 0.83684 0.0051113 0.0058491 0.0015046 0.98539 0.99068 3.2607e-06 1.3043e-05 0.13051 0.78986 0.8262 0.0014584 0.87934 0.5157 0.0019625 0.42284 1.4535 1.4506 16.0089 144.9839 0.00030866 -85.1606 0.24921
0.35323 0.98802 5.5234e-05 3.8182 0.012045 4.6554e-06 0.001154 0.076983 0.00065551 0.077634 0.069616 0 0.042332 0.0389 0 0.85231 0.23008 0.059901 0.0084757 4.1113 0.053225 6.3526e-05 0.83684 0.0051114 0.0058492 0.0015037 0.9854 0.99069 3.2586e-06 1.3035e-05 0.13051 0.79046 0.82662 0.001458 0.88006 0.51586 0.0019619 0.42285 1.455 1.4521 16.0089 144.9839 0.00030798 -85.1642 0.25021
0.35423 0.98802 5.5234e-05 3.8182 0.012045 4.6686e-06 0.001154 0.07711 0.00065552 0.077761 0.069732 0 0.042322 0.0389 0 0.85235 0.2301 0.059907 0.0084764 4.1114 0.053229 6.3531e-05 0.83683 0.0051115 0.0058493 0.0015028 0.98542 0.99069 3.2565e-06 1.3026e-05 0.13051 0.79106 0.82703 0.0014575 0.88079 0.51603 0.0019613 0.42286 1.4565 1.4536 16.0089 144.9839 0.00030731 -85.1678 0.25121
0.35523 0.98802 5.5234e-05 3.8182 0.012045 4.6818e-06 0.001154 0.077237 0.00065553 0.077888 0.069849 0 0.042311 0.0389 0 0.85238 0.23011 0.059913 0.0084772 4.1114 0.053232 6.3536e-05 0.83683 0.0051115 0.0058493 0.001502 0.98543 0.9907 3.2545e-06 1.3018e-05 0.13051 0.79166 0.82744 0.0014571 0.88151 0.51619 0.0019607 0.42287 1.458 1.4551 16.0089 144.9839 0.00030665 -85.1713 0.25221
0.35623 0.98802 5.5234e-05 3.8182 0.012045 4.695e-06 0.001154 0.077364 0.00065554 0.078015 0.069965 0 0.042301 0.0389 0 0.85242 0.23013 0.059919 0.0084779 4.1115 0.053236 6.3541e-05 0.83683 0.0051116 0.0058494 0.0015011 0.98544 0.99071 3.2525e-06 1.301e-05 0.13051 0.79226 0.82785 0.0014566 0.88222 0.51636 0.0019601 0.42288 1.4594 1.4566 16.009 144.9839 0.00030598 -85.1749 0.25321
0.35723 0.98802 5.5234e-05 3.8182 0.012045 4.7081e-06 0.001154 0.077491 0.00065555 0.078142 0.070082 0 0.042291 0.0389 0 0.85246 0.23014 0.059925 0.0084786 4.1115 0.05324 6.3546e-05 0.83682 0.0051117 0.0058495 0.0015002 0.98545 0.99072 3.2505e-06 1.3002e-05 0.13051 0.79285 0.82825 0.0014562 0.88294 0.51653 0.0019595 0.42289 1.4609 1.4581 16.009 144.9839 0.00030532 -85.1784 0.25421
0.35823 0.98802 5.5234e-05 3.8182 0.012045 4.7213e-06 0.001154 0.077618 0.00065556 0.078269 0.070198 0 0.04228 0.0389 0 0.8525 0.23016 0.05993 0.0084794 4.1116 0.053244 6.3551e-05 0.83682 0.0051117 0.0058495 0.0014993 0.98546 0.99073 3.2485e-06 1.2994e-05 0.13051 0.79345 0.82866 0.0014557 0.88364 0.51669 0.0019589 0.4229 1.4624 1.4596 16.009 144.984 0.00030467 -85.1818 0.25521
0.35923 0.98802 5.5234e-05 3.8182 0.012045 4.7345e-06 0.001154 0.077744 0.00065557 0.078395 0.070314 0 0.04227 0.0389 0 0.85253 0.23018 0.059936 0.0084801 4.1116 0.053248 6.3556e-05 0.83682 0.0051118 0.0058496 0.0014985 0.98547 0.99073 3.2465e-06 1.2986e-05 0.13051 0.79404 0.82906 0.0014553 0.88435 0.51686 0.0019584 0.42291 1.4638 1.461 16.009 144.984 0.00030401 -85.1853 0.25621
0.36023 0.98802 5.5234e-05 3.8182 0.012045 4.7476e-06 0.001154 0.077871 0.00065558 0.078522 0.07043 0 0.042259 0.0389 0 0.85257 0.23019 0.059942 0.0084809 4.1117 0.053252 6.3561e-05 0.83681 0.0051119 0.0058496 0.0014976 0.98549 0.99074 3.2445e-06 1.2978e-05 0.13051 0.79463 0.82946 0.0014549 0.88505 0.51702 0.0019578 0.42292 1.4653 1.4625 16.0091 144.984 0.00030336 -85.1887 0.25721
0.36123 0.98802 5.5234e-05 3.8182 0.012045 4.7608e-06 0.001154 0.077997 0.00065559 0.078648 0.070546 0 0.042249 0.0389 0 0.85261 0.23021 0.059948 0.0084816 4.1118 0.053256 6.3566e-05 0.83681 0.0051119 0.0058497 0.0014968 0.9855 0.99075 3.2426e-06 1.2971e-05 0.13051 0.79522 0.82986 0.0014544 0.88574 0.51719 0.0019572 0.42293 1.4667 1.464 16.0091 144.984 0.00030271 -85.1921 0.25821
0.36223 0.98802 5.5234e-05 3.8182 0.012045 4.774e-06 0.001154 0.078124 0.0006556 0.078775 0.070662 0 0.042238 0.0389 0 0.85264 0.23023 0.059954 0.0084824 4.1118 0.05326 6.3571e-05 0.8368 0.005112 0.0058498 0.0014959 0.98551 0.99076 3.2407e-06 1.2963e-05 0.13051 0.7958 0.83026 0.001454 0.88643 0.51735 0.0019567 0.42294 1.4682 1.4654 16.0091 144.984 0.00030207 -85.1954 0.25921
0.36323 0.98802 5.5234e-05 3.8182 0.012045 4.7872e-06 0.001154 0.07825 0.00065561 0.078901 0.070778 0 0.042228 0.0389 0 0.85268 0.23024 0.05996 0.0084831 4.1119 0.053264 6.3576e-05 0.8368 0.0051121 0.0058498 0.0014951 0.98552 0.99076 3.2388e-06 1.2955e-05 0.13051 0.79639 0.83065 0.0014536 0.88712 0.51752 0.0019561 0.42295 1.4696 1.4669 16.0091 144.984 0.00030143 -85.1988 0.26021
0.36423 0.98802 5.5234e-05 3.8182 0.012045 4.8003e-06 0.001154 0.078376 0.00065561 0.079027 0.070894 0 0.042218 0.0389 0 0.85272 0.23026 0.059966 0.0084839 4.1119 0.053268 6.3581e-05 0.8368 0.0051121 0.0058499 0.0014943 0.98553 0.99077 3.2369e-06 1.2948e-05 0.13051 0.79697 0.83105 0.0014532 0.8878 0.51768 0.0019556 0.42296 1.4711 1.4683 16.0091 144.9841 0.00030079 -85.2021 0.26121
0.36523 0.98802 5.5234e-05 3.8182 0.012045 4.8135e-06 0.001154 0.078502 0.00065562 0.079153 0.071009 0 0.042207 0.0389 0 0.85276 0.23028 0.059972 0.0084846 4.112 0.053272 6.3586e-05 0.83679 0.0051122 0.00585 0.0014935 0.98554 0.99078 3.235e-06 1.294e-05 0.13052 0.79755 0.83144 0.0014528 0.88848 0.51785 0.001955 0.42297 1.4725 1.4698 16.0092 144.9841 0.00030015 -85.2054 0.26221
0.36623 0.98802 5.5234e-05 3.8182 0.012045 4.8267e-06 0.001154 0.078628 0.00065563 0.079279 0.071125 0 0.042197 0.0389 0 0.85279 0.23029 0.059978 0.0084854 4.112 0.053276 6.3592e-05 0.83679 0.0051123 0.00585 0.0014927 0.98555 0.99079 3.2331e-06 1.2933e-05 0.13052 0.79813 0.83183 0.0014523 0.88916 0.51802 0.0019545 0.42298 1.474 1.4712 16.0092 144.9841 0.00029952 -85.2086 0.26321
0.36723 0.98802 5.5234e-05 3.8182 0.012045 4.8398e-06 0.001154 0.078754 0.00065564 0.079405 0.07124 0 0.042187 0.0389 0 0.85283 0.23031 0.059984 0.0084861 4.1121 0.05328 6.3597e-05 0.83678 0.0051123 0.0058501 0.0014918 0.98556 0.99079 3.2312e-06 1.2925e-05 0.13052 0.7987 0.83222 0.0014519 0.88983 0.51818 0.0019539 0.42299 1.4754 1.4727 16.0092 144.9841 0.00029889 -85.2119 0.26421
0.36823 0.98802 5.5233e-05 3.8182 0.012045 4.853e-06 0.001154 0.078879 0.00065565 0.079531 0.071356 0 0.042176 0.0389 0 0.85287 0.23033 0.05999 0.0084869 4.1121 0.053284 6.3602e-05 0.83678 0.0051124 0.0058502 0.001491 0.98557 0.9908 3.2294e-06 1.2918e-05 0.13052 0.79928 0.8326 0.0014515 0.89049 0.51835 0.0019534 0.423 1.4768 1.4741 16.0092 144.9841 0.00029826 -85.2151 0.26521
0.36923 0.98802 5.5233e-05 3.8182 0.012045 4.8662e-06 0.001154 0.079005 0.00065566 0.079656 0.071471 0 0.042166 0.0389 0 0.85291 0.23034 0.059996 0.0084876 4.1122 0.053288 6.3607e-05 0.83678 0.0051125 0.0058502 0.0014903 0.98558 0.99081 3.2276e-06 1.291e-05 0.13052 0.79985 0.83299 0.0014511 0.89116 0.51851 0.0019529 0.42301 1.4782 1.4755 16.0092 144.9841 0.00029764 -85.2183 0.26621
0.37023 0.98802 5.5233e-05 3.8182 0.012045 4.8794e-06 0.001154 0.079131 0.00065567 0.079782 0.071586 0 0.042156 0.0389 0 0.85295 0.23036 0.060002 0.0084884 4.1122 0.053292 6.3612e-05 0.83677 0.0051125 0.0058503 0.0014895 0.98559 0.99082 3.2258e-06 1.2903e-05 0.13052 0.80042 0.83337 0.0014507 0.89182 0.51868 0.0019523 0.42302 1.4797 1.477 16.0093 144.9842 0.00029701 -85.2215 0.26721
0.37123 0.98802 5.5233e-05 3.8182 0.012045 4.8925e-06 0.001154 0.079256 0.00065568 0.079907 0.071701 0 0.042145 0.0389 0 0.85298 0.23038 0.060008 0.0084891 4.1123 0.053296 6.3617e-05 0.83677 0.0051126 0.0058504 0.0014887 0.9856 0.99082 3.224e-06 1.2896e-05 0.13052 0.80099 0.83375 0.0014503 0.89247 0.51884 0.0019518 0.42303 1.4811 1.4784 16.0093 144.9842 0.0002964 -85.2246 0.26821
0.37223 0.98802 5.5233e-05 3.8182 0.012045 4.9057e-06 0.001154 0.079381 0.00065569 0.080032 0.071816 0 0.042135 0.0389 0 0.85302 0.23039 0.060014 0.0084899 4.1123 0.053301 6.3622e-05 0.83676 0.0051127 0.0058504 0.0014879 0.98561 0.99083 3.2222e-06 1.2889e-05 0.13052 0.80156 0.83413 0.0014499 0.89312 0.51901 0.0019513 0.42304 1.4825 1.4798 16.0093 144.9842 0.00029578 -85.2277 0.26921
0.37323 0.98802 5.5233e-05 3.8182 0.012045 4.9189e-06 0.001154 0.079507 0.0006557 0.080158 0.071931 0 0.042125 0.0389 0 0.85306 0.23041 0.06002 0.0084907 4.1124 0.053305 6.3628e-05 0.83676 0.0051127 0.0058505 0.0014871 0.98563 0.99084 3.2204e-06 1.2882e-05 0.13052 0.80213 0.83451 0.0014495 0.89377 0.51917 0.0019508 0.42305 1.4839 1.4812 16.0093 144.9842 0.00029517 -85.2308 0.27021
0.37423 0.98802 5.5233e-05 3.8182 0.012045 4.932e-06 0.001154 0.079632 0.0006557 0.080283 0.072046 0 0.042115 0.0389 0 0.8531 0.23043 0.060026 0.0084914 4.1125 0.053309 6.3633e-05 0.83675 0.0051128 0.0058506 0.0014864 0.98564 0.99084 3.2187e-06 1.2875e-05 0.13052 0.80269 0.83489 0.0014491 0.89442 0.51934 0.0019503 0.42306 1.4853 1.4826 16.0093 144.9842 0.00029456 -85.2339 0.27121
0.37523 0.98802 5.5233e-05 3.8182 0.012045 4.9452e-06 0.001154 0.079757 0.00065571 0.080408 0.072161 0 0.042104 0.0389 0 0.85314 0.23044 0.060032 0.0084922 4.1125 0.053313 6.3638e-05 0.83675 0.0051129 0.0058507 0.0014856 0.98565 0.99085 3.2169e-06 1.2868e-05 0.13052 0.80326 0.83526 0.0014487 0.89506 0.5195 0.0019498 0.42308 1.4867 1.4841 16.0094 144.9842 0.00029395 -85.237 0.27221
0.37623 0.98802 5.5233e-05 3.8182 0.012045 4.9584e-06 0.001154 0.079882 0.00065572 0.080533 0.072276 0 0.042094 0.0389 0 0.85318 0.23046 0.060038 0.008493 4.1126 0.053317 6.3643e-05 0.83675 0.0051129 0.0058507 0.0014849 0.98566 0.99086 3.2152e-06 1.2861e-05 0.13052 0.80382 0.83563 0.0014484 0.89569 0.51967 0.0019493 0.42309 1.4881 1.4855 16.0094 144.9843 0.00029334 -85.24 0.27321
0.37723 0.98802 5.5233e-05 3.8182 0.012045 4.9716e-06 0.001154 0.080006 0.00065573 0.080658 0.07239 0 0.042084 0.0389 0 0.85321 0.23048 0.060045 0.0084937 4.1126 0.053321 6.3649e-05 0.83674 0.005113 0.0058508 0.0014841 0.98567 0.99086 3.2135e-06 1.2854e-05 0.13052 0.80438 0.83601 0.001448 0.89632 0.51983 0.0019488 0.4231 1.4895 1.4869 16.0094 144.9843 0.00029274 -85.243 0.27421
0.37823 0.98802 5.5233e-05 3.8182 0.012045 4.9847e-06 0.001154 0.080131 0.00065574 0.080782 0.072505 0 0.042074 0.0389 0 0.85325 0.23049 0.060051 0.0084945 4.1127 0.053325 6.3654e-05 0.83674 0.0051131 0.0058509 0.0014834 0.98567 0.99087 3.2118e-06 1.2847e-05 0.13052 0.80493 0.83637 0.0014476 0.89695 0.52 0.0019483 0.42311 1.4909 1.4883 16.0094 144.9843 0.00029214 -85.246 0.27521
0.37923 0.98802 5.5233e-05 3.8182 0.012045 4.9979e-06 0.001154 0.080256 0.00065575 0.080907 0.072619 0 0.042063 0.0389 0 0.85329 0.23051 0.060057 0.0084953 4.1127 0.053329 6.3659e-05 0.83673 0.0051132 0.0058509 0.0014827 0.98568 0.99088 3.2101e-06 1.284e-05 0.13052 0.80549 0.83674 0.0014472 0.89758 0.52016 0.0019478 0.42312 1.4923 1.4897 16.0094 144.9843 0.00029155 -85.249 0.27621
0.38023 0.98802 5.5233e-05 3.8182 0.012045 5.0111e-06 0.001154 0.08038 0.00065576 0.081031 0.072734 0 0.042053 0.0389 0 0.85333 0.23053 0.060063 0.0084961 4.1128 0.053334 6.3664e-05 0.83673 0.0051132 0.005851 0.0014819 0.98569 0.99088 3.2084e-06 1.2834e-05 0.13052 0.80604 0.83711 0.0014468 0.8982 0.52033 0.0019473 0.42313 1.4936 1.491 16.0095 144.9843 0.00029095 -85.2519 0.27721
0.38123 0.98802 5.5233e-05 3.8182 0.012045 5.0242e-06 0.001154 0.080505 0.00065577 0.081156 0.072848 0 0.042043 0.0389 0 0.85337 0.23055 0.060069 0.0084968 4.1128 0.053338 6.367e-05 0.83673 0.0051133 0.0058511 0.0014812 0.9857 0.99089 3.2068e-06 1.2827e-05 0.13052 0.8066 0.83747 0.0014465 0.89882 0.52049 0.0019468 0.42314 1.495 1.4924 16.0095 144.9843 0.00029036 -85.2548 0.27821
0.38223 0.98802 5.5233e-05 3.8182 0.012045 5.0374e-06 0.001154 0.080629 0.00065577 0.08128 0.072962 0 0.042033 0.0389 0 0.85341 0.23056 0.060075 0.0084976 4.1129 0.053342 6.3675e-05 0.83672 0.0051134 0.0058511 0.0014805 0.98571 0.9909 3.2051e-06 1.2821e-05 0.13053 0.80715 0.83784 0.0014461 0.89943 0.52066 0.0019463 0.42315 1.4964 1.4938 16.0095 144.9844 0.00028977 -85.2577 0.27921
0.38323 0.98802 5.5233e-05 3.8182 0.012045 5.0506e-06 0.001154 0.080753 0.00065578 0.081404 0.073076 0 0.042023 0.0389 0 0.85345 0.23058 0.060081 0.0084984 4.113 0.053346 6.368e-05 0.83672 0.0051135 0.0058512 0.0014798 0.98572 0.9909 3.2035e-06 1.2814e-05 0.13053 0.8077 0.8382 0.0014457 0.90004 0.52082 0.0019459 0.42316 1.4978 1.4952 16.0095 144.9844 0.00028919 -85.2606 0.28021
0.38423 0.98802 5.5232e-05 3.8182 0.012045 5.0638e-06 0.001154 0.080877 0.00065579 0.081529 0.07319 0 0.042013 0.0389 0 0.85349 0.2306 0.060088 0.0084992 4.113 0.05335 6.3686e-05 0.83671 0.0051135 0.0058513 0.0014791 0.98573 0.99091 3.2019e-06 1.2808e-05 0.13053 0.80824 0.83856 0.0014454 0.90065 0.52099 0.0019454 0.42317 1.4991 1.4966 16.0095 144.9844 0.00028861 -85.2635 0.28121
0.38523 0.98802 5.5232e-05 3.8182 0.012045 5.0769e-06 0.001154 0.081001 0.0006558 0.081653 0.073304 0 0.042003 0.0389 0 0.85353 0.23061 0.060094 0.0085 4.1131 0.053355 6.3691e-05 0.83671 0.0051136 0.0058514 0.0014784 0.98574 0.99091 3.2003e-06 1.2801e-05 0.13053 0.80879 0.83892 0.001445 0.90125 0.52115 0.0019449 0.42318 1.5005 1.4979 16.0095 144.9844 0.00028803 -85.2663 0.28221
0.38623 0.98802 5.5232e-05 3.8182 0.012045 5.0901e-06 0.001154 0.081125 0.00065581 0.081777 0.073418 0 0.041993 0.0389 0 0.85356 0.23063 0.0601 0.0085007 4.1131 0.053359 6.3697e-05 0.8367 0.0051137 0.0058514 0.0014777 0.98575 0.99092 3.1987e-06 1.2795e-05 0.13053 0.80933 0.83927 0.0014447 0.90185 0.52131 0.0019444 0.42319 1.5019 1.4993 16.0096 144.9844 0.00028745 -85.2692 0.28321
0.38723 0.98802 5.5232e-05 3.8182 0.012045 5.1033e-06 0.001154 0.081249 0.00065582 0.0819 0.073532 0 0.041982 0.0389 0 0.8536 0.23065 0.060106 0.0085015 4.1132 0.053363 6.3702e-05 0.8367 0.0051138 0.0058515 0.001477 0.98576 0.99093 3.1971e-06 1.2788e-05 0.13053 0.80987 0.83963 0.0014443 0.90245 0.52148 0.001944 0.4232 1.5032 1.5007 16.0096 144.9845 0.00028687 -85.272 0.28421
0.38823 0.98802 5.5232e-05 3.8182 0.012045 5.1164e-06 0.001154 0.081373 0.00065582 0.082024 0.073645 0 0.041972 0.0389 0 0.85364 0.23067 0.060113 0.0085023 4.1133 0.053367 6.3707e-05 0.8367 0.0051138 0.0058516 0.0014763 0.98577 0.99093 3.1955e-06 1.2782e-05 0.13053 0.81042 0.83998 0.001444 0.90304 0.52164 0.0019435 0.42321 1.5046 1.502 16.0096 144.9845 0.0002863 -85.2747 0.28521
0.38923 0.98802 5.5232e-05 3.8182 0.012045 5.1296e-06 0.001154 0.081496 0.00065583 0.082148 0.073759 0 0.041962 0.0389 0 0.85368 0.23068 0.060119 0.0085031 4.1133 0.053372 6.3713e-05 0.83669 0.0051139 0.0058517 0.0014756 0.98578 0.99094 3.1939e-06 1.2776e-05 0.13053 0.81095 0.84033 0.0014436 0.90363 0.52181 0.0019431 0.42323 1.5059 1.5034 16.0096 144.9845 0.00028573 -85.2775 0.28621
0.39023 0.98802 5.5232e-05 3.8182 0.012045 5.1428e-06 0.001154 0.08162 0.00065584 0.082271 0.073872 0 0.041952 0.0389 0 0.85372 0.2307 0.060125 0.0085039 4.1134 0.053376 6.3718e-05 0.83669 0.005114 0.0058517 0.0014749 0.98579 0.99095 3.1924e-06 1.277e-05 0.13053 0.81149 0.84068 0.0014433 0.90421 0.52197 0.0019426 0.42324 1.5073 1.5048 16.0096 144.9845 0.00028516 -85.2802 0.28721
0.39123 0.98802 5.5232e-05 3.8182 0.012045 5.1559e-06 0.001154 0.081743 0.00065585 0.082395 0.073986 0 0.041942 0.0389 0 0.85376 0.23072 0.060131 0.0085047 4.1134 0.05338 6.3724e-05 0.83668 0.0051141 0.0058518 0.0014743 0.9858 0.99095 3.1909e-06 1.2763e-05 0.13053 0.81203 0.84103 0.0014429 0.9048 0.52214 0.0019422 0.42325 1.5086 1.5061 16.0096 144.9845 0.0002846 -85.283 0.28821
0.39223 0.98802 5.5232e-05 3.8182 0.012045 5.1691e-06 0.001154 0.081867 0.00065586 0.082518 0.074099 0 0.041932 0.0389 0 0.8538 0.23074 0.060138 0.0085055 4.1135 0.053385 6.3729e-05 0.83668 0.0051141 0.0058519 0.0014736 0.9858 0.99096 3.1893e-06 1.2757e-05 0.13053 0.81256 0.84138 0.0014426 0.90537 0.5223 0.0019417 0.42326 1.5099 1.5075 16.0096 144.9845 0.00028404 -85.2857 0.28921
0.39323 0.98802 5.5232e-05 3.8182 0.012045 5.1823e-06 0.001154 0.08199 0.00065587 0.082641 0.074212 0 0.041922 0.0389 0 0.85384 0.23075 0.060144 0.0085063 4.1136 0.053389 6.3735e-05 0.83667 0.0051142 0.005852 0.001473 0.98581 0.99096 3.1878e-06 1.2751e-05 0.13053 0.81309 0.84172 0.0014422 0.90595 0.52247 0.0019413 0.42327 1.5113 1.5088 16.0097 144.9846 0.00028348 -85.2883 0.29021
0.39423 0.98802 5.5232e-05 3.8182 0.012045 5.1955e-06 0.001154 0.082113 0.00065587 0.082764 0.074325 0 0.041912 0.0389 0 0.85388 0.23077 0.06015 0.0085071 4.1136 0.053393 6.374e-05 0.83667 0.0051143 0.005852 0.0014723 0.98582 0.99097 3.1863e-06 1.2745e-05 0.13053 0.81362 0.84207 0.0014419 0.90652 0.52263 0.0019408 0.42328 1.5126 1.5101 16.0097 144.9846 0.00028292 -85.291 0.29121
0.39523 0.98802 5.5232e-05 3.8182 0.012045 5.2086e-06 0.001154 0.082236 0.00065588 0.082887 0.074438 0 0.041902 0.0389 0 0.85392 0.23079 0.060157 0.0085079 4.1137 0.053398 6.3746e-05 0.83667 0.0051144 0.0058521 0.0014717 0.98583 0.99097 3.1848e-06 1.2739e-05 0.13053 0.81415 0.84241 0.0014416 0.90709 0.52279 0.0019404 0.42329 1.5139 1.5115 16.0097 144.9846 0.00028237 -85.2936 0.29221
0.39623 0.98802 5.5232e-05 3.8182 0.012045 5.2218e-06 0.001154 0.082359 0.00065589 0.08301 0.074551 0 0.041892 0.0389 0 0.85396 0.23081 0.060163 0.0085087 4.1137 0.053402 6.3751e-05 0.83666 0.0051144 0.0058522 0.001471 0.98584 0.99098 3.1833e-06 1.2733e-05 0.13053 0.81468 0.84275 0.0014412 0.90765 0.52296 0.00194 0.4233 1.5153 1.5128 16.0097 144.9846 0.00028182 -85.2963 0.29321
0.39723 0.98802 5.5232e-05 3.8182 0.012045 5.235e-06 0.001154 0.082482 0.0006559 0.083133 0.074664 0 0.041882 0.0389 0 0.854 0.23082 0.060169 0.0085095 4.1138 0.053406 6.3757e-05 0.83666 0.0051145 0.0058523 0.0014704 0.98585 0.99099 3.1819e-06 1.2728e-05 0.13053 0.81521 0.84309 0.0014409 0.90821 0.52312 0.0019395 0.42331 1.5166 1.5141 16.0097 144.9846 0.00028127 -85.2989 0.29421
0.39823 0.98802 5.5232e-05 3.8182 0.012045 5.2481e-06 0.001154 0.082605 0.00065591 0.083256 0.074777 0 0.041872 0.0389 0 0.85404 0.23084 0.060176 0.0085103 4.1139 0.053411 6.3762e-05 0.83665 0.0051146 0.0058523 0.0014697 0.98586 0.99099 3.1804e-06 1.2722e-05 0.13054 0.81573 0.84343 0.0014406 0.90877 0.52329 0.0019391 0.42333 1.5179 1.5155 16.0097 144.9846 0.00028072 -85.3015 0.29521
0.39923 0.98802 5.5232e-05 3.8182 0.012045 5.2613e-06 0.001154 0.082727 0.00065591 0.083379 0.07489 0 0.041862 0.0389 0 0.85408 0.23086 0.060182 0.0085111 4.1139 0.053415 6.3768e-05 0.83665 0.0051147 0.0058524 0.0014691 0.98586 0.991 3.179e-06 1.2716e-05 0.13054 0.81625 0.84377 0.0014403 0.90933 0.52345 0.0019387 0.42334 1.5192 1.5168 16.0097 144.9847 0.00028017 -85.304 0.29621
0.40023 0.98802 5.5231e-05 3.8182 0.012045 5.2745e-06 0.001154 0.08285 0.00065592 0.083501 0.075002 0 0.041852 0.0389 0 0.85412 0.23088 0.060189 0.0085119 4.114 0.053419 6.3773e-05 0.83664 0.0051147 0.0058525 0.0014685 0.98587 0.991 3.1775e-06 1.271e-05 0.13054 0.81677 0.8441 0.0014399 0.90988 0.52361 0.0019383 0.42335 1.5205 1.5181 16.0098 144.9847 0.00027963 -85.3066 0.29721
0.40123 0.98802 5.5231e-05 3.8182 0.012045 5.2876e-06 0.001154 0.082972 0.00065593 0.083624 0.075115 0 0.041843 0.0389 0 0.85416 0.2309 0.060195 0.0085127 4.114 0.053424 6.3779e-05 0.83664 0.0051148 0.0058526 0.0014679 0.98588 0.99101 3.1761e-06 1.2705e-05 0.13054 0.81729 0.84444 0.0014396 0.91043 0.52378 0.0019379 0.42336 1.5218 1.5194 16.0098 144.9847 0.00027909 -85.3091 0.29821
0.40223 0.98802 5.5231e-05 3.8182 0.012045 5.3008e-06 0.001154 0.083095 0.00065594 0.083746 0.075227 0 0.041833 0.0389 0 0.8542 0.23091 0.060201 0.0085135 4.1141 0.053428 6.3785e-05 0.83664 0.0051149 0.0058526 0.0014672 0.98589 0.99101 3.1747e-06 1.2699e-05 0.13054 0.81781 0.84477 0.0014393 0.91097 0.52394 0.0019374 0.42337 1.5231 1.5207 16.0098 144.9847 0.00027856 -85.3116 0.29921
0.40323 0.98802 5.5231e-05 3.8182 0.012045 5.314e-06 0.001154 0.083217 0.00065595 0.083868 0.07534 0 0.041823 0.0389 0 0.85424 0.23093 0.060208 0.0085143 4.1142 0.053433 6.379e-05 0.83663 0.005115 0.0058527 0.0014666 0.9859 0.99102 3.1733e-06 1.2693e-05 0.13054 0.81833 0.8451 0.001439 0.91151 0.52411 0.001937 0.42338 1.5244 1.522 16.0098 144.9847 0.00027802 -85.3141 0.30021
0.40423 0.98802 5.5231e-05 3.8182 0.012045 5.3272e-06 0.001154 0.083339 0.00065595 0.08399 0.075452 0 0.041813 0.0389 0 0.85428 0.23095 0.060214 0.0085151 4.1142 0.053437 6.3796e-05 0.83663 0.0051151 0.0058528 0.001466 0.9859 0.99102 3.1719e-06 1.2688e-05 0.13054 0.81884 0.84543 0.0014387 0.91205 0.52427 0.0019366 0.42339 1.5257 1.5233 16.0098 144.9847 0.00027749 -85.3166 0.30121
0.40523 0.98802 5.5231e-05 3.8182 0.012045 5.3403e-06 0.001154 0.083461 0.00065596 0.084112 0.075564 0 0.041803 0.0389 0 0.85433 0.23097 0.060221 0.0085159 4.1143 0.053441 6.3801e-05 0.83662 0.0051151 0.0058529 0.0014654 0.98591 0.99103 3.1705e-06 1.2682e-05 0.13054 0.81935 0.84576 0.0014384 0.91258 0.52443 0.0019362 0.4234 1.527 1.5246 16.0098 144.9848 0.00027696 -85.319 0.30221
0.40623 0.98802 5.5231e-05 3.8182 0.012045 5.3535e-06 0.001154 0.083583 0.00065597 0.084234 0.075676 0 0.041793 0.0389 0 0.85437 0.23099 0.060227 0.0085168 4.1144 0.053446 6.3807e-05 0.83662 0.0051152 0.005853 0.0014648 0.98592 0.99103 3.1692e-06 1.2677e-05 0.13054 0.81986 0.84608 0.0014381 0.91312 0.5246 0.0019358 0.42342 1.5283 1.5259 16.0098 144.9848 0.00027643 -85.3215 0.30321
0.40723 0.98802 5.5231e-05 3.8182 0.012045 5.3667e-06 0.001154 0.083705 0.00065598 0.084356 0.075788 0 0.041783 0.0389 0 0.85441 0.231 0.060234 0.0085176 4.1144 0.05345 6.3813e-05 0.83661 0.0051153 0.005853 0.0014642 0.98593 0.99104 3.1678e-06 1.2671e-05 0.13054 0.82037 0.84641 0.0014378 0.91364 0.52476 0.0019354 0.42343 1.5296 1.5272 16.0098 144.9848 0.00027591 -85.3239 0.30421
0.40823 0.98802 5.5231e-05 3.8182 0.012045 5.3798e-06 0.001154 0.083827 0.00065598 0.084478 0.0759 0 0.041773 0.0389 0 0.85445 0.23102 0.06024 0.0085184 4.1145 0.053455 6.3818e-05 0.83661 0.0051154 0.0058531 0.0014637 0.98594 0.99104 3.1665e-06 1.2666e-05 0.13054 0.82088 0.84673 0.0014375 0.91417 0.52492 0.001935 0.42344 1.5309 1.5285 16.0099 144.9848 0.00027538 -85.3263 0.30521
0.40923 0.98802 5.5231e-05 3.8182 0.012045 5.393e-06 0.001154 0.083948 0.00065599 0.0846 0.076012 0 0.041764 0.0389 0 0.85449 0.23104 0.060247 0.0085192 4.1146 0.053459 6.3824e-05 0.8366 0.0051155 0.0058532 0.0014631 0.98594 0.99105 3.1651e-06 1.2661e-05 0.13054 0.82139 0.84705 0.0014372 0.91469 0.52509 0.0019346 0.42345 1.5322 1.5298 16.0099 144.9848 0.00027486 -85.3287 0.30621
0.41023 0.98802 5.5231e-05 3.8182 0.012045 5.4062e-06 0.001154 0.08407 0.000656 0.084721 0.076124 0 0.041754 0.0389 0 0.85453 0.23106 0.060253 0.00852 4.1146 0.053464 6.383e-05 0.8366 0.0051156 0.0058533 0.0014625 0.98595 0.99105 3.1638e-06 1.2655e-05 0.13054 0.82189 0.84737 0.0014369 0.91521 0.52525 0.0019342 0.42346 1.5334 1.5311 16.0099 144.9849 0.00027434 -85.3311 0.30721
0.41123 0.98802 5.5231e-05 3.8182 0.012045 5.4193e-06 0.001154 0.084191 0.00065601 0.084843 0.076235 0 0.041744 0.0389 0 0.85457 0.23108 0.06026 0.0085208 4.1147 0.053468 6.3835e-05 0.8366 0.0051156 0.0058534 0.0014619 0.98596 0.99106 3.1625e-06 1.265e-05 0.13054 0.8224 0.84769 0.0014366 0.91573 0.52542 0.0019339 0.42347 1.5347 1.5324 16.0099 144.9849 0.00027383 -85.3334 0.30821
0.41223 0.98802 5.5231e-05 3.8182 0.012045 5.4325e-06 0.001154 0.084313 0.00065601 0.084964 0.076347 0 0.041734 0.0389 0 0.85461 0.23109 0.060266 0.0085217 4.1147 0.053473 6.3841e-05 0.83659 0.0051157 0.0058534 0.0014614 0.98597 0.99106 3.1612e-06 1.2645e-05 0.13054 0.8229 0.84801 0.0014363 0.91624 0.52558 0.0019335 0.42348 1.536 1.5336 16.0099 144.9849 0.00027331 -85.3358 0.30921
0.41323 0.98802 5.5231e-05 3.8182 0.012045 5.4457e-06 0.001154 0.084434 0.00065602 0.085085 0.076458 0 0.041725 0.0389 0 0.85465 0.23111 0.060273 0.0085225 4.1148 0.053477 6.3847e-05 0.83659 0.0051158 0.0058535 0.0014608 0.98597 0.99107 3.1599e-06 1.264e-05 0.13055 0.8234 0.84833 0.001436 0.91675 0.52574 0.0019331 0.4235 1.5372 1.5349 16.0099 144.9849 0.0002728 -85.3381 0.31021
0.41423 0.98802 5.5231e-05 3.8182 0.012045 5.4588e-06 0.001154 0.084555 0.00065603 0.085207 0.07657 0 0.041715 0.0389 0 0.85469 0.23113 0.060279 0.0085233 4.1149 0.053482 6.3853e-05 0.83658 0.0051159 0.0058536 0.0014602 0.98598 0.99107 3.1586e-06 1.2634e-05 0.13055 0.8239 0.84864 0.0014357 0.91726 0.52591 0.0019327 0.42351 1.5385 1.5362 16.0099 144.9849 0.00027229 -85.3404 0.31121
0.41523 0.98802 5.5231e-05 3.8182 0.012045 5.472e-06 0.001154 0.084676 0.00065604 0.085328 0.076681 0 0.041705 0.0389 0 0.85474 0.23115 0.060286 0.0085241 4.1149 0.053486 6.3858e-05 0.83658 0.005116 0.0058537 0.0014597 0.98599 0.99108 3.1573e-06 1.2629e-05 0.13055 0.8244 0.84896 0.0014354 0.91776 0.52607 0.0019323 0.42352 1.5398 1.5375 16.0099 144.9849 0.00027179 -85.3427 0.31221
0.41623 0.98802 5.523e-05 3.8182 0.012045 5.4852e-06 0.001154 0.084797 0.00065604 0.085449 0.076792 0 0.041695 0.0389 0 0.85478 0.23117 0.060293 0.008525 4.115 0.053491 6.3864e-05 0.83657 0.0051161 0.0058538 0.0014591 0.986 0.99108 3.156e-06 1.2624e-05 0.13055 0.82489 0.84927 0.0014351 0.91826 0.52623 0.001932 0.42353 1.541 1.5387 16.0099 144.985 0.00027128 -85.3449 0.31321
0.41723 0.98802 5.523e-05 3.8182 0.012044 5.4984e-06 0.001154 0.084918 0.00065605 0.085569 0.076904 0 0.041686 0.0389 0 0.85482 0.23118 0.060299 0.0085258 4.1151 0.053496 6.387e-05 0.83657 0.0051161 0.0058538 0.0014586 0.986 0.99109 3.1548e-06 1.2619e-05 0.13055 0.82538 0.84958 0.0014348 0.91876 0.5264 0.0019316 0.42354 1.5423 1.54 16.01 144.985 0.00027078 -85.3472 0.31421
0.41823 0.98802 5.523e-05 3.8182 0.012044 5.5115e-06 0.001154 0.085039 0.00065606 0.08569 0.077015 0 0.041676 0.0389 0 0.85486 0.2312 0.060306 0.0085266 4.1151 0.0535 6.3876e-05 0.83656 0.0051162 0.0058539 0.001458 0.98601 0.99109 3.1535e-06 1.2614e-05 0.13055 0.82588 0.84989 0.0014346 0.91925 0.52656 0.0019312 0.42355 1.5435 1.5412 16.01 144.985 0.00027028 -85.3494 0.31521
0.41923 0.98802 5.523e-05 3.8182 0.012044 5.5247e-06 0.001154 0.085159 0.00065607 0.085811 0.077126 0 0.041666 0.0389 0 0.8549 0.23122 0.060312 0.0085275 4.1152 0.053505 6.3882e-05 0.83656 0.0051163 0.005854 0.0014575 0.98602 0.9911 3.1523e-06 1.2609e-05 0.13055 0.82637 0.8502 0.0014343 0.91974 0.52672 0.0019309 0.42357 1.5448 1.5425 16.01 144.985 0.00026978 -85.3516 0.31621
0.42023 0.98802 5.523e-05 3.8182 0.012044 5.5379e-06 0.001154 0.08528 0.00065607 0.085932 0.077237 0 0.041656 0.0389 0 0.85494 0.23124 0.060319 0.0085283 4.1153 0.053509 6.3888e-05 0.83655 0.0051164 0.0058541 0.001457 0.98602 0.9911 3.1511e-06 1.2604e-05 0.13055 0.82686 0.85051 0.001434 0.92023 0.52689 0.0019305 0.42358 1.546 1.5437 16.01 144.985 0.00026929 -85.3538 0.31721
0.42123 0.98802 5.523e-05 3.8182 0.012044 5.551e-06 0.001154 0.085401 0.00065608 0.086052 0.077347 0 0.041647 0.0389 0 0.85499 0.23126 0.060326 0.0085291 4.1154 0.053514 6.3893e-05 0.83655 0.0051165 0.0058542 0.0014564 0.98603 0.99111 3.1498e-06 1.2599e-05 0.13055 0.82735 0.85082 0.0014337 0.92072 0.52705 0.0019301 0.42359 1.5472 1.545 16.01 144.9851 0.00026879 -85.356 0.31821
0.42223 0.98802 5.523e-05 3.8182 0.012044 5.5642e-06 0.001154 0.085521 0.00065609 0.086172 0.077458 0 0.041637 0.0389 0 0.85503 0.23128 0.060332 0.00853 4.1154 0.053519 6.3899e-05 0.83655 0.0051166 0.0058543 0.0014559 0.98604 0.99111 3.1486e-06 1.2595e-05 0.13055 0.82783 0.85112 0.0014335 0.9212 0.52721 0.0019298 0.4236 1.5485 1.5462 16.01 144.9851 0.0002683 -85.3582 0.31921
0.42323 0.98802 5.523e-05 3.8182 0.012044 5.5774e-06 0.001154 0.085641 0.0006561 0.086293 0.077569 0 0.041628 0.0389 0 0.85507 0.2313 0.060339 0.0085308 4.1155 0.053523 6.3905e-05 0.83654 0.0051166 0.0058544 0.0014554 0.98604 0.99112 3.1474e-06 1.259e-05 0.13055 0.82832 0.85142 0.0014332 0.92168 0.52737 0.0019294 0.42361 1.5497 1.5475 16.01 144.9851 0.00026781 -85.3604 0.32021
0.42423 0.98802 5.523e-05 3.8182 0.012044 5.5905e-06 0.001154 0.085761 0.0006561 0.086413 0.077679 0 0.041618 0.0389 0 0.85511 0.23131 0.060346 0.0085317 4.1156 0.053528 6.3911e-05 0.83654 0.0051167 0.0058544 0.0014548 0.98605 0.99112 3.1462e-06 1.2585e-05 0.13055 0.8288 0.85173 0.0014329 0.92215 0.52754 0.0019291 0.42362 1.5509 1.5487 16.01 144.9851 0.00026733 -85.3625 0.32121
0.42523 0.98802 5.523e-05 3.8182 0.012044 5.6037e-06 0.001154 0.085882 0.00065611 0.086533 0.07779 0 0.041608 0.0389 0 0.85515 0.23133 0.060352 0.0085325 4.1156 0.053532 6.3917e-05 0.83653 0.0051168 0.0058545 0.0014543 0.98606 0.99113 3.1451e-06 1.258e-05 0.13055 0.82928 0.85203 0.0014326 0.92263 0.5277 0.0019287 0.42364 1.5521 1.5499 16.01 144.9851 0.00026684 -85.3646 0.32221
0.42623 0.98802 5.523e-05 3.8182 0.012044 5.6169e-06 0.001154 0.086002 0.00065612 0.086653 0.0779 0 0.041599 0.0389 0 0.8552 0.23135 0.060359 0.0085333 4.1157 0.053537 6.3923e-05 0.83653 0.0051169 0.0058546 0.0014538 0.98607 0.99113 3.1439e-06 1.2576e-05 0.13055 0.82976 0.85233 0.0014324 0.9231 0.52786 0.0019284 0.42365 1.5534 1.5512 16.01 144.9851 0.00026636 -85.3668 0.32321
0.42723 0.98802 5.523e-05 3.8182 0.012044 5.63e-06 0.001154 0.086121 0.00065612 0.086773 0.078011 0 0.041589 0.0389 0 0.85524 0.23137 0.060366 0.0085342 4.1158 0.053542 6.3929e-05 0.83652 0.005117 0.0058547 0.0014533 0.98607 0.99113 3.1427e-06 1.2571e-05 0.13056 0.83024 0.85262 0.0014321 0.92357 0.52803 0.001928 0.42366 1.5546 1.5524 16.01 144.9852 0.00026588 -85.3689 0.32421
0.42823 0.98802 5.523e-05 3.8182 0.012044 5.6432e-06 0.001154 0.086241 0.00065613 0.086893 0.078121 0 0.041579 0.0389 0 0.85528 0.23139 0.060373 0.008535 4.1158 0.053546 6.3935e-05 0.83652 0.0051171 0.0058548 0.0014528 0.98608 0.99114 3.1416e-06 1.2566e-05 0.13056 0.83072 0.85292 0.0014319 0.92403 0.52819 0.0019277 0.42367 1.5558 1.5536 16.0101 144.9852 0.0002654 -85.3709 0.32521
0.42923 0.98802 5.523e-05 3.8182 0.012044 5.6564e-06 0.001154 0.086361 0.00065614 0.087013 0.078231 0 0.04157 0.0389 0 0.85532 0.23141 0.060379 0.0085359 4.1159 0.053551 6.3941e-05 0.83651 0.0051172 0.0058549 0.0014523 0.98609 0.99114 3.1404e-06 1.2562e-05 0.13056 0.8312 0.85322 0.0014316 0.92449 0.52835 0.0019274 0.42368 1.557 1.5548 16.0101 144.9852 0.00026492 -85.373 0.32621
0.43023 0.98802 5.523e-05 3.8182 0.012044 5.6695e-06 0.001154 0.086481 0.00065615 0.087132 0.078341 0 0.04156 0.0389 0 0.85537 0.23143 0.060386 0.0085367 4.116 0.053556 6.3947e-05 0.83651 0.0051173 0.005855 0.0014518 0.98609 0.99115 3.1393e-06 1.2557e-05 0.13056 0.83167 0.85351 0.0014313 0.92495 0.52851 0.001927 0.4237 1.5582 1.556 16.0101 144.9852 0.00026445 -85.3751 0.32721
0.43123 0.98802 5.523e-05 3.8182 0.012044 5.6827e-06 0.001154 0.0866 0.00065615 0.087252 0.078451 0 0.041551 0.0389 0 0.85541 0.23145 0.060393 0.0085376 4.116 0.05356 6.3953e-05 0.8365 0.0051174 0.005855 0.0014513 0.9861 0.99115 3.1381e-06 1.2553e-05 0.13056 0.83214 0.85381 0.0014311 0.92541 0.52868 0.0019267 0.42371 1.5594 1.5572 16.0101 144.9852 0.00026398 -85.3771 0.32821
0.43223 0.98802 5.523e-05 3.8182 0.012044 5.6959e-06 0.001154 0.08672 0.00065616 0.087371 0.078561 0 0.041541 0.0389 0 0.85545 0.23146 0.0604 0.0085384 4.1161 0.053565 6.3959e-05 0.8365 0.0051174 0.0058551 0.0014508 0.9861 0.99116 3.137e-06 1.2548e-05 0.13056 0.83262 0.8541 0.0014308 0.92586 0.52884 0.0019264 0.42372 1.5606 1.5585 16.0101 144.9853 0.00026351 -85.3791 0.32921
0.43323 0.98802 5.5229e-05 3.8182 0.012044 5.7091e-06 0.001154 0.086839 0.00065617 0.087491 0.078671 0 0.041532 0.0389 0 0.85549 0.23148 0.060406 0.0085393 4.1162 0.05357 6.3965e-05 0.83649 0.0051175 0.0058552 0.0014503 0.98611 0.99116 3.1359e-06 1.2544e-05 0.13056 0.83309 0.85439 0.0014306 0.92632 0.529 0.001926 0.42373 1.5618 1.5597 16.0101 144.9853 0.00026304 -85.3811 0.33021
0.43423 0.98802 5.5229e-05 3.8182 0.012044 5.7222e-06 0.001154 0.086958 0.00065617 0.08761 0.07878 0 0.041522 0.0389 0 0.85554 0.2315 0.060413 0.0085402 4.1163 0.053575 6.3971e-05 0.83649 0.0051176 0.0058553 0.0014499 0.98612 0.99116 3.1348e-06 1.2539e-05 0.13056 0.83355 0.85468 0.0014303 0.92676 0.52916 0.0019257 0.42374 1.563 1.5609 16.0101 144.9853 0.00026257 -85.3831 0.33121
0.43523 0.98802 5.5229e-05 3.8182 0.012044 5.7354e-06 0.001154 0.087077 0.00065618 0.087729 0.07889 0 0.041513 0.0389 0 0.85558 0.23152 0.06042 0.008541 4.1163 0.053579 6.3977e-05 0.83648 0.0051177 0.0058554 0.0014494 0.98612 0.99117 3.1337e-06 1.2535e-05 0.13056 0.83402 0.85497 0.0014301 0.92721 0.52933 0.0019254 0.42375 1.5642 1.5621 16.0101 144.9853 0.00026211 -85.3851 0.33221
0.43623 0.98802 5.5229e-05 3.8182 0.012044 5.7486e-06 0.001154 0.087196 0.00065619 0.087848 0.079 0 0.041503 0.0389 0 0.85562 0.23154 0.060427 0.0085419 4.1164 0.053584 6.3983e-05 0.83648 0.0051178 0.0058555 0.0014489 0.98613 0.99117 3.1326e-06 1.253e-05 0.13056 0.83449 0.85525 0.0014298 0.92765 0.52949 0.0019251 0.42377 1.5654 1.5633 16.0101 144.9853 0.00026165 -85.3871 0.33321
0.43723 0.98802 5.5229e-05 3.8182 0.012044 5.7617e-06 0.001154 0.087315 0.00065619 0.087967 0.079109 0 0.041494 0.0389 0 0.85567 0.23156 0.060434 0.0085427 4.1165 0.053589 6.3989e-05 0.83648 0.0051179 0.0058556 0.0014484 0.98614 0.99118 3.1315e-06 1.2526e-05 0.13056 0.83495 0.85554 0.0014296 0.92809 0.52965 0.0019247 0.42378 1.5666 1.5644 16.0101 144.9853 0.00026119 -85.389 0.33421
0.43823 0.98802 5.5229e-05 3.8182 0.012044 5.7749e-06 0.001154 0.087434 0.0006562 0.088086 0.079218 0 0.041484 0.0389 0 0.85571 0.23158 0.060441 0.0085436 4.1166 0.053594 6.3995e-05 0.83647 0.005118 0.0058557 0.001448 0.98614 0.99118 3.1304e-06 1.2522e-05 0.13056 0.83541 0.85582 0.0014293 0.92853 0.52981 0.0019244 0.42379 1.5678 1.5656 16.0101 144.9854 0.00026073 -85.391 0.33521
0.43923 0.98802 5.5229e-05 3.8182 0.012044 5.7881e-06 0.001154 0.087553 0.00065621 0.088205 0.079328 0 0.041475 0.0389 0 0.85575 0.2316 0.060447 0.0085445 4.1166 0.053598 6.4001e-05 0.83647 0.0051181 0.0058558 0.0014475 0.98615 0.99118 3.1294e-06 1.2518e-05 0.13056 0.83588 0.85611 0.0014291 0.92896 0.52998 0.0019241 0.4238 1.5689 1.5668 16.0101 144.9854 0.00026027 -85.3929 0.33621
0.44023 0.98802 5.5229e-05 3.8182 0.012044 5.8012e-06 0.001154 0.087672 0.00065622 0.088323 0.079437 0 0.041465 0.0389 0 0.8558 0.23162 0.060454 0.0085453 4.1167 0.053603 6.4007e-05 0.83646 0.0051182 0.0058558 0.001447 0.98615 0.99119 3.1283e-06 1.2513e-05 0.13057 0.83634 0.85639 0.0014289 0.9294 0.53014 0.0019238 0.42381 1.5701 1.568 16.0101 144.9854 0.00025982 -85.3948 0.33721
0.44123 0.98802 5.5229e-05 3.8182 0.012044 5.8144e-06 0.001154 0.08779 0.00065622 0.088442 0.079546 0 0.041456 0.0389 0 0.85584 0.23163 0.060461 0.0085462 4.1168 0.053608 6.4013e-05 0.83646 0.0051183 0.0058559 0.0014466 0.98616 0.99119 3.1273e-06 1.2509e-05 0.13057 0.83679 0.85667 0.0014286 0.92983 0.5303 0.0019235 0.42383 1.5713 1.5692 16.0101 144.9854 0.00025937 -85.3967 0.33821
0.44223 0.98802 5.5229e-05 3.8182 0.012044 5.8276e-06 0.001154 0.087909 0.00065623 0.08856 0.079655 0 0.041446 0.0389 0 0.85588 0.23165 0.060468 0.008547 4.1168 0.053613 6.4019e-05 0.83645 0.0051184 0.005856 0.0014461 0.98617 0.9912 3.1262e-06 1.2505e-05 0.13057 0.83725 0.85695 0.0014284 0.93025 0.53046 0.0019232 0.42384 1.5725 1.5704 16.0102 144.9854 0.00025892 -85.3986 0.33921
0.44323 0.98802 5.5229e-05 3.8182 0.012044 5.8407e-06 0.001154 0.088027 0.00065624 0.088679 0.079764 0 0.041437 0.0389 0 0.85593 0.23167 0.060475 0.0085479 4.1169 0.053618 6.4025e-05 0.83645 0.0051184 0.0058561 0.0014457 0.98617 0.9912 3.1252e-06 1.2501e-05 0.13057 0.83771 0.85723 0.0014282 0.93068 0.53062 0.0019229 0.42385 1.5736 1.5715 16.0102 144.9855 0.00025847 -85.4005 0.34021
0.44423 0.98802 5.5229e-05 3.8182 0.012044 5.8539e-06 0.001154 0.088145 0.00065624 0.088797 0.079873 0 0.041428 0.0389 0 0.85597 0.23169 0.060482 0.0085488 4.117 0.053623 6.4031e-05 0.83644 0.0051185 0.0058562 0.0014452 0.98618 0.9912 3.1242e-06 1.2497e-05 0.13057 0.83816 0.85751 0.0014279 0.9311 0.53079 0.0019226 0.42386 1.5748 1.5727 16.0102 144.9855 0.00025802 -85.4023 0.34121
0.44523 0.98802 5.5229e-05 3.8182 0.012044 5.8671e-06 0.001154 0.088264 0.00065625 0.088915 0.079982 0 0.041418 0.0389 0 0.85601 0.23171 0.060489 0.0085497 4.1171 0.053627 6.4038e-05 0.83644 0.0051186 0.0058563 0.0014448 0.98618 0.99121 3.1231e-06 1.2493e-05 0.13057 0.83861 0.85778 0.0014277 0.93152 0.53095 0.0019223 0.42388 1.5759 1.5739 16.0102 144.9855 0.00025758 -85.4042 0.34221
0.44623 0.98802 5.5229e-05 3.8182 0.012044 5.8802e-06 0.001154 0.088382 0.00065626 0.089033 0.080091 0 0.041409 0.0389 0 0.85606 0.23173 0.060496 0.0085505 4.1171 0.053632 6.4044e-05 0.83643 0.0051187 0.0058564 0.0014443 0.98619 0.99121 3.1221e-06 1.2489e-05 0.13057 0.83907 0.85806 0.0014275 0.93193 0.53111 0.001922 0.42389 1.5771 1.575 16.0102 144.9855 0.00025714 -85.406 0.34321
0.44723 0.98802 5.5229e-05 3.8182 0.012044 5.8934e-06 0.001154 0.0885 0.00065626 0.089151 0.080199 0 0.041399 0.0389 0 0.8561 0.23175 0.060503 0.0085514 4.1172 0.053637 6.405e-05 0.83643 0.0051188 0.0058565 0.0014439 0.9862 0.99122 3.1211e-06 1.2484e-05 0.13057 0.83952 0.85833 0.0014272 0.93235 0.53127 0.0019217 0.4239 1.5783 1.5762 16.0102 144.9855 0.0002567 -85.4078 0.34421
0.44823 0.98802 5.5229e-05 3.8182 0.012044 5.9066e-06 0.001154 0.088618 0.00065627 0.089269 0.080308 0 0.04139 0.0389 0 0.85615 0.23177 0.06051 0.0085523 4.1173 0.053642 6.4056e-05 0.83642 0.0051189 0.0058566 0.0014435 0.9862 0.99122 3.1201e-06 1.2481e-05 0.13057 0.83997 0.85861 0.001427 0.93276 0.53143 0.0019214 0.42391 1.5794 1.5773 16.0102 144.9855 0.00025626 -85.4096 0.34521
0.44923 0.98802 5.5228e-05 3.8182 0.012044 5.9197e-06 0.001154 0.088735 0.00065628 0.089387 0.080416 0 0.041381 0.0389 0 0.85619 0.23179 0.060517 0.0085532 4.1174 0.053647 6.4062e-05 0.83642 0.005119 0.0058567 0.001443 0.98621 0.99122 3.1191e-06 1.2477e-05 0.13057 0.84041 0.85888 0.0014268 0.93317 0.5316 0.0019211 0.42392 1.5806 1.5785 16.0102 144.9856 0.00025582 -85.4114 0.34621
0.45023 0.98802 5.5228e-05 3.8182 0.012044 5.9329e-06 0.001154 0.088853 0.00065628 0.089505 0.080525 0 0.041371 0.0389 0 0.85623 0.23181 0.060524 0.008554 4.1175 0.053652 6.4068e-05 0.83641 0.0051191 0.0058568 0.0014426 0.98621 0.99123 3.1182e-06 1.2473e-05 0.13057 0.84086 0.85915 0.0014266 0.93357 0.53176 0.0019208 0.42394 1.5817 1.5797 16.0102 144.9856 0.00025539 -85.4132 0.34721
0.45123 0.98802 5.5228e-05 3.8182 0.012044 5.9461e-06 0.001154 0.088971 0.00065629 0.089622 0.080633 0 0.041362 0.0389 0 0.85628 0.23183 0.060531 0.0085549 4.1175 0.053657 6.4075e-05 0.83641 0.0051192 0.0058569 0.0014422 0.98622 0.99123 3.1172e-06 1.2469e-05 0.13057 0.8413 0.85942 0.0014264 0.93398 0.53192 0.0019205 0.42395 1.5828 1.5808 16.0102 144.9856 0.00025495 -85.415 0.34821
0.45223 0.98802 5.5228e-05 3.8182 0.012044 5.9592e-06 0.001154 0.089088 0.0006563 0.08974 0.080741 0 0.041353 0.0389 0 0.85632 0.23185 0.060538 0.0085558 4.1176 0.053662 6.4081e-05 0.8364 0.0051193 0.005857 0.0014418 0.98622 0.99123 3.1162e-06 1.2465e-05 0.13057 0.84175 0.85969 0.0014261 0.93438 0.53208 0.0019202 0.42396 1.584 1.5819 16.0102 144.9856 0.00025452 -85.4167 0.34921
0.45323 0.98802 5.5228e-05 3.8182 0.012044 5.9724e-06 0.001154 0.089206 0.0006563 0.089857 0.080849 0 0.041344 0.0389 0 0.85637 0.23187 0.060545 0.0085567 4.1177 0.053666 6.4087e-05 0.8364 0.0051194 0.005857 0.0014413 0.98623 0.99124 3.1152e-06 1.2461e-05 0.13058 0.84219 0.85996 0.0014259 0.93478 0.53224 0.0019199 0.42397 1.5851 1.5831 16.0102 144.9856 0.00025409 -85.4185 0.35021
0.45423 0.98802 5.5228e-05 3.8182 0.012044 5.9856e-06 0.001154 0.089323 0.00065631 0.089975 0.080957 0 0.041334 0.0389 0 0.85641 0.23189 0.060552 0.0085576 4.1178 0.053671 6.4093e-05 0.83639 0.0051195 0.0058571 0.0014409 0.98623 0.99124 3.1143e-06 1.2457e-05 0.13058 0.84263 0.86022 0.0014257 0.93517 0.53241 0.0019196 0.42398 1.5862 1.5842 16.0102 144.9857 0.00025367 -85.4202 0.35121
0.45523 0.98802 5.5228e-05 3.8182 0.012044 5.9987e-06 0.001154 0.08944 0.00065632 0.090092 0.081065 0 0.041325 0.0389 0 0.85645 0.23191 0.060559 0.0085584 4.1178 0.053676 6.41e-05 0.83639 0.0051196 0.0058572 0.0014405 0.98624 0.99125 3.1133e-06 1.2453e-05 0.13058 0.84307 0.86049 0.0014255 0.93557 0.53257 0.0019194 0.424 1.5874 1.5854 16.0102 144.9857 0.00025324 -85.4219 0.35221
0.45623 0.98802 5.5228e-05 3.8182 0.012044 6.0119e-06 0.001154 0.089557 0.00065632 0.090209 0.081173 0 0.041316 0.0389 0 0.8565 0.23193 0.060566 0.0085593 4.1179 0.053681 6.4106e-05 0.83638 0.0051197 0.0058573 0.0014401 0.98625 0.99125 3.1124e-06 1.245e-05 0.13058 0.84351 0.86075 0.0014253 0.93596 0.53273 0.0019191 0.42401 1.5885 1.5865 16.0102 144.9857 0.00025282 -85.4236 0.35321
0.45723 0.98802 5.5228e-05 3.8182 0.012044 6.0251e-06 0.001154 0.089675 0.00065633 0.090326 0.081281 0 0.041306 0.0389 0 0.85654 0.23194 0.060573 0.0085602 4.118 0.053686 6.4112e-05 0.83638 0.0051198 0.0058574 0.0014397 0.98625 0.99125 3.1115e-06 1.2446e-05 0.13058 0.84394 0.86101 0.0014251 0.93635 0.53289 0.0019188 0.42402 1.5896 1.5876 16.0102 144.9857 0.0002524 -85.4253 0.35421
0.45823 0.98802 5.5228e-05 3.8182 0.012044 6.0382e-06 0.001154 0.089792 0.00065633 0.090443 0.081389 0 0.041297 0.0389 0 0.85659 0.23196 0.06058 0.0085611 4.1181 0.053691 6.4119e-05 0.83637 0.0051199 0.0058575 0.0014393 0.98626 0.99126 3.1105e-06 1.2442e-05 0.13058 0.84438 0.86128 0.0014248 0.93673 0.53305 0.0019185 0.42403 1.5907 1.5887 16.0102 144.9857 0.00025198 -85.427 0.35521
0.45923 0.98802 5.5228e-05 3.8182 0.012044 6.0514e-06 0.001154 0.089908 0.00065634 0.09056 0.081496 0 0.041288 0.0389 0 0.85663 0.23198 0.060587 0.008562 4.1182 0.053696 6.4125e-05 0.83637 0.00512 0.0058576 0.0014389 0.98626 0.99126 3.1096e-06 1.2439e-05 0.13058 0.84481 0.86154 0.0014246 0.93712 0.53321 0.0019183 0.42405 1.5918 1.5899 16.0102 144.9858 0.00025156 -85.4287 0.35621
0.46023 0.98802 5.5228e-05 3.8182 0.012044 6.0646e-06 0.001154 0.090025 0.00065635 0.090677 0.081604 0 0.041279 0.0389 0 0.85668 0.232 0.060594 0.0085629 4.1182 0.053701 6.4131e-05 0.83636 0.0051201 0.0058577 0.0014385 0.98627 0.99126 3.1087e-06 1.2435e-05 0.13058 0.84524 0.8618 0.0014244 0.9375 0.53337 0.001918 0.42406 1.593 1.591 16.0102 144.9858 0.00025114 -85.4303 0.35721
0.46123 0.98802 5.5228e-05 3.8182 0.012044 6.0778e-06 0.001154 0.090142 0.00065635 0.090794 0.081711 0 0.04127 0.0389 0 0.85672 0.23202 0.060601 0.0085638 4.1183 0.053706 6.4138e-05 0.83636 0.0051202 0.0058578 0.0014381 0.98627 0.99127 3.1078e-06 1.2431e-05 0.13058 0.84567 0.86206 0.0014242 0.93788 0.53353 0.0019177 0.42407 1.5941 1.5921 16.0102 144.9858 0.00025073 -85.432 0.35821
0.46223 0.98802 5.5228e-05 3.8182 0.012044 6.0909e-06 0.001154 0.090258 0.00065636 0.09091 0.081819 0 0.04126 0.0389 0 0.85677 0.23204 0.060608 0.0085647 4.1184 0.053711 6.4144e-05 0.83635 0.0051203 0.0058579 0.0014377 0.98628 0.99127 3.1069e-06 1.2428e-05 0.13058 0.8461 0.86231 0.001424 0.93826 0.5337 0.0019175 0.42408 1.5952 1.5932 16.0102 144.9858 0.00025031 -85.4336 0.35921
0.46323 0.98802 5.5228e-05 3.8182 0.012044 6.1041e-06 0.001154 0.090375 0.00065637 0.091027 0.081926 0 0.041251 0.0389 0 0.85681 0.23206 0.060616 0.0085656 4.1185 0.053716 6.415e-05 0.83635 0.0051204 0.005858 0.0014373 0.98628 0.99127 3.106e-06 1.2424e-05 0.13058 0.84653 0.86257 0.0014238 0.93863 0.53386 0.0019172 0.4241 1.5963 1.5943 16.0102 144.9858 0.0002499 -85.4352 0.36021
0.46423 0.98802 5.5228e-05 3.8182 0.012044 6.1173e-06 0.001154 0.090491 0.00065637 0.091143 0.082033 0 0.041242 0.0389 0 0.85686 0.23208 0.060623 0.0085665 4.1186 0.053721 6.4157e-05 0.83634 0.0051205 0.0058581 0.0014369 0.98629 0.99128 3.1051e-06 1.2421e-05 0.13058 0.84696 0.86283 0.0014236 0.939 0.53402 0.0019169 0.42411 1.5974 1.5954 16.0102 144.9858 0.00024949 -85.4368 0.36121
0.46523 0.98802 5.5227e-05 3.8182 0.012044 6.1304e-06 0.001154 0.090608 0.00065638 0.091259 0.08214 0 0.041233 0.0389 0 0.8569 0.2321 0.06063 0.0085674 4.1186 0.053726 6.4163e-05 0.83634 0.0051206 0.0058582 0.0014365 0.98629 0.99128 3.1042e-06 1.2417e-05 0.13059 0.84738 0.86308 0.0014234 0.93938 0.53418 0.0019167 0.42412 1.5985 1.5965 16.0102 144.9859 0.00024909 -85.4384 0.36221
0.46623 0.98802 5.5227e-05 3.8182 0.012044 6.1436e-06 0.001154 0.090724 0.00065638 0.091376 0.082248 0 0.041224 0.0389 0 0.85695 0.23212 0.060637 0.0085683 4.1187 0.053731 6.417e-05 0.83633 0.0051207 0.0058583 0.0014362 0.9863 0.99128 3.1034e-06 1.2414e-05 0.13059 0.84781 0.86333 0.0014232 0.93974 0.53434 0.0019164 0.42413 1.5996 1.5976 16.0102 144.9859 0.00024868 -85.44 0.36321
0.46723 0.98802 5.5227e-05 3.8182 0.012044 6.1568e-06 0.001154 0.09084 0.00065639 0.091492 0.082355 0 0.041214 0.0389 0 0.85699 0.23214 0.060644 0.0085692 4.1188 0.053736 6.4176e-05 0.83633 0.0051208 0.0058584 0.0014358 0.9863 0.99129 3.1025e-06 1.241e-05 0.13059 0.84823 0.86359 0.001423 0.94011 0.5345 0.0019162 0.42414 1.6007 1.5987 16.0102 144.9859 0.00024828 -85.4416 0.36421
0.46823 0.98802 5.5227e-05 3.8182 0.012044 6.1699e-06 0.001154 0.090956 0.0006564 0.091608 0.082461 0 0.041205 0.0389 0 0.85704 0.23216 0.060651 0.0085701 4.1189 0.053741 6.4182e-05 0.83632 0.0051209 0.0058585 0.0014354 0.98631 0.99129 3.1016e-06 1.2407e-05 0.13059 0.84865 0.86384 0.0014228 0.94047 0.53466 0.0019159 0.42416 1.6018 1.5998 16.0103 144.9859 0.00024787 -85.4432 0.36521
0.46923 0.98802 5.5227e-05 3.8182 0.012044 6.1831e-06 0.001154 0.091072 0.0006564 0.091724 0.082568 0 0.041196 0.0389 0 0.85708 0.23218 0.060659 0.008571 4.119 0.053746 6.4189e-05 0.83632 0.005121 0.0058586 0.001435 0.98631 0.99129 3.1008e-06 1.2403e-05 0.13059 0.84907 0.86409 0.0014226 0.94083 0.53482 0.0019156 0.42417 1.6028 1.6009 16.0103 144.9859 0.00024747 -85.4447 0.36621
0.47023 0.98802 5.5227e-05 3.8182 0.012044 6.1963e-06 0.001154 0.091188 0.00065641 0.09184 0.082675 0 0.041187 0.0389 0 0.85713 0.2322 0.060666 0.0085719 4.119 0.053752 6.4195e-05 0.83631 0.0051211 0.0058587 0.0014347 0.98632 0.9913 3.0999e-06 1.24e-05 0.13059 0.84949 0.86434 0.0014224 0.94119 0.53498 0.0019154 0.42418 1.6039 1.602 16.0103 144.986 0.00024707 -85.4463 0.36721
0.47123 0.98802 5.5227e-05 3.8182 0.012044 6.2094e-06 0.001154 0.091304 0.00065642 0.091955 0.082782 0 0.041178 0.0389 0 0.85717 0.23222 0.060673 0.0085728 4.1191 0.053757 6.4202e-05 0.83631 0.0051212 0.0058588 0.0014343 0.98632 0.9913 3.0991e-06 1.2396e-05 0.13059 0.84991 0.86458 0.0014223 0.94155 0.53514 0.0019151 0.42419 1.605 1.6031 16.0103 144.986 0.00024668 -85.4478 0.36821
0.47223 0.98802 5.5227e-05 3.8182 0.012044 6.2226e-06 0.001154 0.091419 0.00065642 0.092071 0.082888 0 0.041169 0.0389 0 0.85722 0.23224 0.06068 0.0085737 4.1192 0.053762 6.4208e-05 0.8363 0.0051213 0.0058589 0.0014339 0.98633 0.9913 3.0983e-06 1.2393e-05 0.13059 0.85033 0.86483 0.0014221 0.9419 0.53531 0.0019149 0.42421 1.6061 1.6042 16.0103 144.986 0.00024628 -85.4493 0.36921
0.47323 0.98802 5.5227e-05 3.8182 0.012044 6.2358e-06 0.001154 0.091535 0.00065643 0.092187 0.082995 0 0.04116 0.0389 0 0.85726 0.23226 0.060687 0.0085746 4.1193 0.053767 6.4215e-05 0.8363 0.0051214 0.005859 0.0014336 0.98633 0.9913 3.0974e-06 1.239e-05 0.13059 0.85074 0.86508 0.0014219 0.94226 0.53547 0.0019146 0.42422 1.6072 1.6053 16.0103 144.986 0.00024589 -85.4509 0.37021
0.47423 0.98802 5.5227e-05 3.8182 0.012044 6.2489e-06 0.001154 0.09165 0.00065643 0.092302 0.083101 0 0.041151 0.0389 0 0.85731 0.23228 0.060695 0.0085755 4.1194 0.053772 6.4221e-05 0.83629 0.0051215 0.0058591 0.0014332 0.98634 0.99131 3.0966e-06 1.2386e-05 0.13059 0.85116 0.86532 0.0014217 0.94261 0.53563 0.0019144 0.42423 1.6082 1.6063 16.0103 144.986 0.0002455 -85.4524 0.37121
0.47523 0.98802 5.5227e-05 3.8182 0.012044 6.2621e-06 0.001154 0.091766 0.00065644 0.092418 0.083207 0 0.041142 0.0389 0 0.85736 0.2323 0.060702 0.0085764 4.1195 0.053777 6.4228e-05 0.83629 0.0051216 0.0058592 0.0014329 0.98634 0.99131 3.0958e-06 1.2383e-05 0.13059 0.85157 0.86557 0.0014215 0.94295 0.53579 0.0019142 0.42424 1.6093 1.6074 16.0103 144.9861 0.0002451 -85.4539 0.37221
0.47623 0.98802 5.5227e-05 3.8182 0.012044 6.2753e-06 0.001154 0.091881 0.00065645 0.092533 0.083314 0 0.041133 0.0389 0 0.8574 0.23232 0.060709 0.0085773 4.1195 0.053782 6.4234e-05 0.83628 0.0051217 0.0058593 0.0014325 0.98634 0.99131 3.095e-06 1.238e-05 0.13059 0.85198 0.86581 0.0014213 0.9433 0.53595 0.0019139 0.42426 1.6104 1.6085 16.0103 144.9861 0.00024472 -85.4553 0.37321
0.47723 0.98802 5.5227e-05 3.8182 0.012044 6.2884e-06 0.001154 0.091996 0.00065645 0.092648 0.08342 0 0.041124 0.0389 0 0.85745 0.23234 0.060717 0.0085783 4.1196 0.053787 6.4241e-05 0.83628 0.0051218 0.0058594 0.0014321 0.98635 0.99132 3.0942e-06 1.2377e-05 0.1306 0.85239 0.86605 0.0014211 0.94364 0.53611 0.0019137 0.42427 1.6114 1.6096 16.0103 144.9861 0.00024433 -85.4568 0.37421
0.47823 0.98802 5.5227e-05 3.8182 0.012044 6.3016e-06 0.001154 0.092111 0.00065646 0.092763 0.083526 0 0.041115 0.0389 0 0.85749 0.23236 0.060724 0.0085792 4.1197 0.053793 6.4247e-05 0.83627 0.0051219 0.0058595 0.0014318 0.98635 0.99132 3.0934e-06 1.2374e-05 0.1306 0.8528 0.86629 0.001421 0.94398 0.53627 0.0019134 0.42428 1.6125 1.6106 16.0103 144.9861 0.00024394 -85.4583 0.37521
0.47923 0.98802 5.5227e-05 3.8182 0.012044 6.3148e-06 0.001154 0.092226 0.00065646 0.092878 0.083632 0 0.041106 0.0389 0 0.85754 0.23238 0.060731 0.0085801 4.1198 0.053798 6.4254e-05 0.83627 0.005122 0.0058596 0.0014315 0.98636 0.99132 3.0926e-06 1.237e-05 0.1306 0.85321 0.86653 0.0014208 0.94432 0.53643 0.0019132 0.42429 1.6135 1.6117 16.0103 144.9861 0.00024356 -85.4597 0.37621
0.48023 0.98802 5.5227e-05 3.8182 0.012044 6.3279e-06 0.001154 0.092341 0.00065647 0.092993 0.083738 0 0.041097 0.0389 0 0.85759 0.2324 0.060738 0.008581 4.1199 0.053803 6.4261e-05 0.83626 0.0051221 0.0058597 0.0014311 0.98636 0.99133 3.0918e-06 1.2367e-05 0.1306 0.85361 0.86677 0.0014206 0.94466 0.53659 0.001913 0.42431 1.6146 1.6128 16.0103 144.9861 0.00024318 -85.4612 0.37721
0.48123 0.98802 5.5226e-05 3.8182 0.012044 6.3411e-06 0.001154 0.092456 0.00065648 0.093108 0.083844 0 0.041088 0.0389 0 0.85763 0.23242 0.060746 0.0085819 4.12 0.053808 6.4267e-05 0.83626 0.0051222 0.0058598 0.0014308 0.98637 0.99133 3.091e-06 1.2364e-05 0.1306 0.85402 0.86701 0.0014204 0.945 0.53675 0.0019127 0.42432 1.6157 1.6138 16.0103 144.9862 0.0002428 -85.4626 0.37821
0.48223 0.98802 5.5226e-05 3.8182 0.012044 6.3543e-06 0.001154 0.092571 0.00065648 0.093223 0.083949 0 0.041079 0.0389 0 0.85768 0.23244 0.060753 0.0085829 4.1201 0.053813 6.4274e-05 0.83625 0.0051224 0.00586 0.0014304 0.98637 0.99133 3.0902e-06 1.2361e-05 0.1306 0.85442 0.86725 0.0014202 0.94533 0.53691 0.0019125 0.42433 1.6167 1.6149 16.0103 144.9862 0.00024242 -85.464 0.37921
0.48323 0.98802 5.5226e-05 3.8182 0.012044 6.3674e-06 0.001154 0.092685 0.00065649 0.093337 0.084055 0 0.04107 0.0389 0 0.85772 0.23247 0.06076 0.0085838 4.1201 0.053818 6.428e-05 0.83625 0.0051225 0.0058601 0.0014301 0.98638 0.99133 3.0895e-06 1.2358e-05 0.1306 0.85482 0.86749 0.0014201 0.94566 0.53707 0.0019123 0.42434 1.6177 1.6159 16.0103 144.9862 0.00024204 -85.4654 0.38021
0.48423 0.98802 5.5226e-05 3.8182 0.012044 6.3806e-06 0.001154 0.0928 0.00065649 0.093452 0.084161 0 0.041061 0.0389 0 0.85777 0.23249 0.060768 0.0085847 4.1202 0.053824 6.4287e-05 0.83624 0.0051226 0.0058602 0.0014298 0.98638 0.99134 3.0887e-06 1.2355e-05 0.1306 0.85523 0.86772 0.0014199 0.94599 0.53723 0.0019121 0.42436 1.6188 1.617 16.0103 144.9862 0.00024166 -85.4668 0.38121
0.48523 0.98802 5.5226e-05 3.8182 0.012044 6.3937e-06 0.001154 0.092914 0.0006565 0.093566 0.084266 0 0.041052 0.0389 0 0.85782 0.23251 0.060775 0.0085856 4.1203 0.053829 6.4294e-05 0.83624 0.0051227 0.0058603 0.0014294 0.98638 0.99134 3.0879e-06 1.2352e-05 0.1306 0.85563 0.86796 0.0014197 0.94631 0.53739 0.0019118 0.42437 1.6198 1.618 16.0103 144.9862 0.00024129 -85.4682 0.38221
0.48623 0.98802 5.5226e-05 3.8182 0.012044 6.4069e-06 0.001154 0.093029 0.0006565 0.093681 0.084372 0 0.041043 0.0389 0 0.85786 0.23253 0.060783 0.0085866 4.1204 0.053834 6.43e-05 0.83623 0.0051228 0.0058604 0.0014291 0.98639 0.99134 3.0872e-06 1.2349e-05 0.1306 0.85603 0.86819 0.0014195 0.94664 0.53755 0.0019116 0.42438 1.6209 1.6191 16.0103 144.9863 0.00024092 -85.4696 0.38321
0.48723 0.98802 5.5226e-05 3.8182 0.012044 6.4201e-06 0.001154 0.093143 0.00065651 0.093795 0.084477 0 0.041034 0.0389 0 0.85791 0.23255 0.06079 0.0085875 4.1205 0.053839 6.4307e-05 0.83622 0.0051229 0.0058605 0.0014288 0.98639 0.99135 3.0864e-06 1.2346e-05 0.1306 0.85642 0.86842 0.0014194 0.94696 0.53771 0.0019114 0.4244 1.6219 1.6201 16.0103 144.9863 0.00024054 -85.471 0.38421
0.48823 0.98802 5.5226e-05 3.8182 0.012044 6.4332e-06 0.001154 0.093257 0.00065652 0.093909 0.084582 0 0.041025 0.0389 0 0.85796 0.23257 0.060797 0.0085884 4.1206 0.053845 6.4314e-05 0.83622 0.005123 0.0058606 0.0014284 0.9864 0.99135 3.0857e-06 1.2343e-05 0.13061 0.85682 0.86865 0.0014192 0.94728 0.53787 0.0019112 0.42441 1.6229 1.6211 16.0103 144.9863 0.00024017 -85.4723 0.38521
0.48923 0.98802 5.5226e-05 3.8182 0.012044 6.4464e-06 0.001154 0.093371 0.00065652 0.094023 0.084688 0 0.041016 0.0389 0 0.858 0.23259 0.060805 0.0085893 4.1207 0.05385 6.432e-05 0.83621 0.0051231 0.0058607 0.0014281 0.9864 0.99135 3.085e-06 1.234e-05 0.13061 0.85721 0.86888 0.001419 0.9476 0.53803 0.0019109 0.42442 1.624 1.6222 16.0103 144.9863 0.00023981 -85.4737 0.38621
0.49023 0.98802 5.5226e-05 3.8182 0.012044 6.4596e-06 0.001154 0.093485 0.00065653 0.094137 0.084793 0 0.041007 0.0389 0 0.85805 0.23261 0.060812 0.0085903 4.1208 0.053855 6.4327e-05 0.83621 0.0051232 0.0058608 0.0014278 0.98641 0.99135 3.0842e-06 1.2337e-05 0.13061 0.85761 0.86911 0.0014189 0.94792 0.53819 0.0019107 0.42443 1.625 1.6232 16.0103 144.9863 0.00023944 -85.475 0.38721
0.49123 0.98802 5.5226e-05 3.8182 0.012044 6.4727e-06 0.001154 0.093599 0.00065653 0.094251 0.084898 0 0.040998 0.0389 0 0.8581 0.23263 0.06082 0.0085912 4.1208 0.05386 6.4334e-05 0.8362 0.0051233 0.0058609 0.0014275 0.98641 0.99136 3.0835e-06 1.2334e-05 0.13061 0.858 0.86934 0.0014187 0.94823 0.53835 0.0019105 0.42445 1.626 1.6242 16.0103 144.9864 0.00023907 -85.4764 0.38821
0.49223 0.98802 5.5226e-05 3.8182 0.012043 6.4859e-06 0.001154 0.093713 0.00065654 0.094365 0.085003 0 0.040989 0.0389 0 0.85814 0.23265 0.060827 0.0085922 4.1209 0.053866 6.434e-05 0.8362 0.0051234 0.005861 0.0014272 0.98641 0.99136 3.0828e-06 1.2331e-05 0.13061 0.85839 0.86957 0.0014185 0.94855 0.53851 0.0019103 0.42446 1.627 1.6253 16.0102 144.9864 0.00023871 -85.4777 0.38921
0.49323 0.98802 5.5226e-05 3.8182 0.012043 6.4991e-06 0.001154 0.093827 0.00065655 0.094479 0.085108 0 0.040981 0.0389 0 0.85819 0.23267 0.060835 0.0085931 4.121 0.053871 6.4347e-05 0.83619 0.0051235 0.0058611 0.0014269 0.98642 0.99136 3.0821e-06 1.2328e-05 0.13061 0.85878 0.8698 0.0014184 0.94886 0.53867 0.0019101 0.42447 1.628 1.6263 16.0102 144.9864 0.00023835 -85.479 0.39021
0.49423 0.98802 5.5226e-05 3.8182 0.012043 6.5122e-06 0.001154 0.093941 0.00065655 0.094593 0.085212 0 0.040972 0.0389 0 0.85824 0.23269 0.060842 0.008594 4.1211 0.053876 6.4354e-05 0.83619 0.0051237 0.0058612 0.0014265 0.98642 0.99136 3.0813e-06 1.2325e-05 0.13061 0.85917 0.87002 0.0014182 0.94917 0.53883 0.0019099 0.42448 1.6291 1.6273 16.0102 144.9864 0.00023799 -85.4803 0.39121
0.49523 0.98802 5.5226e-05 3.8182 0.012043 6.5254e-06 0.001154 0.094054 0.00065656 0.094706 0.085317 0 0.040963 0.0389 0 0.85828 0.23271 0.06085 0.008595 4.1212 0.053882 6.4361e-05 0.83618 0.0051238 0.0058614 0.0014262 0.98643 0.99137 3.0806e-06 1.2322e-05 0.13061 0.85956 0.87025 0.0014181 0.94947 0.53899 0.0019097 0.4245 1.6301 1.6283 16.0102 144.9864 0.00023763 -85.4816 0.39221
0.49623 0.98802 5.5226e-05 3.8182 0.012043 6.5386e-06 0.001154 0.094168 0.00065656 0.09482 0.085422 0 0.040954 0.0389 0 0.85833 0.23273 0.060857 0.0085959 4.1213 0.053887 6.4367e-05 0.83618 0.0051239 0.0058615 0.0014259 0.98643 0.99137 3.0799e-06 1.232e-05 0.13061 0.85995 0.87047 0.0014179 0.94978 0.53915 0.0019094 0.42451 1.6311 1.6293 16.0102 144.9865 0.00023727 -85.4829 0.39321
0.49723 0.98802 5.5225e-05 3.8182 0.012043 6.5517e-06 0.001154 0.094281 0.00065657 0.094933 0.085526 0 0.040945 0.0389 0 0.85838 0.23275 0.060865 0.0085968 4.1214 0.053892 6.4374e-05 0.83617 0.005124 0.0058616 0.0014256 0.98643 0.99137 3.0792e-06 1.2317e-05 0.13061 0.86033 0.8707 0.0014177 0.95008 0.53931 0.0019092 0.42452 1.6321 1.6303 16.0102 144.9865 0.00023692 -85.4842 0.39421
0.49823 0.98802 5.5225e-05 3.8182 0.012043 6.5649e-06 0.001154 0.094394 0.00065657 0.095046 0.085631 0 0.040936 0.0389 0 0.85843 0.23277 0.060872 0.0085978 4.1215 0.053898 6.4381e-05 0.83617 0.0051241 0.0058617 0.0014253 0.98644 0.99138 3.0785e-06 1.2314e-05 0.13061 0.86071 0.87092 0.0014176 0.95038 0.53947 0.001909 0.42453 1.6331 1.6314 16.0102 144.9865 0.00023656 -85.4854 0.39521
0.49923 0.98802 5.5225e-05 3.8182 0.012043 6.5781e-06 0.001154 0.094507 0.00065658 0.095159 0.085735 0 0.040928 0.0389 0 0.85847 0.2328 0.06088 0.0085987 4.1216 0.053903 6.4388e-05 0.83616 0.0051242 0.0058618 0.001425 0.98644 0.99138 3.0779e-06 1.2311e-05 0.13062 0.8611 0.87114 0.0014174 0.95068 0.53963 0.0019088 0.42455 1.6341 1.6324 16.0102 144.9865 0.00023621 -85.4867 0.39621
0.50023 0.98802 5.5225e-05 3.8182 0.012043 6.5912e-06 0.001154 0.09462 0.00065658 0.095272 0.085839 0 0.040919 0.0389 0 0.85852 0.23282 0.060887 0.0085997 4.1217 0.053908 6.4395e-05 0.83616 0.0051243 0.0058619 0.0014247 0.98645 0.99138 3.0772e-06 1.2309e-05 0.13062 0.86148 0.87136 0.0014173 0.95098 0.53979 0.0019086 0.42456 1.6351 1.6334 16.0102 144.9865 0.00023586 -85.488 0.39721
0.50123 0.98802 5.5225e-05 3.8182 0.012043 6.6044e-06 0.001154 0.094734 0.00065659 0.095385 0.085944 0 0.04091 0.0389 0 0.85857 0.23284 0.060895 0.0086006 4.1218 0.053914 6.4401e-05 0.83615 0.0051244 0.005862 0.0014244 0.98645 0.99138 3.0765e-06 1.2306e-05 0.13062 0.86186 0.87158 0.0014171 0.95127 0.53995 0.0019084 0.42457 1.6361 1.6344 16.0102 144.9865 0.00023551 -85.4892 0.39821
0.50223 0.98802 5.5225e-05 3.8182 0.012043 6.6176e-06 0.001154 0.094846 0.0006566 0.095498 0.086048 0 0.040901 0.0389 0 0.85862 0.23286 0.060902 0.0086016 4.1218 0.053919 6.4408e-05 0.83615 0.0051246 0.0058621 0.0014241 0.98645 0.99139 3.0758e-06 1.2303e-05 0.13062 0.86224 0.8718 0.001417 0.95157 0.54011 0.0019082 0.42459 1.6371 1.6354 16.0102 144.9866 0.00023516 -85.4904 0.39921
0.50323 0.98802 5.5225e-05 3.8182 0.012043 6.6307e-06 0.001154 0.094959 0.0006566 0.095611 0.086152 0 0.040893 0.0389 0 0.85866 0.23288 0.06091 0.0086025 4.1219 0.053925 6.4415e-05 0.83614 0.0051247 0.0058622 0.0014238 0.98646 0.99139 3.0752e-06 1.2301e-05 0.13062 0.86262 0.87202 0.0014168 0.95186 0.54027 0.001908 0.4246 1.6381 1.6364 16.0102 144.9866 0.00023481 -85.4917 0.40021
0.50423 0.98802 5.5225e-05 3.8182 0.012043 6.6439e-06 0.001154 0.095072 0.00065661 0.095724 0.086256 0 0.040884 0.0389 0 0.85871 0.2329 0.060917 0.0086035 4.122 0.05393 6.4422e-05 0.83613 0.0051248 0.0058624 0.0014236 0.98646 0.99139 3.0745e-06 1.2298e-05 0.13062 0.86299 0.87223 0.0014167 0.95215 0.54042 0.0019078 0.42461 1.6391 1.6374 16.0102 144.9866 0.00023446 -85.4929 0.40121
0.50523 0.98802 5.5225e-05 3.8182 0.012043 6.6571e-06 0.001154 0.095185 0.00065661 0.095837 0.08636 0 0.040875 0.0389 0 0.85876 0.23292 0.060925 0.0086044 4.1221 0.053935 6.4429e-05 0.83613 0.0051249 0.0058625 0.0014233 0.98646 0.99139 3.0738e-06 1.2295e-05 0.13062 0.86337 0.87245 0.0014165 0.95244 0.54058 0.0019076 0.42462 1.6401 1.6383 16.0102 144.9866 0.00023412 -85.4941 0.40221
0.50623 0.98802 5.5225e-05 3.8182 0.012043 6.6702e-06 0.001154 0.095297 0.00065662 0.095949 0.086464 0 0.040866 0.0389 0 0.85881 0.23294 0.060933 0.0086054 4.1222 0.053941 6.4436e-05 0.83612 0.005125 0.0058626 0.001423 0.98647 0.9914 3.0732e-06 1.2293e-05 0.13062 0.86375 0.87267 0.0014164 0.95272 0.54074 0.0019074 0.42464 1.641 1.6393 16.0102 144.9866 0.00023378 -85.4953 0.40321
0.50723 0.98802 5.5225e-05 3.8182 0.012043 6.6834e-06 0.001154 0.09541 0.00065662 0.096062 0.086567 0 0.040858 0.0389 0 0.85885 0.23296 0.06094 0.0086063 4.1223 0.053946 6.4443e-05 0.83612 0.0051251 0.0058627 0.0014227 0.98647 0.9914 3.0725e-06 1.229e-05 0.13062 0.86412 0.87288 0.0014162 0.95301 0.5409 0.0019072 0.42465 1.642 1.6403 16.0102 144.9867 0.00023343 -85.4965 0.40421
0.50823 0.98802 5.5225e-05 3.8182 0.012043 6.6966e-06 0.001154 0.095522 0.00065663 0.096174 0.086671 0 0.040849 0.0389 0 0.8589 0.23299 0.060948 0.0086073 4.1224 0.053952 6.445e-05 0.83611 0.0051253 0.0058628 0.0014224 0.98648 0.9914 3.0719e-06 1.2288e-05 0.13062 0.86449 0.87309 0.0014161 0.95329 0.54106 0.001907 0.42466 1.643 1.6413 16.0102 144.9867 0.00023309 -85.4977 0.40521
0.50923 0.98802 5.5225e-05 3.8182 0.012043 6.7097e-06 0.001154 0.095634 0.00065663 0.096286 0.086775 0 0.04084 0.0389 0 0.85895 0.23301 0.060955 0.0086083 4.1225 0.053957 6.4457e-05 0.83611 0.0051254 0.0058629 0.0014221 0.98648 0.9914 3.0712e-06 1.2285e-05 0.13062 0.86486 0.87331 0.0014159 0.95357 0.54122 0.0019069 0.42468 1.644 1.6423 16.0102 144.9867 0.00023276 -85.4988 0.40621
0.51023 0.98802 5.5225e-05 3.8182 0.012043 6.7229e-06 0.001154 0.095746 0.00065664 0.096399 0.086878 0 0.040832 0.0389 0 0.859 0.23303 0.060963 0.0086092 4.1226 0.053962 6.4463e-05 0.8361 0.0051255 0.005863 0.0014219 0.98648 0.9914 3.0706e-06 1.2282e-05 0.13063 0.86523 0.87352 0.0014158 0.95385 0.54138 0.0019067 0.42469 1.6449 1.6433 16.0102 144.9867 0.00023242 -85.5 0.40721
0.51123 0.98802 5.5225e-05 3.8182 0.012043 6.7361e-06 0.001154 0.095859 0.00065664 0.096511 0.086981 0 0.040823 0.0389 0 0.85905 0.23305 0.060971 0.0086102 4.1227 0.053968 6.447e-05 0.8361 0.0051256 0.0058632 0.0014216 0.98649 0.99141 3.07e-06 1.228e-05 0.13063 0.8656 0.87373 0.0014156 0.95413 0.54154 0.0019065 0.4247 1.6459 1.6442 16.0102 144.9867 0.00023208 -85.5012 0.40821
0.51223 0.98802 5.5225e-05 3.8182 0.012043 6.7492e-06 0.001154 0.095971 0.00065665 0.096623 0.087085 0 0.040814 0.0389 0 0.8591 0.23307 0.060978 0.0086111 4.1228 0.053973 6.4477e-05 0.83609 0.0051257 0.0058633 0.0014213 0.98649 0.99141 3.0694e-06 1.2277e-05 0.13063 0.86597 0.87394 0.0014155 0.95441 0.5417 0.0019063 0.42471 1.6469 1.6452 16.0102 144.9868 0.00023175 -85.5023 0.40921
0.51323 0.98802 5.5225e-05 3.8182 0.012043 6.7624e-06 0.001154 0.096083 0.00065665 0.096735 0.087188 0 0.040806 0.0389 0 0.85914 0.23309 0.060986 0.0086121 4.1229 0.053979 6.4484e-05 0.83609 0.0051258 0.0058634 0.001421 0.98649 0.99141 3.0687e-06 1.2275e-05 0.13063 0.86634 0.87415 0.0014153 0.95468 0.54185 0.0019061 0.42473 1.6478 1.6462 16.0102 144.9868 0.00023141 -85.5035 0.41021
0.51423 0.98802 5.5224e-05 3.8182 0.012043 6.7755e-06 0.001154 0.096194 0.00065666 0.096846 0.087291 0 0.040797 0.0389 0 0.85919 0.23311 0.060994 0.0086131 4.123 0.053984 6.4491e-05 0.83608 0.005126 0.0058635 0.0014208 0.9865 0.99141 3.0681e-06 1.2272e-05 0.13063 0.8667 0.87436 0.0014152 0.95495 0.54201 0.0019059 0.42474 1.6488 1.6471 16.0102 144.9868 0.00023108 -85.5046 0.41121
0.51523 0.98802 5.5224e-05 3.8182 0.012043 6.7887e-06 0.001154 0.096306 0.00065667 0.096958 0.087394 0 0.040788 0.0389 0 0.85924 0.23313 0.061001 0.008614 4.1231 0.05399 6.4498e-05 0.83607 0.0051261 0.0058636 0.0014205 0.9865 0.99142 3.0675e-06 1.227e-05 0.13063 0.86707 0.87457 0.0014151 0.95522 0.54217 0.0019057 0.42475 1.6498 1.6481 16.0102 144.9868 0.00023075 -85.5057 0.41221
0.51623 0.98802 5.5224e-05 3.8182 0.012043 6.8019e-06 0.001154 0.096418 0.00065667 0.09707 0.087497 0 0.04078 0.0389 0 0.85929 0.23316 0.061009 0.008615 4.1232 0.053995 6.4505e-05 0.83607 0.0051262 0.0058637 0.0014202 0.9865 0.99142 3.0669e-06 1.2268e-05 0.13063 0.86743 0.87477 0.0014149 0.95549 0.54233 0.0019056 0.42477 1.6507 1.6491 16.0102 144.9868 0.00023042 -85.5069 0.41321
0.51723 0.98802 5.5224e-05 3.8182 0.012043 6.815e-06 0.001154 0.096529 0.00065668 0.097181 0.0876 0 0.040771 0.0389 0 0.85934 0.23318 0.061017 0.008616 4.1233 0.054001 6.4512e-05 0.83606 0.0051263 0.0058639 0.00142 0.98651 0.99142 3.0663e-06 1.2265e-05 0.13063 0.86779 0.87498 0.0014148 0.95576 0.54249 0.0019054 0.42478 1.6517 1.65 16.0102 144.9869 0.00023009 -85.508 0.41421
0.51823 0.98802 5.5224e-05 3.8182 0.012043 6.8282e-06 0.001154 0.096641 0.00065668 0.097293 0.087703 0 0.040762 0.0389 0 0.85939 0.2332 0.061025 0.0086169 4.1234 0.054006 6.4519e-05 0.83606 0.0051264 0.005864 0.0014197 0.98651 0.99142 3.0657e-06 1.2263e-05 0.13063 0.86815 0.87519 0.0014147 0.95602 0.54265 0.0019052 0.42479 1.6526 1.651 16.0102 144.9869 0.00022977 -85.5091 0.41521
0.51923 0.98802 5.5224e-05 3.8182 0.012043 6.8414e-06 0.001154 0.096752 0.00065669 0.097404 0.087806 0 0.040754 0.0389 0 0.85943 0.23322 0.061032 0.0086179 4.1235 0.054012 6.4526e-05 0.83605 0.0051266 0.0058641 0.0014195 0.98651 0.99143 3.0651e-06 1.226e-05 0.13063 0.86851 0.87539 0.0014145 0.95629 0.54281 0.001905 0.4248 1.6536 1.6519 16.0102 144.9869 0.00022944 -85.5102 0.41621
0.52023 0.98802 5.5224e-05 3.8182 0.012043 6.8545e-06 0.001154 0.096863 0.00065669 0.097516 0.087909 0 0.040745 0.0389 0 0.85948 0.23324 0.06104 0.0086189 4.1236 0.054017 6.4533e-05 0.83605 0.0051267 0.0058642 0.0014192 0.98652 0.99143 3.0645e-06 1.2258e-05 0.13064 0.86887 0.87559 0.0014144 0.95655 0.54296 0.0019048 0.42482 1.6545 1.6529 16.0102 144.9869 0.00022912 -85.5113 0.41721
0.52123 0.98802 5.5224e-05 3.8182 0.012043 6.8677e-06 0.001154 0.096975 0.0006567 0.097627 0.088011 0 0.040737 0.0389 0 0.85953 0.23326 0.061048 0.0086198 4.1237 0.054023 6.454e-05 0.83604 0.0051268 0.0058643 0.0014189 0.98652 0.99143 3.0639e-06 1.2256e-05 0.13064 0.86923 0.8758 0.0014142 0.95681 0.54312 0.0019047 0.42483 1.6555 1.6538 16.0101 144.9869 0.0002288 -85.5124 0.41821
0.52223 0.98802 5.5224e-05 3.8182 0.012043 6.8809e-06 0.001154 0.097086 0.0006567 0.097738 0.088114 0 0.040728 0.0389 0 0.85958 0.23328 0.061056 0.0086208 4.1238 0.054029 6.4548e-05 0.83604 0.0051269 0.0058645 0.0014187 0.98652 0.99143 3.0633e-06 1.2253e-05 0.13064 0.86959 0.876 0.0014141 0.95707 0.54328 0.0019045 0.42484 1.6564 1.6548 16.0101 144.987 0.00022848 -85.5134 0.41921
0.52323 0.98802 5.5224e-05 3.8182 0.012043 6.894e-06 0.001154 0.097197 0.00065671 0.097849 0.088216 0 0.04072 0.0389 0 0.85963 0.23331 0.061063 0.0086218 4.1239 0.054034 6.4555e-05 0.83603 0.005127 0.0058646 0.0014184 0.98653 0.99143 3.0628e-06 1.2251e-05 0.13064 0.86994 0.8762 0.001414 0.95733 0.54344 0.0019043 0.42486 1.6573 1.6557 16.0101 144.987 0.00022816 -85.5145 0.42021
0.52423 0.98802 5.5224e-05 3.8182 0.012043 6.9072e-06 0.001154 0.097308 0.00065671 0.09796 0.088319 0 0.040711 0.0389 0 0.85968 0.23333 0.061071 0.0086228 4.124 0.05404 6.4562e-05 0.83602 0.0051272 0.0058647 0.0014182 0.98653 0.99144 3.0622e-06 1.2249e-05 0.13064 0.87029 0.8764 0.0014139 0.95758 0.5436 0.0019042 0.42487 1.6583 1.6567 16.0101 144.987 0.00022784 -85.5156 0.42121
0.52523 0.98802 5.5224e-05 3.8182 0.012043 6.9204e-06 0.001154 0.097419 0.00065672 0.098071 0.088421 0 0.040703 0.0389 0 0.85973 0.23335 0.061079 0.0086237 4.1241 0.054045 6.4569e-05 0.83602 0.0051273 0.0058648 0.0014179 0.98653 0.99144 3.0616e-06 1.2246e-05 0.13064 0.87065 0.8766 0.0014137 0.95784 0.54376 0.001904 0.42488 1.6592 1.6576 16.0101 144.987 0.00022752 -85.5166 0.42221
0.52623 0.98802 5.5224e-05 3.8182 0.012043 6.9335e-06 0.001154 0.097529 0.00065672 0.098182 0.088523 0 0.040694 0.0389 0 0.85978 0.23337 0.061087 0.0086247 4.1242 0.054051 6.4576e-05 0.83601 0.0051274 0.0058649 0.0014177 0.98654 0.99144 3.061e-06 1.2244e-05 0.13064 0.871 0.8768 0.0014136 0.95809 0.54391 0.0019038 0.42489 1.6601 1.6586 16.0101 144.987 0.0002272 -85.5177 0.42321
0.52723 0.98802 5.5224e-05 3.8182 0.012043 6.9467e-06 0.001154 0.09764 0.00065673 0.098292 0.088626 0 0.040686 0.0389 0 0.85983 0.23339 0.061095 0.0086257 4.1243 0.054057 6.4583e-05 0.83601 0.0051275 0.0058651 0.0014174 0.98654 0.99144 3.0605e-06 1.2242e-05 0.13064 0.87135 0.877 0.0014135 0.95834 0.54407 0.0019036 0.42491 1.6611 1.6595 16.0101 144.987 0.00022689 -85.5187 0.42421
0.52823 0.98802 5.5224e-05 3.8182 0.012043 6.9599e-06 0.001154 0.097751 0.00065673 0.098403 0.088728 0 0.040677 0.0389 0 0.85988 0.23341 0.061102 0.0086267 4.1244 0.054062 6.459e-05 0.836 0.0051277 0.0058652 0.0014172 0.98654 0.99144 3.0599e-06 1.224e-05 0.13064 0.8717 0.87719 0.0014133 0.95859 0.54423 0.0019035 0.42492 1.662 1.6604 16.0101 144.9871 0.00022658 -85.5197 0.42521
0.52923 0.98802 5.5224e-05 3.8182 0.012043 6.973e-06 0.001154 0.097861 0.00065674 0.098513 0.08883 0 0.040669 0.0389 0 0.85992 0.23344 0.06111 0.0086277 4.1245 0.054068 6.4597e-05 0.836 0.0051278 0.0058653 0.001417 0.98655 0.99145 3.0594e-06 1.2237e-05 0.13064 0.87205 0.87739 0.0014132 0.95884 0.54439 0.0019033 0.42493 1.6629 1.6614 16.0101 144.9871 0.00022626 -85.5207 0.42621
0.53023 0.98802 5.5223e-05 3.8182 0.012043 6.9862e-06 0.001154 0.097972 0.00065674 0.098624 0.088932 0 0.04066 0.0389 0 0.85997 0.23346 0.061118 0.0086287 4.1246 0.054073 6.4604e-05 0.83599 0.0051279 0.0058654 0.0014167 0.98655 0.99145 3.0588e-06 1.2235e-05 0.13065 0.8724 0.87759 0.0014131 0.95908 0.54455 0.0019031 0.42495 1.6639 1.6623 16.0101 144.9871 0.00022595 -85.5218 0.42721
0.53123 0.98802 5.5223e-05 3.8182 0.012043 6.9993e-06 0.001154 0.098082 0.00065675 0.098734 0.089033 0 0.040652 0.0389 0 0.86002 0.23348 0.061126 0.0086296 4.1247 0.054079 6.4612e-05 0.83599 0.005128 0.0058655 0.0014165 0.98655 0.99145 3.0583e-06 1.2233e-05 0.13065 0.87274 0.87778 0.001413 0.95933 0.5447 0.001903 0.42496 1.6648 1.6632 16.0101 144.9871 0.00022564 -85.5228 0.42821
0.53223 0.98802 5.5223e-05 3.8182 0.012043 7.0125e-06 0.001154 0.098192 0.00065675 0.098844 0.089135 0 0.040643 0.0389 0 0.86007 0.2335 0.061134 0.0086306 4.1248 0.054085 6.4619e-05 0.83598 0.0051282 0.0058657 0.0014162 0.98656 0.99145 3.0577e-06 1.2231e-05 0.13065 0.87309 0.87798 0.0014128 0.95957 0.54486 0.0019028 0.42497 1.6657 1.6641 16.0101 144.9871 0.00022533 -85.5238 0.42921
0.53323 0.98802 5.5223e-05 3.8182 0.012043 7.0257e-06 0.001154 0.098302 0.00065676 0.098954 0.089237 0 0.040635 0.0389 0 0.86012 0.23352 0.061142 0.0086316 4.1249 0.05409 6.4626e-05 0.83597 0.0051283 0.0058658 0.001416 0.98656 0.99145 3.0572e-06 1.2229e-05 0.13065 0.87343 0.87817 0.0014127 0.95981 0.54502 0.0019027 0.42498 1.6666 1.665 16.0101 144.9872 0.00022503 -85.5248 0.43021
0.53423 0.98802 5.5223e-05 3.8182 0.012043 7.0388e-06 0.001154 0.098412 0.00065676 0.099064 0.089339 0 0.040626 0.0389 0 0.86017 0.23355 0.06115 0.0086326 4.125 0.054096 6.4633e-05 0.83597 0.0051284 0.0058659 0.0014158 0.98656 0.99146 3.0566e-06 1.2227e-05 0.13065 0.87378 0.87836 0.0014126 0.96005 0.54518 0.0019025 0.425 1.6675 1.666 16.0101 144.9872 0.00022472 -85.5258 0.43121
0.53523 0.98802 5.5223e-05 3.8182 0.012043 7.052e-06 0.001154 0.098522 0.00065677 0.099174 0.08944 0 0.040618 0.0389 0 0.86022 0.23357 0.061158 0.0086336 4.1251 0.054102 6.464e-05 0.83596 0.0051285 0.005866 0.0014155 0.98657 0.99146 3.0561e-06 1.2224e-05 0.13065 0.87412 0.87855 0.0014125 0.96029 0.54534 0.0019023 0.42501 1.6684 1.6669 16.0101 144.9872 0.00022442 -85.5268 0.43221
0.53623 0.98802 5.5223e-05 3.8182 0.012043 7.0652e-06 0.001154 0.098632 0.00065677 0.099284 0.089542 0 0.040609 0.0389 0 0.86027 0.23359 0.061165 0.0086346 4.1252 0.054107 6.4648e-05 0.83596 0.0051287 0.0058662 0.0014153 0.98657 0.99146 3.0556e-06 1.2222e-05 0.13065 0.87446 0.87875 0.0014123 0.96053 0.54549 0.0019022 0.42502 1.6693 1.6678 16.0101 144.9872 0.00022411 -85.5277 0.43321
0.53723 0.98802 5.5223e-05 3.8182 0.012043 7.0783e-06 0.001154 0.098742 0.00065678 0.099394 0.089643 0 0.040601 0.0389 0 0.86032 0.23361 0.061173 0.0086356 4.1253 0.054113 6.4655e-05 0.83595 0.0051288 0.0058663 0.0014151 0.98657 0.99146 3.0551e-06 1.222e-05 0.13065 0.8748 0.87894 0.0014122 0.96076 0.54565 0.001902 0.42504 1.6702 1.6687 16.01 144.9872 0.00022381 -85.5287 0.43421
0.53823 0.98802 5.5223e-05 3.8182 0.012043 7.0915e-06 0.001154 0.098852 0.00065678 0.099504 0.089744 0 0.040593 0.0389 0 0.86037 0.23363 0.061181 0.0086366 4.1254 0.054119 6.4662e-05 0.83595 0.0051289 0.0058664 0.0014148 0.98657 0.99146 3.0545e-06 1.2218e-05 0.13065 0.87514 0.87913 0.0014121 0.961 0.54581 0.0019019 0.42505 1.6711 1.6696 16.01 144.9873 0.00022351 -85.5297 0.43521
0.53923 0.98802 5.5223e-05 3.8182 0.012043 7.1047e-06 0.001154 0.098961 0.00065679 0.099613 0.089845 0 0.040584 0.0389 0 0.86042 0.23365 0.061189 0.0086376 4.1255 0.054124 6.4669e-05 0.83594 0.005129 0.0058665 0.0014146 0.98658 0.99147 3.054e-06 1.2216e-05 0.13066 0.87548 0.87932 0.001412 0.96123 0.54597 0.0019017 0.42506 1.672 1.6705 16.01 144.9873 0.00022321 -85.5306 0.43621
0.54023 0.98802 5.5223e-05 3.8182 0.012043 7.1178e-06 0.001154 0.099071 0.00065679 0.099723 0.089947 0 0.040576 0.0389 0 0.86047 0.23368 0.061197 0.0086386 4.1256 0.05413 6.4677e-05 0.83593 0.0051292 0.0058667 0.0014144 0.98658 0.99147 3.0535e-06 1.2214e-05 0.13066 0.87582 0.8795 0.0014119 0.96146 0.54612 0.0019016 0.42508 1.6729 1.6714 16.01 144.9873 0.00022291 -85.5316 0.43721
0.54123 0.98802 5.5223e-05 3.8182 0.012043 7.131e-06 0.001154 0.09918 0.0006568 0.099832 0.090048 0 0.040567 0.0389 0 0.86052 0.2337 0.061205 0.0086396 4.1257 0.054136 6.4684e-05 0.83593 0.0051293 0.0058668 0.0014142 0.98658 0.99147 3.053e-06 1.2212e-05 0.13066 0.87615 0.87969 0.0014118 0.96169 0.54628 0.0019014 0.42509 1.6738 1.6723 16.01 144.9873 0.00022261 -85.5325 0.43821
0.54223 0.98802 5.5223e-05 3.8182 0.012043 7.1441e-06 0.001154 0.09929 0.0006568 0.099942 0.090149 0 0.040559 0.0389 0 0.86057 0.23372 0.061213 0.0086406 4.1258 0.054142 6.4691e-05 0.83592 0.0051294 0.0058669 0.001414 0.98659 0.99147 3.0525e-06 1.221e-05 0.13066 0.87649 0.87988 0.0014116 0.96192 0.54644 0.0019013 0.4251 1.6747 1.6732 16.01 144.9873 0.00022232 -85.5334 0.43921
0.54323 0.98802 5.5223e-05 3.8182 0.012043 7.1573e-06 0.001154 0.099399 0.00065681 0.10005 0.09025 0 0.040551 0.0389 0 0.86062 0.23374 0.061221 0.0086416 4.1259 0.054147 6.4699e-05 0.83592 0.0051296 0.005867 0.0014137 0.98659 0.99147 3.052e-06 1.2208e-05 0.13066 0.87682 0.88006 0.0014115 0.96215 0.5466 0.0019011 0.42511 1.6756 1.6741 16.01 144.9874 0.00022202 -85.5344 0.44021
0.54423 0.98802 5.5223e-05 3.8182 0.012043 7.1705e-06 0.001154 0.099508 0.00065681 0.10016 0.09035 0 0.040542 0.0389 0 0.86067 0.23377 0.061229 0.0086426 4.126 0.054153 6.4706e-05 0.83591 0.0051297 0.0058672 0.0014135 0.98659 0.99148 3.0515e-06 1.2206e-05 0.13066 0.87715 0.88025 0.0014114 0.96237 0.54675 0.001901 0.42513 1.6765 1.675 16.01 144.9874 0.00022173 -85.5353 0.44121
0.54523 0.98802 5.5223e-05 3.8182 0.012043 7.1836e-06 0.001154 0.099617 0.00065682 0.10027 0.090451 0 0.040534 0.0389 0 0.86072 0.23379 0.061237 0.0086436 4.1261 0.054159 6.4713e-05 0.83591 0.0051298 0.0058673 0.0014133 0.98659 0.99148 3.051e-06 1.2204e-05 0.13066 0.87749 0.88043 0.0014113 0.96259 0.54691 0.0019008 0.42514 1.6774 1.6759 16.01 144.9874 0.00022144 -85.5362 0.44221
0.54623 0.98802 5.5222e-05 3.8182 0.012043 7.1968e-06 0.001154 0.099726 0.00065682 0.10038 0.090552 0 0.040526 0.0389 0 0.86077 0.23381 0.061245 0.0086446 4.1262 0.054165 6.4721e-05 0.8359 0.0051299 0.0058674 0.0014131 0.9866 0.99148 3.0505e-06 1.2202e-05 0.13066 0.87782 0.88062 0.0014112 0.96282 0.54707 0.0019007 0.42515 1.6783 1.6768 16.01 144.9874 0.00022114 -85.5371 0.44321
0.54723 0.98802 5.5222e-05 3.8182 0.012043 7.21e-06 0.001154 0.099835 0.00065683 0.10049 0.090652 0 0.040517 0.0389 0 0.86082 0.23383 0.061253 0.0086456 4.1263 0.05417 6.4728e-05 0.83589 0.0051301 0.0058676 0.0014129 0.9866 0.99148 3.05e-06 1.22e-05 0.13066 0.87815 0.8808 0.0014111 0.96304 0.54722 0.0019005 0.42517 1.6792 1.6777 16.01 144.9874 0.00022085 -85.538 0.44421
0.54823 0.98802 5.5222e-05 3.8182 0.012043 7.2231e-06 0.001154 0.099944 0.00065683 0.1006 0.090753 0 0.040509 0.0389 0 0.86087 0.23385 0.061261 0.0086466 4.1265 0.054176 6.4735e-05 0.83589 0.0051302 0.0058677 0.0014127 0.9866 0.99148 3.0495e-06 1.2198e-05 0.13067 0.87848 0.88098 0.001411 0.96326 0.54738 0.0019004 0.42518 1.68 1.6785 16.01 144.9875 0.00022056 -85.5389 0.44521
0.54923 0.98802 5.5222e-05 3.8182 0.012043 7.2363e-06 0.001154 0.10005 0.00065684 0.1007 0.090853 0 0.040501 0.0389 0 0.86092 0.23388 0.061269 0.0086476 4.1266 0.054182 6.4743e-05 0.83588 0.0051303 0.0058678 0.0014125 0.98661 0.99148 3.0491e-06 1.2196e-05 0.13067 0.8788 0.88117 0.0014109 0.96348 0.54754 0.0019002 0.42519 1.6809 1.6794 16.01 144.9875 0.00022028 -85.5398 0.44621
0.55023 0.98802 5.5222e-05 3.8182 0.012043 7.2495e-06 0.001154 0.10016 0.00065684 0.10081 0.090954 0 0.040493 0.0389 0 0.86098 0.2339 0.061277 0.0086486 4.1267 0.054188 6.475e-05 0.83588 0.0051305 0.0058679 0.0014122 0.98661 0.99149 3.0486e-06 1.2194e-05 0.13067 0.87913 0.88135 0.0014107 0.96369 0.54769 0.0019001 0.42521 1.6818 1.6803 16.0099 144.9875 0.00021999 -85.5407 0.44721
0.55123 0.98802 5.5222e-05 3.8182 0.012043 7.2626e-06 0.001154 0.10027 0.00065685 0.10092 0.091054 0 0.040484 0.0389 0 0.86103 0.23392 0.061285 0.0086496 4.1268 0.054194 6.4757e-05 0.83587 0.0051306 0.0058681 0.001412 0.98661 0.99149 3.0481e-06 1.2192e-05 0.13067 0.87946 0.88153 0.0014106 0.96391 0.54785 0.0018999 0.42522 1.6827 1.6812 16.0099 144.9875 0.0002197 -85.5416 0.44821
0.55223 0.98802 5.5222e-05 3.8182 0.012043 7.2758e-06 0.001154 0.10038 0.00065685 0.10103 0.091154 0 0.040476 0.0389 0 0.86108 0.23394 0.061293 0.0086506 4.1269 0.054199 6.4765e-05 0.83587 0.0051307 0.0058682 0.0014118 0.98661 0.99149 3.0476e-06 1.219e-05 0.13067 0.87978 0.88171 0.0014105 0.96412 0.54801 0.0018998 0.42523 1.6835 1.6821 16.0099 144.9875 0.00021942 -85.5425 0.44921
0.55323 0.98802 5.5222e-05 3.8182 0.012043 7.2889e-06 0.001154 0.10049 0.00065685 0.10114 0.091254 0 0.040468 0.0389 0 0.86113 0.23397 0.061301 0.0086516 4.127 0.054205 6.4772e-05 0.83586 0.0051309 0.0058683 0.0014116 0.98662 0.99149 3.0472e-06 1.2189e-05 0.13067 0.8801 0.88189 0.0014104 0.96434 0.54817 0.0018997 0.42524 1.6844 1.6829 16.0099 144.9876 0.00021914 -85.5433 0.45021
0.55423 0.98802 5.5222e-05 3.8182 0.012043 7.3021e-06 0.001154 0.10059 0.00065686 0.10125 0.091355 0 0.04046 0.0389 0 0.86118 0.23399 0.061309 0.0086527 4.1271 0.054211 6.478e-05 0.83585 0.005131 0.0058685 0.0014114 0.98662 0.99149 3.0467e-06 1.2187e-05 0.13067 0.88043 0.88206 0.0014103 0.96455 0.54832 0.0018995 0.42526 1.6853 1.6838 16.0099 144.9876 0.00021885 -85.5442 0.45121
0.55523 0.98802 5.5222e-05 3.8182 0.012043 7.3153e-06 0.001154 0.1007 0.00065686 0.10136 0.091455 0 0.040451 0.0389 0 0.86123 0.23401 0.061318 0.0086537 4.1272 0.054217 6.4787e-05 0.83585 0.0051311 0.0058686 0.0014112 0.98662 0.99149 3.0462e-06 1.2185e-05 0.13067 0.88075 0.88224 0.0014102 0.96476 0.54848 0.0018994 0.42527 1.6861 1.6847 16.0099 144.9876 0.00021857 -85.5451 0.45221
0.55623 0.98802 5.5222e-05 3.8182 0.012043 7.3284e-06 0.001154 0.10081 0.00065687 0.10146 0.091554 0 0.040443 0.0389 0 0.86128 0.23403 0.061326 0.0086547 4.1273 0.054223 6.4795e-05 0.83584 0.0051313 0.0058687 0.001411 0.98662 0.9915 3.0458e-06 1.2183e-05 0.13067 0.88107 0.88242 0.0014101 0.96497 0.54864 0.0018992 0.42528 1.687 1.6855 16.0099 144.9876 0.00021829 -85.5459 0.45321
0.55723 0.98802 5.5222e-05 3.8182 0.012043 7.3416e-06 0.001154 0.10092 0.00065687 0.10157 0.091654 0 0.040435 0.0389 0 0.86133 0.23406 0.061334 0.0086557 4.1274 0.054229 6.4802e-05 0.83584 0.0051314 0.0058689 0.0014108 0.98663 0.9915 3.0453e-06 1.2181e-05 0.13068 0.88139 0.88259 0.00141 0.96517 0.54879 0.0018991 0.4253 1.6878 1.6864 16.0099 144.9876 0.00021801 -85.5468 0.45421
0.55823 0.98802 5.5222e-05 3.8182 0.012043 7.3548e-06 0.001154 0.10103 0.00065688 0.10168 0.091754 0 0.040427 0.0389 0 0.86138 0.23408 0.061342 0.0086567 4.1275 0.054235 6.4809e-05 0.83583 0.0051315 0.005869 0.0014106 0.98663 0.9915 3.0449e-06 1.2179e-05 0.13068 0.88171 0.88277 0.0014099 0.96538 0.54895 0.001899 0.42531 1.6887 1.6873 16.0099 144.9877 0.00021774 -85.5476 0.45521
0.55923 0.98802 5.5222e-05 3.8182 0.012043 7.3679e-06 0.001154 0.10114 0.00065688 0.10179 0.091854 0 0.040419 0.0389 0 0.86143 0.2341 0.06135 0.0086577 4.1277 0.05424 6.4817e-05 0.83582 0.0051317 0.0058691 0.0014104 0.98663 0.9915 3.0444e-06 1.2178e-05 0.13068 0.88203 0.88294 0.0014098 0.96558 0.5491 0.0018988 0.42532 1.6895 1.6881 16.0099 144.9877 0.00021746 -85.5484 0.45621
0.56023 0.98802 5.5222e-05 3.8182 0.012043 7.3811e-06 0.001154 0.10124 0.00065689 0.1019 0.091953 0 0.04041 0.0389 0 0.86149 0.23412 0.061358 0.0086588 4.1278 0.054246 6.4824e-05 0.83582 0.0051318 0.0058693 0.0014102 0.98663 0.9915 3.044e-06 1.2176e-05 0.13068 0.88234 0.88312 0.0014097 0.96579 0.54926 0.0018987 0.42534 1.6904 1.689 16.0099 144.9877 0.00021718 -85.5493 0.45721
0.56123 0.98802 5.5222e-05 3.8182 0.012043 7.3942e-06 0.001154 0.10135 0.00065689 0.102 0.092053 0 0.040402 0.0389 0 0.86154 0.23415 0.061366 0.0086598 4.1279 0.054252 6.4832e-05 0.83581 0.0051319 0.0058694 0.00141 0.98664 0.9915 3.0435e-06 1.2174e-05 0.13068 0.88266 0.88329 0.0014096 0.96599 0.54942 0.0018986 0.42535 1.6913 1.6898 16.0098 144.9877 0.00021691 -85.5501 0.45821
0.56223 0.98802 5.5221e-05 3.8182 0.012043 7.4074e-06 0.001154 0.10146 0.0006569 0.10211 0.092152 0 0.040394 0.0389 0 0.86159 0.23417 0.061375 0.0086608 4.128 0.054258 6.4839e-05 0.83581 0.0051321 0.0058695 0.0014098 0.98664 0.99151 3.0431e-06 1.2172e-05 0.13068 0.88297 0.88347 0.0014095 0.96619 0.54957 0.0018984 0.42536 1.6921 1.6907 16.0098 144.9877 0.00021664 -85.5509 0.45921
0.56323 0.98802 5.5221e-05 3.8182 0.012043 7.4206e-06 0.001154 0.10157 0.0006569 0.10222 0.092252 0 0.040386 0.0389 0 0.86164 0.23419 0.061383 0.0086618 4.1281 0.054264 6.4847e-05 0.8358 0.0051322 0.0058697 0.0014097 0.98664 0.99151 3.0427e-06 1.2171e-05 0.13068 0.88329 0.88364 0.0014094 0.96639 0.54973 0.0018983 0.42538 1.6929 1.6915 16.0098 144.9878 0.00021636 -85.5517 0.46021
0.56423 0.98802 5.5221e-05 3.8182 0.012043 7.4337e-06 0.001154 0.10167 0.00065691 0.10233 0.092351 0 0.040378 0.0389 0 0.86169 0.23421 0.061391 0.0086629 4.1282 0.05427 6.4854e-05 0.83579 0.0051323 0.0058698 0.0014095 0.98664 0.99151 3.0422e-06 1.2169e-05 0.13068 0.8836 0.88381 0.0014093 0.96659 0.54989 0.0018982 0.42539 1.6938 1.6924 16.0098 144.9878 0.00021609 -85.5525 0.46121
0.56523 0.98802 5.5221e-05 3.8182 0.012043 7.4469e-06 0.001154 0.10178 0.00065691 0.10243 0.09245 0 0.04037 0.0389 0 0.86174 0.23424 0.061399 0.0086639 4.1283 0.054276 6.4862e-05 0.83579 0.0051325 0.0058699 0.0014093 0.98665 0.99151 3.0418e-06 1.2167e-05 0.13068 0.88391 0.88398 0.0014092 0.96678 0.55004 0.0018981 0.4254 1.6946 1.6932 16.0098 144.9878 0.00021582 -85.5533 0.46221
0.56623 0.98802 5.5221e-05 3.8182 0.012043 7.4601e-06 0.001154 0.10189 0.00065691 0.10254 0.092549 0 0.040361 0.0389 0 0.86179 0.23426 0.061407 0.0086649 4.1284 0.054282 6.487e-05 0.83578 0.0051326 0.0058701 0.0014091 0.98665 0.99151 3.0414e-06 1.2165e-05 0.13069 0.88422 0.88415 0.0014091 0.96698 0.5502 0.0018979 0.42541 1.6955 1.6941 16.0098 144.9878 0.00021555 -85.5541 0.46321
0.56723 0.98802 5.5221e-05 3.8182 0.012042 7.4732e-06 0.001154 0.102 0.00065692 0.10265 0.092648 0 0.040353 0.0389 0 0.86185 0.23428 0.061416 0.0086659 4.1286 0.054288 6.4877e-05 0.83578 0.0051328 0.0058702 0.0014089 0.98665 0.99151 3.0409e-06 1.2164e-05 0.13069 0.88453 0.88432 0.001409 0.96718 0.55035 0.0018978 0.42543 1.6963 1.6949 16.0098 144.9878 0.00021528 -85.5549 0.46421
0.56823 0.98802 5.5221e-05 3.8182 0.012042 7.4864e-06 0.001154 0.1021 0.00065692 0.10275 0.092747 0 0.040345 0.0389 0 0.8619 0.23431 0.061424 0.008667 4.1287 0.054294 6.4885e-05 0.83577 0.0051329 0.0058703 0.0014087 0.98665 0.99152 3.0405e-06 1.2162e-05 0.13069 0.88484 0.88449 0.0014089 0.96737 0.55051 0.0018977 0.42544 1.6971 1.6957 16.0098 144.9878 0.00021502 -85.5557 0.46521
0.56923 0.98802 5.5221e-05 3.8182 0.012042 7.4995e-06 0.001154 0.10221 0.00065693 0.10286 0.092846 0 0.040337 0.0389 0 0.86195 0.23433 0.061432 0.008668 4.1288 0.0543 6.4892e-05 0.83577 0.005133 0.0058705 0.0014085 0.98666 0.99152 3.0401e-06 1.216e-05 0.13069 0.88515 0.88466 0.0014088 0.96756 0.55067 0.0018975 0.42545 1.698 1.6966 16.0098 144.9879 0.00021475 -85.5565 0.46621
0.57023 0.98802 5.5221e-05 3.8182 0.012042 7.5127e-06 0.001154 0.10232 0.00065693 0.10297 0.092945 0 0.040329 0.0389 0 0.862 0.23435 0.06144 0.008669 4.1289 0.054306 6.49e-05 0.83576 0.0051332 0.0058706 0.0014084 0.98666 0.99152 3.0397e-06 1.2159e-05 0.13069 0.88546 0.88482 0.0014087 0.96775 0.55082 0.0018974 0.42547 1.6988 1.6974 16.0097 144.9879 0.00021449 -85.5572 0.46721
0.57123 0.98802 5.5221e-05 3.8182 0.012042 7.5259e-06 0.001154 0.10242 0.00065694 0.10308 0.093044 0 0.040321 0.0389 0 0.86205 0.23437 0.061449 0.0086701 4.129 0.054312 6.4907e-05 0.83575 0.0051333 0.0058708 0.0014082 0.98666 0.99152 3.0393e-06 1.2157e-05 0.13069 0.88576 0.88499 0.0014086 0.96794 0.55098 0.0018973 0.42548 1.6996 1.6982 16.0097 144.9879 0.00021422 -85.558 0.46821
0.57223 0.98802 5.5221e-05 3.8182 0.012042 7.539e-06 0.001154 0.10253 0.00065694 0.10318 0.093143 0 0.040313 0.0389 0 0.86211 0.2344 0.061457 0.0086711 4.1291 0.054318 6.4915e-05 0.83575 0.0051335 0.0058709 0.001408 0.98666 0.99152 3.0389e-06 1.2155e-05 0.13069 0.88607 0.88516 0.0014085 0.96813 0.55113 0.0018972 0.42549 1.7004 1.6991 16.0097 144.9879 0.00021396 -85.5588 0.46921
0.57323 0.98802 5.5221e-05 3.8182 0.012042 7.5522e-06 0.001154 0.10264 0.00065695 0.10329 0.093241 0 0.040305 0.0389 0 0.86216 0.23442 0.061465 0.0086722 4.1293 0.054324 6.4923e-05 0.83574 0.0051336 0.005871 0.0014078 0.98667 0.99152 3.0384e-06 1.2154e-05 0.13069 0.88637 0.88532 0.0014084 0.96832 0.55129 0.0018971 0.42551 1.7013 1.6999 16.0097 144.9879 0.0002137 -85.5595 0.47021
0.57423 0.98802 5.5221e-05 3.8182 0.012042 7.5654e-06 0.001154 0.10274 0.00065695 0.1034 0.09334 0 0.040297 0.0389 0 0.86221 0.23444 0.061473 0.0086732 4.1294 0.05433 6.493e-05 0.83574 0.0051337 0.0058712 0.0014076 0.98667 0.99152 3.038e-06 1.2152e-05 0.13069 0.88667 0.88549 0.0014083 0.9685 0.55145 0.0018969 0.42552 1.7021 1.7007 16.0097 144.988 0.00021344 -85.5603 0.47121
0.57523 0.98802 5.5221e-05 3.8182 0.012042 7.5785e-06 0.001154 0.10285 0.00065695 0.1035 0.093438 0 0.040289 0.0389 0 0.86226 0.23447 0.061482 0.0086742 4.1295 0.054336 6.4938e-05 0.83573 0.0051339 0.0058713 0.0014075 0.98667 0.99153 3.0376e-06 1.2151e-05 0.1307 0.88698 0.88565 0.0014082 0.96869 0.5516 0.0018968 0.42553 1.7029 1.7015 16.0097 144.988 0.00021318 -85.561 0.47221
0.57623 0.98802 5.5221e-05 3.8182 0.012042 7.5917e-06 0.001154 0.10296 0.00065696 0.10361 0.093537 0 0.040281 0.0389 0 0.86231 0.23449 0.06149 0.0086753 4.1296 0.054342 6.4946e-05 0.83572 0.005134 0.0058715 0.0014073 0.98667 0.99153 3.0372e-06 1.2149e-05 0.1307 0.88728 0.88582 0.0014081 0.96887 0.55176 0.0018967 0.42555 1.7037 1.7024 16.0097 144.988 0.00021292 -85.5618 0.47321
0.57723 0.98802 5.5221e-05 3.8182 0.012042 7.6048e-06 0.001154 0.10306 0.00065696 0.10371 0.093635 0 0.040273 0.0389 0 0.86237 0.23451 0.061498 0.0086763 4.1297 0.054348 6.4953e-05 0.83572 0.0051342 0.0058716 0.0014071 0.98667 0.99153 3.0368e-06 1.2147e-05 0.1307 0.88758 0.88598 0.0014081 0.96905 0.55191 0.0018966 0.42556 1.7045 1.7032 16.0097 144.988 0.00021266 -85.5625 0.47421
0.57823 0.98802 5.522e-05 3.8182 0.012042 7.618e-06 0.001154 0.10317 0.00065697 0.10382 0.093733 0 0.040265 0.0389 0 0.86242 0.23454 0.061507 0.0086774 4.1298 0.054354 6.4961e-05 0.83571 0.0051343 0.0058717 0.0014069 0.98668 0.99153 3.0365e-06 1.2146e-05 0.1307 0.88788 0.88614 0.001408 0.96924 0.55207 0.0018965 0.42557 1.7054 1.704 16.0097 144.988 0.0002124 -85.5632 0.47521
0.57923 0.98802 5.522e-05 3.8182 0.012042 7.6312e-06 0.001154 0.10327 0.00065697 0.10393 0.093831 0 0.040257 0.0389 0 0.86247 0.23456 0.061515 0.0086784 4.13 0.05436 6.4969e-05 0.83571 0.0051344 0.0058719 0.0014068 0.98668 0.99153 3.0361e-06 1.2144e-05 0.1307 0.88818 0.8863 0.0014079 0.96942 0.55222 0.0018963 0.42559 1.7062 1.7048 16.0096 144.9881 0.00021215 -85.564 0.47621
0.58023 0.98802 5.522e-05 3.8182 0.012042 7.6443e-06 0.001154 0.10338 0.00065698 0.10403 0.093929 0 0.040249 0.0389 0 0.86252 0.23458 0.061523 0.0086794 4.1301 0.054366 6.4976e-05 0.8357 0.0051346 0.005872 0.0014066 0.98668 0.99153 3.0357e-06 1.2143e-05 0.1307 0.88847 0.88646 0.0014078 0.96959 0.55238 0.0018962 0.4256 1.707 1.7056 16.0096 144.9881 0.00021189 -85.5647 0.47721
0.58123 0.98802 5.522e-05 3.8182 0.012042 7.6575e-06 0.001154 0.10349 0.00065698 0.10414 0.094027 0 0.040241 0.0389 0 0.86258 0.23461 0.061532 0.0086805 4.1302 0.054372 6.4984e-05 0.83569 0.0051347 0.0058722 0.0014064 0.98668 0.99153 3.0353e-06 1.2141e-05 0.1307 0.88877 0.88662 0.0014077 0.96977 0.55253 0.0018961 0.42561 1.7078 1.7064 16.0096 144.9881 0.00021164 -85.5654 0.47821
0.58223 0.98802 5.522e-05 3.8182 0.012042 7.6707e-06 0.001154 0.10359 0.00065699 0.10424 0.094125 0 0.040233 0.0389 0 0.86263 0.23463 0.06154 0.0086815 4.1303 0.054378 6.4992e-05 0.83569 0.0051349 0.0058723 0.0014063 0.98669 0.99154 3.0349e-06 1.214e-05 0.1307 0.88907 0.88678 0.0014076 0.96995 0.55269 0.001896 0.42562 1.7086 1.7072 16.0096 144.9881 0.00021139 -85.5661 0.47921
0.58323 0.98802 5.522e-05 3.8182 0.012042 7.6838e-06 0.001154 0.1037 0.00065699 0.10435 0.094223 0 0.040225 0.0389 0 0.86268 0.23465 0.061548 0.0086826 4.1304 0.054384 6.5e-05 0.83568 0.005135 0.0058724 0.0014061 0.98669 0.99154 3.0345e-06 1.2138e-05 0.13071 0.88936 0.88694 0.0014075 0.97012 0.55285 0.0018959 0.42564 1.7094 1.7081 16.0096 144.9881 0.00021114 -85.5668 0.48021
0.58423 0.98802 5.522e-05 3.8182 0.012042 7.697e-06 0.001154 0.1038 0.00065699 0.10446 0.094321 0 0.040217 0.0389 0 0.86273 0.23467 0.061557 0.0086836 4.1306 0.05439 6.5007e-05 0.83567 0.0051352 0.0058726 0.0014059 0.98669 0.99154 3.0341e-06 1.2137e-05 0.13071 0.88965 0.8871 0.0014074 0.9703 0.553 0.0018958 0.42565 1.7102 1.7089 16.0096 144.9882 0.00021088 -85.5675 0.48121
0.58523 0.98802 5.522e-05 3.8182 0.012042 7.7101e-06 0.001154 0.10391 0.000657 0.10456 0.094419 0 0.040209 0.0389 0 0.86279 0.2347 0.061565 0.0086847 4.1307 0.054396 6.5015e-05 0.83567 0.0051353 0.0058727 0.0014058 0.98669 0.99154 3.0338e-06 1.2135e-05 0.13071 0.88995 0.88726 0.0014074 0.97047 0.55316 0.0018957 0.42566 1.711 1.7097 16.0096 144.9882 0.00021063 -85.5682 0.48221
0.58623 0.98802 5.522e-05 3.8182 0.012042 7.7233e-06 0.001154 0.10402 0.000657 0.10467 0.094516 0 0.040201 0.0389 0 0.86284 0.23472 0.061574 0.0086857 4.1308 0.054402 6.5023e-05 0.83566 0.0051355 0.0058729 0.0014056 0.98669 0.99154 3.0334e-06 1.2134e-05 0.13071 0.89024 0.88742 0.0014073 0.97065 0.55331 0.0018955 0.42568 1.7118 1.7105 16.0096 144.9882 0.00021039 -85.5689 0.48321
0.58723 0.98802 5.522e-05 3.8182 0.012042 7.7365e-06 0.001154 0.10412 0.00065701 0.10477 0.094614 0 0.040193 0.0389 0 0.86289 0.23475 0.061582 0.0086868 4.1309 0.054408 6.5031e-05 0.83566 0.0051356 0.005873 0.0014055 0.9867 0.99154 3.033e-06 1.2132e-05 0.13071 0.89053 0.88758 0.0014072 0.97082 0.55347 0.0018954 0.42569 1.7126 1.7113 16.0096 144.9882 0.00021014 -85.5696 0.48421
0.58823 0.98802 5.522e-05 3.8182 0.012042 7.7496e-06 0.001154 0.10423 0.00065701 0.10488 0.094711 0 0.040185 0.0389 0 0.86295 0.23477 0.06159 0.0086878 4.131 0.054414 6.5038e-05 0.83565 0.0051357 0.0058732 0.0014053 0.9867 0.99154 3.0327e-06 1.2131e-05 0.13071 0.89082 0.88773 0.0014071 0.97099 0.55362 0.0018953 0.4257 1.7134 1.7121 16.0095 144.9882 0.00020989 -85.5703 0.48521
0.58923 0.98802 5.522e-05 3.8182 0.012042 7.7628e-06 0.001154 0.10433 0.00065702 0.10498 0.094809 0 0.040177 0.0389 0 0.863 0.23479 0.061599 0.0086889 4.1312 0.054421 6.5046e-05 0.83564 0.0051359 0.0058733 0.0014051 0.9867 0.99155 3.0323e-06 1.2129e-05 0.13071 0.89111 0.88789 0.001407 0.97116 0.55378 0.0018952 0.42572 1.7142 1.7128 16.0095 144.9883 0.00020964 -85.571 0.48621
0.59023 0.98802 5.522e-05 3.8182 0.012042 7.776e-06 0.001154 0.10444 0.00065702 0.10509 0.094906 0 0.040169 0.0389 0 0.86305 0.23482 0.061607 0.00869 4.1313 0.054427 6.5054e-05 0.83564 0.005136 0.0058735 0.001405 0.9867 0.99155 3.0319e-06 1.2128e-05 0.13071 0.8914 0.88804 0.0014069 0.97132 0.55393 0.0018951 0.42573 1.7149 1.7136 16.0095 144.9883 0.0002094 -85.5716 0.48721
0.59123 0.98802 5.522e-05 3.8182 0.012042 7.7891e-06 0.001154 0.10454 0.00065702 0.10519 0.095003 0 0.040161 0.0389 0 0.8631 0.23484 0.061616 0.008691 4.1314 0.054433 6.5062e-05 0.83563 0.0051362 0.0058736 0.0014048 0.9867 0.99155 3.0316e-06 1.2126e-05 0.13071 0.89169 0.8882 0.0014068 0.97149 0.55409 0.001895 0.42574 1.7157 1.7144 16.0095 144.9883 0.00020916 -85.5723 0.48821
0.59223 0.98802 5.522e-05 3.8182 0.012042 7.8023e-06 0.001154 0.10465 0.00065703 0.1053 0.0951 0 0.040153 0.0389 0 0.86316 0.23486 0.061624 0.0086921 4.1315 0.054439 6.507e-05 0.83563 0.0051363 0.0058737 0.0014047 0.98671 0.99155 3.0312e-06 1.2125e-05 0.13072 0.89197 0.88835 0.0014068 0.97166 0.55424 0.0018949 0.42576 1.7165 1.7152 16.0095 144.9883 0.00020891 -85.573 0.48921
0.59323 0.98802 5.522e-05 3.8182 0.012042 7.8154e-06 0.001154 0.10475 0.00065703 0.1054 0.095197 0 0.040146 0.0389 0 0.86321 0.23489 0.061633 0.0086931 4.1316 0.054445 6.5077e-05 0.83562 0.0051365 0.0058739 0.0014045 0.98671 0.99155 3.0309e-06 1.2123e-05 0.13072 0.89226 0.8885 0.0014067 0.97182 0.5544 0.0018948 0.42577 1.7173 1.716 16.0095 144.9883 0.00020867 -85.5736 0.49021
0.59423 0.98802 5.522e-05 3.8182 0.012042 7.8286e-06 0.001154 0.10486 0.00065704 0.10551 0.095294 0 0.040138 0.0389 0 0.86326 0.23491 0.061641 0.0086942 4.1318 0.054451 6.5085e-05 0.83561 0.0051366 0.005874 0.0014044 0.98671 0.99155 3.0305e-06 1.2122e-05 0.13072 0.89254 0.88866 0.0014066 0.97198 0.55455 0.0018947 0.42578 1.7181 1.7168 16.0095 144.9884 0.00020843 -85.5743 0.49121
0.59523 0.98802 5.5219e-05 3.8182 0.012042 7.8418e-06 0.001154 0.10496 0.00065704 0.10561 0.095391 0 0.04013 0.0389 0 0.86332 0.23493 0.06165 0.0086953 4.1319 0.054457 6.5093e-05 0.83561 0.0051368 0.0058742 0.0014042 0.98671 0.99155 3.0302e-06 1.2121e-05 0.13072 0.89283 0.88881 0.0014065 0.97215 0.5547 0.0018946 0.4258 1.7189 1.7176 16.0095 144.9884 0.00020819 -85.5749 0.49221
0.59623 0.98802 5.5219e-05 3.8182 0.012042 7.8549e-06 0.001154 0.10507 0.00065704 0.10572 0.095488 0 0.040122 0.0389 0 0.86337 0.23496 0.061658 0.0086963 4.132 0.054464 6.5101e-05 0.8356 0.0051369 0.0058743 0.001404 0.98671 0.99156 3.0298e-06 1.2119e-05 0.13072 0.89311 0.88896 0.0014064 0.97231 0.55486 0.0018945 0.42581 1.7196 1.7183 16.0094 144.9884 0.00020795 -85.5756 0.49321
0.59723 0.98802 5.5219e-05 3.8182 0.012042 7.8681e-06 0.001154 0.10517 0.00065705 0.10582 0.095585 0 0.040114 0.0389 0 0.86342 0.23498 0.061667 0.0086974 4.1321 0.05447 6.5109e-05 0.8356 0.0051371 0.0058745 0.0014039 0.98672 0.99156 3.0295e-06 1.2118e-05 0.13072 0.89339 0.88911 0.0014064 0.97247 0.55501 0.0018944 0.42582 1.7204 1.7191 16.0094 144.9884 0.00020771 -85.5762 0.49421
0.59823 0.98802 5.5219e-05 3.8182 0.012042 7.8812e-06 0.001154 0.10528 0.00065705 0.10593 0.095682 0 0.040106 0.0389 0 0.86348 0.235 0.061675 0.0086985 4.1323 0.054476 6.5117e-05 0.83559 0.0051372 0.0058746 0.0014037 0.98672 0.99156 3.0291e-06 1.2116e-05 0.13072 0.89367 0.88926 0.0014063 0.97263 0.55517 0.0018943 0.42583 1.7212 1.7199 16.0094 144.9884 0.00020747 -85.5769 0.49521
0.59923 0.98802 5.5219e-05 3.8182 0.012042 7.8944e-06 0.001154 0.10538 0.00065706 0.10603 0.095778 0 0.040099 0.0389 0 0.86353 0.23503 0.061684 0.0086995 4.1324 0.054482 6.5125e-05 0.83558 0.0051374 0.0058748 0.0014036 0.98672 0.99156 3.0288e-06 1.2115e-05 0.13072 0.89395 0.88941 0.0014062 0.97279 0.55532 0.0018942 0.42585 1.7219 1.7207 16.0094 144.9885 0.00020724 -85.5775 0.49621
0.60023 0.98802 5.5219e-05 3.8182 0.012042 7.9076e-06 0.001154 0.10548 0.00065706 0.10614 0.095875 0 0.040091 0.0389 0 0.86359 0.23505 0.061692 0.0087006 4.1325 0.054488 6.5133e-05 0.83558 0.0051375 0.0058749 0.0014034 0.98672 0.99156 3.0284e-06 1.2114e-05 0.13073 0.89423 0.88956 0.0014061 0.97294 0.55548 0.0018941 0.42586 1.7227 1.7214 16.0094 144.9885 0.000207 -85.5781 0.49721
0.60123 0.98802 5.5219e-05 3.8182 0.012042 7.9207e-06 0.001154 0.10559 0.00065706 0.10624 0.095971 0 0.040083 0.0389 0 0.86364 0.23507 0.061701 0.0087017 4.1326 0.054495 6.5141e-05 0.83557 0.0051377 0.0058751 0.0014033 0.98672 0.99156 3.0281e-06 1.2112e-05 0.13073 0.89451 0.88971 0.0014061 0.9731 0.55563 0.001894 0.42587 1.7235 1.7222 16.0094 144.9885 0.00020677 -85.5788 0.49821
0.60223 0.98802 5.5219e-05 3.8182 0.012042 7.9339e-06 0.001154 0.10569 0.00065707 0.10635 0.096068 0 0.040075 0.0389 0 0.86369 0.2351 0.061709 0.0087027 4.1328 0.054501 6.5148e-05 0.83556 0.0051378 0.0058752 0.0014032 0.98673 0.99156 3.0278e-06 1.2111e-05 0.13073 0.89479 0.88986 0.001406 0.97326 0.55579 0.0018939 0.42589 1.7242 1.723 16.0094 144.9885 0.00020653 -85.5794 0.49921
0.60323 0.98802 5.5219e-05 3.8182 0.012042 7.947e-06 0.001154 0.1058 0.00065707 0.10645 0.096164 0 0.040067 0.0389 0 0.86375 0.23512 0.061718 0.0087038 4.1329 0.054507 6.5156e-05 0.83556 0.005138 0.0058754 0.001403 0.98673 0.99156 3.0274e-06 1.211e-05 0.13073 0.89507 0.89001 0.0014059 0.97341 0.55594 0.0018938 0.4259 1.725 1.7238 16.0093 144.9885 0.0002063 -85.58 0.50021
0.60423 0.98802 5.5219e-05 3.8182 0.012042 7.9602e-06 0.001154 0.1059 0.00065708 0.10655 0.09626 0 0.04006 0.0389 0 0.8638 0.23515 0.061727 0.0087049 4.133 0.054513 6.5164e-05 0.83555 0.0051381 0.0058755 0.0014029 0.98673 0.99156 3.0271e-06 1.2108e-05 0.13073 0.89534 0.89015 0.0014058 0.97357 0.55609 0.0018937 0.42591 1.7258 1.7245 16.0093 144.9886 0.00020607 -85.5806 0.50121
0.60523 0.98802 5.5219e-05 3.8182 0.012042 7.9734e-06 0.001154 0.106 0.00065708 0.10666 0.096357 0 0.040052 0.0389 0 0.86386 0.23517 0.061735 0.008706 4.1331 0.05452 6.5172e-05 0.83555 0.0051383 0.0058757 0.0014027 0.98673 0.99157 3.0268e-06 1.2107e-05 0.13073 0.89562 0.8903 0.0014058 0.97372 0.55625 0.0018936 0.42593 1.7265 1.7253 16.0093 144.9886 0.00020584 -85.5812 0.50221
0.60623 0.98802 5.5219e-05 3.8182 0.012042 7.9865e-06 0.001154 0.10611 0.00065709 0.10676 0.096453 0 0.040044 0.0389 0 0.86391 0.23519 0.061744 0.008707 4.1333 0.054526 6.518e-05 0.83554 0.0051384 0.0058758 0.0014026 0.98673 0.99157 3.0265e-06 1.2106e-05 0.13073 0.89589 0.89045 0.0014057 0.97387 0.5564 0.0018935 0.42594 1.7273 1.726 16.0093 144.9886 0.00020561 -85.5818 0.50321
0.60723 0.98802 5.5219e-05 3.8182 0.012042 7.9997e-06 0.001154 0.10621 0.00065709 0.10687 0.096549 0 0.040036 0.0389 0 0.86396 0.23522 0.061752 0.0087081 4.1334 0.054532 6.5188e-05 0.83553 0.0051386 0.005876 0.0014024 0.98673 0.99157 3.0261e-06 1.2105e-05 0.13074 0.89617 0.89059 0.0014056 0.97402 0.55656 0.0018934 0.42595 1.728 1.7268 16.0093 144.9886 0.00020538 -85.5824 0.50421
0.60823 0.98802 5.5219e-05 3.8182 0.012042 8.0129e-06 0.001154 0.10632 0.00065709 0.10697 0.096645 0 0.040029 0.0389 0 0.86402 0.23524 0.061761 0.0087092 4.1335 0.054538 6.5196e-05 0.83553 0.0051388 0.0058761 0.0014023 0.98674 0.99157 3.0258e-06 1.2103e-05 0.13074 0.89644 0.89074 0.0014055 0.97417 0.55671 0.0018933 0.42597 1.7288 1.7276 16.0093 144.9886 0.00020515 -85.583 0.50521
0.60923 0.98802 5.5219e-05 3.8182 0.012042 8.026e-06 0.001154 0.10642 0.0006571 0.10707 0.096741 0 0.040021 0.0389 0 0.86407 0.23527 0.06177 0.0087103 4.1337 0.054545 6.5204e-05 0.83552 0.0051389 0.0058763 0.0014022 0.98674 0.99157 3.0255e-06 1.2102e-05 0.13074 0.89671 0.89088 0.0014055 0.97432 0.55687 0.0018932 0.42598 1.7295 1.7283 16.0093 144.9887 0.00020492 -85.5836 0.50621
0.61023 0.98802 5.5219e-05 3.8182 0.012042 8.0392e-06 0.001154 0.10652 0.0006571 0.10718 0.096837 0 0.040013 0.0389 0 0.86413 0.23529 0.061778 0.0087113 4.1338 0.054551 6.5212e-05 0.83551 0.0051391 0.0058764 0.001402 0.98674 0.99157 3.0252e-06 1.2101e-05 0.13074 0.89698 0.89103 0.0014054 0.97447 0.55702 0.0018931 0.42599 1.7303 1.7291 16.0092 144.9887 0.00020469 -85.5842 0.50721
0.61123 0.98802 5.5218e-05 3.8182 0.012042 8.0523e-06 0.001154 0.10663 0.00065711 0.10728 0.096932 0 0.040005 0.0389 0 0.86418 0.23531 0.061787 0.0087124 4.1339 0.054557 6.522e-05 0.83551 0.0051392 0.0058766 0.0014019 0.98674 0.99157 3.0249e-06 1.2099e-05 0.13074 0.89725 0.89117 0.0014053 0.97461 0.55717 0.001893 0.42601 1.731 1.7298 16.0092 144.9887 0.00020447 -85.5848 0.50821
0.61223 0.98802 5.5218e-05 3.8182 0.012042 8.0655e-06 0.001154 0.10673 0.00065711 0.10738 0.097028 0 0.039998 0.0389 0 0.86423 0.23534 0.061795 0.0087135 4.134 0.054564 6.5228e-05 0.8355 0.0051394 0.0058767 0.0014018 0.98674 0.99157 3.0246e-06 1.2098e-05 0.13074 0.89752 0.89131 0.0014052 0.97476 0.55733 0.0018929 0.42602 1.7318 1.7306 16.0092 144.9887 0.00020424 -85.5854 0.50921
0.61323 0.98802 5.5218e-05 3.8182 0.012042 8.0787e-06 0.001154 0.10683 0.00065711 0.10749 0.097124 0 0.03999 0.0389 0 0.86429 0.23536 0.061804 0.0087146 4.1342 0.05457 6.5236e-05 0.8355 0.0051395 0.0058769 0.0014016 0.98675 0.99158 3.0243e-06 1.2097e-05 0.13074 0.89779 0.89145 0.0014052 0.9749 0.55748 0.0018928 0.42603 1.7325 1.7313 16.0092 144.9887 0.00020402 -85.586 0.51021
0.61423 0.98802 5.5218e-05 3.8182 0.012042 8.0918e-06 0.001154 0.10694 0.00065712 0.10759 0.097219 0 0.039982 0.0389 0 0.86434 0.23539 0.061813 0.0087157 4.1343 0.054576 6.5244e-05 0.83549 0.0051397 0.0058771 0.0014015 0.98675 0.99158 3.024e-06 1.2096e-05 0.13074 0.89806 0.8916 0.0014051 0.97505 0.55763 0.0018927 0.42605 1.7333 1.732 16.0092 144.9888 0.0002038 -85.5865 0.51121
0.61523 0.98802 5.5218e-05 3.8182 0.012042 8.105e-06 0.001154 0.10704 0.00065712 0.10769 0.097315 0 0.039975 0.0389 0 0.8644 0.23541 0.061821 0.0087168 4.1344 0.054583 6.5252e-05 0.83548 0.0051398 0.0058772 0.0014014 0.98675 0.99158 3.0236e-06 1.2095e-05 0.13075 0.89833 0.89174 0.001405 0.97519 0.55779 0.0018926 0.42606 1.734 1.7328 16.0092 144.9888 0.00020357 -85.5871 0.51221
0.61623 0.98802 5.5218e-05 3.8182 0.012042 8.1181e-06 0.001154 0.10714 0.00065712 0.1078 0.09741 0 0.039967 0.0389 0 0.86445 0.23543 0.06183 0.0087178 4.1346 0.054589 6.5261e-05 0.83548 0.00514 0.0058774 0.0014012 0.98675 0.99158 3.0233e-06 1.2093e-05 0.13075 0.89859 0.89188 0.001405 0.97533 0.55794 0.0018925 0.42607 1.7347 1.7335 16.0092 144.9888 0.00020335 -85.5877 0.51321
0.61723 0.98802 5.5218e-05 3.8182 0.012042 8.1313e-06 0.001154 0.10725 0.00065713 0.1079 0.097505 0 0.039959 0.0389 0 0.86451 0.23546 0.061839 0.0087189 4.1347 0.054595 6.5269e-05 0.83547 0.0051402 0.0058775 0.0014011 0.98675 0.99158 3.023e-06 1.2092e-05 0.13075 0.89886 0.89202 0.0014049 0.97547 0.55809 0.0018924 0.42608 1.7355 1.7343 16.0091 144.9888 0.00020313 -85.5882 0.51421
0.61823 0.98802 5.5218e-05 3.8182 0.012042 8.1445e-06 0.001154 0.10735 0.00065713 0.108 0.097601 0 0.039952 0.0389 0 0.86456 0.23548 0.061848 0.00872 4.1348 0.054602 6.5277e-05 0.83546 0.0051403 0.0058777 0.001401 0.98675 0.99158 3.0227e-06 1.2091e-05 0.13075 0.89912 0.89216 0.0014048 0.97561 0.55825 0.0018923 0.4261 1.7362 1.735 16.0091 144.9888 0.00020291 -85.5888 0.51521
0.61923 0.98802 5.5218e-05 3.8182 0.012042 8.1576e-06 0.001154 0.10745 0.00065714 0.1081 0.097696 0 0.039944 0.0389 0 0.86462 0.23551 0.061856 0.0087211 4.135 0.054608 6.5285e-05 0.83546 0.0051405 0.0058778 0.0014008 0.98676 0.99158 3.0225e-06 1.209e-05 0.13075 0.89938 0.8923 0.0014048 0.97575 0.5584 0.0018923 0.42611 1.7369 1.7357 16.0091 144.9889 0.00020269 -85.5893 0.51621
0.62023 0.98802 5.5218e-05 3.8182 0.012042 8.1708e-06 0.001154 0.10755 0.00065714 0.10821 0.097791 0 0.039936 0.0389 0 0.86467 0.23553 0.061865 0.0087222 4.1351 0.054614 6.5293e-05 0.83545 0.0051406 0.005878 0.0014007 0.98676 0.99158 3.0222e-06 1.2089e-05 0.13075 0.89965 0.89243 0.0014047 0.97589 0.55856 0.0018922 0.42612 1.7377 1.7365 16.0091 144.9889 0.00020247 -85.5899 0.51721
0.62123 0.98802 5.5218e-05 3.8182 0.012042 8.1839e-06 0.001154 0.10766 0.00065714 0.10831 0.097886 0 0.039929 0.0389 0 0.86473 0.23555 0.061874 0.0087233 4.1352 0.054621 6.5301e-05 0.83544 0.0051408 0.0058781 0.0014006 0.98676 0.99158 3.0219e-06 1.2087e-05 0.13075 0.89991 0.89257 0.0014046 0.97603 0.55871 0.0018921 0.42614 1.7384 1.7372 16.0091 144.9889 0.00020226 -85.5904 0.51821
0.62223 0.98802 5.5218e-05 3.8182 0.012042 8.1971e-06 0.001154 0.10776 0.00065715 0.10841 0.097981 0 0.039921 0.0389 0 0.86478 0.23558 0.061883 0.0087244 4.1354 0.054627 6.5309e-05 0.83544 0.0051409 0.0058783 0.0014004 0.98676 0.99159 3.0216e-06 1.2086e-05 0.13075 0.90017 0.89271 0.0014046 0.97617 0.55886 0.001892 0.42615 1.7391 1.7379 16.0091 144.9889 0.00020204 -85.591 0.51921
0.62323 0.98802 5.5218e-05 3.8182 0.012042 8.2103e-06 0.001154 0.10786 0.00065715 0.10851 0.098076 0 0.039914 0.0389 0 0.86484 0.2356 0.061891 0.0087255 4.1355 0.054633 6.5317e-05 0.83543 0.0051411 0.0058785 0.0014003 0.98676 0.99159 3.0213e-06 1.2085e-05 0.13076 0.90043 0.89285 0.0014045 0.9763 0.55902 0.0018919 0.42616 1.7399 1.7387 16.0091 144.9889 0.00020182 -85.5915 0.52021
0.62423 0.98802 5.5218e-05 3.8182 0.012042 8.2234e-06 0.001154 0.10796 0.00065716 0.10862 0.09817 0 0.039906 0.0389 0 0.86489 0.23563 0.0619 0.0087266 4.1356 0.05464 6.5325e-05 0.83543 0.0051413 0.0058786 0.0014002 0.98676 0.99159 3.021e-06 1.2084e-05 0.13076 0.90069 0.89298 0.0014044 0.97644 0.55917 0.0018918 0.42618 1.7406 1.7394 16.009 144.989 0.00020161 -85.5921 0.52121
0.62523 0.98802 5.5218e-05 3.8182 0.012042 8.2366e-06 0.001154 0.10807 0.00065716 0.10872 0.098265 0 0.039898 0.0389 0 0.86495 0.23565 0.061909 0.0087277 4.1358 0.054646 6.5334e-05 0.83542 0.0051414 0.0058788 0.0014001 0.98677 0.99159 3.0207e-06 1.2083e-05 0.13076 0.90095 0.89312 0.0014044 0.97657 0.55932 0.0018917 0.42619 1.7413 1.7401 16.009 144.989 0.00020139 -85.5926 0.52221
0.62623 0.98802 5.5218e-05 3.8182 0.012042 8.2497e-06 0.001154 0.10817 0.00065716 0.10882 0.09836 0 0.039891 0.0389 0 0.865 0.23568 0.061918 0.0087288 4.1359 0.054653 6.5342e-05 0.83541 0.0051416 0.0058789 0.0013999 0.98677 0.99159 3.0204e-06 1.2082e-05 0.13076 0.90121 0.89326 0.0014043 0.9767 0.55947 0.0018916 0.4262 1.742 1.7408 16.009 144.989 0.00020118 -85.5931 0.52321
0.62723 0.98802 5.5217e-05 3.8182 0.012042 8.2629e-06 0.001154 0.10827 0.00065717 0.10892 0.098454 0 0.039883 0.0389 0 0.86506 0.2357 0.061926 0.0087299 4.136 0.054659 6.535e-05 0.83541 0.0051417 0.0058791 0.0013998 0.98677 0.99159 3.0201e-06 1.2081e-05 0.13076 0.90146 0.89339 0.0014042 0.97684 0.55963 0.0018916 0.42622 1.7427 1.7416 16.009 144.989 0.00020097 -85.5937 0.52421
0.62823 0.98802 5.5217e-05 3.8182 0.012042 8.2761e-06 0.001154 0.10837 0.00065717 0.10903 0.098549 0 0.039876 0.0389 0 0.86511 0.23572 0.061935 0.008731 4.1362 0.054666 6.5358e-05 0.8354 0.0051419 0.0058793 0.0013997 0.98677 0.99159 3.0199e-06 1.2079e-05 0.13076 0.90172 0.89352 0.0014042 0.97697 0.55978 0.0018915 0.42623 1.7435 1.7423 16.009 144.989 0.00020076 -85.5942 0.52521
0.62923 0.98802 5.5217e-05 3.8182 0.012042 8.2892e-06 0.001154 0.10848 0.00065717 0.10913 0.098643 0 0.039868 0.0389 0 0.86517 0.23575 0.061944 0.0087321 4.1363 0.054672 6.5366e-05 0.83539 0.0051421 0.0058794 0.0013996 0.98677 0.99159 3.0196e-06 1.2078e-05 0.13076 0.90197 0.89366 0.0014041 0.9771 0.55993 0.0018914 0.42624 1.7442 1.743 16.009 144.9891 0.00020055 -85.5947 0.52621
0.63023 0.98802 5.5217e-05 3.8182 0.012042 8.3024e-06 0.001154 0.10858 0.00065718 0.10923 0.098738 0 0.039861 0.0389 0 0.86522 0.23577 0.061953 0.0087332 4.1364 0.054678 6.5375e-05 0.83539 0.0051422 0.0058796 0.0013995 0.98677 0.99159 3.0193e-06 1.2077e-05 0.13077 0.90223 0.89379 0.001404 0.97723 0.56009 0.0018913 0.42626 1.7449 1.7437 16.0089 144.9891 0.00020034 -85.5952 0.52721
0.63123 0.98802 5.5217e-05 3.8182 0.012042 8.3155e-06 0.001154 0.10868 0.00065718 0.10933 0.098832 0 0.039853 0.0389 0 0.86528 0.2358 0.061962 0.0087343 4.1366 0.054685 6.5383e-05 0.83538 0.0051424 0.0058797 0.0013993 0.98678 0.99159 3.019e-06 1.2076e-05 0.13077 0.90248 0.89392 0.001404 0.97736 0.56024 0.0018912 0.42627 1.7456 1.7444 16.0089 144.9891 0.00020013 -85.5957 0.52821
0.63223 0.98802 5.5217e-05 3.8182 0.012042 8.3287e-06 0.001154 0.10878 0.00065719 0.10943 0.098926 0 0.039846 0.0389 0 0.86533 0.23582 0.06197 0.0087354 4.1367 0.054691 6.5391e-05 0.83537 0.0051426 0.0058799 0.0013992 0.98678 0.9916 3.0188e-06 1.2075e-05 0.13077 0.90274 0.89406 0.0014039 0.97749 0.56039 0.0018911 0.42628 1.7463 1.7451 16.0089 144.9891 0.00019992 -85.5962 0.52921
0.63323 0.98802 5.5217e-05 3.8182 0.012042 8.3419e-06 0.001154 0.10888 0.00065719 0.10953 0.09902 0 0.039838 0.0389 0 0.86539 0.23585 0.061979 0.0087365 4.1368 0.054698 6.5399e-05 0.83537 0.0051427 0.0058801 0.0013991 0.98678 0.9916 3.0185e-06 1.2074e-05 0.13077 0.90299 0.89419 0.0014038 0.97761 0.56055 0.0018911 0.4263 1.747 1.7459 16.0089 144.9891 0.00019971 -85.5967 0.53021
0.63423 0.98802 5.5217e-05 3.8182 0.012042 8.355e-06 0.001154 0.10898 0.00065719 0.10964 0.099114 0 0.039831 0.0389 0 0.86545 0.23587 0.061988 0.0087376 4.137 0.054704 6.5408e-05 0.83536 0.0051429 0.0058802 0.001399 0.98678 0.9916 3.0182e-06 1.2073e-05 0.13077 0.90324 0.89432 0.0014038 0.97774 0.5607 0.001891 0.42631 1.7477 1.7466 16.0089 144.9892 0.0001995 -85.5972 0.53121
0.63523 0.98802 5.5217e-05 3.8182 0.012042 8.3682e-06 0.001154 0.10909 0.0006572 0.10974 0.099208 0 0.039823 0.0389 0 0.8655 0.2359 0.061997 0.0087387 4.1371 0.054711 6.5416e-05 0.83535 0.0051431 0.0058804 0.0013989 0.98678 0.9916 3.018e-06 1.2072e-05 0.13077 0.90349 0.89445 0.0014037 0.97787 0.56085 0.0018909 0.42632 1.7484 1.7473 16.0089 144.9892 0.0001993 -85.5977 0.53221
0.63623 0.98802 5.5217e-05 3.8182 0.012042 8.3813e-06 0.001154 0.10919 0.0006572 0.10984 0.099302 0 0.039816 0.0389 0 0.86556 0.23592 0.062006 0.0087398 4.1373 0.054717 6.5424e-05 0.83535 0.0051432 0.0058805 0.0013988 0.98678 0.9916 3.0177e-06 1.2071e-05 0.13077 0.90374 0.89458 0.0014037 0.97799 0.561 0.0018908 0.42633 1.7491 1.748 16.0088 144.9892 0.00019909 -85.5982 0.53321
0.63723 0.98802 5.5217e-05 3.8182 0.012042 8.3945e-06 0.001154 0.10929 0.0006572 0.10994 0.099396 0 0.039808 0.0389 0 0.86561 0.23595 0.062015 0.0087409 4.1374 0.054724 6.5432e-05 0.83534 0.0051434 0.0058807 0.0013986 0.98678 0.9916 3.0174e-06 1.207e-05 0.13077 0.90399 0.89471 0.0014036 0.97812 0.56116 0.0018907 0.42635 1.7498 1.7487 16.0088 144.9892 0.00019889 -85.5987 0.53421
0.63823 0.98802 5.5217e-05 3.8182 0.012042 8.4077e-06 0.001154 0.10939 0.00065721 0.11004 0.09949 0 0.039801 0.0389 0 0.86567 0.23597 0.062024 0.008742 4.1375 0.05473 6.5441e-05 0.83534 0.0051435 0.0058809 0.0013985 0.98679 0.9916 3.0172e-06 1.2069e-05 0.13078 0.90424 0.89484 0.0014035 0.97824 0.56131 0.0018907 0.42636 1.7505 1.7494 16.0088 144.9892 0.00019868 -85.5992 0.53521
0.63923 0.98802 5.5217e-05 3.8182 0.012042 8.4208e-06 0.001154 0.10949 0.00065721 0.11014 0.099584 0 0.039793 0.0389 0 0.86572 0.23599 0.062033 0.0087431 4.1377 0.054737 6.5449e-05 0.83533 0.0051437 0.005881 0.0013984 0.98679 0.9916 3.0169e-06 1.2068e-05 0.13078 0.90449 0.89497 0.0014035 0.97836 0.56146 0.0018906 0.42637 1.7512 1.7501 16.0088 144.9893 0.00019848 -85.5997 0.53621
0.64023 0.98802 5.5217e-05 3.8182 0.012042 8.434e-06 0.001154 0.10959 0.00065722 0.11024 0.099677 0 0.039786 0.0389 0 0.86578 0.23602 0.062041 0.0087442 4.1378 0.054743 6.5457e-05 0.83532 0.0051439 0.0058812 0.0013983 0.98679 0.9916 3.0167e-06 1.2067e-05 0.13078 0.90473 0.8951 0.0014034 0.97848 0.56161 0.0018905 0.42639 1.7519 1.7508 16.0088 144.9893 0.00019828 -85.6002 0.53721
0.64123 0.98802 5.5217e-05 3.8182 0.012042 8.4471e-06 0.001154 0.10969 0.00065722 0.11035 0.099771 0 0.039778 0.0389 0 0.86584 0.23604 0.06205 0.0087454 4.138 0.05475 6.5466e-05 0.83532 0.005144 0.0058814 0.0013982 0.98679 0.9916 3.0164e-06 1.2066e-05 0.13078 0.90498 0.89523 0.0014034 0.9786 0.56177 0.0018904 0.4264 1.7526 1.7515 16.0088 144.9893 0.00019808 -85.6006 0.53821
0.64223 0.98802 5.5217e-05 3.8182 0.012042 8.4603e-06 0.001154 0.10979 0.00065722 0.11045 0.099864 0 0.039771 0.0389 0 0.86589 0.23607 0.062059 0.0087465 4.1381 0.054756 6.5474e-05 0.83531 0.0051442 0.0058815 0.0013981 0.98679 0.99161 3.0162e-06 1.2065e-05 0.13078 0.90522 0.89535 0.0014033 0.97872 0.56192 0.0018904 0.42641 1.7533 1.7522 16.0087 144.9893 0.00019787 -85.6011 0.53921
0.64323 0.98802 5.5216e-05 3.8182 0.012041 8.4735e-06 0.001154 0.10989 0.00065723 0.11055 0.099958 0 0.039763 0.0389 0 0.86595 0.23609 0.062068 0.0087476 4.1382 0.054763 6.5482e-05 0.8353 0.0051444 0.0058817 0.001398 0.98679 0.99161 3.0159e-06 1.2064e-05 0.13078 0.90547 0.89548 0.0014032 0.97884 0.56207 0.0018903 0.42643 1.754 1.7529 16.0087 144.9893 0.00019767 -85.6016 0.54021
0.64423 0.98802 5.5216e-05 3.8182 0.012041 8.4866e-06 0.001154 0.11 0.00065723 0.11065 0.10005 0 0.039756 0.0389 0 0.866 0.23612 0.062077 0.0087487 4.1384 0.054769 6.5491e-05 0.8353 0.0051445 0.0058819 0.0013979 0.98679 0.99161 3.0157e-06 1.2063e-05 0.13078 0.90571 0.89561 0.0014032 0.97896 0.56222 0.0018902 0.42644 1.7547 1.7535 16.0087 144.9894 0.00019748 -85.6021 0.54121
0.64523 0.98802 5.5216e-05 3.8182 0.012041 8.4998e-06 0.001154 0.1101 0.00065723 0.11075 0.10014 0 0.039749 0.0389 0 0.86606 0.23614 0.062086 0.0087498 4.1385 0.054776 6.5499e-05 0.83529 0.0051447 0.005882 0.0013978 0.9868 0.99161 3.0154e-06 1.2062e-05 0.13079 0.90596 0.89573 0.0014031 0.97908 0.56237 0.0018901 0.42645 1.7554 1.7542 16.0087 144.9894 0.00019728 -85.6025 0.54221
0.64623 0.98802 5.5216e-05 3.8182 0.012041 8.5129e-06 0.001154 0.1102 0.00065724 0.11085 0.10024 0 0.039741 0.0389 0 0.86612 0.23617 0.062095 0.0087509 4.1387 0.054783 6.5507e-05 0.83528 0.0051449 0.0058822 0.0013976 0.9868 0.99161 3.0152e-06 1.2061e-05 0.13079 0.9062 0.89586 0.0014031 0.9792 0.56253 0.0018901 0.42647 1.756 1.7549 16.0087 144.9894 0.00019708 -85.603 0.54321
0.64723 0.98802 5.5216e-05 3.8182 0.012041 8.5261e-06 0.001154 0.1103 0.00065724 0.11095 0.10033 0 0.039734 0.0389 0 0.86617 0.23619 0.062104 0.0087521 4.1388 0.054789 6.5516e-05 0.83528 0.0051451 0.0058824 0.0013975 0.9868 0.99161 3.0149e-06 1.206e-05 0.13079 0.90644 0.89599 0.001403 0.97931 0.56268 0.00189 0.42648 1.7567 1.7556 16.0087 144.9894 0.00019688 -85.6034 0.54421
0.64823 0.98802 5.5216e-05 3.8182 0.012041 8.5392e-06 0.001154 0.1104 0.00065724 0.11105 0.10042 0 0.039726 0.0389 0 0.86623 0.23622 0.062113 0.0087532 4.1389 0.054796 6.5524e-05 0.83527 0.0051452 0.0058825 0.0013974 0.9868 0.99161 3.0147e-06 1.2059e-05 0.13079 0.90668 0.89611 0.001403 0.97943 0.56283 0.0018899 0.42649 1.7574 1.7563 16.0086 144.9894 0.00019669 -85.6039 0.54521
0.64923 0.98802 5.5216e-05 3.8182 0.012041 8.5524e-06 0.001154 0.1105 0.00065725 0.11115 0.10052 0 0.039719 0.0389 0 0.86629 0.23624 0.062122 0.0087543 4.1391 0.054802 6.5532e-05 0.83526 0.0051454 0.0058827 0.0013973 0.9868 0.99161 3.0144e-06 1.2058e-05 0.13079 0.90692 0.89623 0.0014029 0.97955 0.56298 0.0018898 0.42651 1.7581 1.757 16.0086 144.9895 0.00019649 -85.6044 0.54621
0.65023 0.98802 5.5216e-05 3.8182 0.012041 8.5656e-06 0.001154 0.1106 0.00065725 0.11125 0.10061 0 0.039712 0.0389 0 0.86634 0.23627 0.062131 0.0087554 4.1392 0.054809 6.5541e-05 0.83526 0.0051456 0.0058829 0.0013972 0.9868 0.99161 3.0142e-06 1.2057e-05 0.13079 0.90716 0.89636 0.0014029 0.97966 0.56313 0.0018898 0.42652 1.7588 1.7577 16.0086 144.9895 0.0001963 -85.6048 0.54721
0.65123 0.98802 5.5216e-05 3.8182 0.012041 8.5787e-06 0.001154 0.1107 0.00065726 0.11135 0.1007 0 0.039704 0.0389 0 0.8664 0.23629 0.06214 0.0087566 4.1394 0.054816 6.5549e-05 0.83525 0.0051457 0.005883 0.0013971 0.9868 0.99161 3.014e-06 1.2056e-05 0.13079 0.9074 0.89648 0.0014028 0.97977 0.56329 0.0018897 0.42653 1.7594 1.7583 16.0086 144.9895 0.0001961 -85.6053 0.54821
0.65223 0.98802 5.5216e-05 3.8182 0.012041 8.5919e-06 0.001154 0.1108 0.00065726 0.11145 0.1008 0 0.039697 0.0389 0 0.86646 0.23632 0.062149 0.0087577 4.1395 0.054822 6.5558e-05 0.83524 0.0051459 0.0058832 0.001397 0.98681 0.99161 3.0137e-06 1.2055e-05 0.1308 0.90763 0.8966 0.0014027 0.97989 0.56344 0.0018896 0.42655 1.7601 1.759 16.0086 144.9895 0.00019591 -85.6057 0.54921
0.65323 0.98802 5.5216e-05 3.8182 0.012041 8.605e-06 0.001154 0.1109 0.00065726 0.11155 0.10089 0 0.03969 0.0389 0 0.86651 0.23634 0.062158 0.0087588 4.1397 0.054829 6.5566e-05 0.83524 0.0051461 0.0058834 0.0013969 0.98681 0.99161 3.0135e-06 1.2054e-05 0.1308 0.90787 0.89673 0.0014027 0.98 0.56359 0.0018896 0.42656 1.7608 1.7597 16.0086 144.9895 0.00019571 -85.6061 0.55021
0.65423 0.98802 5.5216e-05 3.8182 0.012041 8.6182e-06 0.001154 0.111 0.00065727 0.11165 0.10098 0 0.039682 0.0389 0 0.86657 0.23637 0.062167 0.0087599 4.1398 0.054835 6.5575e-05 0.83523 0.0051462 0.0058835 0.0013968 0.98681 0.99162 3.0132e-06 1.2053e-05 0.1308 0.90811 0.89685 0.0014026 0.98011 0.56374 0.0018895 0.42657 1.7615 1.7604 16.0085 144.9896 0.00019552 -85.6066 0.55121
0.65523 0.98802 5.5216e-05 3.8182 0.012041 8.6314e-06 0.001154 0.1111 0.00065727 0.11175 0.10107 0 0.039675 0.0389 0 0.86663 0.23639 0.062176 0.0087611 4.14 0.054842 6.5583e-05 0.83522 0.0051464 0.0058837 0.0013967 0.98681 0.99162 3.013e-06 1.2052e-05 0.1308 0.90834 0.89697 0.0014026 0.98022 0.56389 0.0018894 0.42658 1.7621 1.761 16.0085 144.9896 0.00019533 -85.607 0.55221
0.65623 0.98802 5.5216e-05 3.8182 0.012041 8.6445e-06 0.001154 0.1112 0.00065727 0.11185 0.10117 0 0.039668 0.0389 0 0.86668 0.23642 0.062185 0.0087622 4.1401 0.054849 6.5591e-05 0.83522 0.0051466 0.0058839 0.0013966 0.98681 0.99162 3.0128e-06 1.2051e-05 0.1308 0.90858 0.89709 0.0014025 0.98033 0.56404 0.0018893 0.4266 1.7628 1.7617 16.0085 144.9896 0.00019514 -85.6074 0.55321
0.65723 0.98802 5.5216e-05 3.8182 0.012041 8.6577e-06 0.001154 0.1113 0.00065728 0.11195 0.10126 0 0.03966 0.0389 0 0.86674 0.23644 0.062194 0.0087633 4.1402 0.054855 6.56e-05 0.83521 0.0051468 0.0058841 0.0013965 0.98681 0.99162 3.0126e-06 1.205e-05 0.1308 0.90881 0.89721 0.0014025 0.98044 0.5642 0.0018893 0.42661 1.7635 1.7624 16.0085 144.9896 0.00019495 -85.6079 0.55421
0.65823 0.98802 5.5216e-05 3.8182 0.012041 8.6708e-06 0.001154 0.1114 0.00065728 0.11205 0.10135 0 0.039653 0.0389 0 0.8668 0.23647 0.062203 0.0087645 4.1404 0.054862 6.5608e-05 0.8352 0.0051469 0.0058842 0.0013964 0.98681 0.99162 3.0123e-06 1.2049e-05 0.1308 0.90905 0.89733 0.0014024 0.98055 0.56435 0.0018892 0.42662 1.7641 1.763 16.0085 144.9896 0.00019476 -85.6083 0.55521
0.65923 0.98802 5.5215e-05 3.8182 0.012041 8.684e-06 0.001154 0.1115 0.00065728 0.11215 0.10144 0 0.039646 0.0389 0 0.86685 0.23649 0.062212 0.0087656 4.1405 0.054869 6.5617e-05 0.8352 0.0051471 0.0058844 0.0013963 0.98681 0.99162 3.0121e-06 1.2048e-05 0.13081 0.90928 0.89745 0.0014024 0.98065 0.5645 0.0018891 0.42664 1.7648 1.7637 16.0084 144.9897 0.00019457 -85.6087 0.55621
0.66023 0.98802 5.5215e-05 3.8182 0.012041 8.6972e-06 0.001154 0.1116 0.00065729 0.11225 0.10153 0 0.039638 0.0389 0 0.86691 0.23652 0.062221 0.0087667 4.1407 0.054875 6.5625e-05 0.83519 0.0051473 0.0058846 0.0013962 0.98682 0.99162 3.0119e-06 1.2047e-05 0.13081 0.90951 0.89757 0.0014023 0.98076 0.56465 0.0018891 0.42665 1.7654 1.7644 16.0084 144.9897 0.00019439 -85.6091 0.55721
0.66123 0.98802 5.5215e-05 3.8182 0.012041 8.7103e-06 0.001154 0.1117 0.00065729 0.11235 0.10163 0 0.039631 0.0389 0 0.86697 0.23654 0.062231 0.0087679 4.1408 0.054882 6.5634e-05 0.83518 0.0051475 0.0058847 0.0013961 0.98682 0.99162 3.0117e-06 1.2047e-05 0.13081 0.90974 0.89769 0.0014023 0.98087 0.5648 0.001889 0.42666 1.7661 1.765 16.0084 144.9897 0.0001942 -85.6096 0.55821
0.66223 0.98802 5.5215e-05 3.8182 0.012041 8.7235e-06 0.001154 0.1118 0.00065729 0.11245 0.10172 0 0.039624 0.0389 0 0.86703 0.23657 0.06224 0.008769 4.141 0.054889 6.5642e-05 0.83518 0.0051476 0.0058849 0.001396 0.98682 0.99162 3.0114e-06 1.2046e-05 0.13081 0.90997 0.89781 0.0014022 0.98097 0.56495 0.0018889 0.42668 1.7668 1.7657 16.0084 144.9897 0.00019401 -85.61 0.55921
0.66323 0.98802 5.5215e-05 3.8182 0.012041 8.7366e-06 0.001154 0.11189 0.0006573 0.11255 0.10181 0 0.039617 0.0389 0 0.86708 0.23659 0.062249 0.0087701 4.1411 0.054895 6.5651e-05 0.83517 0.0051478 0.0058851 0.0013959 0.98682 0.99162 3.0112e-06 1.2045e-05 0.13081 0.9102 0.89793 0.0014022 0.98108 0.5651 0.0018889 0.42669 1.7674 1.7664 16.0084 144.9897 0.00019383 -85.6104 0.56021
0.66423 0.98802 5.5215e-05 3.8182 0.012041 8.7498e-06 0.001154 0.11199 0.0006573 0.11265 0.1019 0 0.039609 0.0389 0 0.86714 0.23662 0.062258 0.0087713 4.1413 0.054902 6.5659e-05 0.83516 0.005148 0.0058853 0.0013958 0.98682 0.99162 3.011e-06 1.2044e-05 0.13081 0.91043 0.89805 0.0014021 0.98118 0.56526 0.0018888 0.4267 1.7681 1.767 16.0084 144.9898 0.00019364 -85.6108 0.56121
0.66523 0.98802 5.5215e-05 3.8182 0.012041 8.7629e-06 0.001154 0.11209 0.0006573 0.11275 0.10199 0 0.039602 0.0389 0 0.8672 0.23665 0.062267 0.0087724 4.1414 0.054909 6.5668e-05 0.83516 0.0051482 0.0058854 0.0013957 0.98682 0.99162 3.0108e-06 1.2043e-05 0.13081 0.91066 0.89816 0.0014021 0.98129 0.56541 0.0018887 0.42672 1.7687 1.7677 16.0083 144.9898 0.00019346 -85.6112 0.56221
0.66623 0.98802 5.5215e-05 3.8182 0.012041 8.7761e-06 0.001154 0.11219 0.00065731 0.11284 0.10209 0 0.039595 0.0389 0 0.86725 0.23667 0.062276 0.0087736 4.1416 0.054915 6.5677e-05 0.83515 0.0051483 0.0058856 0.0013956 0.98682 0.99163 3.0106e-06 1.2042e-05 0.13082 0.91089 0.89828 0.001402 0.98139 0.56556 0.0018887 0.42673 1.7694 1.7683 16.0083 144.9898 0.00019327 -85.6116 0.56321
0.66723 0.98802 5.5215e-05 3.8182 0.012041 8.7893e-06 0.001154 0.11229 0.00065731 0.11294 0.10218 0 0.039588 0.0389 0 0.86731 0.2367 0.062285 0.0087747 4.1417 0.054922 6.5685e-05 0.83514 0.0051485 0.0058858 0.0013955 0.98682 0.99163 3.0103e-06 1.2041e-05 0.13082 0.91111 0.8984 0.001402 0.98149 0.56571 0.0018886 0.42674 1.77 1.769 16.0083 144.9898 0.00019309 -85.612 0.56421
0.66823 0.98802 5.5215e-05 3.8182 0.012041 8.8024e-06 0.001154 0.11239 0.00065731 0.11304 0.10227 0 0.03958 0.0389 0 0.86737 0.23672 0.062294 0.0087758 4.1419 0.054929 6.5694e-05 0.83514 0.0051487 0.005886 0.0013954 0.98683 0.99163 3.0101e-06 1.204e-05 0.13082 0.91134 0.89851 0.0014019 0.98159 0.56586 0.0018885 0.42676 1.7707 1.7696 16.0083 144.9898 0.00019291 -85.6124 0.56521
0.66923 0.98802 5.5215e-05 3.8182 0.012041 8.8156e-06 0.001154 0.11249 0.00065732 0.11314 0.10236 0 0.039573 0.0389 0 0.86743 0.23675 0.062304 0.008777 4.142 0.054936 6.5702e-05 0.83513 0.0051489 0.0058861 0.0013954 0.98683 0.99163 3.0099e-06 1.204e-05 0.13082 0.91156 0.89863 0.0014019 0.98169 0.56601 0.0018885 0.42677 1.7713 1.7703 16.0083 144.9899 0.00019273 -85.6128 0.56621
0.67023 0.98802 5.5215e-05 3.8182 0.012041 8.8287e-06 0.001154 0.11259 0.00065732 0.11324 0.10245 0 0.039566 0.0389 0 0.86748 0.23677 0.062313 0.0087781 4.1422 0.054942 6.5711e-05 0.83512 0.005149 0.0058863 0.0013953 0.98683 0.99163 3.0097e-06 1.2039e-05 0.13082 0.91179 0.89874 0.0014018 0.9818 0.56616 0.0018884 0.42678 1.772 1.7709 16.0082 144.9899 0.00019255 -85.6132 0.56721
0.67123 0.98802 5.5215e-05 3.8182 0.012041 8.8419e-06 0.001154 0.11269 0.00065732 0.11334 0.10254 0 0.039559 0.0389 0 0.86754 0.2368 0.062322 0.0087793 4.1423 0.054949 6.572e-05 0.83512 0.0051492 0.0058865 0.0013952 0.98683 0.99163 3.0095e-06 1.2038e-05 0.13082 0.91201 0.89886 0.0014018 0.98189 0.56631 0.0018884 0.42679 1.7726 1.7716 16.0082 144.9899 0.00019237 -85.6136 0.56821
0.67223 0.98802 5.5215e-05 3.8182 0.012041 8.8551e-06 0.001154 0.11278 0.00065733 0.11344 0.10264 0 0.039552 0.0389 0 0.8676 0.23682 0.062331 0.0087804 4.1425 0.054956 6.5728e-05 0.83511 0.0051494 0.0058867 0.0013951 0.98683 0.99163 3.0093e-06 1.2037e-05 0.13082 0.91224 0.89897 0.0014017 0.98199 0.56646 0.0018883 0.42681 1.7733 1.7722 16.0082 144.9899 0.00019219 -85.614 0.56921
0.67323 0.98802 5.5215e-05 3.8182 0.012041 8.8682e-06 0.001154 0.11288 0.00065733 0.11354 0.10273 0 0.039544 0.0389 0 0.86766 0.23685 0.06234 0.0087816 4.1426 0.054963 6.5737e-05 0.8351 0.0051496 0.0058869 0.001395 0.98683 0.99163 3.0091e-06 1.2036e-05 0.13083 0.91246 0.89908 0.0014017 0.98209 0.56661 0.0018882 0.42682 1.7739 1.7729 16.0082 144.9899 0.00019201 -85.6144 0.57021
0.67423 0.98802 5.5215e-05 3.8182 0.012041 8.8814e-06 0.001154 0.11298 0.00065733 0.11363 0.10282 0 0.039537 0.0389 0 0.86772 0.23687 0.06235 0.0087827 4.1428 0.054969 6.5745e-05 0.8351 0.0051498 0.005887 0.0013949 0.98683 0.99163 3.0089e-06 1.2035e-05 0.13083 0.91268 0.8992 0.0014016 0.98219 0.56676 0.0018882 0.42683 1.7745 1.7735 16.0082 144.99 0.00019183 -85.6148 0.57121
0.67523 0.98802 5.5214e-05 3.8182 0.012041 8.8945e-06 0.001154 0.11308 0.00065734 0.11373 0.10291 0 0.03953 0.0389 0 0.86777 0.2369 0.062359 0.0087839 4.1429 0.054976 6.5754e-05 0.83509 0.0051499 0.0058872 0.0013948 0.98683 0.99163 3.0087e-06 1.2035e-05 0.13083 0.9129 0.89931 0.0014016 0.98229 0.56691 0.0018881 0.42685 1.7752 1.7741 16.0081 144.99 0.00019165 -85.6151 0.57221
0.67623 0.98802 5.5214e-05 3.8182 0.012041 8.9077e-06 0.001154 0.11318 0.00065734 0.11383 0.103 0 0.039523 0.0389 0 0.86783 0.23693 0.062368 0.008785 4.1431 0.054983 6.5763e-05 0.83508 0.0051501 0.0058874 0.0013947 0.98683 0.99163 3.0085e-06 1.2034e-05 0.13083 0.91312 0.89942 0.0014015 0.98238 0.56707 0.0018881 0.42686 1.7758 1.7748 16.0081 144.99 0.00019147 -85.6155 0.57321
0.67723 0.98802 5.5214e-05 3.8182 0.012041 8.9208e-06 0.001154 0.11328 0.00065734 0.11393 0.10309 0 0.039516 0.0389 0 0.86789 0.23695 0.062377 0.0087862 4.1432 0.05499 6.5771e-05 0.83508 0.0051503 0.0058876 0.0013946 0.98684 0.99163 3.0083e-06 1.2033e-05 0.13083 0.91334 0.89954 0.0014015 0.98248 0.56722 0.001888 0.42687 1.7764 1.7754 16.0081 144.99 0.0001913 -85.6159 0.57421
0.67823 0.98802 5.5214e-05 3.8182 0.012041 8.934e-06 0.001154 0.11337 0.00065735 0.11403 0.10318 0 0.039509 0.0389 0 0.86795 0.23698 0.062386 0.0087873 4.1434 0.054997 6.578e-05 0.83507 0.0051505 0.0058877 0.0013946 0.98684 0.99163 3.0081e-06 1.2032e-05 0.13083 0.91356 0.89965 0.0014014 0.98258 0.56737 0.0018879 0.42689 1.7771 1.7761 16.0081 144.99 0.00019112 -85.6163 0.57521
0.67923 0.98802 5.5214e-05 3.8182 0.012041 8.9472e-06 0.001154 0.11347 0.00065735 0.11412 0.10327 0 0.039501 0.0389 0 0.86801 0.237 0.062396 0.0087885 4.1435 0.055003 6.5789e-05 0.83506 0.0051507 0.0058879 0.0013945 0.98684 0.99164 3.0079e-06 1.2031e-05 0.13084 0.91378 0.89976 0.0014014 0.98267 0.56752 0.0018879 0.4269 1.7777 1.7767 16.0081 144.9901 0.00019095 -85.6166 0.57621
0.68023 0.98802 5.5214e-05 3.8182 0.012041 8.9603e-06 0.001154 0.11357 0.00065735 0.11422 0.10336 0 0.039494 0.0389 0 0.86806 0.23703 0.062405 0.0087896 4.1437 0.05501 6.5797e-05 0.83506 0.0051508 0.0058881 0.0013944 0.98684 0.99164 3.0077e-06 1.2031e-05 0.13084 0.914 0.89987 0.0014014 0.98276 0.56767 0.0018878 0.42691 1.7783 1.7773 16.0081 144.9901 0.00019077 -85.617 0.57721
0.68123 0.98802 5.5214e-05 3.8182 0.012041 8.9735e-06 0.001154 0.11367 0.00065736 0.11432 0.10345 0 0.039487 0.0389 0 0.86812 0.23705 0.062414 0.0087908 4.1439 0.055017 6.5806e-05 0.83505 0.005151 0.0058883 0.0013943 0.98684 0.99164 3.0075e-06 1.203e-05 0.13084 0.91422 0.89998 0.0014013 0.98286 0.56782 0.0018878 0.42693 1.779 1.778 16.008 144.9901 0.0001906 -85.6174 0.57821
0.68223 0.98802 5.5214e-05 3.8182 0.012041 8.9866e-06 0.001154 0.11376 0.00065736 0.11442 0.10354 0 0.03948 0.0389 0 0.86818 0.23708 0.062423 0.008792 4.144 0.055024 6.5815e-05 0.83504 0.0051512 0.0058885 0.0013942 0.98684 0.99164 3.0073e-06 1.2029e-05 0.13084 0.91443 0.90009 0.0014013 0.98295 0.56797 0.0018877 0.42694 1.7796 1.7786 16.008 144.9901 0.00019043 -85.6177 0.57921
0.68323 0.98802 5.5214e-05 3.8182 0.012041 8.9998e-06 0.001154 0.11386 0.00065736 0.11452 0.10364 0 0.039473 0.0389 0 0.86824 0.2371 0.062433 0.0087931 4.1442 0.055031 6.5823e-05 0.83504 0.0051514 0.0058887 0.0013941 0.98684 0.99164 3.0071e-06 1.2028e-05 0.13084 0.91465 0.9002 0.0014012 0.98304 0.56812 0.0018876 0.42695 1.7802 1.7792 16.008 144.9901 0.00019025 -85.6181 0.58021
0.68423 0.98802 5.5214e-05 3.8182 0.012041 9.0129e-06 0.001154 0.11396 0.00065737 0.11461 0.10373 0 0.039466 0.0389 0 0.8683 0.23713 0.062442 0.0087943 4.1443 0.055038 6.5832e-05 0.83503 0.0051516 0.0058888 0.001394 0.98684 0.99164 3.0069e-06 1.2028e-05 0.13084 0.91486 0.90031 0.0014012 0.98313 0.56827 0.0018876 0.42697 1.7808 1.7798 16.008 144.9902 0.00019008 -85.6184 0.58121
0.68523 0.98802 5.5214e-05 3.8182 0.012041 9.0261e-06 0.001154 0.11406 0.00065737 0.11471 0.10382 0 0.039459 0.0389 0 0.86835 0.23716 0.062451 0.0087954 4.1445 0.055044 6.5841e-05 0.83502 0.0051518 0.005889 0.001394 0.98684 0.99164 3.0067e-06 1.2027e-05 0.13084 0.91508 0.90042 0.0014011 0.98323 0.56842 0.0018875 0.42698 1.7815 1.7805 16.008 144.9902 0.00018991 -85.6188 0.58221
0.68623 0.98802 5.5214e-05 3.8182 0.012041 9.0393e-06 0.001154 0.11415 0.00065737 0.11481 0.10391 0 0.039452 0.0389 0 0.86841 0.23718 0.062461 0.0087966 4.1446 0.055051 6.585e-05 0.83501 0.0051519 0.0058892 0.0013939 0.98685 0.99164 3.0065e-06 1.2026e-05 0.13085 0.91529 0.90053 0.0014011 0.98332 0.56857 0.0018875 0.42699 1.7821 1.7811 16.0079 144.9902 0.00018974 -85.6192 0.58321
0.68723 0.98802 5.5214e-05 3.8182 0.012041 9.0524e-06 0.001154 0.11425 0.00065738 0.11491 0.104 0 0.039445 0.0389 0 0.86847 0.23721 0.06247 0.0087978 4.1448 0.055058 6.5858e-05 0.83501 0.0051521 0.0058894 0.0013938 0.98685 0.99164 3.0064e-06 1.2025e-05 0.13085 0.9155 0.90064 0.0014011 0.98341 0.56872 0.0018874 0.427 1.7827 1.7817 16.0079 144.9902 0.00018957 -85.6195 0.58421
0.68823 0.98802 5.5214e-05 3.8182 0.012041 9.0656e-06 0.001154 0.11435 0.00065738 0.115 0.10409 0 0.039438 0.0389 0 0.86853 0.23723 0.062479 0.0087989 4.145 0.055065 6.5867e-05 0.835 0.0051523 0.0058896 0.0013937 0.98685 0.99164 3.0062e-06 1.2025e-05 0.13085 0.91572 0.90074 0.001401 0.98349 0.56887 0.0018874 0.42702 1.7833 1.7823 16.0079 144.9902 0.0001894 -85.6199 0.58521
0.68923 0.98802 5.5214e-05 3.8182 0.012041 9.0787e-06 0.001154 0.11445 0.00065738 0.1151 0.10418 0 0.039431 0.0389 0 0.86859 0.23726 0.062489 0.0088001 4.1451 0.055072 6.5876e-05 0.83499 0.0051525 0.0058898 0.0013936 0.98685 0.99164 3.006e-06 1.2024e-05 0.13085 0.91593 0.90085 0.001401 0.98358 0.56902 0.0018873 0.42703 1.7839 1.783 16.0079 144.9903 0.00018923 -85.6202 0.58621
0.69023 0.98802 5.5214e-05 3.8182 0.012041 9.0919e-06 0.001154 0.11454 0.00065739 0.1152 0.10427 0 0.039424 0.0389 0 0.86865 0.23729 0.062498 0.0088012 4.1453 0.055079 6.5885e-05 0.83499 0.0051527 0.0058899 0.0013936 0.98685 0.99164 3.0058e-06 1.2023e-05 0.13085 0.91614 0.90096 0.0014009 0.98367 0.56917 0.0018872 0.42704 1.7846 1.7836 16.0079 144.9903 0.00018906 -85.6205 0.58721
0.69123 0.98802 5.5213e-05 3.8182 0.012041 9.105e-06 0.001154 0.11464 0.00065739 0.11529 0.10436 0 0.039416 0.0389 0 0.86871 0.23731 0.062507 0.0088024 4.1454 0.055086 6.5894e-05 0.83498 0.0051529 0.0058901 0.0013935 0.98685 0.99164 3.0056e-06 1.2022e-05 0.13085 0.91635 0.90106 0.0014009 0.98376 0.56932 0.0018872 0.42706 1.7852 1.7842 16.0078 144.9903 0.0001889 -85.6209 0.58821
0.69223 0.98802 5.5213e-05 3.8182 0.012041 9.1182e-06 0.001154 0.11474 0.00065739 0.11539 0.10445 0 0.039409 0.0389 0 0.86877 0.23734 0.062517 0.0088036 4.1456 0.055093 6.5902e-05 0.83497 0.0051531 0.0058903 0.0013934 0.98685 0.99164 3.0054e-06 1.2022e-05 0.13086 0.91656 0.90117 0.0014008 0.98385 0.56947 0.0018871 0.42707 1.7858 1.7848 16.0078 144.9903 0.00018873 -85.6212 0.58921
0.69323 0.98802 5.5213e-05 3.8182 0.012041 9.1314e-06 0.001154 0.11483 0.0006574 0.11549 0.10454 0 0.039402 0.0389 0 0.86882 0.23736 0.062526 0.0088048 4.1457 0.055099 6.5911e-05 0.83497 0.0051533 0.0058905 0.0013933 0.98685 0.99164 3.0053e-06 1.2021e-05 0.13086 0.91677 0.90128 0.0014008 0.98393 0.56962 0.0018871 0.42708 1.7864 1.7854 16.0078 144.9903 0.00018856 -85.6216 0.59021
0.69423 0.98802 5.5213e-05 3.8182 0.012041 9.1445e-06 0.001154 0.11493 0.0006574 0.11558 0.10463 0 0.039395 0.0389 0 0.86888 0.23739 0.062535 0.0088059 4.1459 0.055106 6.592e-05 0.83496 0.0051534 0.0058907 0.0013932 0.98685 0.99165 3.0051e-06 1.202e-05 0.13086 0.91698 0.90138 0.0014008 0.98402 0.56977 0.001887 0.4271 1.787 1.786 16.0078 144.9904 0.0001884 -85.6219 0.59121
0.69523 0.98802 5.5213e-05 3.8182 0.012041 9.1577e-06 0.001154 0.11503 0.0006574 0.11568 0.10472 0 0.039388 0.0389 0 0.86894 0.23742 0.062545 0.0088071 4.1461 0.055113 6.5929e-05 0.83495 0.0051536 0.0058909 0.0013932 0.98685 0.99165 3.0049e-06 1.202e-05 0.13086 0.91719 0.90149 0.0014007 0.9841 0.56992 0.001887 0.42711 1.7876 1.7866 16.0077 144.9904 0.00018823 -85.6222 0.59221
0.69623 0.98802 5.5213e-05 3.8182 0.012041 9.1708e-06 0.001154 0.11512 0.00065741 0.11578 0.10481 0 0.039381 0.0389 0 0.869 0.23744 0.062554 0.0088083 4.1462 0.05512 6.5938e-05 0.83495 0.0051538 0.0058911 0.0013931 0.98686 0.99165 3.0047e-06 1.2019e-05 0.13086 0.91739 0.90159 0.0014007 0.98419 0.57007 0.0018869 0.42712 1.7882 1.7873 16.0077 144.9904 0.00018807 -85.6226 0.59321
0.69723 0.98802 5.5213e-05 3.8182 0.012041 9.184e-06 0.001154 0.11522 0.00065741 0.11587 0.1049 0 0.039374 0.0389 0 0.86906 0.23747 0.062564 0.0088094 4.1464 0.055127 6.5946e-05 0.83494 0.005154 0.0058912 0.001393 0.98686 0.99165 3.0046e-06 1.2018e-05 0.13086 0.9176 0.9017 0.0014006 0.98427 0.57022 0.0018869 0.42714 1.7888 1.7879 16.0077 144.9904 0.0001879 -85.6229 0.59421
0.69823 0.98802 5.5213e-05 3.8182 0.012041 9.1971e-06 0.001154 0.11532 0.00065741 0.11597 0.10499 0 0.039367 0.0389 0 0.86912 0.23749 0.062573 0.0088106 4.1465 0.055134 6.5955e-05 0.83493 0.0051542 0.0058914 0.0013929 0.98686 0.99165 3.0044e-06 1.2017e-05 0.13086 0.91781 0.9018 0.0014006 0.98436 0.57036 0.0018868 0.42715 1.7894 1.7885 16.0077 144.9904 0.00018774 -85.6232 0.59521
0.69923 0.98802 5.5213e-05 3.8182 0.012041 9.2103e-06 0.001154 0.11541 0.00065742 0.11607 0.10507 0 0.039361 0.0389 0 0.86918 0.23752 0.062582 0.0088118 4.1467 0.055141 6.5964e-05 0.83492 0.0051544 0.0058916 0.0013929 0.98686 0.99165 3.0042e-06 1.2017e-05 0.13087 0.91801 0.9019 0.0014006 0.98444 0.57051 0.0018868 0.42716 1.79 1.7891 16.0077 144.9905 0.00018758 -85.6235 0.59621
0.70023 0.98802 5.5213e-05 3.8182 0.012041 9.2235e-06 0.001154 0.11551 0.00065742 0.11616 0.10516 0 0.039354 0.0389 0 0.86924 0.23755 0.062592 0.008813 4.1469 0.055148 6.5973e-05 0.83492 0.0051546 0.0058918 0.0013928 0.98686 0.99165 3.004e-06 1.2016e-05 0.13087 0.91822 0.90201 0.0014005 0.98452 0.57066 0.0018867 0.42717 1.7906 1.7897 16.0076 144.9905 0.00018742 -85.6239 0.59721
0.70123 0.98802 5.5213e-05 3.8182 0.012041 9.2366e-06 0.001154 0.11561 0.00065742 0.11626 0.10525 0 0.039347 0.0389 0 0.8693 0.23757 0.062601 0.0088141 4.147 0.055155 6.5982e-05 0.83491 0.0051548 0.005892 0.0013927 0.98686 0.99165 3.0039e-06 1.2015e-05 0.13087 0.91842 0.90211 0.0014005 0.98461 0.57081 0.0018867 0.42719 1.7912 1.7903 16.0076 144.9905 0.00018725 -85.6242 0.59821
0.70223 0.98802 5.5213e-05 3.8182 0.012041 9.2498e-06 0.001154 0.1157 0.00065743 0.11636 0.10534 0 0.03934 0.0389 0 0.86936 0.2376 0.062611 0.0088153 4.1472 0.055162 6.5991e-05 0.8349 0.005155 0.0058922 0.0013926 0.98686 0.99165 3.0037e-06 1.2015e-05 0.13087 0.91862 0.90221 0.0014004 0.98469 0.57096 0.0018866 0.4272 1.7918 1.7909 16.0076 144.9905 0.00018709 -85.6245 0.59921
0.70323 0.98802 5.5213e-05 3.8182 0.012041 9.2629e-06 0.001154 0.1158 0.00065743 0.11645 0.10543 0 0.039333 0.0389 0 0.86942 0.23762 0.06262 0.0088165 4.1474 0.055169 6.6e-05 0.8349 0.0051551 0.0058924 0.0013926 0.98686 0.99165 3.0035e-06 1.2014e-05 0.13087 0.91883 0.90231 0.0014004 0.98477 0.57111 0.0018866 0.42721 1.7924 1.7915 16.0076 144.9905 0.00018693 -85.6248 0.60021
0.70423 0.98802 5.5213e-05 3.8182 0.012041 9.2761e-06 0.001154 0.1159 0.00065743 0.11655 0.10552 0 0.039326 0.0389 0 0.86947 0.23765 0.06263 0.0088177 4.1475 0.055176 6.6009e-05 0.83489 0.0051553 0.0058926 0.0013925 0.98686 0.99165 3.0034e-06 1.2013e-05 0.13087 0.91903 0.90241 0.0014004 0.98485 0.57126 0.0018865 0.42723 1.793 1.7921 16.0076 144.9906 0.00018677 -85.6251 0.60121
0.70523 0.98802 5.5213e-05 3.8182 0.012041 9.2892e-06 0.001154 0.11599 0.00065743 0.11664 0.10561 0 0.039319 0.0389 0 0.86953 0.23768 0.062639 0.0088189 4.1477 0.055183 6.6017e-05 0.83488 0.0051555 0.0058927 0.0013924 0.98686 0.99165 3.0032e-06 1.2013e-05 0.13088 0.91923 0.90252 0.0014003 0.98493 0.57141 0.0018865 0.42724 1.7936 1.7927 16.0075 144.9906 0.00018661 -85.6254 0.60221
0.70623 0.98802 5.5213e-05 3.8182 0.012041 9.3024e-06 0.001154 0.11609 0.00065744 0.11674 0.1057 0 0.039312 0.0389 0 0.86959 0.2377 0.062649 0.00882 4.1478 0.05519 6.6026e-05 0.83488 0.0051557 0.0058929 0.0013923 0.98687 0.99165 3.003e-06 1.2012e-05 0.13088 0.91943 0.90262 0.0014003 0.98501 0.57156 0.0018864 0.42725 1.7942 1.7933 16.0075 144.9906 0.00018646 -85.6258 0.60321
0.70723 0.98802 5.5212e-05 3.8182 0.012041 9.3156e-06 0.001154 0.11618 0.00065744 0.11684 0.10579 0 0.039305 0.0389 0 0.86965 0.23773 0.062658 0.0088212 4.148 0.055197 6.6035e-05 0.83487 0.0051559 0.0058931 0.0013923 0.98687 0.99165 3.0029e-06 1.2011e-05 0.13088 0.91963 0.90272 0.0014002 0.98509 0.57171 0.0018864 0.42727 1.7948 1.7939 16.0075 144.9906 0.0001863 -85.6261 0.60421
0.70823 0.98802 5.5212e-05 3.8182 0.012041 9.3287e-06 0.0011541 0.11628 0.00065744 0.11693 0.10588 0 0.039298 0.0389 0 0.86971 0.23776 0.062668 0.0088224 4.1482 0.055204 6.6044e-05 0.83486 0.0051561 0.0058933 0.0013922 0.98687 0.99165 3.0027e-06 1.2011e-05 0.13088 0.91983 0.90282 0.0014002 0.98517 0.57186 0.0018863 0.42728 1.7954 1.7945 16.0075 144.9906 0.00018614 -85.6264 0.60521
0.70923 0.98802 5.5212e-05 3.8182 0.012041 9.3419e-06 0.0011541 0.11637 0.00065745 0.11703 0.10597 0 0.039291 0.0389 0 0.86977 0.23778 0.062677 0.0088236 4.1483 0.055211 6.6053e-05 0.83486 0.0051563 0.0058935 0.0013921 0.98687 0.99165 3.0026e-06 1.201e-05 0.13088 0.92003 0.90292 0.0014002 0.98524 0.57201 0.0018863 0.42729 1.796 1.7951 16.0075 144.9907 0.00018598 -85.6267 0.60621
0.71023 0.98802 5.5212e-05 3.8182 0.012041 9.355e-06 0.0011541 0.11647 0.00065745 0.11712 0.10605 0 0.039284 0.0389 0 0.86983 0.23781 0.062687 0.0088248 4.1485 0.055218 6.6062e-05 0.83485 0.0051565 0.0058937 0.0013921 0.98687 0.99166 3.0024e-06 1.2009e-05 0.13088 0.92023 0.90302 0.0014001 0.98532 0.57215 0.0018862 0.4273 1.7966 1.7956 16.0074 144.9907 0.00018583 -85.627 0.60721
0.71123 0.98802 5.5212e-05 3.8182 0.012041 9.3682e-06 0.0011541 0.11657 0.00065745 0.11722 0.10614 0 0.039277 0.0389 0 0.86989 0.23784 0.062696 0.008826 4.1487 0.055225 6.6071e-05 0.83484 0.0051567 0.0058939 0.001392 0.98687 0.99166 3.0022e-06 1.2009e-05 0.13089 0.92043 0.90312 0.0014001 0.9854 0.5723 0.0018862 0.42732 1.7972 1.7962 16.0074 144.9907 0.00018567 -85.6273 0.60821
0.71223 0.98802 5.5212e-05 3.8182 0.012041 9.3813e-06 0.0011541 0.11666 0.00065746 0.11731 0.10623 0 0.039271 0.0389 0 0.86995 0.23786 0.062706 0.0088271 4.1488 0.055232 6.608e-05 0.83483 0.0051569 0.0058941 0.0013919 0.98687 0.99166 3.0021e-06 1.2008e-05 0.13089 0.92062 0.90321 0.0014001 0.98547 0.57245 0.0018861 0.42733 1.7977 1.7968 16.0074 144.9907 0.00018552 -85.6276 0.60921
0.71323 0.98802 5.5212e-05 3.8182 0.012041 9.3945e-06 0.0011541 0.11676 0.00065746 0.11741 0.10632 0 0.039264 0.0389 0 0.87001 0.23789 0.062715 0.0088283 4.149 0.055239 6.6089e-05 0.83483 0.0051571 0.0058943 0.0013919 0.98687 0.99166 3.0019e-06 1.2008e-05 0.13089 0.92082 0.90331 0.0014 0.98555 0.5726 0.0018861 0.42734 1.7983 1.7974 16.0074 144.9907 0.00018536 -85.6279 0.61021
0.71423 0.98802 5.5212e-05 3.8182 0.012041 9.4076e-06 0.0011541 0.11685 0.00065746 0.1175 0.10641 0 0.039257 0.0389 0 0.87007 0.23791 0.062725 0.0088295 4.1492 0.055246 6.6098e-05 0.83482 0.0051573 0.0058945 0.0013918 0.98687 0.99166 3.0018e-06 1.2007e-05 0.13089 0.92101 0.90341 0.0014 0.98563 0.57275 0.001886 0.42736 1.7989 1.798 16.0073 144.9908 0.00018521 -85.6282 0.61121
0.71523 0.98802 5.5212e-05 3.8182 0.012041 9.4208e-06 0.0011541 0.11695 0.00065747 0.1176 0.1065 0 0.03925 0.0389 0 0.87013 0.23794 0.062734 0.0088307 4.1493 0.055253 6.6107e-05 0.83481 0.0051575 0.0058947 0.0013917 0.98687 0.99166 3.0016e-06 1.2006e-05 0.13089 0.92121 0.90351 0.0014 0.9857 0.5729 0.001886 0.42737 1.7995 1.7986 16.0073 144.9908 0.00018505 -85.6284 0.61221
0.71623 0.98802 5.5212e-05 3.8182 0.012041 9.434e-06 0.0011541 0.11704 0.00065747 0.11769 0.10658 0 0.039243 0.0389 0 0.87019 0.23797 0.062744 0.0088319 4.1495 0.05526 6.6116e-05 0.83481 0.0051577 0.0058949 0.0013917 0.98687 0.99166 3.0015e-06 1.2006e-05 0.13089 0.9214 0.90361 0.0013999 0.98577 0.57305 0.0018859 0.42738 1.8001 1.7992 16.0073 144.9908 0.0001849 -85.6287 0.61321
0.71723 0.98802 5.5212e-05 3.8182 0.012041 9.4471e-06 0.0011541 0.11714 0.00065747 0.11779 0.10667 0 0.039236 0.0389 0 0.87025 0.23799 0.062753 0.0088331 4.1497 0.055267 6.6125e-05 0.8348 0.0051579 0.0058951 0.0013916 0.98688 0.99166 3.0013e-06 1.2005e-05 0.1309 0.9216 0.9037 0.0013999 0.98585 0.5732 0.0018859 0.4274 1.8006 1.7997 16.0073 144.9908 0.00018475 -85.629 0.61421
0.71823 0.98802 5.5212e-05 3.8182 0.01204 9.4603e-06 0.0011541 0.11723 0.00065747 0.11788 0.10676 0 0.03923 0.0389 0 0.87031 0.23802 0.062763 0.0088343 4.1498 0.055274 6.6134e-05 0.83479 0.0051581 0.0058953 0.0013915 0.98688 0.99166 3.0012e-06 1.2005e-05 0.1309 0.92179 0.9038 0.0013998 0.98592 0.57334 0.0018858 0.42741 1.8012 1.8003 16.0073 144.9909 0.0001846 -85.6293 0.61521
0.71923 0.98802 5.5212e-05 3.8182 0.01204 9.4734e-06 0.0011541 0.11733 0.00065748 0.11798 0.10685 0 0.039223 0.0389 0 0.87037 0.23805 0.062773 0.0088355 4.15 0.055281 6.6143e-05 0.83478 0.0051583 0.0058955 0.0013915 0.98688 0.99166 3.001e-06 1.2004e-05 0.1309 0.92198 0.9039 0.0013998 0.986 0.57349 0.0018858 0.42742 1.8018 1.8009 16.0072 144.9909 0.00018445 -85.6296 0.61621
0.72023 0.98802 5.5212e-05 3.8182 0.01204 9.4866e-06 0.0011541 0.11742 0.00065748 0.11807 0.10694 0 0.039216 0.0389 0 0.87043 0.23807 0.062782 0.0088367 4.1502 0.055289 6.6152e-05 0.83478 0.0051585 0.0058957 0.0013914 0.98688 0.99166 3.0009e-06 1.2003e-05 0.1309 0.92218 0.90399 0.0013998 0.98607 0.57364 0.0018857 0.42744 1.8024 1.8015 16.0072 144.9909 0.00018429 -85.6299 0.61721
0.72123 0.98802 5.5212e-05 3.8182 0.01204 9.4997e-06 0.0011541 0.11752 0.00065748 0.11817 0.10703 0 0.039209 0.0389 0 0.87049 0.2381 0.062792 0.0088379 4.1504 0.055296 6.6161e-05 0.83477 0.0051587 0.0058959 0.0013913 0.98688 0.99166 3.0007e-06 1.2003e-05 0.1309 0.92237 0.90409 0.0013997 0.98614 0.57379 0.0018857 0.42745 1.8029 1.802 16.0072 144.9909 0.00018414 -85.6302 0.61821
0.72223 0.98802 5.5212e-05 3.8182 0.01204 9.5129e-06 0.0011541 0.11761 0.00065749 0.11826 0.10711 0 0.039202 0.0389 0 0.87055 0.23813 0.062801 0.0088391 4.1505 0.055303 6.617e-05 0.83476 0.0051589 0.005896 0.0013913 0.98688 0.99166 3.0006e-06 1.2002e-05 0.1309 0.92256 0.90418 0.0013997 0.98621 0.57394 0.0018857 0.42746 1.8035 1.8026 16.0072 144.9909 0.000184 -85.6304 0.61921
0.72323 0.98802 5.5212e-05 3.8182 0.01204 9.5261e-06 0.0011541 0.11771 0.00065749 0.11836 0.1072 0 0.039196 0.0389 0 0.87061 0.23815 0.062811 0.0088403 4.1507 0.05531 6.6179e-05 0.83476 0.005159 0.0058962 0.0013912 0.98688 0.99166 3.0004e-06 1.2002e-05 0.13091 0.92275 0.90428 0.0013997 0.98628 0.57408 0.0018856 0.42747 1.8041 1.8032 16.0072 144.991 0.00018385 -85.6307 0.62021
0.72423 0.98802 5.5211e-05 3.8182 0.01204 9.5392e-06 0.0011541 0.1178 0.00065749 0.11845 0.10729 0 0.039189 0.0389 0 0.87067 0.23818 0.062821 0.0088415 4.1509 0.055317 6.6188e-05 0.83475 0.0051592 0.0058964 0.0013911 0.98688 0.99166 3.0003e-06 1.2001e-05 0.13091 0.92294 0.90437 0.0013996 0.98635 0.57423 0.0018856 0.42749 1.8047 1.8038 16.0071 144.991 0.0001837 -85.631 0.62121
0.72523 0.98802 5.5211e-05 3.8182 0.01204 9.5524e-06 0.0011541 0.11789 0.0006575 0.11855 0.10738 0 0.039182 0.0389 0 0.87073 0.23821 0.06283 0.0088427 4.151 0.055324 6.6198e-05 0.83474 0.0051594 0.0058966 0.0013911 0.98688 0.99166 3.0001e-06 1.2e-05 0.13091 0.92313 0.90447 0.0013996 0.98642 0.57438 0.0018855 0.4275 1.8052 1.8043 16.0071 144.991 0.00018355 -85.6313 0.62221
0.72623 0.98802 5.5211e-05 3.8182 0.01204 9.5655e-06 0.0011541 0.11799 0.0006575 0.11864 0.10746 0 0.039175 0.0389 0 0.87079 0.23823 0.06284 0.0088439 4.1512 0.055331 6.6207e-05 0.83473 0.0051596 0.0058968 0.001391 0.98688 0.99166 3e-06 1.2e-05 0.13091 0.92332 0.90456 0.0013996 0.98649 0.57453 0.0018855 0.42751 1.8058 1.8049 16.0071 144.991 0.0001834 -85.6315 0.62321
0.72723 0.98802 5.5211e-05 3.8182 0.01204 9.5787e-06 0.0011541 0.11808 0.0006575 0.11874 0.10755 0 0.039168 0.0389 0 0.87085 0.23826 0.062849 0.0088451 4.1514 0.055338 6.6216e-05 0.83473 0.0051598 0.005897 0.0013909 0.98688 0.99166 2.9998e-06 1.1999e-05 0.13091 0.92351 0.90465 0.0013995 0.98656 0.57468 0.0018854 0.42753 1.8064 1.8055 16.0071 144.991 0.00018325 -85.6318 0.62421
0.72823 0.98802 5.5211e-05 3.8182 0.01204 9.5918e-06 0.0011541 0.11818 0.0006575 0.11883 0.10764 0 0.039162 0.0389 0 0.87092 0.23829 0.062859 0.0088463 4.1516 0.055346 6.6225e-05 0.83472 0.0051601 0.0058972 0.0013909 0.98688 0.99167 2.9997e-06 1.1999e-05 0.13091 0.92369 0.90475 0.0013995 0.98663 0.57483 0.0018854 0.42754 1.8069 1.806 16.007 144.9911 0.00018311 -85.6321 0.62521
0.72923 0.98802 5.5211e-05 3.8182 0.01204 9.605e-06 0.0011541 0.11827 0.00065751 0.11892 0.10773 0 0.039155 0.0389 0 0.87098 0.23831 0.062869 0.0088475 4.1517 0.055353 6.6234e-05 0.83471 0.0051603 0.0058974 0.0013908 0.98688 0.99167 2.9996e-06 1.1998e-05 0.13092 0.92388 0.90484 0.0013995 0.9867 0.57497 0.0018854 0.42755 1.8075 1.8066 16.007 144.9911 0.00018296 -85.6323 0.62621
0.73023 0.98802 5.5211e-05 3.8182 0.01204 9.6181e-06 0.0011541 0.11837 0.00065751 0.11902 0.10781 0 0.039148 0.0389 0 0.87104 0.23834 0.062878 0.0088487 4.1519 0.05536 6.6243e-05 0.83471 0.0051605 0.0058976 0.0013908 0.98689 0.99167 2.9994e-06 1.1998e-05 0.13092 0.92407 0.90493 0.0013994 0.98677 0.57512 0.0018853 0.42756 1.808 1.8072 16.007 144.9911 0.00018282 -85.6326 0.62721
0.73123 0.98802 5.5211e-05 3.8182 0.01204 9.6313e-06 0.0011541 0.11846 0.00065751 0.11911 0.1079 0 0.039142 0.0389 0 0.8711 0.23837 0.062888 0.0088499 4.1521 0.055367 6.6252e-05 0.8347 0.0051607 0.0058978 0.0013907 0.98689 0.99167 2.9993e-06 1.1997e-05 0.13092 0.92425 0.90503 0.0013994 0.98684 0.57527 0.0018853 0.42758 1.8086 1.8077 16.007 144.9911 0.00018267 -85.6328 0.62821
0.73223 0.98802 5.5211e-05 3.8182 0.01204 9.6444e-06 0.0011541 0.11855 0.00065752 0.11921 0.10799 0 0.039135 0.0389 0 0.87116 0.23839 0.062898 0.0088511 4.1522 0.055374 6.6261e-05 0.83469 0.0051609 0.005898 0.0013906 0.98689 0.99167 2.9991e-06 1.1996e-05 0.13092 0.92444 0.90512 0.0013994 0.9869 0.57542 0.0018852 0.42759 1.8092 1.8083 16.007 144.9911 0.00018253 -85.6331 0.62921
0.73323 0.98802 5.5211e-05 3.8182 0.01204 9.6576e-06 0.0011541 0.11865 0.00065752 0.1193 0.10807 0 0.039128 0.0389 0 0.87122 0.23842 0.062908 0.0088523 4.1524 0.055381 6.6271e-05 0.83468 0.0051611 0.0058982 0.0013906 0.98689 0.99167 2.999e-06 1.1996e-05 0.13092 0.92462 0.90521 0.0013994 0.98697 0.57556 0.0018852 0.4276 1.8097 1.8088 16.0069 144.9912 0.00018238 -85.6334 0.63021
0.73423 0.98802 5.5211e-05 3.8182 0.01204 9.6708e-06 0.0011541 0.11874 0.00065752 0.11939 0.10816 0 0.039121 0.0389 0 0.87128 0.23845 0.062917 0.0088535 4.1526 0.055389 6.628e-05 0.83468 0.0051613 0.0058984 0.0013905 0.98689 0.99167 2.9989e-06 1.1995e-05 0.13092 0.92481 0.9053 0.0013993 0.98704 0.57571 0.0018851 0.42762 1.8103 1.8094 16.0069 144.9912 0.00018224 -85.6336 0.63121
0.73523 0.98802 5.5211e-05 3.8182 0.01204 9.6839e-06 0.0011541 0.11883 0.00065752 0.11949 0.10825 0 0.039115 0.0389 0 0.87134 0.23848 0.062927 0.0088547 4.1528 0.055396 6.6289e-05 0.83467 0.0051615 0.0058987 0.0013905 0.98689 0.99167 2.9987e-06 1.1995e-05 0.13093 0.92499 0.90539 0.0013993 0.9871 0.57586 0.0018851 0.42763 1.8108 1.81 16.0069 144.9912 0.0001821 -85.6339 0.63221
0.73623 0.98802 5.5211e-05 3.8182 0.01204 9.6971e-06 0.0011541 0.11893 0.00065753 0.11958 0.10834 0 0.039108 0.0389 0 0.8714 0.2385 0.062937 0.0088559 4.1529 0.055403 6.6298e-05 0.83466 0.0051617 0.0058989 0.0013904 0.98689 0.99167 2.9986e-06 1.1994e-05 0.13093 0.92517 0.90548 0.0013993 0.98717 0.57601 0.0018851 0.42764 1.8114 1.8105 16.0069 144.9912 0.00018195 -85.6341 0.63321
0.73723 0.98802 5.5211e-05 3.8182 0.01204 9.7102e-06 0.0011541 0.11902 0.00065753 0.11967 0.10842 0 0.039101 0.0389 0 0.87146 0.23853 0.062946 0.0088571 4.1531 0.05541 6.6307e-05 0.83466 0.0051619 0.0058991 0.0013903 0.98689 0.99167 2.9985e-06 1.1994e-05 0.13093 0.92536 0.90557 0.0013992 0.98723 0.57615 0.001885 0.42766 1.8119 1.8111 16.0068 144.9912 0.00018181 -85.6344 0.63421
0.73823 0.98802 5.5211e-05 3.8182 0.01204 9.7234e-06 0.0011541 0.11911 0.00065753 0.11977 0.10851 0 0.039095 0.0389 0 0.87152 0.23856 0.062956 0.0088584 4.1533 0.055417 6.6317e-05 0.83465 0.0051621 0.0058993 0.0013903 0.98689 0.99167 2.9983e-06 1.1993e-05 0.13093 0.92554 0.90566 0.0013992 0.9873 0.5763 0.001885 0.42767 1.8125 1.8116 16.0068 144.9913 0.00018167 -85.6346 0.63521
0.73923 0.98802 5.5211e-05 3.8182 0.01204 9.7365e-06 0.0011541 0.11921 0.00065754 0.11986 0.1086 0 0.039088 0.0389 0 0.87159 0.23858 0.062966 0.0088596 4.1535 0.055425 6.6326e-05 0.83464 0.0051623 0.0058995 0.0013902 0.98689 0.99167 2.9982e-06 1.1993e-05 0.13093 0.92572 0.90575 0.0013992 0.98736 0.57645 0.0018849 0.42768 1.813 1.8122 16.0068 144.9913 0.00018153 -85.6349 0.63621
0.74023 0.98802 5.521e-05 3.8182 0.01204 9.7497e-06 0.0011541 0.1193 0.00065754 0.11995 0.10868 0 0.039081 0.0389 0 0.87165 0.23861 0.062976 0.0088608 4.1537 0.055432 6.6335e-05 0.83463 0.0051625 0.0058997 0.0013902 0.98689 0.99167 2.9981e-06 1.1992e-05 0.13093 0.9259 0.90584 0.0013991 0.98743 0.5766 0.0018849 0.42769 1.8136 1.8127 16.0068 144.9913 0.00018139 -85.6351 0.63721
0.74123 0.98802 5.521e-05 3.8182 0.01204 9.7628e-06 0.0011541 0.11939 0.00065754 0.12005 0.10877 0 0.039075 0.0389 0 0.87171 0.23864 0.062985 0.008862 4.1538 0.055439 6.6344e-05 0.83463 0.0051627 0.0058999 0.0013901 0.98689 0.99167 2.9979e-06 1.1992e-05 0.13094 0.92608 0.90593 0.0013991 0.98749 0.57674 0.0018849 0.42771 1.8141 1.8133 16.0067 144.9913 0.00018125 -85.6354 0.63821
0.74223 0.98802 5.521e-05 3.8182 0.01204 9.776e-06 0.0011541 0.11949 0.00065754 0.12014 0.10886 0 0.039068 0.0389 0 0.87177 0.23866 0.062995 0.0088632 4.154 0.055446 6.6353e-05 0.83462 0.0051629 0.0059001 0.0013901 0.98689 0.99167 2.9978e-06 1.1991e-05 0.13094 0.92626 0.90602 0.0013991 0.98755 0.57689 0.0018848 0.42772 1.8147 1.8138 16.0067 144.9913 0.00018111 -85.6356 0.63921
0.74323 0.98802 5.521e-05 3.8182 0.01204 9.7892e-06 0.0011541 0.11958 0.00065755 0.12023 0.10894 0 0.039061 0.0389 0 0.87183 0.23869 0.063005 0.0088644 4.1542 0.055454 6.6363e-05 0.83461 0.0051631 0.0059003 0.00139 0.9869 0.99167 2.9977e-06 1.1991e-05 0.13094 0.92644 0.90611 0.001399 0.98761 0.57704 0.0018848 0.42773 1.8152 1.8144 16.0067 144.9914 0.00018097 -85.6359 0.64021
0.74423 0.98802 5.521e-05 3.8182 0.01204 9.8023e-06 0.0011541 0.11967 0.00065755 0.12033 0.10903 0 0.039055 0.0389 0 0.87189 0.23872 0.063015 0.0088656 4.1544 0.055461 6.6372e-05 0.83461 0.0051633 0.0059005 0.0013899 0.9869 0.99167 2.9975e-06 1.199e-05 0.13094 0.92662 0.9062 0.001399 0.98768 0.57719 0.0018848 0.42775 1.8158 1.8149 16.0067 144.9914 0.00018083 -85.6361 0.64121
0.74523 0.98802 5.521e-05 3.8182 0.01204 9.8155e-06 0.0011541 0.11977 0.00065755 0.12042 0.10911 0 0.039048 0.0389 0 0.87195 0.23875 0.063025 0.0088669 4.1545 0.055468 6.6381e-05 0.8346 0.0051635 0.0059007 0.0013899 0.9869 0.99167 2.9974e-06 1.199e-05 0.13094 0.92679 0.90628 0.001399 0.98774 0.57733 0.0018847 0.42776 1.8163 1.8155 16.0067 144.9914 0.0001807 -85.6363 0.64221
0.74623 0.98802 5.521e-05 3.8182 0.01204 9.8286e-06 0.0011541 0.11986 0.00065756 0.12051 0.1092 0 0.039042 0.0389 0 0.87201 0.23877 0.063034 0.0088681 4.1547 0.055475 6.639e-05 0.83459 0.0051637 0.0059009 0.0013898 0.9869 0.99167 2.9973e-06 1.1989e-05 0.13094 0.92697 0.90637 0.001399 0.9878 0.57748 0.0018847 0.42777 1.8168 1.816 16.0066 144.9914 0.00018056 -85.6366 0.64321
0.74723 0.98802 5.521e-05 3.8182 0.01204 9.8418e-06 0.0011541 0.11995 0.00065756 0.12061 0.10929 0 0.039035 0.0389 0 0.87208 0.2388 0.063044 0.0088693 4.1549 0.055483 6.64e-05 0.83458 0.0051639 0.0059011 0.0013898 0.9869 0.99167 2.9972e-06 1.1989e-05 0.13095 0.92715 0.90646 0.0013989 0.98786 0.57763 0.0018846 0.42778 1.8174 1.8165 16.0066 144.9914 0.00018042 -85.6368 0.64421
0.74823 0.98802 5.521e-05 3.8182 0.01204 9.8549e-06 0.0011541 0.12005 0.00065756 0.1207 0.10937 0 0.039028 0.0389 0 0.87214 0.23883 0.063054 0.0088705 4.1551 0.05549 6.6409e-05 0.83458 0.0051642 0.0059013 0.0013897 0.9869 0.99167 2.997e-06 1.1988e-05 0.13095 0.92732 0.90654 0.0013989 0.98792 0.57777 0.0018846 0.4278 1.8179 1.8171 16.0066 144.9915 0.00018029 -85.637 0.64521
0.74923 0.98802 5.521e-05 3.8182 0.01204 9.8681e-06 0.0011541 0.12014 0.00065756 0.12079 0.10946 0 0.039022 0.0389 0 0.8722 0.23885 0.063064 0.0088718 4.1553 0.055497 6.6418e-05 0.83457 0.0051644 0.0059015 0.0013897 0.9869 0.99168 2.9969e-06 1.1988e-05 0.13095 0.9275 0.90663 0.0013989 0.98798 0.57792 0.0018846 0.42781 1.8185 1.8176 16.0066 144.9915 0.00018015 -85.6373 0.64621
0.75023 0.98802 5.521e-05 3.8182 0.01204 9.8812e-06 0.0011541 0.12023 0.00065757 0.12088 0.10955 0 0.039015 0.0389 0 0.87226 0.23888 0.063074 0.008873 4.1554 0.055504 6.6428e-05 0.83456 0.0051646 0.0059017 0.0013896 0.9869 0.99168 2.9968e-06 1.1987e-05 0.13095 0.92767 0.90672 0.0013988 0.98804 0.57807 0.0018845 0.42782 1.819 1.8182 16.0065 144.9915 0.00018001 -85.6375 0.64721
0.75123 0.98802 5.521e-05 3.8182 0.01204 9.8944e-06 0.0011541 0.12032 0.00065757 0.12098 0.10963 0 0.039009 0.0389 0 0.87232 0.23891 0.063083 0.0088742 4.1556 0.055512 6.6437e-05 0.83455 0.0051648 0.0059019 0.0013896 0.9869 0.99168 2.9967e-06 1.1987e-05 0.13095 0.92785 0.9068 0.0013988 0.9881 0.57821 0.0018845 0.42784 1.8195 1.8187 16.0065 144.9915 0.00017988 -85.6377 0.64821
0.75223 0.98802 5.521e-05 3.8182 0.01204 9.9075e-06 0.0011541 0.12042 0.00065757 0.12107 0.10972 0 0.039002 0.0389 0 0.87238 0.23894 0.063093 0.0088754 4.1558 0.055519 6.6446e-05 0.83455 0.005165 0.0059022 0.0013895 0.9869 0.99168 2.9966e-06 1.1986e-05 0.13095 0.92802 0.90689 0.0013988 0.98816 0.57836 0.0018845 0.42785 1.8201 1.8192 16.0065 144.9915 0.00017974 -85.638 0.64921
0.75323 0.98802 5.521e-05 3.8182 0.01204 9.9207e-06 0.0011541 0.12051 0.00065758 0.12116 0.1098 0 0.038995 0.0389 0 0.87245 0.23896 0.063103 0.0088767 4.156 0.055526 6.6456e-05 0.83454 0.0051652 0.0059024 0.0013895 0.9869 0.99168 2.9964e-06 1.1986e-05 0.13096 0.9282 0.90697 0.0013988 0.98822 0.57851 0.0018844 0.42786 1.8206 1.8198 16.0065 144.9916 0.00017961 -85.6382 0.65021
0.75423 0.98802 5.521e-05 3.8182 0.01204 9.9339e-06 0.0011541 0.1206 0.00065758 0.12125 0.10989 0 0.038989 0.0389 0 0.87251 0.23899 0.063113 0.0088779 4.1562 0.055534 6.6465e-05 0.83453 0.0051654 0.0059026 0.0013894 0.9869 0.99168 2.9963e-06 1.1985e-05 0.13096 0.92837 0.90706 0.0013987 0.98828 0.57865 0.0018844 0.42788 1.8211 1.8203 16.0064 144.9916 0.00017948 -85.6384 0.65121
0.75523 0.98802 5.521e-05 3.8182 0.01204 9.947e-06 0.0011541 0.12069 0.00065758 0.12134 0.10997 0 0.038982 0.0389 0 0.87257 0.23902 0.063123 0.0088791 4.1564 0.055541 6.6474e-05 0.83453 0.0051656 0.0059028 0.0013894 0.9869 0.99168 2.9962e-06 1.1985e-05 0.13096 0.92854 0.90714 0.0013987 0.98833 0.5788 0.0018843 0.42789 1.8217 1.8208 16.0064 144.9916 0.00017934 -85.6386 0.65221
0.75623 0.98802 5.5209e-05 3.8182 0.01204 9.9602e-06 0.0011541 0.12078 0.00065758 0.12144 0.11006 0 0.038976 0.0389 0 0.87263 0.23905 0.063133 0.0088803 4.1565 0.055548 6.6484e-05 0.83452 0.0051658 0.005903 0.0013893 0.9869 0.99168 2.9961e-06 1.1984e-05 0.13096 0.92871 0.90723 0.0013987 0.98839 0.57895 0.0018843 0.4279 1.8222 1.8214 16.0064 144.9916 0.00017921 -85.6389 0.65321
0.75723 0.98802 5.5209e-05 3.8182 0.01204 9.9733e-06 0.0011541 0.12088 0.00065759 0.12153 0.11015 0 0.038969 0.0389 0 0.87269 0.23907 0.063143 0.0088816 4.1567 0.055556 6.6493e-05 0.83451 0.0051661 0.0059032 0.0013893 0.98691 0.99168 2.996e-06 1.1984e-05 0.13096 0.92888 0.90731 0.0013987 0.98845 0.57909 0.0018843 0.42791 1.8227 1.8219 16.0064 144.9916 0.00017908 -85.6391 0.65421
0.75823 0.98802 5.5209e-05 3.8182 0.01204 9.9865e-06 0.0011541 0.12097 0.00065759 0.12162 0.11023 0 0.038963 0.0389 0 0.87276 0.2391 0.063153 0.0088828 4.1569 0.055563 6.6502e-05 0.8345 0.0051663 0.0059034 0.0013892 0.98691 0.99168 2.9959e-06 1.1983e-05 0.13097 0.92906 0.9074 0.0013986 0.9885 0.57924 0.0018842 0.42793 1.8232 1.8224 16.0063 144.9917 0.00017895 -85.6393 0.65521
0.75923 0.98802 5.5209e-05 3.8182 0.01204 9.9996e-06 0.0011541 0.12106 0.00065759 0.12171 0.11032 0 0.038956 0.0389 0 0.87282 0.23913 0.063162 0.008884 4.1571 0.05557 6.6512e-05 0.8345 0.0051665 0.0059036 0.0013892 0.98691 0.99168 2.9957e-06 1.1983e-05 0.13097 0.92923 0.90748 0.0013986 0.98856 0.57939 0.0018842 0.42794 1.8238 1.8229 16.0063 144.9917 0.00017882 -85.6395 0.65621
0.76023 0.98802 5.5209e-05 3.8182 0.01204 1.0013e-05 0.0011541 0.12115 0.00065759 0.1218 0.1104 0 0.03895 0.0389 0 0.87288 0.23916 0.063172 0.0088853 4.1573 0.055578 6.6521e-05 0.83449 0.0051667 0.0059038 0.0013891 0.98691 0.99168 2.9956e-06 1.1982e-05 0.13097 0.9294 0.90756 0.0013986 0.98862 0.57953 0.0018842 0.42795 1.8243 1.8235 16.0063 144.9917 0.00017869 -85.6397 0.65721
0.76123 0.98802 5.5209e-05 3.8182 0.01204 1.0026e-05 0.0011541 0.12124 0.0006576 0.1219 0.11049 0 0.038943 0.0389 0 0.87294 0.23918 0.063182 0.0088865 4.1575 0.055585 6.6531e-05 0.83448 0.0051669 0.0059041 0.0013891 0.98691 0.99168 2.9955e-06 1.1982e-05 0.13097 0.92956 0.90765 0.0013985 0.98867 0.57968 0.0018841 0.42797 1.8248 1.824 16.0063 144.9917 0.00017856 -85.6399 0.65821
0.76223 0.98802 5.5209e-05 3.8182 0.01204 1.0039e-05 0.0011541 0.12134 0.0006576 0.12199 0.11057 0 0.038937 0.0389 0 0.87301 0.23921 0.063192 0.0088877 4.1577 0.055592 6.654e-05 0.83447 0.0051671 0.0059043 0.001389 0.98691 0.99168 2.9954e-06 1.1982e-05 0.13097 0.92973 0.90773 0.0013985 0.98873 0.57983 0.0018841 0.42798 1.8253 1.8245 16.0062 144.9917 0.00017843 -85.6402 0.65921
0.76323 0.98802 5.5209e-05 3.8182 0.01204 1.0052e-05 0.0011541 0.12143 0.0006576 0.12208 0.11066 0 0.03893 0.0389 0 0.87307 0.23924 0.063202 0.008889 4.1578 0.0556 6.6549e-05 0.83447 0.0051673 0.0059045 0.001389 0.98691 0.99168 2.9953e-06 1.1981e-05 0.13097 0.9299 0.90781 0.0013985 0.98878 0.57997 0.0018841 0.42799 1.8259 1.825 16.0062 144.9918 0.0001783 -85.6404 0.66021
0.76423 0.98802 5.5209e-05 3.8182 0.01204 1.0065e-05 0.0011541 0.12152 0.0006576 0.12217 0.11074 0 0.038924 0.0389 0 0.87313 0.23927 0.063212 0.0088902 4.158 0.055607 6.6559e-05 0.83446 0.0051676 0.0059047 0.0013889 0.98691 0.99168 2.9952e-06 1.1981e-05 0.13098 0.93007 0.90789 0.0013985 0.98884 0.58012 0.001884 0.428 1.8264 1.8256 16.0062 144.9918 0.00017817 -85.6406 0.66121
0.76523 0.98802 5.5209e-05 3.8182 0.01204 1.0079e-05 0.0011541 0.12161 0.00065761 0.12226 0.11083 0 0.038917 0.0389 0 0.87319 0.23929 0.063222 0.0088914 4.1582 0.055615 6.6568e-05 0.83445 0.0051678 0.0059049 0.0013889 0.98691 0.99168 2.9951e-06 1.198e-05 0.13098 0.93024 0.90797 0.0013984 0.98889 0.58026 0.001884 0.42802 1.8269 1.8261 16.0062 144.9918 0.00017804 -85.6408 0.66221
0.76623 0.98802 5.5209e-05 3.8182 0.01204 1.0092e-05 0.0011541 0.1217 0.00065761 0.12235 0.11091 0 0.038911 0.0389 0 0.87325 0.23932 0.063232 0.0088927 4.1584 0.055622 6.6578e-05 0.83444 0.005168 0.0059051 0.0013888 0.98691 0.99168 2.995e-06 1.198e-05 0.13098 0.9304 0.90806 0.0013984 0.98895 0.58041 0.001884 0.42803 1.8274 1.8266 16.0061 144.9918 0.00017791 -85.641 0.66321
0.76723 0.98802 5.5209e-05 3.8182 0.01204 1.0105e-05 0.0011541 0.12179 0.00065761 0.12245 0.111 0 0.038904 0.0389 0 0.87332 0.23935 0.063242 0.0088939 4.1586 0.055629 6.6587e-05 0.83444 0.0051682 0.0059053 0.0013888 0.98691 0.99168 2.9948e-06 1.1979e-05 0.13098 0.93057 0.90814 0.0013984 0.989 0.58056 0.0018839 0.42804 1.8279 1.8271 16.0061 144.9918 0.00017778 -85.6412 0.66421
0.76823 0.98802 5.5209e-05 3.8182 0.01204 1.0118e-05 0.0011541 0.12188 0.00065762 0.12254 0.11108 0 0.038898 0.0389 0 0.87338 0.23938 0.063252 0.0088952 4.1588 0.055637 6.6596e-05 0.83443 0.0051684 0.0059056 0.0013887 0.98691 0.99168 2.9947e-06 1.1979e-05 0.13098 0.93073 0.90822 0.0013984 0.98905 0.5807 0.0018839 0.42806 1.8285 1.8276 16.0061 144.9919 0.00017766 -85.6414 0.66521
0.76923 0.98802 5.5209e-05 3.8182 0.01204 1.0131e-05 0.0011541 0.12197 0.00065762 0.12263 0.11117 0 0.038891 0.0389 0 0.87344 0.2394 0.063262 0.0088964 4.159 0.055644 6.6606e-05 0.83442 0.0051686 0.0059058 0.0013887 0.98691 0.99168 2.9946e-06 1.1978e-05 0.13098 0.9309 0.9083 0.0013983 0.98911 0.58085 0.0018839 0.42807 1.829 1.8282 16.0061 144.9919 0.00017753 -85.6416 0.66621
0.77023 0.98802 5.5209e-05 3.8182 0.01204 1.0144e-05 0.0011541 0.12207 0.00065762 0.12272 0.11125 0 0.038885 0.0389 0 0.8735 0.23943 0.063272 0.0088976 4.1592 0.055652 6.6616e-05 0.83442 0.0051689 0.005906 0.0013886 0.98691 0.99168 2.9945e-06 1.1978e-05 0.13099 0.93106 0.90838 0.0013983 0.98916 0.58099 0.0018838 0.42808 1.8295 1.8287 16.0061 144.9919 0.0001774 -85.6418 0.66721
0.77123 0.98802 5.5209e-05 3.8182 0.01204 1.0157e-05 0.0011541 0.12216 0.00065762 0.12281 0.11134 0 0.038879 0.0389 0 0.87357 0.23946 0.063282 0.0088989 4.1593 0.055659 6.6625e-05 0.83441 0.0051691 0.0059062 0.0013886 0.98691 0.99168 2.9944e-06 1.1978e-05 0.13099 0.93123 0.90846 0.0013983 0.98921 0.58114 0.0018838 0.42809 1.83 1.8292 16.006 144.9919 0.00017728 -85.642 0.66821
0.77223 0.98802 5.5208e-05 3.8182 0.01204 1.0171e-05 0.0011541 0.12225 0.00065763 0.1229 0.11142 0 0.038872 0.0389 0 0.87363 0.23949 0.063292 0.0089001 4.1595 0.055666 6.6634e-05 0.8344 0.0051693 0.0059064 0.0013885 0.98691 0.99168 2.9943e-06 1.1977e-05 0.13099 0.93139 0.90854 0.0013983 0.98926 0.58128 0.0018838 0.42811 1.8305 1.8297 16.006 144.9919 0.00017715 -85.6422 0.66921
0.77323 0.98802 5.5208e-05 3.8182 0.01204 1.0184e-05 0.0011541 0.12234 0.00065763 0.12299 0.1115 0 0.038866 0.0389 0 0.87369 0.23952 0.063302 0.0089014 4.1597 0.055674 6.6644e-05 0.83439 0.0051695 0.0059066 0.0013885 0.98692 0.99169 2.9942e-06 1.1977e-05 0.13099 0.93155 0.90862 0.0013982 0.98931 0.58143 0.0018837 0.42812 1.831 1.8302 16.006 144.992 0.00017703 -85.6424 0.67021
0.77423 0.98802 5.5208e-05 3.8182 0.01204 1.0197e-05 0.0011541 0.12243 0.00065763 0.12308 0.11159 0 0.038859 0.0389 0 0.87376 0.23954 0.063312 0.0089026 4.1599 0.055681 6.6653e-05 0.83439 0.0051697 0.0059069 0.0013884 0.98692 0.99169 2.9941e-06 1.1976e-05 0.13099 0.93172 0.9087 0.0013982 0.98936 0.58158 0.0018837 0.42813 1.8315 1.8307 16.006 144.992 0.0001769 -85.6426 0.67121
0.77523 0.98802 5.5208e-05 3.8182 0.01204 1.021e-05 0.0011541 0.12252 0.00065763 0.12317 0.11167 0 0.038853 0.0389 0 0.87382 0.23957 0.063322 0.0089039 4.1601 0.055689 6.6663e-05 0.83438 0.00517 0.0059071 0.0013884 0.98692 0.99169 2.994e-06 1.1976e-05 0.131 0.93188 0.90878 0.0013982 0.98941 0.58172 0.0018837 0.42814 1.832 1.8312 16.0059 144.992 0.00017678 -85.6428 0.67221
0.77623 0.98802 5.5208e-05 3.8182 0.01204 1.0223e-05 0.0011541 0.12261 0.00065764 0.12326 0.11176 0 0.038847 0.0389 0 0.87388 0.2396 0.063332 0.0089051 4.1603 0.055696 6.6672e-05 0.83437 0.0051702 0.0059073 0.0013883 0.98692 0.99169 2.9939e-06 1.1975e-05 0.131 0.93204 0.90886 0.0013982 0.98947 0.58187 0.0018837 0.42816 1.8325 1.8317 16.0059 144.992 0.00017666 -85.643 0.67321
0.77723 0.98802 5.5208e-05 3.8182 0.01204 1.0236e-05 0.0011541 0.1227 0.00065764 0.12335 0.11184 0 0.03884 0.0389 0 0.87394 0.23963 0.063342 0.0089064 4.1605 0.055704 6.6682e-05 0.83436 0.0051704 0.0059075 0.0013883 0.98692 0.99169 2.9938e-06 1.1975e-05 0.131 0.9322 0.90893 0.0013982 0.98952 0.58201 0.0018836 0.42817 1.833 1.8323 16.0059 144.992 0.00017653 -85.6432 0.67421
0.77823 0.98802 5.5208e-05 3.8182 0.01204 1.025e-05 0.0011541 0.12279 0.00065764 0.12344 0.11193 0 0.038834 0.0389 0 0.87401 0.23965 0.063352 0.0089076 4.1607 0.055711 6.6691e-05 0.83436 0.0051706 0.0059077 0.0013883 0.98692 0.99169 2.9937e-06 1.1975e-05 0.131 0.93236 0.90901 0.0013981 0.98957 0.58216 0.0018836 0.42818 1.8335 1.8328 16.0059 144.9921 0.00017641 -85.6434 0.67521
0.77923 0.98802 5.5208e-05 3.8182 0.01204 1.0263e-05 0.0011541 0.12288 0.00065764 0.12354 0.11201 0 0.038827 0.0389 0 0.87407 0.23968 0.063362 0.0089089 4.1609 0.055719 6.6701e-05 0.83435 0.0051708 0.005908 0.0013882 0.98692 0.99169 2.9936e-06 1.1974e-05 0.131 0.93252 0.90909 0.0013981 0.98961 0.5823 0.0018836 0.4282 1.834 1.8333 16.0058 144.9921 0.00017629 -85.6436 0.67621
0.78023 0.98802 5.5208e-05 3.8182 0.01204 1.0276e-05 0.0011541 0.12297 0.00065765 0.12363 0.11209 0 0.038821 0.0389 0 0.87413 0.23971 0.063372 0.0089101 4.1611 0.055726 6.6711e-05 0.83434 0.0051711 0.0059082 0.0013882 0.98692 0.99169 2.9935e-06 1.1974e-05 0.13101 0.93268 0.90917 0.0013981 0.98966 0.58245 0.0018835 0.42821 1.8346 1.8338 16.0058 144.9921 0.00017617 -85.6437 0.67721
0.78123 0.98802 5.5208e-05 3.8182 0.01204 1.0289e-05 0.0011541 0.12306 0.00065765 0.12372 0.11218 0 0.038815 0.0389 0 0.8742 0.23974 0.063382 0.0089114 4.1613 0.055734 6.672e-05 0.83433 0.0051713 0.0059084 0.0013881 0.98692 0.99169 2.9934e-06 1.1973e-05 0.13101 0.93284 0.90924 0.0013981 0.98971 0.58259 0.0018835 0.42822 1.8351 1.8343 16.0058 144.9921 0.00017604 -85.6439 0.67821
0.78223 0.98802 5.5208e-05 3.8182 0.01204 1.0302e-05 0.0011541 0.12315 0.00065765 0.12381 0.11226 0 0.038808 0.0389 0 0.87426 0.23977 0.063392 0.0089126 4.1615 0.055741 6.673e-05 0.83433 0.0051715 0.0059086 0.0013881 0.98692 0.99169 2.9933e-06 1.1973e-05 0.13101 0.933 0.90932 0.001398 0.98976 0.58274 0.0018835 0.42823 1.8356 1.8348 16.0058 144.9922 0.00017592 -85.6441 0.67921
0.78323 0.98802 5.5208e-05 3.8182 0.01204 1.0315e-05 0.0011541 0.12324 0.00065765 0.1239 0.11235 0 0.038802 0.0389 0 0.87432 0.23979 0.063402 0.0089139 4.1616 0.055749 6.674e-05 0.83432 0.0051717 0.0059089 0.001388 0.98692 0.99169 2.9932e-06 1.1973e-05 0.13101 0.93315 0.9094 0.001398 0.98981 0.58288 0.0018834 0.42825 1.8361 1.8353 16.0057 144.9922 0.0001758 -85.6443 0.68021
0.78423 0.98802 5.5208e-05 3.8182 0.01204 1.0328e-05 0.0011541 0.12333 0.00065766 0.12399 0.11243 0 0.038796 0.0389 0 0.87439 0.23982 0.063413 0.0089151 4.1618 0.055756 6.6748e-05 0.83431 0.0051719 0.0059091 0.001388 0.98692 0.99169 2.9931e-06 1.1972e-05 0.13101 0.93331 0.90948 0.001398 0.98986 0.58303 0.0018834 0.42826 1.8365 1.8358 16.0057 144.9922 0.00017568 -85.6445 0.68121
0.78523 0.98802 5.5208e-05 3.8182 0.01204 1.0342e-05 0.0011541 0.12342 0.00065766 0.12408 0.11251 0 0.038789 0.0389 0 0.87445 0.23985 0.063423 0.0089164 4.162 0.055764 6.6758e-05 0.8343 0.0051722 0.0059093 0.001388 0.98692 0.99169 2.993e-06 1.1972e-05 0.13101 0.93347 0.90955 0.001398 0.9899 0.58317 0.0018834 0.42827 1.837 1.8363 16.0057 144.9922 0.00017556 -85.6447 0.68221
0.78623 0.98802 5.5208e-05 3.8182 0.01204 1.0355e-05 0.0011541 0.12351 0.00065766 0.12417 0.1126 0 0.038783 0.0389 0 0.87451 0.23988 0.063433 0.0089176 4.1622 0.055771 6.6769e-05 0.8343 0.0051724 0.0059095 0.0013879 0.98692 0.99169 2.9929e-06 1.1972e-05 0.13102 0.93363 0.90963 0.0013979 0.98995 0.58332 0.0018834 0.42829 1.8375 1.8368 16.0057 144.9922 0.00017544 -85.6448 0.68321
0.78723 0.98802 5.5208e-05 3.8182 0.01204 1.0368e-05 0.0011541 0.1236 0.00065767 0.12426 0.11268 0 0.038777 0.0389 0 0.87458 0.23991 0.063443 0.0089189 4.1624 0.055779 6.6777e-05 0.83429 0.0051726 0.0059097 0.0013879 0.98692 0.99169 2.9928e-06 1.1971e-05 0.13102 0.93378 0.9097 0.0013979 0.99 0.58346 0.0018833 0.4283 1.838 1.8373 16.0056 144.9923 0.00017532 -85.645 0.68421
0.78823 0.98802 5.5207e-05 3.8182 0.01204 1.0381e-05 0.0011541 0.12369 0.00065767 0.12435 0.11276 0 0.03877 0.0389 0 0.87464 0.23993 0.063453 0.0089202 4.1626 0.055786 6.6785e-05 0.83428 0.0051728 0.00591 0.0013878 0.98692 0.99169 2.9927e-06 1.1971e-05 0.13102 0.93394 0.90978 0.0013979 0.99005 0.58361 0.0018833 0.42831 1.8385 1.8378 16.0056 144.9923 0.00017521 -85.6452 0.68521
0.78923 0.98802 5.5207e-05 3.8182 0.01204 1.0394e-05 0.0011541 0.12378 0.00065767 0.12444 0.11285 0 0.038764 0.0389 0 0.8747 0.23996 0.063463 0.0089214 4.1628 0.055794 6.6797e-05 0.83427 0.0051731 0.0059102 0.0013878 0.98692 0.99169 2.9926e-06 1.197e-05 0.13102 0.93409 0.90985 0.0013979 0.99009 0.58375 0.0018833 0.42832 1.839 1.8383 16.0056 144.9923 0.00017509 -85.6454 0.68621
0.79023 0.98802 5.5207e-05 3.8182 0.01204 1.0407e-05 0.0011541 0.12387 0.00065767 0.12453 0.11293 0 0.038758 0.0389 0 0.87477 0.23999 0.063473 0.0089227 4.163 0.055801 6.6807e-05 0.83427 0.0051733 0.0059104 0.0013877 0.98692 0.99169 2.9925e-06 1.197e-05 0.13102 0.93425 0.90993 0.0013979 0.99014 0.5839 0.0018832 0.42834 1.8395 1.8387 16.0056 144.9923 0.00017497 -85.6456 0.68721
0.79123 0.98802 5.5207e-05 3.8182 0.01204 1.0421e-05 0.0011541 0.12396 0.00065768 0.12461 0.11301 0 0.038751 0.0389 0 0.87483 0.24002 0.063483 0.0089239 4.1632 0.055809 6.6815e-05 0.83426 0.0051735 0.0059106 0.0013877 0.98692 0.99169 2.9924e-06 1.197e-05 0.13103 0.9344 0.91 0.0013978 0.99018 0.58404 0.0018832 0.42835 1.84 1.8392 16.0055 144.9923 0.00017485 -85.6457 0.68821
0.79223 0.98802 5.5207e-05 3.8182 0.012039 1.0434e-05 0.0011541 0.12405 0.00065768 0.1247 0.1131 0 0.038745 0.0389 0 0.8749 0.24005 0.063494 0.0089252 4.1634 0.055816 6.6826e-05 0.83425 0.0051738 0.0059109 0.0013877 0.98693 0.99169 2.9923e-06 1.1969e-05 0.13103 0.93455 0.91008 0.0013978 0.99023 0.58419 0.0018832 0.42836 1.8405 1.8397 16.0055 144.9924 0.00017474 -85.6459 0.68921
0.79323 0.98802 5.5207e-05 3.8182 0.012039 1.0447e-05 0.0011541 0.12414 0.00065768 0.12479 0.11318 0 0.038739 0.0389 0 0.87496 0.24007 0.063504 0.0089265 4.1636 0.055824 6.6836e-05 0.83424 0.005174 0.0059111 0.0013876 0.98693 0.99169 2.9923e-06 1.1969e-05 0.13103 0.93471 0.91015 0.0013978 0.99027 0.58433 0.0018832 0.42837 1.841 1.8402 16.0055 144.9924 0.00017462 -85.6461 0.69021
0.79423 0.98802 5.5207e-05 3.8182 0.012039 1.046e-05 0.0011541 0.12423 0.00065768 0.12488 0.11326 0 0.038733 0.0389 0 0.87502 0.2401 0.063514 0.0089277 4.1638 0.055831 6.6845e-05 0.83424 0.0051742 0.0059113 0.0013876 0.98693 0.99169 2.9922e-06 1.1969e-05 0.13103 0.93486 0.91023 0.0013978 0.99032 0.58448 0.0018831 0.42839 1.8415 1.8407 16.0054 144.9924 0.0001745 -85.6463 0.69121
0.79523 0.98802 5.5207e-05 3.8182 0.012039 1.0473e-05 0.0011541 0.12432 0.00065769 0.12497 0.11335 0 0.038726 0.0389 0 0.87509 0.24013 0.063524 0.008929 4.164 0.055839 6.6855e-05 0.83423 0.0051744 0.0059115 0.0013875 0.98693 0.99169 2.9921e-06 1.1968e-05 0.13103 0.93501 0.9103 0.0013978 0.99036 0.58462 0.0018831 0.4284 1.842 1.8412 16.0054 144.9924 0.00017439 -85.6464 0.69221
0.79623 0.98802 5.5207e-05 3.8182 0.012039 1.0486e-05 0.0011541 0.12441 0.00065769 0.12506 0.11343 0 0.03872 0.0389 0 0.87515 0.24016 0.063534 0.0089303 4.1642 0.055847 6.6865e-05 0.83422 0.0051747 0.0059118 0.0013875 0.98693 0.99169 2.992e-06 1.1968e-05 0.13104 0.93516 0.91037 0.0013977 0.99041 0.58477 0.0018831 0.42841 1.8424 1.8417 16.0054 144.9924 0.00017427 -85.6466 0.69321
0.79723 0.98802 5.5207e-05 3.8182 0.012039 1.0499e-05 0.0011541 0.1245 0.00065769 0.12515 0.11351 0 0.038714 0.0389 0 0.87521 0.24019 0.063544 0.0089315 4.1644 0.055854 6.6874e-05 0.83421 0.0051749 0.005912 0.0013875 0.98693 0.99169 2.9919e-06 1.1967e-05 0.13104 0.93531 0.91045 0.0013977 0.99045 0.58491 0.001883 0.42843 1.8429 1.8422 16.0054 144.9925 0.00017416 -85.6468 0.69421
0.79823 0.98802 5.5207e-05 3.8182 0.012039 1.0513e-05 0.0011541 0.12459 0.00065769 0.12524 0.11359 0 0.038708 0.0389 0 0.87528 0.24022 0.063555 0.0089328 4.1646 0.055862 6.6884e-05 0.83421 0.0051751 0.0059122 0.0013874 0.98693 0.99169 2.9918e-06 1.1967e-05 0.13104 0.93546 0.91052 0.0013977 0.9905 0.58506 0.001883 0.42844 1.8434 1.8427 16.0053 144.9925 0.00017404 -85.6469 0.69521
0.79923 0.98802 5.5207e-05 3.8182 0.012039 1.0526e-05 0.0011541 0.12468 0.0006577 0.12533 0.11368 0 0.038701 0.0389 0 0.87534 0.24024 0.063565 0.0089341 4.1648 0.055869 6.6894e-05 0.8342 0.0051753 0.0059125 0.0013874 0.98693 0.99169 2.9917e-06 1.1967e-05 0.13104 0.93562 0.91059 0.0013977 0.99054 0.5852 0.001883 0.42845 1.8439 1.8431 16.0053 144.9925 0.00017393 -85.6471 0.69621
0.80023 0.98802 5.5207e-05 3.8182 0.012039 1.0539e-05 0.0011541 0.12476 0.0006577 0.12542 0.11376 0 0.038695 0.0389 0 0.87541 0.24027 0.063575 0.0089353 4.165 0.055877 6.6903e-05 0.83419 0.0051756 0.0059127 0.0013874 0.98693 0.99169 2.9916e-06 1.1966e-05 0.13104 0.93576 0.91066 0.0013977 0.99058 0.58534 0.001883 0.42846 1.8444 1.8436 16.0053 144.9925 0.00017382 -85.6473 0.69721
0.80123 0.98802 5.5207e-05 3.8182 0.012039 1.0552e-05 0.0011541 0.12485 0.0006577 0.12551 0.11384 0 0.038689 0.0389 0 0.87547 0.2403 0.063585 0.0089366 4.1652 0.055885 6.6913e-05 0.83418 0.0051758 0.0059129 0.0013873 0.98693 0.99169 2.9915e-06 1.1966e-05 0.13104 0.93591 0.91074 0.0013976 0.99063 0.58549 0.0018829 0.42848 1.8449 1.8441 16.0053 144.9925 0.0001737 -85.6474 0.69821
0.80223 0.98802 5.5207e-05 3.8182 0.012039 1.0565e-05 0.0011541 0.12494 0.0006577 0.12559 0.11392 0 0.038683 0.0389 0 0.87553 0.24033 0.063596 0.0089379 4.1654 0.055892 6.6923e-05 0.83417 0.005176 0.0059131 0.0013873 0.98693 0.9917 2.9915e-06 1.1966e-05 0.13105 0.93606 0.91081 0.0013976 0.99067 0.58563 0.0018829 0.42849 1.8453 1.8446 16.0052 144.9926 0.00017359 -85.6476 0.69921
0.80323 0.98802 5.5207e-05 3.8182 0.012039 1.0578e-05 0.0011541 0.12503 0.00065771 0.12568 0.11401 0 0.038677 0.0389 0 0.8756 0.24036 0.063606 0.0089391 4.1656 0.0559 6.6932e-05 0.83417 0.0051763 0.0059134 0.0013872 0.98693 0.9917 2.9914e-06 1.1965e-05 0.13105 0.93621 0.91088 0.0013976 0.99071 0.58578 0.0018829 0.4285 1.8458 1.8451 16.0052 144.9926 0.00017348 -85.6477 0.70021
0.80423 0.98802 5.5206e-05 3.8182 0.012039 1.0592e-05 0.0011541 0.12512 0.00065771 0.12577 0.11409 0 0.03867 0.0389 0 0.87566 0.24039 0.063616 0.0089404 4.1658 0.055907 6.6942e-05 0.83416 0.0051765 0.0059136 0.0013872 0.98693 0.9917 2.9913e-06 1.1965e-05 0.13105 0.93636 0.91095 0.0013976 0.99075 0.58592 0.0018829 0.42851 1.8463 1.8455 16.0052 144.9926 0.00017336 -85.6479 0.70121
0.80523 0.98802 5.5206e-05 3.8182 0.012039 1.0605e-05 0.0011541 0.12521 0.00065771 0.12586 0.11417 0 0.038664 0.0389 0 0.87573 0.24041 0.063626 0.0089417 4.166 0.055915 6.6952e-05 0.83415 0.0051767 0.0059138 0.0013872 0.98693 0.9917 2.9912e-06 1.1965e-05 0.13105 0.93651 0.91102 0.0013976 0.99079 0.58607 0.0018828 0.42853 1.8468 1.846 16.0052 144.9926 0.00017325 -85.6481 0.70221
0.80623 0.98802 5.5206e-05 3.8182 0.012039 1.0618e-05 0.0011541 0.1253 0.00065771 0.12595 0.11425 0 0.038658 0.0389 0 0.87579 0.24044 0.063637 0.008943 4.1662 0.055923 6.6962e-05 0.83414 0.005177 0.0059141 0.0013871 0.98693 0.9917 2.9911e-06 1.1964e-05 0.13105 0.93665 0.91109 0.0013975 0.99084 0.58621 0.0018828 0.42854 1.8472 1.8465 16.0051 144.9926 0.00017314 -85.6482 0.70321
0.80723 0.98802 5.5206e-05 3.8182 0.012039 1.0631e-05 0.0011541 0.12538 0.00065771 0.12604 0.11434 0 0.038652 0.0389 0 0.87586 0.24047 0.063647 0.0089442 4.1664 0.05593 6.6971e-05 0.83414 0.0051772 0.0059143 0.0013871 0.98693 0.9917 2.991e-06 1.1964e-05 0.13106 0.9368 0.91116 0.0013975 0.99088 0.58635 0.0018828 0.42855 1.8477 1.847 16.0051 144.9927 0.00017303 -85.6484 0.70421
0.80823 0.98802 5.5206e-05 3.8182 0.012039 1.0644e-05 0.0011541 0.12547 0.00065772 0.12613 0.11442 0 0.038646 0.0389 0 0.87592 0.2405 0.063657 0.0089455 4.1666 0.055938 6.6981e-05 0.83413 0.0051774 0.0059145 0.0013871 0.98693 0.9917 2.991e-06 1.1964e-05 0.13106 0.93695 0.91123 0.0013975 0.99092 0.5865 0.0018828 0.42857 1.8482 1.8475 16.0051 144.9927 0.00017292 -85.6485 0.70521
0.80923 0.98802 5.5206e-05 3.8182 0.012039 1.0657e-05 0.0011541 0.12556 0.00065772 0.12621 0.1145 0 0.038639 0.0389 0 0.87598 0.24053 0.063667 0.0089468 4.1668 0.055946 6.6991e-05 0.83412 0.0051777 0.0059148 0.001387 0.98693 0.9917 2.9909e-06 1.1963e-05 0.13106 0.93709 0.9113 0.0013975 0.99096 0.58664 0.0018827 0.42858 1.8487 1.8479 16.0051 144.9927 0.00017281 -85.6487 0.70621
0.81023 0.98802 5.5206e-05 3.8182 0.012039 1.067e-05 0.0011541 0.12565 0.00065772 0.1263 0.11458 0 0.038633 0.0389 0 0.87605 0.24056 0.063678 0.0089481 4.167 0.055953 6.7001e-05 0.83411 0.0051779 0.005915 0.001387 0.98693 0.9917 2.9908e-06 1.1963e-05 0.13106 0.93724 0.91137 0.0013975 0.991 0.58679 0.0018827 0.42859 1.8491 1.8484 16.005 144.9927 0.0001727 -85.6488 0.70721
0.81123 0.98802 5.5206e-05 3.8182 0.012039 1.0684e-05 0.0011541 0.12574 0.00065772 0.12639 0.11466 0 0.038627 0.0389 0 0.87611 0.24059 0.063688 0.0089494 4.1672 0.055961 6.7011e-05 0.83411 0.0051781 0.0059152 0.001387 0.98693 0.9917 2.9907e-06 1.1963e-05 0.13106 0.93738 0.91144 0.0013974 0.99104 0.58693 0.0018827 0.4286 1.8496 1.8489 16.005 144.9927 0.00017259 -85.649 0.70821
0.81223 0.98802 5.5206e-05 3.8182 0.012039 1.0697e-05 0.0011541 0.12583 0.00065773 0.12648 0.11475 0 0.038621 0.0389 0 0.87618 0.24061 0.063698 0.0089506 4.1674 0.055969 6.702e-05 0.8341 0.0051784 0.0059155 0.0013869 0.98694 0.9917 2.9906e-06 1.1962e-05 0.13107 0.93753 0.91151 0.0013974 0.99108 0.58707 0.0018827 0.42862 1.8501 1.8493 16.005 144.9928 0.00017248 -85.6492 0.70921
0.81323 0.98802 5.5206e-05 3.8182 0.012039 1.071e-05 0.0011541 0.12591 0.00065773 0.12657 0.11483 0 0.038615 0.0389 0 0.87624 0.24064 0.063709 0.0089519 4.1677 0.055976 6.703e-05 0.83409 0.0051786 0.0059157 0.0013869 0.98694 0.9917 2.9906e-06 1.1962e-05 0.13107 0.93767 0.91158 0.0013974 0.99112 0.58722 0.0018826 0.42863 1.8505 1.8498 16.005 144.9928 0.00017237 -85.6493 0.71021
0.81423 0.98802 5.5206e-05 3.8182 0.012039 1.0723e-05 0.0011541 0.126 0.00065773 0.12665 0.11491 0 0.038609 0.0389 0 0.87631 0.24067 0.063719 0.0089532 4.1679 0.055984 6.704e-05 0.83408 0.0051788 0.0059159 0.0013868 0.98694 0.9917 2.9905e-06 1.1962e-05 0.13107 0.93781 0.91165 0.0013974 0.99116 0.58736 0.0018826 0.42864 1.851 1.8503 16.0049 144.9928 0.00017227 -85.6495 0.71121
0.81523 0.98802 5.5206e-05 3.8182 0.012039 1.0736e-05 0.0011541 0.12609 0.00065773 0.12674 0.11499 0 0.038603 0.0389 0 0.87637 0.2407 0.063729 0.0089545 4.1681 0.055992 6.705e-05 0.83408 0.0051791 0.0059162 0.0013868 0.98694 0.9917 2.9904e-06 1.1961e-05 0.13107 0.93796 0.91172 0.0013974 0.9912 0.5875 0.0018826 0.42865 1.8515 1.8507 16.0049 144.9928 0.00017216 -85.6496 0.71221
0.81623 0.98802 5.5206e-05 3.8182 0.012039 1.0749e-05 0.0011541 0.12618 0.00065774 0.12683 0.11507 0 0.038596 0.0389 0 0.87644 0.24073 0.06374 0.0089558 4.1683 0.055999 6.706e-05 0.83407 0.0051793 0.0059164 0.0013868 0.98694 0.9917 2.9903e-06 1.1961e-05 0.13107 0.9381 0.91179 0.0013973 0.99124 0.58765 0.0018826 0.42867 1.8519 1.8512 16.0049 144.9928 0.00017205 -85.6497 0.71321
0.81723 0.98802 5.5206e-05 3.8182 0.012039 1.0762e-05 0.0011541 0.12626 0.00065774 0.12692 0.11516 0 0.03859 0.0389 0 0.8765 0.24076 0.06375 0.008957 4.1685 0.056007 6.707e-05 0.83406 0.0051796 0.0059166 0.0013867 0.98694 0.9917 2.9902e-06 1.1961e-05 0.13108 0.93824 0.91186 0.0013973 0.99127 0.58779 0.0018825 0.42868 1.8524 1.8517 16.0048 144.9929 0.00017194 -85.6499 0.71421
0.81823 0.98802 5.5206e-05 3.8182 0.012039 1.0776e-05 0.0011541 0.12635 0.00065774 0.12701 0.11524 0 0.038584 0.0389 0 0.87657 0.24079 0.06376 0.0089583 4.1687 0.056015 6.7079e-05 0.83405 0.0051798 0.0059169 0.0013867 0.98694 0.9917 2.9902e-06 1.1961e-05 0.13108 0.93838 0.91192 0.0013973 0.99131 0.58793 0.0018825 0.42869 1.8529 1.8521 16.0048 144.9929 0.00017184 -85.65 0.71521
0.81923 0.98802 5.5206e-05 3.8182 0.012039 1.0789e-05 0.0011541 0.12644 0.00065774 0.12709 0.11532 0 0.038578 0.0389 0 0.87663 0.24081 0.063771 0.0089596 4.1689 0.056023 6.7089e-05 0.83404 0.00518 0.0059171 0.0013867 0.98694 0.9917 2.9901e-06 1.196e-05 0.13108 0.93852 0.91199 0.0013973 0.99135 0.58808 0.0018825 0.4287 1.8533 1.8526 16.0048 144.9929 0.00017173 -85.6502 0.71621
0.82023 0.98802 5.5205e-05 3.8182 0.012039 1.0802e-05 0.0011541 0.12653 0.00065775 0.12718 0.1154 0 0.038572 0.0389 0 0.8767 0.24084 0.063781 0.0089609 4.1691 0.05603 6.71e-05 0.83404 0.0051803 0.0059174 0.0013866 0.98694 0.9917 2.99e-06 1.196e-05 0.13108 0.93866 0.91206 0.0013973 0.99139 0.58822 0.0018825 0.42872 1.8538 1.8531 16.0048 144.9929 0.00017162 -85.6503 0.71721
0.82123 0.98802 5.5205e-05 3.8182 0.012039 1.0815e-05 0.0011541 0.12661 0.00065775 0.12727 0.11548 0 0.038566 0.0389 0 0.87676 0.24087 0.063791 0.0089622 4.1693 0.056038 6.711e-05 0.83403 0.0051805 0.0059176 0.0013866 0.98694 0.9917 2.9899e-06 1.196e-05 0.13108 0.9388 0.91213 0.0013973 0.99143 0.58836 0.0018825 0.42873 1.8542 1.8535 16.0047 144.9929 0.00017152 -85.6505 0.71821
0.82223 0.98802 5.5205e-05 3.8182 0.012039 1.0828e-05 0.0011541 0.1267 0.00065775 0.12736 0.11556 0 0.03856 0.0389 0 0.87683 0.2409 0.063802 0.0089635 4.1695 0.056046 6.7118e-05 0.83402 0.0051807 0.0059178 0.0013866 0.98694 0.9917 2.9899e-06 1.1959e-05 0.13109 0.93894 0.91219 0.0013972 0.99146 0.58851 0.0018824 0.42874 1.8547 1.854 16.0047 144.993 0.00017141 -85.6506 0.71921
0.82323 0.98802 5.5205e-05 3.8182 0.012039 1.0841e-05 0.0011541 0.12679 0.00065775 0.12744 0.11564 0 0.038554 0.0389 0 0.87689 0.24093 0.063812 0.0089648 4.1697 0.056053 6.7129e-05 0.83401 0.005181 0.0059181 0.0013865 0.98694 0.9917 2.9898e-06 1.1959e-05 0.13109 0.93908 0.91226 0.0013972 0.9915 0.58865 0.0018824 0.42876 1.8552 1.8545 16.0047 144.993 0.00017131 -85.6508 0.72021
0.82423 0.98802 5.5205e-05 3.8182 0.012039 1.0855e-05 0.0011541 0.12688 0.00065776 0.12753 0.11572 0 0.038548 0.0389 0 0.87696 0.24096 0.063822 0.0089661 4.1699 0.056061 6.7141e-05 0.83401 0.0051812 0.0059183 0.0013865 0.98694 0.9917 2.9897e-06 1.1959e-05 0.13109 0.93922 0.91233 0.0013972 0.99154 0.58879 0.0018824 0.42877 1.8556 1.8549 16.0047 144.993 0.0001712 -85.6509 0.72121
0.82523 0.98802 5.5205e-05 3.8182 0.012039 1.0868e-05 0.0011541 0.12696 0.00065776 0.12762 0.11581 0 0.038542 0.0389 0 0.87702 0.24099 0.063833 0.0089673 4.1702 0.056069 6.7147e-05 0.834 0.0051815 0.0059185 0.0013865 0.98694 0.9917 2.9896e-06 1.1958e-05 0.13109 0.93936 0.91239 0.0013972 0.99158 0.58894 0.0018824 0.42878 1.8561 1.8554 16.0046 144.993 0.0001711 -85.651 0.72221
0.82623 0.98802 5.5205e-05 3.8182 0.012039 1.0881e-05 0.0011541 0.12705 0.00065776 0.1277 0.11589 0 0.038536 0.0389 0 0.87709 0.24102 0.063843 0.0089686 4.1704 0.056077 6.7158e-05 0.83399 0.0051817 0.0059188 0.0013864 0.98694 0.9917 2.9896e-06 1.1958e-05 0.13109 0.9395 0.91246 0.0013972 0.99161 0.58908 0.0018823 0.42879 1.8565 1.8558 16.0046 144.993 0.00017099 -85.6512 0.72321
0.82723 0.98802 5.5205e-05 3.8182 0.012039 1.0894e-05 0.0011541 0.12714 0.00065776 0.12779 0.11597 0 0.03853 0.0389 0 0.87715 0.24105 0.063854 0.0089699 4.1706 0.056085 6.7171e-05 0.83398 0.0051819 0.005919 0.0013864 0.98694 0.9917 2.9895e-06 1.1958e-05 0.1311 0.93964 0.91252 0.0013972 0.99165 0.58922 0.0018823 0.42881 1.857 1.8563 16.0046 144.9931 0.00017089 -85.6513 0.72421
0.82823 0.98802 5.5205e-05 3.8182 0.012039 1.0907e-05 0.0011541 0.12722 0.00065776 0.12788 0.11605 0 0.038524 0.0389 0 0.87722 0.24107 0.063864 0.0089712 4.1708 0.056092 6.7177e-05 0.83397 0.0051822 0.0059193 0.0013864 0.98694 0.9917 2.9894e-06 1.1958e-05 0.1311 0.93977 0.91259 0.0013971 0.99168 0.58937 0.0018823 0.42882 1.8574 1.8567 16.0046 144.9931 0.00017079 -85.6514 0.72521
0.82923 0.98802 5.5205e-05 3.8182 0.012039 1.092e-05 0.0011541 0.12731 0.00065777 0.12796 0.11613 0 0.038517 0.0389 0 0.87728 0.2411 0.063874 0.0089725 4.171 0.0561 6.7187e-05 0.83397 0.0051824 0.0059195 0.0013864 0.98694 0.9917 2.9893e-06 1.1957e-05 0.1311 0.93991 0.91266 0.0013971 0.99172 0.58951 0.0018823 0.42883 1.8579 1.8572 16.0045 144.9931 0.00017068 -85.6516 0.72621
0.83023 0.98802 5.5205e-05 3.8182 0.012039 1.0933e-05 0.0011541 0.1274 0.00065777 0.12805 0.11621 0 0.038511 0.0389 0 0.87735 0.24113 0.063885 0.0089738 4.1712 0.056108 6.72e-05 0.83396 0.0051827 0.0059197 0.0013863 0.98694 0.9917 2.9893e-06 1.1957e-05 0.1311 0.94005 0.91272 0.0013971 0.99175 0.58965 0.0018823 0.42884 1.8583 1.8577 16.0045 144.9931 0.00017058 -85.6517 0.72721
0.83123 0.98802 5.5205e-05 3.8182 0.012039 1.0947e-05 0.0011541 0.12749 0.00065777 0.12814 0.11629 0 0.038505 0.0389 0 0.87741 0.24116 0.063895 0.0089751 4.1714 0.056116 6.7208e-05 0.83395 0.0051829 0.00592 0.0013863 0.98694 0.9917 2.9892e-06 1.1957e-05 0.1311 0.94018 0.91279 0.0013971 0.99179 0.58979 0.0018822 0.42886 1.8588 1.8581 16.0045 144.9932 0.00017048 -85.6518 0.72821
0.83223 0.98802 5.5205e-05 3.8182 0.012039 1.096e-05 0.0011541 0.12757 0.00065777 0.12823 0.11637 0 0.038499 0.0389 0 0.87748 0.24119 0.063906 0.0089764 4.1716 0.056123 6.7218e-05 0.83394 0.0051832 0.0059202 0.0013863 0.98694 0.9917 2.9891e-06 1.1956e-05 0.13111 0.94032 0.91285 0.0013971 0.99183 0.58994 0.0018822 0.42887 1.8593 1.8586 16.0044 144.9932 0.00017038 -85.652 0.72921
0.83323 0.98802 5.5205e-05 3.8182 0.012039 1.0973e-05 0.0011541 0.12766 0.00065778 0.12831 0.11645 0 0.038493 0.0389 0 0.87755 0.24122 0.063916 0.0089777 4.1719 0.056131 6.7228e-05 0.83394 0.0051834 0.0059205 0.0013862 0.98694 0.9917 2.9891e-06 1.1956e-05 0.13111 0.94045 0.91292 0.0013971 0.99186 0.59008 0.0018822 0.42888 1.8597 1.859 16.0044 144.9932 0.00017028 -85.6521 0.73021
0.83423 0.98802 5.5205e-05 3.8182 0.012039 1.0986e-05 0.0011541 0.12775 0.00065778 0.1284 0.11653 0 0.038487 0.0389 0 0.87761 0.24125 0.063927 0.008979 4.1721 0.056139 6.7238e-05 0.83393 0.0051836 0.0059207 0.0013862 0.98694 0.9917 2.989e-06 1.1956e-05 0.13111 0.94059 0.91298 0.001397 0.99189 0.59022 0.0018822 0.42889 1.8601 1.8595 16.0044 144.9932 0.00017018 -85.6522 0.73121
0.83523 0.98802 5.5205e-05 3.8182 0.012039 1.0999e-05 0.0011541 0.12783 0.00065778 0.12848 0.11661 0 0.038481 0.0389 0 0.87768 0.24128 0.063937 0.0089803 4.1723 0.056147 6.7248e-05 0.83392 0.0051839 0.005921 0.0013862 0.98694 0.9917 2.9889e-06 1.1956e-05 0.13111 0.94072 0.91304 0.001397 0.99193 0.59037 0.0018821 0.42891 1.8606 1.8599 16.0044 144.9932 0.00017008 -85.6524 0.73221
0.83623 0.98802 5.5204e-05 3.8182 0.012039 1.1012e-05 0.0011541 0.12792 0.00065778 0.12857 0.11669 0 0.038475 0.0389 0 0.87774 0.24131 0.063948 0.0089816 4.1725 0.056155 6.7258e-05 0.83391 0.0051841 0.0059212 0.0013861 0.98695 0.9917 2.9889e-06 1.1955e-05 0.13111 0.94085 0.91311 0.001397 0.99196 0.59051 0.0018821 0.42892 1.861 1.8604 16.0043 144.9933 0.00016997 -85.6525 0.73321
0.83723 0.98802 5.5204e-05 3.8182 0.012039 1.1026e-05 0.0011541 0.128 0.00065779 0.12866 0.11677 0 0.038469 0.0389 0 0.87781 0.24133 0.063958 0.0089829 4.1727 0.056162 6.7268e-05 0.8339 0.0051844 0.0059215 0.0013861 0.98695 0.9917 2.9888e-06 1.1955e-05 0.13112 0.94099 0.91317 0.001397 0.992 0.59065 0.0018821 0.42893 1.8615 1.8608 16.0043 144.9933 0.00016987 -85.6526 0.73421
0.83823 0.98802 5.5204e-05 3.8182 0.012039 1.1039e-05 0.0011541 0.12809 0.00065779 0.12874 0.11685 0 0.038463 0.0389 0 0.87787 0.24136 0.063969 0.0089842 4.1729 0.05617 6.7278e-05 0.8339 0.0051846 0.0059217 0.0013861 0.98695 0.99171 2.9887e-06 1.1955e-05 0.13112 0.94112 0.91323 0.001397 0.99203 0.59079 0.0018821 0.42894 1.8619 1.8612 16.0043 144.9933 0.00016978 -85.6528 0.73521
0.83923 0.98802 5.5204e-05 3.8182 0.012039 1.1052e-05 0.0011541 0.12818 0.00065779 0.12883 0.11693 0 0.038458 0.0389 0 0.87794 0.24139 0.063979 0.0089855 4.1732 0.056178 6.7288e-05 0.83389 0.0051849 0.0059219 0.0013861 0.98695 0.99171 2.9887e-06 1.1955e-05 0.13112 0.94125 0.9133 0.001397 0.99206 0.59094 0.0018821 0.42896 1.8624 1.8617 16.0043 144.9933 0.00016968 -85.6529 0.73621
0.84023 0.98802 5.5204e-05 3.8182 0.012039 1.1065e-05 0.0011541 0.12826 0.00065779 0.12892 0.11701 0 0.038452 0.0389 0 0.87801 0.24142 0.06399 0.0089868 4.1734 0.056186 6.7298e-05 0.83388 0.0051851 0.0059222 0.001386 0.98695 0.99171 2.9886e-06 1.1954e-05 0.13112 0.94139 0.91336 0.0013969 0.9921 0.59108 0.001882 0.42897 1.8628 1.8621 16.0042 144.9933 0.00016958 -85.653 0.73721
0.84123 0.98802 5.5204e-05 3.8182 0.012039 1.1078e-05 0.0011541 0.12835 0.00065779 0.129 0.11709 0 0.038446 0.0389 0 0.87807 0.24145 0.064 0.0089881 4.1736 0.056194 6.7308e-05 0.83387 0.0051854 0.0059224 0.001386 0.98695 0.99171 2.9885e-06 1.1954e-05 0.13112 0.94152 0.91342 0.0013969 0.99213 0.59122 0.001882 0.42898 1.8633 1.8626 16.0042 144.9934 0.00016948 -85.6531 0.73821
0.84223 0.98802 5.5204e-05 3.8182 0.012039 1.1091e-05 0.0011541 0.12843 0.0006578 0.12909 0.11717 0 0.03844 0.0389 0 0.87814 0.24148 0.064011 0.0089894 4.1738 0.056202 6.7318e-05 0.83387 0.0051856 0.0059227 0.001386 0.98695 0.99171 2.9885e-06 1.1954e-05 0.13113 0.94165 0.91349 0.0013969 0.99216 0.59136 0.001882 0.42899 1.8637 1.863 16.0042 144.9934 0.00016938 -85.6533 0.73921
0.84323 0.98802 5.5204e-05 3.8182 0.012039 1.1104e-05 0.0011541 0.12852 0.0006578 0.12917 0.11725 0 0.038434 0.0389 0 0.8782 0.24151 0.064021 0.0089907 4.174 0.05621 6.7328e-05 0.83386 0.0051858 0.0059229 0.0013859 0.98695 0.99171 2.9884e-06 1.1953e-05 0.13113 0.94178 0.91355 0.0013969 0.9922 0.5915 0.001882 0.42901 1.8641 1.8635 16.0041 144.9934 0.00016928 -85.6534 0.74021
0.84423 0.98802 5.5204e-05 3.8182 0.012039 1.1118e-05 0.0011541 0.12861 0.0006578 0.12926 0.11733 0 0.038428 0.0389 0 0.87827 0.24154 0.064032 0.008992 4.1742 0.056217 6.7338e-05 0.83385 0.0051861 0.0059232 0.0013859 0.98695 0.99171 2.9883e-06 1.1953e-05 0.13113 0.94191 0.91361 0.0013969 0.99223 0.59165 0.001882 0.42902 1.8646 1.8639 16.0041 144.9934 0.00016918 -85.6535 0.74121
0.84523 0.98802 5.5204e-05 3.8182 0.012039 1.1131e-05 0.0011541 0.12869 0.0006578 0.12935 0.11741 0 0.038422 0.0389 0 0.87834 0.24157 0.064042 0.0089933 4.1745 0.056225 6.7348e-05 0.83384 0.0051863 0.0059234 0.0013859 0.98695 0.99171 2.9883e-06 1.1953e-05 0.13113 0.94204 0.91367 0.0013969 0.99226 0.59179 0.0018819 0.42903 1.865 1.8643 16.0041 144.9934 0.00016909 -85.6536 0.74221
0.84623 0.98802 5.5204e-05 3.8182 0.012039 1.1144e-05 0.0011541 0.12878 0.00065781 0.12943 0.11749 0 0.038416 0.0389 0 0.8784 0.2416 0.064053 0.0089946 4.1747 0.056233 6.7358e-05 0.83383 0.0051866 0.0059237 0.0013859 0.98695 0.99171 2.9882e-06 1.1953e-05 0.13113 0.94217 0.91373 0.0013969 0.99229 0.59193 0.0018819 0.42904 1.8655 1.8648 16.0041 144.9935 0.00016899 -85.6537 0.74321
0.84723 0.98802 5.5204e-05 3.8182 0.012039 1.1157e-05 0.0011541 0.12886 0.00065781 0.12952 0.11757 0 0.03841 0.0389 0 0.87847 0.24163 0.064063 0.0089959 4.1749 0.056241 6.7368e-05 0.83383 0.0051868 0.0059239 0.0013858 0.98695 0.99171 2.9881e-06 1.1952e-05 0.13114 0.9423 0.9138 0.0013968 0.99232 0.59207 0.0018819 0.42906 1.8659 1.8652 16.004 144.9935 0.00016889 -85.6539 0.74421
0.84823 0.98802 5.5204e-05 3.8182 0.012039 1.117e-05 0.0011541 0.12895 0.00065781 0.1296 0.11765 0 0.038404 0.0389 0 0.87853 0.24166 0.064074 0.0089973 4.1751 0.056249 6.7379e-05 0.83382 0.0051871 0.0059242 0.0013858 0.98695 0.99171 2.9881e-06 1.1952e-05 0.13114 0.94243 0.91386 0.0013968 0.99236 0.59221 0.0018819 0.42907 1.8663 1.8657 16.004 144.9935 0.0001688 -85.654 0.74521
0.84923 0.98802 5.5204e-05 3.8182 0.012039 1.1183e-05 0.0011541 0.12903 0.00065781 0.12969 0.11773 0 0.038398 0.0389 0 0.8786 0.24169 0.064085 0.0089986 4.1753 0.056257 6.7389e-05 0.83381 0.0051873 0.0059244 0.0013858 0.98695 0.99171 2.988e-06 1.1952e-05 0.13114 0.94256 0.91392 0.0013968 0.99239 0.59236 0.0018819 0.42908 1.8668 1.8661 16.004 144.9935 0.0001687 -85.6541 0.74621
0.85023 0.98802 5.5204e-05 3.8182 0.012039 1.1196e-05 0.0011541 0.12912 0.00065781 0.12977 0.11781 0 0.038392 0.0389 0 0.87867 0.24171 0.064095 0.0089999 4.1756 0.056265 6.7399e-05 0.8338 0.0051876 0.0059247 0.0013857 0.98695 0.99171 2.988e-06 1.1952e-05 0.13114 0.94268 0.91398 0.0013968 0.99242 0.5925 0.0018819 0.42909 1.8672 1.8665 16.0039 144.9935 0.0001686 -85.6542 0.74721
0.85123 0.98802 5.5204e-05 3.8182 0.012039 1.121e-05 0.0011541 0.12921 0.00065782 0.12986 0.11789 0 0.038386 0.0389 0 0.87873 0.24174 0.064106 0.0090012 4.1758 0.056273 6.7409e-05 0.83379 0.0051878 0.0059249 0.0013857 0.98695 0.99171 2.9879e-06 1.1951e-05 0.13114 0.94281 0.91404 0.0013968 0.99245 0.59264 0.0018818 0.42911 1.8676 1.867 16.0039 144.9936 0.00016851 -85.6543 0.74821
0.85223 0.98802 5.5203e-05 3.8182 0.012039 1.1223e-05 0.0011541 0.12929 0.00065782 0.12994 0.11797 0 0.038381 0.0389 0 0.8788 0.24177 0.064116 0.0090025 4.176 0.05628 6.7419e-05 0.83379 0.0051881 0.0059252 0.0013857 0.98695 0.99171 2.9878e-06 1.1951e-05 0.13115 0.94294 0.9141 0.0013968 0.99248 0.59278 0.0018818 0.42912 1.8681 1.8674 16.0039 144.9936 0.00016841 -85.6545 0.74921
0.85323 0.98802 5.5203e-05 3.8182 0.012039 1.1236e-05 0.0011541 0.12938 0.00065782 0.13003 0.11805 0 0.038375 0.0389 0 0.87887 0.2418 0.064127 0.0090038 4.1762 0.056288 6.7429e-05 0.83378 0.0051883 0.0059254 0.0013857 0.98695 0.99171 2.9878e-06 1.1951e-05 0.13115 0.94307 0.91416 0.0013968 0.99251 0.59292 0.0018818 0.42913 1.8685 1.8678 16.0039 144.9936 0.00016832 -85.6546 0.75021
0.85423 0.98802 5.5203e-05 3.8182 0.012039 1.1249e-05 0.0011541 0.12946 0.00065782 0.13011 0.11813 0 0.038369 0.0389 0 0.87893 0.24183 0.064137 0.0090051 4.1765 0.056296 6.7439e-05 0.83377 0.0051886 0.0059257 0.0013856 0.98695 0.99171 2.9877e-06 1.1951e-05 0.13115 0.94319 0.91422 0.0013967 0.99254 0.59307 0.0018818 0.42914 1.8689 1.8683 16.0038 144.9936 0.00016823 -85.6547 0.75121
0.85523 0.98802 5.5203e-05 3.8182 0.012039 1.1262e-05 0.0011541 0.12955 0.00065783 0.1302 0.11821 0 0.038363 0.0389 0 0.879 0.24186 0.064148 0.0090064 4.1767 0.056304 6.7449e-05 0.83376 0.0051888 0.0059259 0.0013856 0.98695 0.99171 2.9876e-06 1.195e-05 0.13115 0.94332 0.91428 0.0013967 0.99257 0.59321 0.0018818 0.42916 1.8694 1.8687 16.0038 144.9936 0.00016813 -85.6548 0.75221
0.85623 0.98802 5.5203e-05 3.8182 0.012039 1.1275e-05 0.0011541 0.12963 0.00065783 0.13028 0.11829 0 0.038357 0.0389 0 0.87906 0.24189 0.064159 0.0090078 4.1769 0.056312 6.7459e-05 0.83376 0.0051891 0.0059262 0.0013856 0.98695 0.99171 2.9876e-06 1.195e-05 0.13116 0.94344 0.91434 0.0013967 0.9926 0.59335 0.0018817 0.42917 1.8698 1.8691 16.0038 144.9937 0.00016804 -85.6549 0.75321
0.85723 0.98802 5.5203e-05 3.8182 0.012039 1.1289e-05 0.0011541 0.12972 0.00065783 0.13037 0.11837 0 0.038351 0.0389 0 0.87913 0.24192 0.064169 0.0090091 4.1771 0.05632 6.7469e-05 0.83375 0.0051894 0.0059264 0.0013856 0.98695 0.99171 2.9875e-06 1.195e-05 0.13116 0.94357 0.9144 0.0013967 0.99263 0.59349 0.0018817 0.42918 1.8702 1.8696 16.0038 144.9937 0.00016794 -85.655 0.75421
0.85823 0.98802 5.5203e-05 3.8182 0.012039 1.1302e-05 0.0011541 0.1298 0.00065783 0.13045 0.11845 0 0.038345 0.0389 0 0.8792 0.24195 0.06418 0.0090104 4.1773 0.056328 6.748e-05 0.83374 0.0051896 0.0059267 0.0013855 0.98695 0.99171 2.9875e-06 1.195e-05 0.13116 0.9437 0.91446 0.0013967 0.99266 0.59363 0.0018817 0.42919 1.8706 1.87 16.0037 144.9937 0.00016785 -85.6551 0.75521
0.85923 0.98802 5.5203e-05 3.8182 0.012039 1.1315e-05 0.0011541 0.12989 0.00065783 0.13054 0.11853 0 0.03834 0.0389 0 0.87926 0.24198 0.064191 0.0090117 4.1776 0.056336 6.749e-05 0.83373 0.0051899 0.0059269 0.0013855 0.98695 0.99171 2.9874e-06 1.195e-05 0.13116 0.94382 0.91452 0.0013967 0.99269 0.59377 0.0018817 0.42921 1.8711 1.8704 16.0037 144.9937 0.00016776 -85.6552 0.75621
0.86023 0.98802 5.5203e-05 3.8182 0.012039 1.1328e-05 0.0011541 0.12997 0.00065784 0.13062 0.1186 0 0.038334 0.0389 0 0.87933 0.24201 0.064201 0.009013 4.1778 0.056344 6.75e-05 0.83372 0.0051901 0.0059272 0.0013855 0.98695 0.99171 2.9874e-06 1.1949e-05 0.13116 0.94394 0.91458 0.0013967 0.99272 0.59391 0.0018817 0.42922 1.8715 1.8708 16.0037 144.9937 0.00016767 -85.6553 0.75721
0.86123 0.98802 5.5203e-05 3.8182 0.012039 1.1341e-05 0.0011541 0.13005 0.00065784 0.13071 0.11868 0 0.038328 0.0389 0 0.8794 0.24204 0.064212 0.0090144 4.178 0.056352 6.7511e-05 0.83372 0.0051904 0.0059274 0.0013855 0.98695 0.99171 2.9873e-06 1.1949e-05 0.13117 0.94407 0.91464 0.0013967 0.99275 0.59406 0.0018817 0.42923 1.8719 1.8713 16.0036 144.9938 0.00016757 -85.6555 0.75821
0.86223 0.98802 5.5203e-05 3.8182 0.012039 1.1354e-05 0.0011541 0.13014 0.00065784 0.13079 0.11876 0 0.038322 0.0389 0 0.87946 0.24207 0.064223 0.0090157 4.1782 0.05636 6.7521e-05 0.83371 0.0051906 0.0059277 0.0013854 0.98695 0.99171 2.9872e-06 1.1949e-05 0.13117 0.94419 0.91469 0.0013966 0.99278 0.5942 0.0018816 0.42924 1.8723 1.8717 16.0036 144.9938 0.00016748 -85.6556 0.75921
0.86323 0.98802 5.5203e-05 3.8182 0.012039 1.1367e-05 0.0011541 0.13022 0.00065784 0.13088 0.11884 0 0.038316 0.0389 0 0.87953 0.2421 0.064233 0.009017 4.1785 0.056368 6.753e-05 0.8337 0.0051909 0.0059279 0.0013854 0.98695 0.99171 2.9872e-06 1.1949e-05 0.13117 0.94431 0.91475 0.0013966 0.99281 0.59434 0.0018816 0.42926 1.8728 1.8721 16.0036 144.9938 0.00016739 -85.6557 0.76021
0.86423 0.98802 5.5203e-05 3.8182 0.012039 1.1381e-05 0.0011541 0.13031 0.00065785 0.13096 0.11892 0 0.03831 0.0389 0 0.8796 0.24213 0.064244 0.0090183 4.1787 0.056376 6.7541e-05 0.83369 0.0051911 0.0059282 0.0013854 0.98695 0.99171 2.9871e-06 1.1948e-05 0.13117 0.94444 0.91481 0.0013966 0.99283 0.59448 0.0018816 0.42927 1.8732 1.8725 16.0036 144.9938 0.0001673 -85.6558 0.76121
0.86523 0.98802 5.5203e-05 3.8182 0.012039 1.1394e-05 0.0011541 0.13039 0.00065785 0.13105 0.119 0 0.038305 0.0389 0 0.87967 0.24216 0.064255 0.0090196 4.1789 0.056384 6.7552e-05 0.83368 0.0051914 0.0059285 0.0013854 0.98696 0.99171 2.9871e-06 1.1948e-05 0.13117 0.94456 0.91487 0.0013966 0.99286 0.59462 0.0018816 0.42928 1.8736 1.873 16.0035 144.9938 0.00016721 -85.6559 0.76221
0.86623 0.98802 5.5203e-05 3.8182 0.012039 1.1407e-05 0.0011541 0.13048 0.00065785 0.13113 0.11908 0 0.038299 0.0389 0 0.87973 0.24219 0.064265 0.009021 4.1792 0.056392 6.756e-05 0.83368 0.0051916 0.0059287 0.0013853 0.98696 0.99171 2.987e-06 1.1948e-05 0.13118 0.94468 0.91493 0.0013966 0.99289 0.59476 0.0018816 0.42929 1.874 1.8734 16.0035 144.9939 0.00016712 -85.656 0.76321
0.86723 0.98802 5.5203e-05 3.8182 0.012038 1.142e-05 0.0011541 0.13056 0.00065785 0.13121 0.11915 0 0.038293 0.0389 0 0.8798 0.24222 0.064276 0.0090223 4.1794 0.0564 6.757e-05 0.83367 0.0051919 0.005929 0.0013853 0.98696 0.99171 2.987e-06 1.1948e-05 0.13118 0.9448 0.91498 0.0013966 0.99292 0.5949 0.0018816 0.42931 1.8745 1.8738 16.0035 144.9939 0.00016703 -85.6561 0.76421
0.86823 0.98802 5.5202e-05 3.8182 0.012038 1.1433e-05 0.0011541 0.13065 0.00065785 0.1313 0.11923 0 0.038287 0.0389 0 0.87987 0.24225 0.064287 0.0090236 4.1796 0.056408 6.7585e-05 0.83366 0.0051922 0.0059292 0.0013853 0.98696 0.99171 2.9869e-06 1.1948e-05 0.13118 0.94492 0.91504 0.0013966 0.99295 0.59504 0.0018815 0.42932 1.8749 1.8742 16.0034 144.9939 0.00016694 -85.6562 0.76521
0.86923 0.98802 5.5202e-05 3.8182 0.012038 1.1446e-05 0.0011541 0.13073 0.00065786 0.13138 0.11931 0 0.038281 0.0389 0 0.87993 0.24228 0.064297 0.0090249 4.1798 0.056416 6.7593e-05 0.83365 0.0051924 0.0059295 0.0013853 0.98696 0.99171 2.9869e-06 1.1947e-05 0.13118 0.94504 0.9151 0.0013965 0.99297 0.59518 0.0018815 0.42933 1.8753 1.8747 16.0034 144.9939 0.00016685 -85.6563 0.76621
0.87023 0.98802 5.5202e-05 3.8182 0.012038 1.1459e-05 0.0011541 0.13081 0.00065786 0.13147 0.11939 0 0.038276 0.0389 0 0.88 0.2423 0.064308 0.0090263 4.1801 0.056424 6.7602e-05 0.83364 0.0051927 0.0059297 0.0013852 0.98696 0.99171 2.9868e-06 1.1947e-05 0.13118 0.94516 0.91515 0.0013965 0.993 0.59533 0.0018815 0.42934 1.8757 1.8751 16.0034 144.9939 0.00016676 -85.6564 0.76721
0.87123 0.98802 5.5202e-05 3.8182 0.012038 1.1473e-05 0.0011541 0.1309 0.00065786 0.13155 0.11947 0 0.03827 0.0389 0 0.88007 0.24233 0.064319 0.0090276 4.1803 0.056432 6.7614e-05 0.83364 0.0051929 0.00593 0.0013852 0.98696 0.99171 2.9867e-06 1.1947e-05 0.13119 0.94528 0.91521 0.0013965 0.99303 0.59547 0.0018815 0.42936 1.8761 1.8755 16.0034 144.994 0.00016667 -85.6565 0.76821
0.87223 0.98802 5.5202e-05 3.8182 0.012038 1.1486e-05 0.0011541 0.13098 0.00065786 0.13164 0.11955 0 0.038264 0.0389 0 0.88013 0.24236 0.06433 0.0090289 4.1805 0.05644 6.7623e-05 0.83363 0.0051932 0.0059303 0.0013852 0.98696 0.99171 2.9867e-06 1.1947e-05 0.13119 0.9454 0.91527 0.0013965 0.99305 0.59561 0.0018815 0.42937 1.8765 1.8759 16.0033 144.994 0.00016658 -85.6566 0.76921
0.87323 0.98802 5.5202e-05 3.8182 0.012038 1.1499e-05 0.0011541 0.13107 0.00065786 0.13172 0.11962 0 0.038258 0.0389 0 0.8802 0.24239 0.06434 0.0090303 4.1808 0.056448 6.7632e-05 0.83362 0.0051935 0.0059305 0.0013852 0.98696 0.99171 2.9866e-06 1.1946e-05 0.13119 0.94552 0.91532 0.0013965 0.99308 0.59575 0.0018815 0.42938 1.877 1.8763 16.0033 144.994 0.00016649 -85.6567 0.77021
0.87423 0.98802 5.5202e-05 3.8182 0.012038 1.1512e-05 0.0011541 0.13115 0.00065787 0.1318 0.1197 0 0.038253 0.0389 0 0.88027 0.24242 0.064351 0.0090316 4.181 0.056456 6.7644e-05 0.83361 0.0051937 0.0059308 0.0013851 0.98696 0.99171 2.9866e-06 1.1946e-05 0.13119 0.94564 0.91538 0.0013965 0.99311 0.59589 0.0018814 0.42939 1.8774 1.8767 16.0033 144.994 0.0001664 -85.6568 0.77121
0.87523 0.98802 5.5202e-05 3.8182 0.012038 1.1525e-05 0.0011541 0.13123 0.00065787 0.13189 0.11978 0 0.038247 0.0389 0 0.88034 0.24245 0.064362 0.0090329 4.1812 0.056464 6.7654e-05 0.8336 0.005194 0.005931 0.0013851 0.98696 0.99171 2.9865e-06 1.1946e-05 0.1312 0.94576 0.91544 0.0013965 0.99313 0.59603 0.0018814 0.4294 1.8778 1.8772 16.0032 144.9941 0.00016632 -85.6569 0.77221
0.87623 0.98802 5.5202e-05 3.8182 0.012038 1.1538e-05 0.0011541 0.13132 0.00065787 0.13197 0.11986 0 0.038241 0.0389 0 0.8804 0.24248 0.064373 0.0090343 4.1815 0.056472 6.7663e-05 0.8336 0.0051942 0.0059313 0.0013851 0.98696 0.99171 2.9865e-06 1.1946e-05 0.1312 0.94588 0.91549 0.0013965 0.99316 0.59617 0.0018814 0.42942 1.8782 1.8776 16.0032 144.9941 0.00016623 -85.657 0.77321
0.87723 0.98802 5.5202e-05 3.8182 0.012038 1.1552e-05 0.0011541 0.1314 0.00065787 0.13205 0.11994 0 0.038235 0.0389 0 0.88047 0.24251 0.064383 0.0090356 4.1817 0.05648 6.7674e-05 0.83359 0.0051945 0.0059316 0.0013851 0.98696 0.99171 2.9864e-06 1.1946e-05 0.1312 0.946 0.91555 0.0013964 0.99319 0.59631 0.0018814 0.42943 1.8786 1.878 16.0032 144.9941 0.00016614 -85.6571 0.77421
0.87823 0.98802 5.5202e-05 3.8182 0.012038 1.1565e-05 0.0011541 0.13148 0.00065788 0.13214 0.12001 0 0.03823 0.0389 0 0.88054 0.24254 0.064394 0.0090369 4.1819 0.056488 6.7685e-05 0.83358 0.0051948 0.0059318 0.0013851 0.98696 0.99171 2.9864e-06 1.1945e-05 0.1312 0.94611 0.9156 0.0013964 0.99321 0.59645 0.0018814 0.42944 1.879 1.8784 16.0032 144.9941 0.00016605 -85.6572 0.77521
0.87923 0.98802 5.5202e-05 3.8182 0.012038 1.1578e-05 0.0011541 0.13157 0.00065788 0.13222 0.12009 0 0.038224 0.0389 0 0.88061 0.24257 0.064405 0.0090383 4.1822 0.056496 6.7694e-05 0.83357 0.005195 0.0059321 0.001385 0.98696 0.99171 2.9863e-06 1.1945e-05 0.1312 0.94623 0.91566 0.0013964 0.99324 0.59659 0.0018814 0.42945 1.8794 1.8788 16.0031 144.9941 0.00016597 -85.6573 0.77621
0.88023 0.98802 5.5202e-05 3.8182 0.012038 1.1591e-05 0.0011541 0.13165 0.00065788 0.1323 0.12017 0 0.038218 0.0389 0 0.88067 0.2426 0.064416 0.0090396 4.1824 0.056504 6.7705e-05 0.83356 0.0051953 0.0059323 0.001385 0.98696 0.99171 2.9863e-06 1.1945e-05 0.13121 0.94635 0.91571 0.0013964 0.99326 0.59673 0.0018813 0.42947 1.8798 1.8792 16.0031 144.9942 0.00016588 -85.6574 0.77721
0.88123 0.98802 5.5202e-05 3.8182 0.012038 1.1604e-05 0.0011541 0.13173 0.00065788 0.13239 0.12025 0 0.038213 0.0389 0 0.88074 0.24263 0.064426 0.0090409 4.1826 0.056512 6.7716e-05 0.83356 0.0051955 0.0059326 0.001385 0.98696 0.99171 2.9862e-06 1.1945e-05 0.13121 0.94646 0.91577 0.0013964 0.99329 0.59687 0.0018813 0.42948 1.8802 1.8796 16.0031 144.9942 0.00016579 -85.6575 0.77821
0.88223 0.98802 5.5202e-05 3.8182 0.012038 1.1617e-05 0.0011541 0.13182 0.00065788 0.13247 0.12032 0 0.038207 0.0389 0 0.88081 0.24266 0.064437 0.0090423 4.1829 0.05652 6.7726e-05 0.83355 0.0051958 0.0059329 0.001385 0.98696 0.99171 2.9862e-06 1.1945e-05 0.13121 0.94658 0.91582 0.0013964 0.99332 0.59701 0.0018813 0.42949 1.8807 1.88 16.003 144.9942 0.00016571 -85.6576 0.77921
0.88323 0.98802 5.5202e-05 3.8182 0.012038 1.163e-05 0.0011541 0.1319 0.00065789 0.13255 0.1204 0 0.038201 0.0389 0 0.88088 0.24269 0.064448 0.0090436 4.1831 0.056528 6.7736e-05 0.83354 0.0051961 0.0059331 0.0013849 0.98696 0.99171 2.9861e-06 1.1944e-05 0.13121 0.94669 0.91588 0.0013964 0.99334 0.59715 0.0018813 0.4295 1.8811 1.8804 16.003 144.9942 0.00016562 -85.6577 0.78021
0.88423 0.98802 5.5201e-05 3.8182 0.012038 1.1644e-05 0.0011541 0.13198 0.00065789 0.13264 0.12048 0 0.038196 0.0389 0 0.88094 0.24272 0.064459 0.0090449 4.1833 0.056536 6.7747e-05 0.83353 0.0051963 0.0059334 0.0013849 0.98696 0.99171 2.9861e-06 1.1944e-05 0.13122 0.94681 0.91593 0.0013964 0.99337 0.59729 0.0018813 0.42952 1.8815 1.8809 16.003 144.9942 0.00016554 -85.6578 0.78121
0.88523 0.98802 5.5201e-05 3.8182 0.012038 1.1657e-05 0.0011541 0.13207 0.00065789 0.13272 0.12056 0 0.03819 0.0389 0 0.88101 0.24275 0.06447 0.0090463 4.1836 0.056545 6.7757e-05 0.83352 0.0051966 0.0059337 0.0013849 0.98696 0.99171 2.986e-06 1.1944e-05 0.13122 0.94692 0.91598 0.0013964 0.99339 0.59743 0.0018813 0.42953 1.8819 1.8813 16.0029 144.9943 0.00016545 -85.6579 0.78221
0.88623 0.98802 5.5201e-05 3.8182 0.012038 1.167e-05 0.0011541 0.13215 0.00065789 0.1328 0.12063 0 0.038184 0.0389 0 0.88108 0.24278 0.06448 0.0090476 4.1838 0.056553 6.7767e-05 0.83352 0.0051969 0.0059339 0.0013849 0.98696 0.99171 2.986e-06 1.1944e-05 0.13122 0.94704 0.91604 0.0013963 0.99341 0.59757 0.0018813 0.42954 1.8823 1.8817 16.0029 144.9943 0.00016537 -85.6579 0.78321
0.88723 0.98802 5.5201e-05 3.8182 0.012038 1.1683e-05 0.0011541 0.13223 0.00065789 0.13289 0.12071 0 0.038179 0.0389 0 0.88115 0.24281 0.064491 0.009049 4.184 0.056561 6.7778e-05 0.83351 0.0051971 0.0059342 0.0013849 0.98696 0.99172 2.9859e-06 1.1944e-05 0.13122 0.94715 0.91609 0.0013963 0.99344 0.59771 0.0018812 0.42955 1.8827 1.8821 16.0029 144.9943 0.00016528 -85.658 0.78421
0.88823 0.98802 5.5201e-05 3.8182 0.012038 1.1696e-05 0.0011541 0.13232 0.0006579 0.13297 0.12079 0 0.038173 0.0389 0 0.88122 0.24284 0.064502 0.0090503 4.1843 0.056569 6.7788e-05 0.8335 0.0051974 0.0059344 0.0013848 0.98696 0.99172 2.9859e-06 1.1943e-05 0.13122 0.94727 0.91615 0.0013963 0.99346 0.59785 0.0018812 0.42957 1.8831 1.8825 16.0029 144.9943 0.0001652 -85.6581 0.78521
0.88923 0.98802 5.5201e-05 3.8182 0.012038 1.1709e-05 0.0011541 0.1324 0.0006579 0.13305 0.12087 0 0.038167 0.0389 0 0.88128 0.24287 0.064513 0.0090516 4.1845 0.056577 6.7798e-05 0.83349 0.0051977 0.0059347 0.0013848 0.98696 0.99172 2.9858e-06 1.1943e-05 0.13123 0.94738 0.9162 0.0013963 0.99349 0.59799 0.0018812 0.42958 1.8835 1.8829 16.0028 144.9943 0.00016512 -85.6582 0.78621
0.89023 0.98802 5.5201e-05 3.8182 0.012038 1.1722e-05 0.0011541 0.13248 0.0006579 0.13313 0.12094 0 0.038162 0.0389 0 0.88135 0.2429 0.064524 0.009053 4.1847 0.056585 6.7809e-05 0.83348 0.0051979 0.005935 0.0013848 0.98696 0.99172 2.9858e-06 1.1943e-05 0.13123 0.94749 0.91625 0.0013963 0.99351 0.59813 0.0018812 0.42959 1.8839 1.8833 16.0028 144.9944 0.00016503 -85.6583 0.78721
0.89123 0.98802 5.5201e-05 3.8182 0.012038 1.1736e-05 0.0011541 0.13256 0.0006579 0.13322 0.12102 0 0.038156 0.0389 0 0.88142 0.24293 0.064535 0.0090543 4.185 0.056593 6.7819e-05 0.83347 0.0051982 0.0059352 0.0013848 0.98696 0.99172 2.9857e-06 1.1943e-05 0.13123 0.9476 0.9163 0.0013963 0.99354 0.59827 0.0018812 0.4296 1.8843 1.8837 16.0028 144.9944 0.00016495 -85.6584 0.78821
0.89223 0.98802 5.5201e-05 3.8182 0.012038 1.1749e-05 0.0011541 0.13265 0.0006579 0.1333 0.1211 0 0.03815 0.0389 0 0.88149 0.24296 0.064546 0.0090557 4.1852 0.056601 6.7829e-05 0.83347 0.0051985 0.0059355 0.0013848 0.98696 0.99172 2.9857e-06 1.1943e-05 0.13123 0.94772 0.91636 0.0013963 0.99356 0.59841 0.0018812 0.42961 1.8847 1.8841 16.0027 144.9944 0.00016487 -85.6585 0.78921
0.89323 0.98802 5.5201e-05 3.8182 0.012038 1.1762e-05 0.0011541 0.13273 0.00065791 0.13338 0.12117 0 0.038145 0.0389 0 0.88156 0.24299 0.064556 0.009057 4.1855 0.056609 6.784e-05 0.83346 0.0051987 0.0059358 0.0013847 0.98696 0.99172 2.9857e-06 1.1943e-05 0.13124 0.94783 0.91641 0.0013963 0.99358 0.59855 0.0018812 0.42963 1.8851 1.8845 16.0027 144.9944 0.00016478 -85.6586 0.79021
0.89423 0.98802 5.5201e-05 3.8182 0.012038 1.1775e-05 0.0011541 0.13281 0.00065791 0.13346 0.12125 0 0.038139 0.0389 0 0.88162 0.24302 0.064567 0.0090584 4.1857 0.056618 6.785e-05 0.83345 0.005199 0.005936 0.0013847 0.98696 0.99172 2.9856e-06 1.1942e-05 0.13124 0.94794 0.91646 0.0013963 0.99361 0.59869 0.0018811 0.42964 1.8855 1.8849 16.0027 144.9944 0.0001647 -85.6587 0.79121
0.89523 0.98802 5.5201e-05 3.8182 0.012038 1.1788e-05 0.0011541 0.13289 0.00065791 0.13355 0.12133 0 0.038133 0.0389 0 0.88169 0.24305 0.064578 0.0090597 4.1859 0.056626 6.786e-05 0.83344 0.0051993 0.0059363 0.0013847 0.98696 0.99172 2.9856e-06 1.1942e-05 0.13124 0.94805 0.91651 0.0013962 0.99363 0.59883 0.0018811 0.42965 1.8859 1.8853 16.0027 144.9945 0.00016462 -85.6587 0.79221
0.89623 0.98802 5.5201e-05 3.8182 0.012038 1.1801e-05 0.0011541 0.13298 0.00065791 0.13363 0.1214 0 0.038128 0.0389 0 0.88176 0.24308 0.064589 0.0090611 4.1862 0.056634 6.7871e-05 0.83343 0.0051995 0.0059366 0.0013847 0.98696 0.99172 2.9855e-06 1.1942e-05 0.13124 0.94816 0.91657 0.0013962 0.99365 0.59897 0.0018811 0.42966 1.8863 1.8857 16.0026 144.9945 0.00016454 -85.6588 0.79321
0.89723 0.98802 5.5201e-05 3.8182 0.012038 1.1814e-05 0.0011541 0.13306 0.00065791 0.13371 0.12148 0 0.038122 0.0389 0 0.88183 0.24311 0.0646 0.0090624 4.1864 0.056642 6.7881e-05 0.83343 0.0051998 0.0059369 0.0013847 0.98696 0.99172 2.9855e-06 1.1942e-05 0.13124 0.94827 0.91662 0.0013962 0.99368 0.59911 0.0018811 0.42968 1.8867 1.8861 16.0026 144.9945 0.00016445 -85.6589 0.79421
0.89823 0.98802 5.5201e-05 3.8182 0.012038 1.1828e-05 0.0011541 0.13314 0.00065792 0.13379 0.12156 0 0.038117 0.0389 0 0.8819 0.24314 0.064611 0.0090638 4.1867 0.05665 6.7891e-05 0.83342 0.0052001 0.0059371 0.0013846 0.98696 0.99172 2.9854e-06 1.1942e-05 0.13125 0.94838 0.91667 0.0013962 0.9937 0.59925 0.0018811 0.42969 1.8871 1.8865 16.0026 144.9945 0.00016437 -85.659 0.79521
0.89923 0.98802 5.5201e-05 3.8182 0.012038 1.1841e-05 0.0011541 0.13322 0.00065792 0.13388 0.12163 0 0.038111 0.0389 0 0.88196 0.24317 0.064622 0.0090651 4.1869 0.056658 6.7902e-05 0.83341 0.0052003 0.0059374 0.0013846 0.98696 0.99172 2.9854e-06 1.1941e-05 0.13125 0.94849 0.91672 0.0013962 0.99372 0.59939 0.0018811 0.4297 1.8875 1.8869 16.0025 144.9945 0.00016429 -85.6591 0.79621
0.90023 0.98802 5.52e-05 3.8182 0.012038 1.1854e-05 0.0011541 0.1333 0.00065792 0.13396 0.12171 0 0.038105 0.0389 0 0.88203 0.2432 0.064633 0.0090665 4.1871 0.056666 6.7914e-05 0.8334 0.0052006 0.0059377 0.0013846 0.98696 0.99172 2.9853e-06 1.1941e-05 0.13125 0.9486 0.91677 0.0013962 0.99374 0.59953 0.0018811 0.42971 1.8879 1.8873 16.0025 144.9946 0.00016421 -85.6592 0.79721
0.90123 0.98802 5.52e-05 3.8182 0.012038 1.1867e-05 0.0011541 0.13339 0.00065792 0.13404 0.12179 0 0.0381 0.0389 0 0.8821 0.24324 0.064644 0.0090678 4.1874 0.056675 6.7922e-05 0.83339 0.0052009 0.0059379 0.0013846 0.98697 0.99172 2.9853e-06 1.1941e-05 0.13125 0.94871 0.91682 0.0013962 0.99377 0.59967 0.0018811 0.42972 1.8883 1.8877 16.0025 144.9946 0.00016413 -85.6592 0.79821
0.90223 0.98802 5.52e-05 3.8182 0.012038 1.188e-05 0.0011541 0.13347 0.00065792 0.13412 0.12186 0 0.038094 0.0389 0 0.88217 0.24327 0.064655 0.0090692 4.1876 0.056683 6.7933e-05 0.83339 0.0052011 0.0059382 0.0013846 0.98697 0.99172 2.9853e-06 1.1941e-05 0.13126 0.94882 0.91688 0.0013962 0.99379 0.59981 0.001881 0.42974 1.8887 1.8881 16.0024 144.9946 0.00016405 -85.6593 0.79921
0.90323 0.98802 5.52e-05 3.8182 0.012038 1.1893e-05 0.0011541 0.13355 0.00065793 0.1342 0.12194 0 0.038089 0.0389 0 0.88224 0.2433 0.064665 0.0090705 4.1879 0.056691 6.7947e-05 0.83338 0.0052014 0.0059385 0.0013845 0.98697 0.99172 2.9852e-06 1.1941e-05 0.13126 0.94893 0.91693 0.0013962 0.99381 0.59995 0.001881 0.42975 1.889 1.8885 16.0024 144.9946 0.00016397 -85.6594 0.80021
0.90423 0.98802 5.52e-05 3.8182 0.012038 1.1907e-05 0.0011541 0.13363 0.00065793 0.13429 0.12202 0 0.038083 0.0389 0 0.88231 0.24333 0.064676 0.0090719 4.1881 0.056699 6.7954e-05 0.83337 0.0052017 0.0059387 0.0013845 0.98697 0.99172 2.9852e-06 1.1941e-05 0.13126 0.94904 0.91698 0.0013962 0.99383 0.60009 0.001881 0.42976 1.8894 1.8888 16.0024 144.9946 0.00016389 -85.6595 0.80121
0.90523 0.98802 5.52e-05 3.8182 0.012038 1.192e-05 0.0011541 0.13371 0.00065793 0.13437 0.12209 0 0.038078 0.0389 0 0.88238 0.24336 0.064687 0.0090732 4.1884 0.056707 6.7965e-05 0.83336 0.005202 0.005939 0.0013845 0.98697 0.99172 2.9851e-06 1.194e-05 0.13126 0.94915 0.91703 0.0013961 0.99385 0.60023 0.001881 0.42977 1.8898 1.8892 16.0024 144.9947 0.00016381 -85.6596 0.80221
0.90623 0.98802 5.52e-05 3.8182 0.012038 1.1933e-05 0.0011541 0.1338 0.00065793 0.13445 0.12217 0 0.038072 0.0389 0 0.88244 0.24339 0.064698 0.0090746 4.1886 0.056716 6.7978e-05 0.83335 0.0052022 0.0059393 0.0013845 0.98697 0.99172 2.9851e-06 1.194e-05 0.13126 0.94925 0.91708 0.0013961 0.99387 0.60036 0.001881 0.42979 1.8902 1.8896 16.0023 144.9947 0.00016373 -85.6596 0.80321
0.90723 0.98802 5.52e-05 3.8182 0.012038 1.1946e-05 0.0011541 0.13388 0.00065793 0.13453 0.12224 0 0.038067 0.0389 0 0.88251 0.24342 0.064709 0.0090759 4.1888 0.056724 6.7986e-05 0.83334 0.0052025 0.0059396 0.0013845 0.98697 0.99172 2.985e-06 1.194e-05 0.13127 0.94936 0.91713 0.0013961 0.9939 0.6005 0.001881 0.4298 1.8906 1.89 16.0023 144.9947 0.00016365 -85.6597 0.80421
0.90823 0.98802 5.52e-05 3.8182 0.012038 1.1959e-05 0.0011541 0.13396 0.00065794 0.13461 0.12232 0 0.038061 0.0389 0 0.88258 0.24345 0.06472 0.0090773 4.1891 0.056732 6.7995e-05 0.83334 0.0052028 0.0059398 0.0013845 0.98697 0.99172 2.985e-06 1.194e-05 0.13127 0.94947 0.91718 0.0013961 0.99392 0.60064 0.001881 0.42981 1.891 1.8904 16.0023 144.9947 0.00016357 -85.6598 0.80521
0.90923 0.98802 5.52e-05 3.8182 0.012038 1.1972e-05 0.0011541 0.13404 0.00065794 0.13469 0.1224 0 0.038055 0.0389 0 0.88265 0.24348 0.064731 0.0090786 4.1893 0.05674 6.8008e-05 0.83333 0.0052031 0.0059401 0.0013844 0.98697 0.99172 2.985e-06 1.194e-05 0.13127 0.94957 0.91723 0.0013961 0.99394 0.60078 0.0018809 0.42982 1.8914 1.8908 16.0022 144.9947 0.0001635 -85.6599 0.80621
0.91023 0.98802 5.52e-05 3.8182 0.012038 1.1985e-05 0.0011541 0.13412 0.00065794 0.13477 0.12247 0 0.03805 0.0389 0 0.88272 0.24351 0.064742 0.00908 4.1896 0.056748 6.8018e-05 0.83332 0.0052033 0.0059404 0.0013844 0.98697 0.99172 2.9849e-06 1.194e-05 0.13127 0.94968 0.91728 0.0013961 0.99396 0.60092 0.0018809 0.42983 1.8918 1.8912 16.0022 144.9948 0.00016342 -85.66 0.80721
0.91123 0.98802 5.52e-05 3.8182 0.012038 1.1999e-05 0.0011541 0.1342 0.00065794 0.13486 0.12255 0 0.038044 0.0389 0 0.88279 0.24354 0.064753 0.0090814 4.1898 0.056757 6.8028e-05 0.83331 0.0052036 0.0059407 0.0013844 0.98697 0.99172 2.9849e-06 1.1939e-05 0.13128 0.94979 0.91733 0.0013961 0.99398 0.60106 0.0018809 0.42985 1.8922 1.8916 16.0022 144.9948 0.00016334 -85.66 0.80821
0.91223 0.98802 5.52e-05 3.8182 0.012038 1.2012e-05 0.0011541 0.13428 0.00065794 0.13494 0.12262 0 0.038039 0.0389 0 0.88286 0.24357 0.064764 0.0090827 4.1901 0.056765 6.8039e-05 0.8333 0.0052039 0.0059409 0.0013844 0.98697 0.99172 2.9848e-06 1.1939e-05 0.13128 0.94989 0.91738 0.0013961 0.994 0.6012 0.0018809 0.42986 1.8925 1.892 16.0022 144.9948 0.00016326 -85.6601 0.80921
0.91323 0.98802 5.52e-05 3.8182 0.012038 1.2025e-05 0.0011541 0.13437 0.00065795 0.13502 0.1227 0 0.038033 0.0389 0 0.88293 0.2436 0.064775 0.0090841 4.1903 0.056773 6.8049e-05 0.83329 0.0052042 0.0059412 0.0013844 0.98697 0.99172 2.9848e-06 1.1939e-05 0.13128 0.95 0.91743 0.0013961 0.99402 0.60134 0.0018809 0.42987 1.8929 1.8923 16.0021 144.9948 0.00016318 -85.6602 0.81021
0.91423 0.98802 5.52e-05 3.8182 0.012038 1.2038e-05 0.0011541 0.13445 0.00065795 0.1351 0.12277 0 0.038028 0.0389 0 0.88299 0.24363 0.064786 0.0090854 4.1906 0.056781 6.806e-05 0.83329 0.0052044 0.0059415 0.0013843 0.98697 0.99172 2.9848e-06 1.1939e-05 0.13128 0.9501 0.91747 0.0013961 0.99404 0.60148 0.0018809 0.42988 1.8933 1.8927 16.0021 144.9949 0.00016311 -85.6603 0.81121
0.91523 0.98802 5.52e-05 3.8182 0.012038 1.2051e-05 0.0011541 0.13453 0.00065795 0.13518 0.12285 0 0.038022 0.0389 0 0.88306 0.24366 0.064797 0.0090868 4.1908 0.05679 6.807e-05 0.83328 0.0052047 0.0059418 0.0013843 0.98697 0.99172 2.9847e-06 1.1939e-05 0.13128 0.95021 0.91752 0.0013961 0.99406 0.60161 0.0018809 0.4299 1.8937 1.8931 16.0021 144.9949 0.00016303 -85.6603 0.81221
0.91623 0.98802 5.5199e-05 3.8182 0.012038 1.2064e-05 0.0011541 0.13461 0.00065795 0.13526 0.12293 0 0.038017 0.0389 0 0.88313 0.24369 0.064808 0.0090882 4.1911 0.056798 6.8081e-05 0.83327 0.005205 0.005942 0.0013843 0.98697 0.99172 2.9847e-06 1.1939e-05 0.13129 0.95031 0.91757 0.001396 0.99408 0.60175 0.0018809 0.42991 1.8941 1.8935 16.002 144.9949 0.00016295 -85.6604 0.81321
0.91723 0.98802 5.5199e-05 3.8182 0.012038 1.2077e-05 0.0011541 0.13469 0.00065795 0.13534 0.123 0 0.038011 0.0389 0 0.8832 0.24372 0.064819 0.0090895 4.1913 0.056806 6.8092e-05 0.83326 0.0052053 0.0059423 0.0013843 0.98697 0.99172 2.9846e-06 1.1938e-05 0.13129 0.95041 0.91762 0.001396 0.9941 0.60189 0.0018809 0.42992 1.8945 1.8939 16.002 144.9949 0.00016288 -85.6605 0.81421
0.91823 0.98802 5.5199e-05 3.8182 0.012038 1.2091e-05 0.0011541 0.13477 0.00065796 0.13542 0.12308 0 0.038006 0.0389 0 0.88327 0.24375 0.06483 0.0090909 4.1916 0.056814 6.8102e-05 0.83325 0.0052055 0.0059426 0.0013843 0.98697 0.99172 2.9846e-06 1.1938e-05 0.13129 0.95052 0.91767 0.001396 0.99412 0.60203 0.0018808 0.42993 1.8948 1.8943 16.002 144.9949 0.0001628 -85.6606 0.81521
0.91923 0.98802 5.5199e-05 3.8182 0.012038 1.2104e-05 0.0011541 0.13485 0.00065796 0.1355 0.12315 0 0.038 0.0389 0 0.88334 0.24378 0.064841 0.0090923 4.1918 0.056823 6.8113e-05 0.83325 0.0052058 0.0059429 0.0013843 0.98697 0.99172 2.9846e-06 1.1938e-05 0.13129 0.95062 0.91772 0.001396 0.99414 0.60217 0.0018808 0.42994 1.8952 1.8946 16.0019 144.995 0.00016273 -85.6606 0.81621
0.92023 0.98802 5.5199e-05 3.8182 0.012038 1.2117e-05 0.0011541 0.13493 0.00065796 0.13559 0.12323 0 0.037995 0.0389 0 0.88341 0.24381 0.064852 0.0090936 4.1921 0.056831 6.8123e-05 0.83324 0.0052061 0.0059431 0.0013842 0.98697 0.99172 2.9845e-06 1.1938e-05 0.1313 0.95072 0.91777 0.001396 0.99416 0.60231 0.0018808 0.42996 1.8956 1.895 16.0019 144.995 0.00016265 -85.6607 0.81721
0.92123 0.98802 5.5199e-05 3.8182 0.012038 1.213e-05 0.0011541 0.13501 0.00065796 0.13567 0.1233 0 0.03799 0.0389 0 0.88348 0.24384 0.064863 0.009095 4.1923 0.056839 6.8134e-05 0.83323 0.0052064 0.0059434 0.0013842 0.98697 0.99172 2.9845e-06 1.1938e-05 0.1313 0.95083 0.91781 0.001396 0.99418 0.60245 0.0018808 0.42997 1.896 1.8954 16.0019 144.995 0.00016258 -85.6608 0.81821
0.92223 0.98802 5.5199e-05 3.8182 0.012038 1.2143e-05 0.0011541 0.13509 0.00065796 0.13575 0.12338 0 0.037984 0.0389 0 0.88355 0.24388 0.064874 0.0090964 4.1926 0.056848 6.8144e-05 0.83322 0.0052066 0.0059437 0.0013842 0.98697 0.99172 2.9844e-06 1.1938e-05 0.1313 0.95093 0.91786 0.001396 0.9942 0.60258 0.0018808 0.42998 1.8964 1.8958 16.0019 144.995 0.0001625 -85.6608 0.81921
0.92323 0.98802 5.5199e-05 3.8182 0.012038 1.2156e-05 0.0011541 0.13517 0.00065797 0.13583 0.12345 0 0.037979 0.0389 0 0.88362 0.24391 0.064886 0.0090977 4.1928 0.056856 6.8155e-05 0.83321 0.0052069 0.005944 0.0013842 0.98697 0.99172 2.9844e-06 1.1938e-05 0.1313 0.95103 0.91791 0.001396 0.99422 0.60272 0.0018808 0.42999 1.8967 1.8962 16.0018 144.995 0.00016243 -85.6609 0.82021
0.92423 0.98802 5.5199e-05 3.8182 0.012038 1.2169e-05 0.0011541 0.13525 0.00065797 0.13591 0.12353 0 0.037973 0.0389 0 0.88369 0.24394 0.064897 0.0090991 4.1931 0.056864 6.8166e-05 0.8332 0.0052072 0.0059443 0.0013842 0.98697 0.99172 2.9844e-06 1.1937e-05 0.13131 0.95113 0.91796 0.001396 0.99424 0.60286 0.0018808 0.43001 1.8971 1.8965 16.0018 144.9951 0.00016235 -85.661 0.82121
0.92523 0.98802 5.5199e-05 3.8182 0.012038 1.2183e-05 0.0011541 0.13533 0.00065797 0.13599 0.1236 0 0.037968 0.0389 0 0.88376 0.24397 0.064908 0.0091005 4.1933 0.056872 6.8176e-05 0.8332 0.0052075 0.0059445 0.0013842 0.98697 0.99172 2.9843e-06 1.1937e-05 0.13131 0.95123 0.918 0.001396 0.99426 0.603 0.0018808 0.43002 1.8975 1.8969 16.0018 144.9951 0.00016228 -85.6611 0.82221
0.92623 0.98802 5.5199e-05 3.8182 0.012038 1.2196e-05 0.0011541 0.13541 0.00065797 0.13607 0.12368 0 0.037962 0.0389 0 0.88382 0.244 0.064919 0.0091018 4.1936 0.056881 6.8187e-05 0.83319 0.0052078 0.0059448 0.0013841 0.98697 0.99172 2.9843e-06 1.1937e-05 0.13131 0.95133 0.91805 0.001396 0.99428 0.60314 0.0018808 0.43003 1.8979 1.8973 16.0017 144.9951 0.0001622 -85.6611 0.82321
0.92723 0.98802 5.5199e-05 3.8182 0.012038 1.2209e-05 0.0011541 0.1355 0.00065797 0.13615 0.12375 0 0.037957 0.0389 0 0.88389 0.24403 0.06493 0.0091032 4.1938 0.056889 6.8198e-05 0.83318 0.005208 0.0059451 0.0013841 0.98697 0.99172 2.9843e-06 1.1937e-05 0.13131 0.95143 0.9181 0.0013959 0.9943 0.60327 0.0018807 0.43004 1.8982 1.8977 16.0017 144.9951 0.00016213 -85.6612 0.82421
0.92823 0.98802 5.5199e-05 3.8182 0.012038 1.2222e-05 0.0011541 0.13558 0.00065797 0.13623 0.12383 0 0.037951 0.0389 0 0.88396 0.24406 0.064941 0.0091046 4.1941 0.056897 6.8208e-05 0.83317 0.0052083 0.0059454 0.0013841 0.98697 0.99172 2.9842e-06 1.1937e-05 0.13132 0.95153 0.91814 0.0013959 0.99432 0.60341 0.0018807 0.43005 1.8986 1.8981 16.0017 144.9951 0.00016206 -85.6613 0.82521
0.92923 0.98802 5.5199e-05 3.8182 0.012038 1.2235e-05 0.0011541 0.13566 0.00065798 0.13631 0.1239 0 0.037946 0.0389 0 0.88403 0.24409 0.064952 0.009106 4.1943 0.056906 6.8219e-05 0.83316 0.0052086 0.0059457 0.0013841 0.98697 0.99172 2.9842e-06 1.1937e-05 0.13132 0.95163 0.91819 0.0013959 0.99434 0.60355 0.0018807 0.43007 1.899 1.8984 16.0016 144.9952 0.00016198 -85.6613 0.82621
0.93023 0.98802 5.5199e-05 3.8182 0.012038 1.2248e-05 0.0011541 0.13574 0.00065798 0.13639 0.12398 0 0.037941 0.0389 0 0.8841 0.24412 0.064963 0.0091073 4.1946 0.056914 6.823e-05 0.83315 0.0052089 0.005946 0.0013841 0.98697 0.99172 2.9842e-06 1.1937e-05 0.13132 0.95173 0.91824 0.0013959 0.99435 0.60369 0.0018807 0.43008 1.8994 1.8988 16.0016 144.9952 0.00016191 -85.6614 0.82721
0.93123 0.98802 5.5199e-05 3.8182 0.012038 1.2262e-05 0.0011541 0.13582 0.00065798 0.13647 0.12405 0 0.037935 0.0389 0 0.88417 0.24415 0.064974 0.0091087 4.1948 0.056922 6.824e-05 0.83315 0.0052092 0.0059462 0.0013841 0.98697 0.99172 2.9841e-06 1.1936e-05 0.13132 0.95183 0.91828 0.0013959 0.99437 0.60383 0.0018807 0.43009 1.8997 1.8992 16.0016 144.9952 0.00016184 -85.6615 0.82821
0.93223 0.98802 5.5198e-05 3.8182 0.012038 1.2275e-05 0.0011541 0.1359 0.00065798 0.13655 0.12413 0 0.03793 0.0389 0 0.88424 0.24418 0.064985 0.0091101 4.1951 0.056931 6.8251e-05 0.83314 0.0052095 0.0059465 0.0013841 0.98697 0.99172 2.9841e-06 1.1936e-05 0.13132 0.95193 0.91833 0.0013959 0.99439 0.60396 0.0018807 0.4301 1.9001 1.8995 16.0015 144.9952 0.00016176 -85.6615 0.82921
0.93323 0.98802 5.5198e-05 3.8182 0.012038 1.2288e-05 0.0011541 0.13598 0.00065798 0.13663 0.1242 0 0.037924 0.0389 0 0.88431 0.24421 0.064997 0.0091115 4.1954 0.056939 6.8261e-05 0.83313 0.0052097 0.0059468 0.001384 0.98697 0.99172 2.9841e-06 1.1936e-05 0.13133 0.95203 0.91838 0.0013959 0.99441 0.6041 0.0018807 0.43011 1.9005 1.8999 16.0015 144.9952 0.00016169 -85.6616 0.83021
0.93423 0.98802 5.5198e-05 3.8182 0.012038 1.2301e-05 0.0011541 0.13606 0.00065799 0.13671 0.12427 0 0.037919 0.0389 0 0.88438 0.24424 0.065008 0.0091128 4.1956 0.056947 6.8272e-05 0.83312 0.00521 0.0059471 0.001384 0.98697 0.99172 2.984e-06 1.1936e-05 0.13133 0.95213 0.91842 0.0013959 0.99443 0.60424 0.0018807 0.43013 1.9009 1.9003 16.0015 144.9953 0.00016162 -85.6617 0.83121
0.93523 0.98802 5.5198e-05 3.8182 0.012038 1.2314e-05 0.0011541 0.13614 0.00065799 0.13679 0.12435 0 0.037914 0.0389 0 0.88445 0.24428 0.065019 0.0091142 4.1959 0.056956 6.8283e-05 0.83311 0.0052103 0.0059474 0.001384 0.98697 0.99172 2.984e-06 1.1936e-05 0.13133 0.95223 0.91847 0.0013959 0.99444 0.60438 0.0018807 0.43014 1.9012 1.9007 16.0015 144.9953 0.00016155 -85.6617 0.83221
0.93623 0.98802 5.5198e-05 3.8182 0.012038 1.2327e-05 0.0011541 0.13621 0.00065799 0.13687 0.12442 0 0.037908 0.0389 0 0.88452 0.24431 0.06503 0.0091156 4.1961 0.056964 6.8294e-05 0.8331 0.0052106 0.0059477 0.001384 0.98697 0.99172 2.984e-06 1.1936e-05 0.13133 0.95233 0.91851 0.0013959 0.99446 0.60452 0.0018806 0.43015 1.9016 1.901 16.0014 144.9953 0.00016148 -85.6618 0.83321
0.93723 0.98802 5.5198e-05 3.8182 0.012038 1.234e-05 0.0011541 0.13629 0.00065799 0.13695 0.1245 0 0.037903 0.0389 0 0.88459 0.24434 0.065041 0.009117 4.1964 0.056972 6.8304e-05 0.8331 0.0052109 0.0059479 0.001384 0.98697 0.99172 2.9839e-06 1.1936e-05 0.13134 0.95242 0.91856 0.0013959 0.99448 0.60465 0.0018806 0.43016 1.902 1.9014 16.0014 144.9953 0.0001614 -85.6619 0.83421
0.93823 0.98802 5.5198e-05 3.8182 0.012038 1.2354e-05 0.0011541 0.13637 0.00065799 0.13703 0.12457 0 0.037898 0.0389 0 0.88466 0.24437 0.065052 0.0091183 4.1966 0.056981 6.8315e-05 0.83309 0.0052112 0.0059482 0.001384 0.98697 0.99172 2.9839e-06 1.1935e-05 0.13134 0.95252 0.9186 0.0013959 0.9945 0.60479 0.0018806 0.43017 1.9023 1.9018 16.0014 144.9953 0.00016133 -85.6619 0.83521
0.93923 0.98802 5.5198e-05 3.8182 0.012038 1.2367e-05 0.0011541 0.13645 0.000658 0.13711 0.12465 0 0.037892 0.0389 0 0.88473 0.2444 0.065063 0.0091197 4.1969 0.056989 6.8326e-05 0.83308 0.0052114 0.0059485 0.001384 0.98697 0.99172 2.9839e-06 1.1935e-05 0.13134 0.95262 0.91865 0.0013959 0.99451 0.60493 0.0018806 0.43019 1.9027 1.9021 16.0013 144.9954 0.00016126 -85.662 0.83621
0.94023 0.98802 5.5198e-05 3.8182 0.012038 1.238e-05 0.0011541 0.13653 0.000658 0.13719 0.12472 0 0.037887 0.0389 0 0.8848 0.24443 0.065075 0.0091211 4.1972 0.056997 6.8336e-05 0.83307 0.0052117 0.0059488 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13134 0.95271 0.91869 0.0013958 0.99453 0.60507 0.0018806 0.4302 1.9031 1.9025 16.0013 144.9954 0.00016119 -85.662 0.83721
0.94123 0.98802 5.5198e-05 3.8182 0.012038 1.2393e-05 0.0011541 0.13661 0.000658 0.13727 0.12479 0 0.037882 0.0389 0 0.88487 0.24446 0.065086 0.0091225 4.1974 0.057006 6.8348e-05 0.83306 0.005212 0.0059491 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13135 0.95281 0.91874 0.0013958 0.99455 0.6052 0.0018806 0.43021 1.9034 1.9029 16.0013 144.9954 0.00016112 -85.6621 0.83821
0.94223 0.98802 5.5198e-05 3.8182 0.012037 1.2406e-05 0.0011541 0.13669 0.000658 0.13735 0.12487 0 0.037876 0.0389 0 0.88494 0.24449 0.065097 0.0091239 4.1977 0.057014 6.8358e-05 0.83305 0.0052123 0.0059494 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13135 0.95291 0.91878 0.0013958 0.99457 0.60534 0.0018806 0.43022 1.9038 1.9032 16.0012 144.9954 0.00016105 -85.6622 0.83921
0.94323 0.98802 5.5198e-05 3.8182 0.012037 1.2419e-05 0.0011541 0.13677 0.000658 0.13742 0.12494 0 0.037871 0.0389 0 0.88501 0.24452 0.065108 0.0091252 4.1979 0.057023 6.8368e-05 0.83305 0.0052126 0.0059497 0.0013839 0.98697 0.99172 2.9837e-06 1.1935e-05 0.13135 0.953 0.91883 0.0013958 0.99458 0.60548 0.0018806 0.43023 1.9042 1.9036 16.0012 144.9954 0.00016098 -85.6622 0.84021
0.94423 0.98802 5.5198e-05 3.8182 0.012037 1.2432e-05 0.0011541 0.13685 0.000658 0.1375 0.12502 0 0.037866 0.0389 0 0.88508 0.24455 0.065119 0.0091266 4.1982 0.057031 6.838e-05 0.83304 0.0052129 0.0059499 0.0013839 0.98697 0.99172 2.9837e-06 1.1935e-05 0.13135 0.9531 0.91887 0.0013958 0.9946 0.60562 0.0018806 0.43025 1.9045 1.904 16.0012 144.9955 0.00016091 -85.6623 0.84121
0.94523 0.98802 5.5198e-05 3.8182 0.012037 1.2446e-05 0.0011541 0.13693 0.00065801 0.13758 0.12509 0 0.03786 0.0389 0 0.88515 0.24459 0.065131 0.009128 4.1985 0.057039 6.839e-05 0.83303 0.0052132 0.0059502 0.0013839 0.98697 0.99172 2.9837e-06 1.1935e-05 0.13136 0.95319 0.91892 0.0013958 0.99462 0.60575 0.0018806 0.43026 1.9049 1.9043 16.0011 144.9955 0.00016084 -85.6623 0.84221
0.94623 0.98802 5.5198e-05 3.8182 0.012037 1.2459e-05 0.0011541 0.13701 0.00065801 0.13766 0.12516 0 0.037855 0.0389 0 0.88522 0.24462 0.065142 0.0091294 4.1987 0.057048 6.8401e-05 0.83302 0.0052135 0.0059505 0.0013839 0.98697 0.99172 2.9836e-06 1.1934e-05 0.13136 0.95329 0.91896 0.0013958 0.99463 0.60589 0.0018805 0.43027 1.9052 1.9047 16.0011 144.9955 0.00016077 -85.6624 0.84321
0.94723 0.98802 5.5198e-05 3.8182 0.012037 1.2472e-05 0.0011541 0.13709 0.00065801 0.13774 0.12524 0 0.03785 0.0389 0 0.88529 0.24465 0.065153 0.0091308 4.199 0.057056 6.8412e-05 0.83301 0.0052137 0.0059508 0.0013838 0.98697 0.99172 2.9836e-06 1.1934e-05 0.13136 0.95338 0.919 0.0013958 0.99465 0.60603 0.0018805 0.43028 1.9056 1.9051 16.0011 144.9955 0.0001607 -85.6625 0.84421
0.94823 0.98802 5.5197e-05 3.8182 0.012037 1.2485e-05 0.0011541 0.13717 0.00065801 0.13782 0.12531 0 0.037844 0.0389 0 0.88536 0.24468 0.065164 0.0091322 4.1992 0.057065 6.8423e-05 0.833 0.005214 0.0059511 0.0013838 0.98697 0.99172 2.9836e-06 1.1934e-05 0.13136 0.95348 0.91905 0.0013958 0.99467 0.60616 0.0018805 0.43029 1.906 1.9054 16.0011 144.9955 0.00016063 -85.6625 0.84521
0.94923 0.98802 5.5197e-05 3.8182 0.012037 1.2498e-05 0.0011541 0.13725 0.00065801 0.1379 0.12538 0 0.037839 0.0389 0 0.88543 0.24471 0.065176 0.0091336 4.1995 0.057073 6.8433e-05 0.833 0.0052143 0.0059514 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13136 0.95357 0.91909 0.0013958 0.99468 0.6063 0.0018805 0.43031 1.9063 1.9058 16.001 144.9956 0.00016057 -85.6626 0.84621
0.95023 0.98802 5.5197e-05 3.8182 0.012037 1.2511e-05 0.0011541 0.13732 0.00065802 0.13798 0.12546 0 0.037834 0.0389 0 0.8855 0.24474 0.065187 0.0091349 4.1998 0.057081 6.8444e-05 0.83299 0.0052146 0.0059517 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13137 0.95366 0.91913 0.0013958 0.9947 0.60644 0.0018805 0.43032 1.9067 1.9061 16.001 144.9956 0.0001605 -85.6626 0.84721
0.95123 0.98802 5.5197e-05 3.8182 0.012037 1.2524e-05 0.0011541 0.1374 0.00065802 0.13806 0.12553 0 0.037828 0.0389 0 0.88557 0.24477 0.065198 0.0091363 4.2 0.05709 6.8455e-05 0.83298 0.0052149 0.005952 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13137 0.95376 0.91918 0.0013958 0.99471 0.60658 0.0018805 0.43033 1.9071 1.9065 16.001 144.9956 0.00016043 -85.6627 0.84821
0.95223 0.98802 5.5197e-05 3.8182 0.012037 1.2538e-05 0.0011541 0.13748 0.00065802 0.13814 0.1256 0 0.037823 0.0389 0 0.88564 0.2448 0.065209 0.0091377 4.2003 0.057098 6.8466e-05 0.83297 0.0052152 0.0059523 0.0013838 0.98698 0.99172 2.9834e-06 1.1934e-05 0.13137 0.95385 0.91922 0.0013958 0.99473 0.60671 0.0018805 0.43034 1.9074 1.9069 16.0009 144.9956 0.00016036 -85.6628 0.84921
0.95323 0.98802 5.5197e-05 3.8182 0.012037 1.2551e-05 0.0011541 0.13756 0.00065802 0.13821 0.12568 0 0.037818 0.0389 0 0.88571 0.24483 0.065221 0.0091391 4.2006 0.057107 6.8477e-05 0.83296 0.0052155 0.0059526 0.0013838 0.98698 0.99172 2.9834e-06 1.1934e-05 0.13137 0.95394 0.91926 0.0013958 0.99475 0.60685 0.0018805 0.43035 1.9078 1.9072 16.0009 144.9957 0.00016029 -85.6628 0.85021
0.95423 0.98802 5.5197e-05 3.8182 0.012037 1.2564e-05 0.0011541 0.13764 0.00065802 0.13829 0.12575 0 0.037813 0.0389 0 0.88578 0.24487 0.065232 0.0091405 4.2008 0.057115 6.8487e-05 0.83295 0.0052158 0.0059529 0.0013837 0.98698 0.99172 2.9834e-06 1.1933e-05 0.13138 0.95404 0.91931 0.0013957 0.99476 0.60699 0.0018805 0.43037 1.9081 1.9076 16.0009 144.9957 0.00016023 -85.6629 0.85121
0.95523 0.98802 5.5197e-05 3.8182 0.012037 1.2577e-05 0.0011541 0.13772 0.00065802 0.13837 0.12582 0 0.037807 0.0389 0 0.88585 0.2449 0.065243 0.0091419 4.2011 0.057124 6.8498e-05 0.83294 0.0052161 0.0059531 0.0013837 0.98698 0.99172 2.9834e-06 1.1933e-05 0.13138 0.95413 0.91935 0.0013957 0.99478 0.60712 0.0018805 0.43038 1.9085 1.9079 16.0008 144.9957 0.00016016 -85.6629 0.85221
0.95623 0.98802 5.5197e-05 3.8182 0.012037 1.259e-05 0.0011541 0.1378 0.00065803 0.13845 0.1259 0 0.037802 0.0389 0 0.88592 0.24493 0.065254 0.0091433 4.2014 0.057132 6.8509e-05 0.83294 0.0052164 0.0059534 0.0013837 0.98698 0.99172 2.9833e-06 1.1933e-05 0.13138 0.95422 0.91939 0.0013957 0.99479 0.60726 0.0018805 0.43039 1.9088 1.9083 16.0008 144.9957 0.00016009 -85.663 0.85321
0.95723 0.98802 5.5197e-05 3.8182 0.012037 1.2603e-05 0.0011541 0.13787 0.00065803 0.13853 0.12597 0 0.037797 0.0389 0 0.886 0.24496 0.065266 0.0091447 4.2016 0.057141 6.852e-05 0.83293 0.0052167 0.0059537 0.0013837 0.98698 0.99172 2.9833e-06 1.1933e-05 0.13138 0.95431 0.91943 0.0013957 0.99481 0.6074 0.0018804 0.4304 1.9092 1.9087 16.0008 144.9957 0.00016002 -85.663 0.85421
0.95823 0.98802 5.5197e-05 3.8182 0.012037 1.2616e-05 0.0011541 0.13795 0.00065803 0.13861 0.12604 0 0.037792 0.0389 0 0.88607 0.24499 0.065277 0.0091461 4.2019 0.057149 6.8531e-05 0.83292 0.0052169 0.005954 0.0013837 0.98698 0.99172 2.9833e-06 1.1933e-05 0.13139 0.9544 0.91948 0.0013957 0.99482 0.60753 0.0018804 0.43041 1.9096 1.909 16.0007 144.9958 0.00015996 -85.6631 0.85521
0.95923 0.98802 5.5197e-05 3.8182 0.012037 1.263e-05 0.0011541 0.13803 0.00065803 0.13868 0.12612 0 0.037786 0.0389 0 0.88614 0.24502 0.065288 0.0091475 4.2022 0.057158 6.8542e-05 0.83291 0.0052172 0.0059543 0.0013837 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13139 0.95449 0.91952 0.0013957 0.99484 0.60767 0.0018804 0.43043 1.9099 1.9094 16.0007 144.9958 0.00015989 -85.6631 0.85621
0.96023 0.98802 5.5197e-05 3.8182 0.012037 1.2643e-05 0.0011541 0.13811 0.00065803 0.13876 0.12619 0 0.037781 0.0389 0 0.88621 0.24505 0.065299 0.0091489 4.2024 0.057166 6.8552e-05 0.8329 0.0052175 0.0059546 0.0013837 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13139 0.95459 0.91956 0.0013957 0.99486 0.60781 0.0018804 0.43044 1.9103 1.9097 16.0007 144.9958 0.00015983 -85.6632 0.85721
0.96123 0.98802 5.5197e-05 3.8182 0.012037 1.2656e-05 0.0011541 0.13819 0.00065803 0.13884 0.12626 0 0.037776 0.0389 0 0.88628 0.24508 0.065311 0.0091503 4.2027 0.057174 6.8563e-05 0.83289 0.0052178 0.0059549 0.0013837 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13139 0.95468 0.9196 0.0013957 0.99487 0.60794 0.0018804 0.43045 1.9106 1.9101 16.0007 144.9958 0.00015976 -85.6632 0.85821
0.96223 0.98802 5.5197e-05 3.8182 0.012037 1.2669e-05 0.0011541 0.13827 0.00065804 0.13892 0.12634 0 0.037771 0.0389 0 0.88635 0.24512 0.065322 0.0091517 4.203 0.057183 6.8574e-05 0.83289 0.0052181 0.0059552 0.0013836 0.98698 0.99173 2.9832e-06 1.1933e-05 0.1314 0.95477 0.91964 0.0013957 0.99489 0.60808 0.0018804 0.43046 1.911 1.9104 16.0006 144.9958 0.00015969 -85.6633 0.85921
0.96323 0.98802 5.5197e-05 3.8182 0.012037 1.2682e-05 0.0011541 0.13834 0.00065804 0.139 0.12641 0 0.037765 0.0389 0 0.88642 0.24515 0.065333 0.0091531 4.2032 0.057191 6.8585e-05 0.83288 0.0052184 0.0059555 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.1314 0.95486 0.91969 0.0013957 0.9949 0.60822 0.0018804 0.43047 1.9113 1.9108 16.0006 144.9959 0.00015963 -85.6634 0.86021
0.96423 0.98802 5.5196e-05 3.8182 0.012037 1.2695e-05 0.0011541 0.13842 0.00065804 0.13907 0.12648 0 0.03776 0.0389 0 0.88649 0.24518 0.065345 0.0091544 4.2035 0.0572 6.8596e-05 0.83287 0.0052187 0.0059558 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.1314 0.95495 0.91973 0.0013957 0.99492 0.60835 0.0018804 0.43049 1.9117 1.9111 16.0006 144.9959 0.00015956 -85.6634 0.86121
0.96523 0.98802 5.5196e-05 3.8182 0.012037 1.2708e-05 0.0011541 0.1385 0.00065804 0.13915 0.12655 0 0.037755 0.0389 0 0.88656 0.24521 0.065356 0.0091558 4.2038 0.057208 6.8607e-05 0.83286 0.005219 0.0059561 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.1314 0.95503 0.91977 0.0013957 0.99493 0.60849 0.0018804 0.4305 1.912 1.9115 16.0005 144.9959 0.0001595 -85.6635 0.86221
0.96623 0.98802 5.5196e-05 3.8182 0.012037 1.2722e-05 0.0011541 0.13858 0.00065804 0.13923 0.12663 0 0.03775 0.0389 0 0.88663 0.24524 0.065367 0.0091572 4.204 0.057217 6.8618e-05 0.83285 0.0052193 0.0059564 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13141 0.95512 0.91981 0.0013957 0.99494 0.60862 0.0018804 0.43051 1.9124 1.9118 16.0005 144.9959 0.00015943 -85.6635 0.86321
0.96723 0.98802 5.5196e-05 3.8182 0.012037 1.2735e-05 0.0011541 0.13865 0.00065805 0.13931 0.1267 0 0.037745 0.0389 0 0.8867 0.24527 0.065379 0.0091586 4.2043 0.057225 6.8629e-05 0.83284 0.0052196 0.0059567 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13141 0.95521 0.91985 0.0013957 0.99496 0.60876 0.0018804 0.43052 1.9127 1.9122 16.0005 144.9959 0.00015937 -85.6636 0.86421
0.96823 0.98802 5.5196e-05 3.8182 0.012037 1.2748e-05 0.0011541 0.13873 0.00065805 0.13939 0.12677 0 0.037739 0.0389 0 0.88677 0.2453 0.06539 0.00916 4.2046 0.057234 6.8639e-05 0.83283 0.0052199 0.005957 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13141 0.9553 0.91989 0.0013957 0.99497 0.6089 0.0018804 0.43053 1.9131 1.9125 16.0004 144.996 0.0001593 -85.6636 0.86521
0.96923 0.98802 5.5196e-05 3.8182 0.012037 1.2761e-05 0.0011541 0.13881 0.00065805 0.13946 0.12684 0 0.037734 0.0389 0 0.88685 0.24534 0.065401 0.0091614 4.2048 0.057242 6.865e-05 0.83283 0.0052202 0.0059573 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13141 0.95539 0.91993 0.0013956 0.99499 0.60903 0.0018803 0.43055 1.9134 1.9129 16.0004 144.996 0.00015924 -85.6637 0.86621
0.97023 0.98802 5.5196e-05 3.8182 0.012037 1.2774e-05 0.0011541 0.13889 0.00065805 0.13954 0.12692 0 0.037729 0.0389 0 0.88692 0.24537 0.065413 0.0091628 4.2051 0.057251 6.8661e-05 0.83282 0.0052205 0.0059576 0.0013836 0.98698 0.99173 2.9829e-06 1.1932e-05 0.13142 0.95548 0.91997 0.0013956 0.995 0.60917 0.0018803 0.43056 1.9138 1.9132 16.0004 144.996 0.00015918 -85.6637 0.86721
0.97123 0.98802 5.5196e-05 3.8182 0.012037 1.2787e-05 0.0011541 0.13896 0.00065805 0.13962 0.12699 0 0.037724 0.0389 0 0.88699 0.2454 0.065424 0.0091642 4.2054 0.05726 6.8672e-05 0.83281 0.0052208 0.0059579 0.0013835 0.98698 0.99173 2.9829e-06 1.1932e-05 0.13142 0.95557 0.92001 0.0013956 0.99502 0.6093 0.0018803 0.43057 1.9141 1.9136 16.0003 144.996 0.00015911 -85.6638 0.86821
0.97223 0.98802 5.5196e-05 3.8182 0.012037 1.28e-05 0.0011541 0.13904 0.00065805 0.1397 0.12706 0 0.037719 0.0389 0 0.88706 0.24543 0.065436 0.0091657 4.2057 0.057268 6.8683e-05 0.8328 0.0052211 0.0059582 0.0013835 0.98698 0.99173 2.9829e-06 1.1931e-05 0.13142 0.95565 0.92005 0.0013956 0.99503 0.60944 0.0018803 0.43058 1.9145 1.9139 16.0003 144.996 0.00015905 -85.6638 0.86921
0.97323 0.98802 5.5196e-05 3.8182 0.012037 1.2814e-05 0.0011541 0.13912 0.00065806 0.13977 0.12713 0 0.037713 0.0389 0 0.88713 0.24546 0.065447 0.0091671 4.2059 0.057277 6.8694e-05 0.83279 0.0052214 0.0059585 0.0013835 0.98698 0.99173 2.9829e-06 1.1931e-05 0.13142 0.95574 0.92009 0.0013956 0.99504 0.60958 0.0018803 0.43059 1.9148 1.9143 16.0003 144.9961 0.00015898 -85.6639 0.87021
0.97423 0.98802 5.5196e-05 3.8182 0.012037 1.2827e-05 0.0011541 0.1392 0.00065806 0.13985 0.12721 0 0.037708 0.0389 0 0.8872 0.24549 0.065458 0.0091685 4.2062 0.057285 6.8705e-05 0.83278 0.0052217 0.0059588 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13143 0.95583 0.92013 0.0013956 0.99506 0.60971 0.0018803 0.43061 1.9152 1.9146 16.0002 144.9961 0.00015892 -85.6639 0.87121
0.97523 0.98802 5.5196e-05 3.8182 0.012037 1.284e-05 0.0011541 0.13927 0.00065806 0.13993 0.12728 0 0.037703 0.0389 0 0.88727 0.24553 0.06547 0.0091699 4.2065 0.057294 6.8716e-05 0.83278 0.005222 0.0059591 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13143 0.95591 0.92017 0.0013956 0.99507 0.60985 0.0018803 0.43062 1.9155 1.915 16.0002 144.9961 0.00015886 -85.664 0.87221
0.97623 0.98802 5.5196e-05 3.8182 0.012037 1.2853e-05 0.0011541 0.13935 0.00065806 0.14001 0.12735 0 0.037698 0.0389 0 0.88734 0.24556 0.065481 0.0091713 4.2068 0.057302 6.8726e-05 0.83277 0.0052223 0.0059594 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13143 0.956 0.92021 0.0013956 0.99509 0.60998 0.0018803 0.43063 1.9158 1.9153 16.0002 144.9961 0.0001588 -85.664 0.87321
0.97723 0.98802 5.5196e-05 3.8182 0.012037 1.2866e-05 0.0011541 0.13943 0.00065806 0.14008 0.12742 0 0.037693 0.0389 0 0.88741 0.24559 0.065493 0.0091727 4.207 0.057311 6.8739e-05 0.83276 0.0052226 0.0059597 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13143 0.95609 0.92025 0.0013956 0.9951 0.61012 0.0018803 0.43064 1.9162 1.9157 16.0002 144.9961 0.00015873 -85.6641 0.87421
0.97823 0.98802 5.5196e-05 3.8182 0.012037 1.2879e-05 0.0011541 0.13951 0.00065806 0.14016 0.12749 0 0.037688 0.0389 0 0.88749 0.24562 0.065504 0.0091741 4.2073 0.057319 6.8749e-05 0.83275 0.0052229 0.00596 0.0013835 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13144 0.95617 0.92029 0.0013956 0.99511 0.61026 0.0018803 0.43065 1.9165 1.916 16.0001 144.9962 0.00015867 -85.6641 0.87521
0.97923 0.98802 5.5196e-05 3.8182 0.012037 1.2892e-05 0.0011541 0.13958 0.00065807 0.14024 0.12757 0 0.037683 0.0389 0 0.88756 0.24565 0.065515 0.0091755 4.2076 0.057328 6.8758e-05 0.83274 0.0052232 0.0059603 0.0013835 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13144 0.95626 0.92033 0.0013956 0.99513 0.61039 0.0018803 0.43066 1.9169 1.9164 16.0001 144.9962 0.00015861 -85.6641 0.87621
0.98023 0.98802 5.5195e-05 3.8182 0.012037 1.2906e-05 0.0011541 0.13966 0.00065807 0.14031 0.12764 0 0.037677 0.0389 0 0.88763 0.24568 0.065527 0.0091769 4.2079 0.057336 6.8771e-05 0.83273 0.0052235 0.0059606 0.0013834 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13144 0.95634 0.92037 0.0013956 0.99514 0.61053 0.0018803 0.43068 1.9172 1.9167 16.0001 144.9962 0.00015855 -85.6642 0.87721
0.98123 0.98802 5.5195e-05 3.8182 0.012037 1.2919e-05 0.0011541 0.13974 0.00065807 0.14039 0.12771 0 0.037672 0.0389 0 0.8877 0.24571 0.065538 0.0091783 4.2081 0.057345 6.8784e-05 0.83272 0.0052238 0.0059609 0.0013834 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13144 0.95643 0.92041 0.0013956 0.99515 0.61066 0.0018803 0.43069 1.9176 1.917 16 144.9962 0.00015849 -85.6642 0.87821
0.98223 0.98802 5.5195e-05 3.8182 0.012037 1.2932e-05 0.0011541 0.13981 0.00065807 0.14047 0.12778 0 0.037667 0.0389 0 0.88777 0.24575 0.06555 0.0091797 4.2084 0.057354 6.879e-05 0.83272 0.0052241 0.0059612 0.0013834 0.98698 0.99173 2.9826e-06 1.193e-05 0.13145 0.95651 0.92045 0.0013956 0.99517 0.6108 0.0018802 0.4307 1.9179 1.9174 16 144.9962 0.00015842 -85.6643 0.87921
0.98323 0.98802 5.5195e-05 3.8182 0.012037 1.2945e-05 0.0011541 0.13989 0.00065807 0.14054 0.12785 0 0.037662 0.0389 0 0.88784 0.24578 0.065561 0.0091811 4.2087 0.057362 6.8804e-05 0.83271 0.0052244 0.0059615 0.0013834 0.98698 0.99173 2.9826e-06 1.193e-05 0.13145 0.9566 0.92049 0.0013956 0.99518 0.61093 0.0018802 0.43071 1.9182 1.9177 16 144.9963 0.00015836 -85.6643 0.88021
0.98423 0.98802 5.5195e-05 3.8182 0.012037 1.2958e-05 0.0011541 0.13997 0.00065807 0.14062 0.12792 0 0.037657 0.0389 0 0.88792 0.24581 0.065573 0.0091825 4.209 0.057371 6.8818e-05 0.8327 0.0052247 0.0059618 0.0013834 0.98698 0.99173 2.9826e-06 1.193e-05 0.13145 0.95668 0.92053 0.0013956 0.99519 0.61107 0.0018802 0.43072 1.9186 1.9181 15.9999 144.9963 0.0001583 -85.6644 0.88121
0.98523 0.98802 5.5195e-05 3.8182 0.012037 1.2971e-05 0.0011541 0.14004 0.00065808 0.1407 0.128 0 0.037652 0.0389 0 0.88799 0.24584 0.065584 0.009184 4.2092 0.057379 6.8824e-05 0.83269 0.005225 0.0059621 0.0013834 0.98698 0.99173 2.9826e-06 1.193e-05 0.13145 0.95676 0.92057 0.0013956 0.9952 0.6112 0.0018802 0.43074 1.9189 1.9184 15.9999 144.9963 0.00015824 -85.6644 0.88221
0.98623 0.98802 5.5195e-05 3.8182 0.012037 1.2985e-05 0.0011541 0.14012 0.00065808 0.14077 0.12807 0 0.037647 0.0389 0 0.88806 0.24587 0.065595 0.0091854 4.2095 0.057388 6.8835e-05 0.83268 0.0052253 0.0059624 0.0013834 0.98698 0.99173 2.9825e-06 1.193e-05 0.13146 0.95685 0.92061 0.0013956 0.99522 0.61134 0.0018802 0.43075 1.9193 1.9187 15.9999 144.9963 0.00015818 -85.6645 0.88321
0.98723 0.98802 5.5195e-05 3.8182 0.012037 1.2998e-05 0.0011541 0.1402 0.00065808 0.14085 0.12814 0 0.037642 0.0389 0 0.88813 0.24591 0.065607 0.0091868 4.2098 0.057397 6.885e-05 0.83267 0.0052256 0.0059627 0.0013834 0.98698 0.99173 2.9825e-06 1.193e-05 0.13146 0.95693 0.92064 0.0013955 0.99523 0.61147 0.0018802 0.43076 1.9196 1.9191 15.9998 144.9963 0.00015812 -85.6645 0.88421
0.98823 0.98802 5.5195e-05 3.8182 0.012037 1.3011e-05 0.0011541 0.14027 0.00065808 0.14093 0.12821 0 0.037637 0.0389 0 0.8882 0.24594 0.065618 0.0091882 4.2101 0.057405 6.8859e-05 0.83266 0.0052259 0.005963 0.0013834 0.98698 0.99173 2.9825e-06 1.193e-05 0.13146 0.95701 0.92068 0.0013955 0.99524 0.61161 0.0018802 0.43077 1.9199 1.9194 15.9998 144.9964 0.00015806 -85.6645 0.88521
0.98923 0.98802 5.5195e-05 3.8182 0.012037 1.3024e-05 0.0011541 0.14035 0.00065808 0.141 0.12828 0 0.037631 0.0389 0 0.88827 0.24597 0.06563 0.0091896 4.2104 0.057414 6.887e-05 0.83266 0.0052262 0.0059633 0.0013833 0.98698 0.99173 2.9825e-06 1.193e-05 0.13146 0.9571 0.92072 0.0013955 0.99526 0.61174 0.0018802 0.43078 1.9203 1.9198 15.9998 144.9964 0.000158 -85.6646 0.88621
0.99023 0.98802 5.5195e-05 3.8182 0.012037 1.3037e-05 0.0011541 0.14043 0.00065808 0.14108 0.12835 0 0.037626 0.0389 0 0.88835 0.246 0.065641 0.009191 4.2106 0.057422 6.8881e-05 0.83265 0.0052265 0.0059636 0.0013833 0.98698 0.99173 2.9824e-06 1.193e-05 0.13147 0.95718 0.92076 0.0013955 0.99527 0.61188 0.0018802 0.43079 1.9206 1.9201 15.9997 144.9964 0.00015794 -85.6646 0.88721
0.99123 0.98802 5.5195e-05 3.8182 0.012037 1.305e-05 0.0011541 0.1405 0.00065809 0.14116 0.12842 0 0.037621 0.0389 0 0.88842 0.24603 0.065653 0.0091924 4.2109 0.057431 6.8892e-05 0.83264 0.0052268 0.0059639 0.0013833 0.98698 0.99173 2.9824e-06 1.193e-05 0.13147 0.95726 0.9208 0.0013955 0.99528 0.61201 0.0018802 0.43081 1.9209 1.9204 15.9997 144.9964 0.00015788 -85.6647 0.88821
0.99223 0.98802 5.5195e-05 3.8182 0.012037 1.3063e-05 0.0011541 0.14058 0.00065809 0.14123 0.12849 0 0.037616 0.0389 0 0.88849 0.24606 0.065664 0.0091939 4.2112 0.05744 6.8903e-05 0.83263 0.0052272 0.0059643 0.0013833 0.98698 0.99173 2.9824e-06 1.193e-05 0.13147 0.95734 0.92083 0.0013955 0.99529 0.61215 0.0018802 0.43082 1.9213 1.9208 15.9997 144.9965 0.00015782 -85.6647 0.88921
0.99323 0.98802 5.5195e-05 3.8182 0.012037 1.3077e-05 0.0011541 0.14065 0.00065809 0.14131 0.12857 0 0.037611 0.0389 0 0.88856 0.2461 0.065676 0.0091953 4.2115 0.057448 6.8914e-05 0.83262 0.0052275 0.0059646 0.0013833 0.98698 0.99173 2.9824e-06 1.1929e-05 0.13147 0.95743 0.92087 0.0013955 0.9953 0.61228 0.0018802 0.43083 1.9216 1.9211 15.9996 144.9965 0.00015776 -85.6648 0.89021
0.99423 0.98802 5.5195e-05 3.8182 0.012037 1.309e-05 0.0011541 0.14073 0.00065809 0.14138 0.12864 0 0.037606 0.0389 0 0.88863 0.24613 0.065687 0.0091967 4.2118 0.057457 6.8925e-05 0.83261 0.0052278 0.0059649 0.0013833 0.98698 0.99173 2.9824e-06 1.1929e-05 0.13148 0.95751 0.92091 0.0013955 0.99532 0.61242 0.0018802 0.43084 1.9219 1.9214 15.9996 144.9965 0.0001577 -85.6648 0.89121
0.99523 0.98802 5.5195e-05 3.8182 0.012037 1.3103e-05 0.0011541 0.14081 0.00065809 0.14146 0.12871 0 0.037601 0.0389 0 0.88871 0.24616 0.065699 0.0091981 4.212 0.057466 6.8936e-05 0.8326 0.0052281 0.0059652 0.0013833 0.98698 0.99173 2.9823e-06 1.1929e-05 0.13148 0.95759 0.92095 0.0013955 0.99533 0.61255 0.0018802 0.43085 1.9223 1.9218 15.9996 144.9965 0.00015764 -85.6648 0.89221
0.99623 0.98802 5.5194e-05 3.8182 0.012037 1.3116e-05 0.0011541 0.14088 0.00065809 0.14154 0.12878 0 0.037596 0.0389 0 0.88878 0.24619 0.06571 0.0091995 4.2123 0.057474 6.8947e-05 0.83259 0.0052284 0.0059655 0.0013833 0.98698 0.99173 2.9823e-06 1.1929e-05 0.13148 0.95767 0.92098 0.0013955 0.99534 0.61269 0.0018801 0.43087 1.9226 1.9221 15.9995 144.9965 0.00015758 -85.6649 0.89321
0.99723 0.98802 5.5194e-05 3.8182 0.012037 1.3129e-05 0.0011541 0.14096 0.0006581 0.14161 0.12885 0 0.037591 0.0389 0 0.88885 0.24622 0.065722 0.009201 4.2126 0.057483 6.8958e-05 0.83259 0.0052287 0.0059658 0.0013833 0.98698 0.99173 2.9823e-06 1.1929e-05 0.13148 0.95775 0.92102 0.0013955 0.99535 0.61282 0.0018801 0.43088 1.9229 1.9224 15.9995 144.9966 0.00015753 -85.6649 0.89421
0.99823 0.98802 5.5194e-05 3.8182 0.012037 1.3142e-05 0.0011541 0.14103 0.0006581 0.14169 0.12892 0 0.037586 0.0389 0 0.88892 0.24626 0.065733 0.0092024 4.2129 0.057491 6.897e-05 0.83258 0.005229 0.0059661 0.0013833 0.98698 0.99173 2.9823e-06 1.1929e-05 0.13149 0.95783 0.92106 0.0013955 0.99536 0.61296 0.0018801 0.43089 1.9233 1.9228 15.9995 144.9966 0.00015747 -85.665 0.89521
0.99923 0.98802 5.5194e-05 3.8182 0.012037 1.3155e-05 0.0011541 0.14111 0.0006581 0.14176 0.12899 0 0.037581 0.0389 0 0.88899 0.24629 0.065745 0.0092038 4.2132 0.0575 6.8981e-05 0.83257 0.0052293 0.0059664 0.0013833 0.98698 0.99173 2.9823e-06 1.1929e-05 0.13149 0.95791 0.9211 0.0013955 0.99538 0.61309 0.0018801 0.4309 1.9236 1.9231 15.9994 144.9966 0.00015741 -85.665 0.89621
1.0002 0.98802 5.5194e-05 3.8182 0.012037 1.3169e-05 0.0011541 0.14119 0.0006581 0.14184 0.12906 0 0.037576 0.0389 0 0.88907 0.24632 0.065757 0.0092052 4.2135 0.057509 6.8992e-05 0.83256 0.0052296 0.0059667 0.0013832 0.98698 0.99173 2.9822e-06 1.1929e-05 0.13149 0.95799 0.92113 0.0013955 0.99539 0.61323 0.0018801 0.43091 1.9239 1.9234 15.9994 144.9966 0.00015735 -85.665 0.89721
1.0012 0.98802 5.5194e-05 3.8182 0.012037 1.3182e-05 0.0011541 0.14126 0.0006581 0.14192 0.12913 0 0.037571 0.0389 0 0.88914 0.24635 0.065768 0.0092066 4.2137 0.057517 6.9003e-05 0.83255 0.0052299 0.005967 0.0013832 0.98698 0.99173 2.9822e-06 1.1929e-05 0.13149 0.95807 0.92117 0.0013955 0.9954 0.61336 0.0018801 0.43092 1.9243 1.9238 15.9994 144.9966 0.00015729 -85.6651 0.89821
1.0022 0.98802 5.5194e-05 3.8182 0.012037 1.3195e-05 0.0011541 0.14134 0.0006581 0.14199 0.1292 0 0.037566 0.0389 0 0.88921 0.24638 0.06578 0.0092081 4.214 0.057526 6.9014e-05 0.83254 0.0052302 0.0059674 0.0013832 0.98698 0.99173 2.9822e-06 1.1929e-05 0.1315 0.95815 0.92121 0.0013955 0.99541 0.6135 0.0018801 0.43094 1.9246 1.9241 15.9994 144.9967 0.00015724 -85.6651 0.89921
1.0032 0.98802 5.5194e-05 3.8182 0.012037 1.3208e-05 0.0011541 0.14141 0.00065811 0.14207 0.12927 0 0.037561 0.0389 0 0.88928 0.24642 0.065791 0.0092095 4.2143 0.057535 6.9025e-05 0.83253 0.0052306 0.0059677 0.0013832 0.98698 0.99173 2.9822e-06 1.1929e-05 0.1315 0.95823 0.92124 0.0013955 0.99542 0.61363 0.0018801 0.43095 1.9249 1.9244 15.9993 144.9967 0.00015718 -85.6652 0.90021
1.0042 0.98802 5.5194e-05 3.8182 0.012037 1.3221e-05 0.0011541 0.14149 0.00065811 0.14214 0.12934 0 0.037556 0.0389 0 0.88935 0.24645 0.065803 0.0092109 4.2146 0.057544 6.9036e-05 0.83253 0.0052309 0.005968 0.0013832 0.98698 0.99173 2.9821e-06 1.1928e-05 0.1315 0.95831 0.92128 0.0013955 0.99543 0.61377 0.0018801 0.43096 1.9253 1.9248 15.9993 144.9967 0.00015712 -85.6652 0.90121
1.0052 0.98802 5.5194e-05 3.8182 0.012037 1.3234e-05 0.0011541 0.14156 0.00065811 0.14222 0.12941 0 0.037551 0.0389 0 0.88943 0.24648 0.065814 0.0092123 4.2149 0.057552 6.9047e-05 0.83252 0.0052312 0.0059683 0.0013832 0.98698 0.99173 2.9821e-06 1.1928e-05 0.1315 0.95839 0.92132 0.0013955 0.99545 0.6139 0.0018801 0.43097 1.9256 1.9251 15.9993 144.9967 0.00015706 -85.6652 0.90221
1.0062 0.98802 5.5194e-05 3.8182 0.012037 1.3247e-05 0.0011541 0.14164 0.00065811 0.14229 0.12948 0 0.037546 0.0389 0 0.8895 0.24651 0.065826 0.0092138 4.2152 0.057561 6.9059e-05 0.83251 0.0052315 0.0059686 0.0013832 0.98698 0.99173 2.9821e-06 1.1928e-05 0.13151 0.95847 0.92135 0.0013955 0.99546 0.61404 0.0018801 0.43098 1.9259 1.9254 15.9992 144.9967 0.00015701 -85.6653 0.90321
1.0072 0.98802 5.5194e-05 3.8182 0.012037 1.3261e-05 0.0011541 0.14171 0.00065811 0.14237 0.12956 0 0.037541 0.0389 0 0.88957 0.24654 0.065837 0.0092152 4.2155 0.05757 6.907e-05 0.8325 0.0052318 0.0059689 0.0013832 0.98698 0.99173 2.9821e-06 1.1928e-05 0.13151 0.95855 0.92139 0.0013954 0.99547 0.61417 0.0018801 0.43099 1.9262 1.9257 15.9992 144.9968 0.00015695 -85.6653 0.90421
1.0082 0.98802 5.5194e-05 3.8182 0.012037 1.3274e-05 0.0011541 0.14179 0.00065811 0.14244 0.12963 0 0.037536 0.0389 0 0.88964 0.24658 0.065849 0.0092166 4.2157 0.057578 6.9081e-05 0.83249 0.0052321 0.0059692 0.0013832 0.98698 0.99173 2.9821e-06 1.1928e-05 0.13151 0.95862 0.92142 0.0013954 0.99548 0.6143 0.0018801 0.43101 1.9266 1.9261 15.9992 144.9968 0.00015689 -85.6654 0.90521
1.0092 0.98802 5.5194e-05 3.8182 0.012037 1.3287e-05 0.0011541 0.14186 0.00065812 0.14252 0.1297 0 0.037531 0.0389 0 0.88972 0.24661 0.065861 0.009218 4.216 0.057587 6.9092e-05 0.83248 0.0052324 0.0059695 0.0013832 0.98698 0.99173 2.982e-06 1.1928e-05 0.13152 0.9587 0.92146 0.0013954 0.99549 0.61444 0.0018801 0.43102 1.9269 1.9264 15.9991 144.9968 0.00015684 -85.6654 0.90621
1.0102 0.98803 5.5194e-05 3.8182 0.012037 1.33e-05 0.0011541 0.14194 0.00065812 0.14259 0.12977 0 0.037526 0.0389 0 0.88979 0.24664 0.065872 0.0092195 4.2163 0.057596 6.9103e-05 0.83247 0.0052327 0.0059699 0.0013832 0.98698 0.99173 2.982e-06 1.1928e-05 0.13152 0.95878 0.92149 0.0013954 0.9955 0.61457 0.0018801 0.43103 1.9272 1.9267 15.9991 144.9968 0.00015678 -85.6654 0.90721
1.0112 0.98803 5.5194e-05 3.8182 0.012037 1.3313e-05 0.0011541 0.14201 0.00065812 0.14267 0.12984 0 0.037521 0.0389 0 0.88986 0.24667 0.065884 0.0092209 4.2166 0.057604 6.9114e-05 0.83246 0.0052331 0.0059702 0.0013831 0.98698 0.99173 2.982e-06 1.1928e-05 0.13152 0.95886 0.92153 0.0013954 0.99551 0.61471 0.0018801 0.43104 1.9275 1.9271 15.9991 144.9968 0.00015673 -85.6655 0.90821
1.0122 0.98803 5.5193e-05 3.8182 0.012037 1.3326e-05 0.0011541 0.14209 0.00065812 0.14274 0.12991 0 0.037516 0.0389 0 0.88993 0.24671 0.065895 0.0092223 4.2169 0.057613 6.9126e-05 0.83246 0.0052334 0.0059705 0.0013831 0.98698 0.99173 2.982e-06 1.1928e-05 0.13152 0.95893 0.92157 0.0013954 0.99552 0.61484 0.0018801 0.43105 1.9279 1.9274 15.999 144.9969 0.00015667 -85.6655 0.90921
1.0132 0.98803 5.5193e-05 3.8182 0.012037 1.3339e-05 0.0011541 0.14216 0.00065812 0.14282 0.12998 0 0.037511 0.0389 0 0.89001 0.24674 0.065907 0.0092238 4.2172 0.057622 6.9137e-05 0.83245 0.0052337 0.0059708 0.0013831 0.98698 0.99173 2.982e-06 1.1928e-05 0.13153 0.95901 0.9216 0.0013954 0.99553 0.61497 0.00188 0.43106 1.9282 1.9277 15.999 144.9969 0.00015661 -85.6655 0.91021
1.0142 0.98803 5.5193e-05 3.8182 0.012037 1.3353e-05 0.0011541 0.14224 0.00065812 0.14289 0.13005 0 0.037506 0.0389 0 0.89008 0.24677 0.065919 0.0092252 4.2175 0.057631 6.9147e-05 0.83244 0.005234 0.0059711 0.0013831 0.98698 0.99173 2.982e-06 1.1928e-05 0.13153 0.95909 0.92164 0.0013954 0.99554 0.61511 0.00188 0.43108 1.9285 1.928 15.999 144.9969 0.00015656 -85.6656 0.91121
1.0152 0.98803 5.5193e-05 3.8182 0.012037 1.3366e-05 0.0011541 0.14231 0.00065813 0.14297 0.13012 0 0.037501 0.0389 0 0.89015 0.2468 0.06593 0.0092266 4.2178 0.057639 6.9159e-05 0.83243 0.0052343 0.0059714 0.0013831 0.98698 0.99173 2.9819e-06 1.1928e-05 0.13153 0.95916 0.92167 0.0013954 0.99555 0.61524 0.00188 0.43109 1.9288 1.9284 15.9989 144.9969 0.0001565 -85.6656 0.91221
1.0162 0.98803 5.5193e-05 3.8182 0.012036 1.3379e-05 0.0011541 0.14239 0.00065813 0.14304 0.13019 0 0.037496 0.0389 0 0.89023 0.24683 0.065942 0.0092281 4.2181 0.057648 6.9171e-05 0.83242 0.0052346 0.0059718 0.0013831 0.98698 0.99173 2.9819e-06 1.1928e-05 0.13153 0.95924 0.92171 0.0013954 0.99557 0.61538 0.00188 0.4311 1.9292 1.9287 15.9989 144.9969 0.00015645 -85.6656 0.91321
1.0172 0.98803 5.5193e-05 3.8182 0.012036 1.3392e-05 0.0011541 0.14246 0.00065813 0.14312 0.13026 0 0.037491 0.0389 0 0.8903 0.24687 0.065954 0.0092295 4.2184 0.057657 6.918e-05 0.83241 0.0052349 0.0059721 0.0013831 0.98698 0.99173 2.9819e-06 1.1927e-05 0.13154 0.95932 0.92174 0.0013954 0.99558 0.61551 0.00188 0.43111 1.9295 1.929 15.9989 144.997 0.00015639 -85.6657 0.91421
1.0182 0.98803 5.5193e-05 3.8182 0.012036 1.3405e-05 0.0011541 0.14254 0.00065813 0.14319 0.13033 0 0.037486 0.0389 0 0.89037 0.2469 0.065965 0.0092309 4.2186 0.057665 6.9192e-05 0.8324 0.0052353 0.0059724 0.0013831 0.98698 0.99173 2.9819e-06 1.1927e-05 0.13154 0.95939 0.92178 0.0013954 0.99559 0.61564 0.00188 0.43112 1.9298 1.9293 15.9988 144.997 0.00015634 -85.6657 0.91521
1.0192 0.98803 5.5193e-05 3.8182 0.012036 1.3418e-05 0.0011541 0.14261 0.00065813 0.14327 0.13039 0 0.037482 0.0389 0 0.89044 0.24693 0.065977 0.0092324 4.2189 0.057674 6.9204e-05 0.83239 0.0052356 0.0059727 0.0013831 0.98698 0.99173 2.9819e-06 1.1927e-05 0.13154 0.95947 0.92181 0.0013954 0.9956 0.61578 0.00188 0.43113 1.9301 1.9296 15.9988 144.997 0.00015628 -85.6657 0.91621
1.0202 0.98803 5.5193e-05 3.8182 0.012036 1.3431e-05 0.0011541 0.14269 0.00065813 0.14334 0.13046 0 0.037477 0.0389 0 0.89052 0.24696 0.065989 0.0092338 4.2192 0.057683 6.9213e-05 0.83239 0.0052359 0.005973 0.0013831 0.98698 0.99173 2.9818e-06 1.1927e-05 0.13154 0.95954 0.92184 0.0013954 0.99561 0.61591 0.00188 0.43115 1.9304 1.93 15.9988 144.997 0.00015623 -85.6658 0.91721
1.0212 0.98803 5.5193e-05 3.8182 0.012036 1.3445e-05 0.0011541 0.14276 0.00065814 0.14342 0.13053 0 0.037472 0.0389 0 0.89059 0.247 0.066 0.0092352 4.2195 0.057692 6.9225e-05 0.83238 0.0052362 0.0059734 0.0013831 0.98698 0.99173 2.9818e-06 1.1927e-05 0.13155 0.95962 0.92188 0.0013954 0.99562 0.61605 0.00188 0.43116 1.9308 1.9303 15.9987 144.997 0.00015618 -85.6658 0.91821
1.0222 0.98803 5.5193e-05 3.8182 0.012036 1.3458e-05 0.0011541 0.14284 0.00065814 0.14349 0.1306 0 0.037467 0.0389 0 0.89066 0.24703 0.066012 0.0092367 4.2198 0.057701 6.9242e-05 0.83237 0.0052365 0.0059737 0.0013831 0.98698 0.99173 2.9818e-06 1.1927e-05 0.13155 0.95969 0.92191 0.0013954 0.99563 0.61618 0.00188 0.43117 1.9311 1.9306 15.9987 144.9971 0.00015612 -85.6658 0.91921
1.0232 0.98803 5.5193e-05 3.8182 0.012036 1.3471e-05 0.0011541 0.14291 0.00065814 0.14356 0.13067 0 0.037462 0.0389 0 0.89074 0.24706 0.066024 0.0092381 4.2201 0.057709 6.9248e-05 0.83236 0.0052369 0.005974 0.0013831 0.98698 0.99173 2.9818e-06 1.1927e-05 0.13155 0.95977 0.92195 0.0013954 0.99564 0.61631 0.00188 0.43118 1.9314 1.9309 15.9987 144.9971 0.00015607 -85.6659 0.92021
1.0242 0.98803 5.5193e-05 3.8182 0.012036 1.3484e-05 0.0011541 0.14299 0.00065814 0.14364 0.13074 0 0.037457 0.0389 0 0.89081 0.24709 0.066035 0.0092395 4.2204 0.057718 6.9253e-05 0.83235 0.0052372 0.0059743 0.001383 0.98699 0.99173 2.9818e-06 1.1927e-05 0.13155 0.95984 0.92198 0.0013954 0.99565 0.61645 0.00188 0.43119 1.9317 1.9312 15.9986 144.9971 0.00015602 -85.6659 0.92121
1.0252 0.98803 5.5193e-05 3.8182 0.012036 1.3497e-05 0.0011541 0.14306 0.00065814 0.14371 0.13081 0 0.037452 0.0389 0 0.89088 0.24712 0.066047 0.009241 4.2207 0.057727 6.928e-05 0.83234 0.0052375 0.0059746 0.001383 0.98699 0.99173 2.9818e-06 1.1927e-05 0.13156 0.95992 0.92202 0.0013954 0.99566 0.61658 0.00188 0.4312 1.932 1.9316 15.9986 144.9971 0.00015596 -85.6659 0.92221
1.0262 0.98803 5.5193e-05 3.8182 0.012036 1.351e-05 0.0011541 0.14313 0.00065814 0.14379 0.13088 0 0.037447 0.0389 0 0.89095 0.24716 0.066059 0.0092424 4.221 0.057736 6.9283e-05 0.83233 0.0052378 0.005975 0.001383 0.98699 0.99173 2.9817e-06 1.1927e-05 0.13156 0.95999 0.92205 0.0013954 0.99567 0.61671 0.00188 0.43122 1.9324 1.9319 15.9986 144.9971 0.00015591 -85.666 0.92321
1.0272 0.98803 5.5193e-05 3.8182 0.012036 1.3523e-05 0.0011541 0.14321 0.00065814 0.14386 0.13095 0 0.037442 0.0389 0 0.89103 0.24719 0.06607 0.0092439 4.2213 0.057744 6.9284e-05 0.83232 0.0052381 0.0059753 0.001383 0.98699 0.99173 2.9817e-06 1.1927e-05 0.13156 0.96006 0.92208 0.0013954 0.99568 0.61685 0.00188 0.43123 1.9327 1.9322 15.9985 144.9972 0.00015586 -85.666 0.92421
1.0282 0.98803 5.5192e-05 3.8182 0.012036 1.3537e-05 0.0011541 0.14328 0.00065815 0.14394 0.13102 0 0.037437 0.0389 0 0.8911 0.24722 0.066082 0.0092453 4.2216 0.057753 6.931e-05 0.83232 0.0052385 0.0059756 0.001383 0.98699 0.99173 2.9817e-06 1.1927e-05 0.13157 0.96014 0.92212 0.0013954 0.99569 0.61698 0.00188 0.43124 1.933 1.9325 15.9985 144.9972 0.0001558 -85.666 0.92521
1.0292 0.98803 5.5192e-05 3.8182 0.012036 1.355e-05 0.0011541 0.14336 0.00065815 0.14401 0.13109 0 0.037433 0.0389 0 0.89117 0.24725 0.066094 0.0092467 4.2219 0.057762 6.9322e-05 0.83231 0.0052388 0.0059759 0.001383 0.98699 0.99173 2.9817e-06 1.1927e-05 0.13157 0.96021 0.92215 0.0013954 0.9957 0.61711 0.00188 0.43125 1.9333 1.9328 15.9985 144.9972 0.00015575 -85.6661 0.92621
1.0302 0.98803 5.5192e-05 3.8182 0.012036 1.3563e-05 0.0011541 0.14343 0.00065815 0.14408 0.13116 0 0.037428 0.0389 0 0.89125 0.24729 0.066105 0.0092482 4.2222 0.057771 6.932e-05 0.8323 0.0052391 0.0059762 0.001383 0.98699 0.99173 2.9817e-06 1.1927e-05 0.13157 0.96028 0.92218 0.0013953 0.99571 0.61725 0.00188 0.43126 1.9336 1.9331 15.9984 144.9972 0.0001557 -85.6661 0.92721
1.0312 0.98803 5.5192e-05 3.8182 0.012036 1.3576e-05 0.0011541 0.1435 0.00065815 0.14416 0.13123 0 0.037423 0.0389 0 0.89132 0.24732 0.066117 0.0092496 4.2225 0.05778 6.9339e-05 0.83229 0.0052394 0.0059766 0.001383 0.98699 0.99173 2.9817e-06 1.1927e-05 0.13157 0.96036 0.92222 0.0013953 0.99572 0.61738 0.0018799 0.43127 1.9339 1.9335 15.9984 144.9973 0.00015564 -85.6661 0.92821
1.0322 0.98803 5.5192e-05 3.8182 0.012036 1.3589e-05 0.0011541 0.14358 0.00065815 0.14423 0.1313 0 0.037418 0.0389 0 0.89139 0.24735 0.066129 0.0092511 4.2228 0.057788 6.9352e-05 0.83228 0.0052397 0.0059769 0.001383 0.98699 0.99173 2.9816e-06 1.1926e-05 0.13158 0.96043 0.92225 0.0013953 0.99572 0.61751 0.0018799 0.43129 1.9342 1.9338 15.9984 144.9973 0.00015559 -85.6662 0.92921
1.0332 0.98803 5.5192e-05 3.8182 0.012036 1.3602e-05 0.0011541 0.14365 0.00065815 0.1443 0.13136 0 0.037413 0.0389 0 0.89147 0.24738 0.066141 0.0092525 4.2231 0.057797 6.9361e-05 0.83227 0.0052401 0.0059772 0.001383 0.98699 0.99173 2.9816e-06 1.1926e-05 0.13158 0.9605 0.92228 0.0013953 0.99573 0.61765 0.0018799 0.4313 1.9346 1.9341 15.9983 144.9973 0.00015554 -85.6662 0.93021
1.0342 0.98803 5.5192e-05 3.8182 0.012036 1.3615e-05 0.0011541 0.14372 0.00065816 0.14438 0.13143 0 0.037408 0.0389 0 0.89154 0.24742 0.066152 0.009254 4.2234 0.057806 6.9375e-05 0.83226 0.0052404 0.0059775 0.001383 0.98699 0.99173 2.9816e-06 1.1926e-05 0.13158 0.96057 0.92232 0.0013953 0.99574 0.61778 0.0018799 0.43131 1.9349 1.9344 15.9983 144.9973 0.00015549 -85.6662 0.93121
1.0352 0.98803 5.5192e-05 3.8182 0.012036 1.3629e-05 0.0011541 0.1438 0.00065816 0.14445 0.1315 0 0.037403 0.0389 0 0.89161 0.24745 0.066164 0.0092554 4.2237 0.057815 6.9386e-05 0.83225 0.0052407 0.0059779 0.001383 0.98699 0.99173 2.9816e-06 1.1926e-05 0.13158 0.96064 0.92235 0.0013953 0.99575 0.61791 0.0018799 0.43132 1.9352 1.9347 15.9983 144.9973 0.00015544 -85.6663 0.93221
1.0362 0.98803 5.5192e-05 3.8182 0.012036 1.3642e-05 0.0011541 0.14387 0.00065816 0.14453 0.13157 0 0.037399 0.0389 0 0.89169 0.24748 0.066176 0.0092568 4.224 0.057824 6.9394e-05 0.83225 0.005241 0.0059782 0.001383 0.98699 0.99173 2.9816e-06 1.1926e-05 0.13159 0.96072 0.92238 0.0013953 0.99576 0.61804 0.0018799 0.43133 1.9355 1.935 15.9982 144.9974 0.00015539 -85.6663 0.93321
1.0372 0.98803 5.5192e-05 3.8182 0.012036 1.3655e-05 0.0011541 0.14395 0.00065816 0.1446 0.13164 0 0.037394 0.0389 0 0.89176 0.24751 0.066188 0.0092583 4.2243 0.057832 6.9407e-05 0.83224 0.0052414 0.0059785 0.0013829 0.98699 0.99173 2.9816e-06 1.1926e-05 0.13159 0.96079 0.92241 0.0013953 0.99577 0.61818 0.0018799 0.43134 1.9358 1.9353 15.9982 144.9974 0.00015533 -85.6663 0.93421
1.0382 0.98803 5.5192e-05 3.8182 0.012036 1.3668e-05 0.0011541 0.14402 0.00065816 0.14467 0.13171 0 0.037389 0.0389 0 0.89183 0.24755 0.066199 0.0092597 4.2246 0.057841 6.942e-05 0.83223 0.0052417 0.0059788 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.13159 0.96086 0.92245 0.0013953 0.99578 0.61831 0.0018799 0.43136 1.9361 1.9357 15.9982 144.9974 0.00015528 -85.6663 0.93521
1.0392 0.98803 5.5192e-05 3.8182 0.012036 1.3681e-05 0.0011541 0.14409 0.00065816 0.14475 0.13178 0 0.037384 0.0389 0 0.89191 0.24758 0.066211 0.0092612 4.2249 0.05785 6.9429e-05 0.83222 0.005242 0.0059792 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.13159 0.96093 0.92248 0.0013953 0.99579 0.61844 0.0018799 0.43137 1.9364 1.936 15.9981 144.9974 0.00015523 -85.6664 0.93621
1.0402 0.98803 5.5192e-05 3.8182 0.012036 1.3694e-05 0.0011541 0.14417 0.00065816 0.14482 0.13184 0 0.037379 0.0389 0 0.89198 0.24761 0.066223 0.0092626 4.2252 0.057859 6.944e-05 0.83221 0.0052423 0.0059795 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.1316 0.961 0.92251 0.0013953 0.9958 0.61858 0.0018799 0.43138 1.9367 1.9363 15.9981 144.9974 0.00015518 -85.6664 0.93721
1.0412 0.98803 5.5192e-05 3.8182 0.012036 1.3707e-05 0.0011541 0.14424 0.00065817 0.14489 0.13191 0 0.037375 0.0389 0 0.89206 0.24765 0.066235 0.0092641 4.2255 0.057868 6.9454e-05 0.8322 0.0052427 0.0059798 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.1316 0.96107 0.92254 0.0013953 0.99581 0.61871 0.0018799 0.43139 1.9371 1.9366 15.9981 144.9975 0.00015513 -85.6664 0.93821
1.0422 0.98803 5.5192e-05 3.8182 0.012036 1.3721e-05 0.0011541 0.14431 0.00065817 0.14497 0.13198 0 0.03737 0.0389 0 0.89213 0.24768 0.066247 0.0092655 4.2258 0.057877 6.9463e-05 0.83219 0.005243 0.0059802 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.1316 0.96114 0.92258 0.0013953 0.99582 0.61884 0.0018799 0.4314 1.9374 1.9369 15.998 144.9975 0.00015508 -85.6665 0.93921
1.0432 0.98803 5.5192e-05 3.8182 0.012036 1.3734e-05 0.0011541 0.14439 0.00065817 0.14504 0.13205 0 0.037365 0.0389 0 0.8922 0.24771 0.066258 0.009267 4.2261 0.057886 6.9474e-05 0.83218 0.0052433 0.0059805 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.13161 0.96121 0.92261 0.0013953 0.99583 0.61897 0.0018799 0.43141 1.9377 1.9372 15.998 144.9975 0.00015503 -85.6665 0.94021
1.0442 0.98803 5.5191e-05 3.8182 0.012036 1.3747e-05 0.0011541 0.14446 0.00065817 0.14511 0.13212 0 0.03736 0.0389 0 0.89228 0.24774 0.06627 0.0092684 4.2264 0.057894 6.9487e-05 0.83218 0.0052436 0.0059808 0.0013829 0.98699 0.99173 2.9815e-06 1.1926e-05 0.13161 0.96128 0.92264 0.0013953 0.99583 0.61911 0.0018799 0.43142 1.938 1.9375 15.998 144.9975 0.00015498 -85.6665 0.94121
1.0452 0.98803 5.5191e-05 3.8182 0.012036 1.376e-05 0.0011541 0.14453 0.00065817 0.14518 0.13219 0 0.037355 0.0389 0 0.89235 0.24778 0.066282 0.0092699 4.2267 0.057903 6.9498e-05 0.83217 0.005244 0.0059811 0.0013829 0.98699 0.99173 2.9814e-06 1.1926e-05 0.13161 0.96135 0.92267 0.0013953 0.99584 0.61924 0.0018799 0.43144 1.9383 1.9378 15.998 144.9975 0.00015493 -85.6665 0.94221
1.0462 0.98803 5.5191e-05 3.8182 0.012036 1.3773e-05 0.0011541 0.1446 0.00065817 0.14526 0.13225 0 0.037351 0.0389 0 0.89242 0.24781 0.066294 0.0092713 4.227 0.057912 6.9509e-05 0.83216 0.0052443 0.0059815 0.0013829 0.98699 0.99173 2.9814e-06 1.1926e-05 0.13161 0.96142 0.9227 0.0013953 0.99585 0.61937 0.0018799 0.43145 1.9386 1.9381 15.9979 144.9976 0.00015488 -85.6666 0.94321
1.0472 0.98803 5.5191e-05 3.8182 0.012036 1.3786e-05 0.0011541 0.14468 0.00065818 0.14533 0.13232 0 0.037346 0.0389 0 0.8925 0.24784 0.066306 0.0092728 4.2273 0.057921 6.9521e-05 0.83215 0.0052446 0.0059818 0.0013829 0.98699 0.99173 2.9814e-06 1.1926e-05 0.13162 0.96149 0.92273 0.0013953 0.99586 0.6195 0.0018799 0.43146 1.9389 1.9384 15.9979 144.9976 0.00015483 -85.6666 0.94421
1.0482 0.98803 5.5191e-05 3.8182 0.012036 1.3799e-05 0.0011541 0.14475 0.00065818 0.1454 0.13239 0 0.037341 0.0389 0 0.89257 0.24787 0.066317 0.0092742 4.2276 0.05793 6.9532e-05 0.83214 0.0052449 0.0059821 0.0013829 0.98699 0.99173 2.9814e-06 1.1925e-05 0.13162 0.96156 0.92277 0.0013953 0.99587 0.61964 0.0018799 0.43147 1.9392 1.9388 15.9979 144.9976 0.00015478 -85.6666 0.94521
1.0492 0.98803 5.5191e-05 3.8182 0.012036 1.3813e-05 0.0011541 0.14482 0.00065818 0.14548 0.13246 0 0.037336 0.0389 0 0.89265 0.24791 0.066329 0.0092757 4.2279 0.057939 6.9543e-05 0.83213 0.0052453 0.0059825 0.0013829 0.98699 0.99173 2.9814e-06 1.1925e-05 0.13162 0.96163 0.9228 0.0013953 0.99588 0.61977 0.0018799 0.43148 1.9395 1.9391 15.9978 144.9976 0.00015473 -85.6667 0.94621
1.0502 0.98803 5.5191e-05 3.8182 0.012036 1.3826e-05 0.0011541 0.1449 0.00065818 0.14555 0.13253 0 0.037331 0.0389 0 0.89272 0.24794 0.066341 0.0092771 4.2282 0.057948 6.9555e-05 0.83212 0.0052456 0.0059828 0.0013829 0.98699 0.99173 2.9814e-06 1.1925e-05 0.13162 0.96169 0.92283 0.0013953 0.99589 0.6199 0.0018799 0.43149 1.9398 1.9394 15.9978 144.9976 0.00015468 -85.6667 0.94721
1.0512 0.98803 5.5191e-05 3.8182 0.012036 1.3839e-05 0.0011541 0.14497 0.00065818 0.14562 0.13259 0 0.037327 0.0389 0 0.89279 0.24797 0.066353 0.0092786 4.2285 0.057956 6.9567e-05 0.83211 0.0052459 0.0059831 0.0013829 0.98699 0.99173 2.9814e-06 1.1925e-05 0.13163 0.96176 0.92286 0.0013953 0.99589 0.62003 0.0018799 0.4315 1.9401 1.9397 15.9978 144.9977 0.00015463 -85.6667 0.94821
1.0522 0.98803 5.5191e-05 3.8182 0.012036 1.3852e-05 0.0011541 0.14504 0.00065818 0.14569 0.13266 0 0.037322 0.0389 0 0.89287 0.24801 0.066365 0.0092801 4.2288 0.057965 6.9577e-05 0.8321 0.0052463 0.0059835 0.0013829 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13163 0.96183 0.92289 0.0013953 0.9959 0.62017 0.0018799 0.43152 1.9404 1.94 15.9977 144.9977 0.00015458 -85.6667 0.94921
1.0532 0.98803 5.5191e-05 3.8182 0.012036 1.3865e-05 0.0011541 0.14511 0.00065818 0.14577 0.13273 0 0.037317 0.0389 0 0.89294 0.24804 0.066377 0.0092815 4.2291 0.057974 6.9589e-05 0.8321 0.0052466 0.0059838 0.0013828 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13163 0.9619 0.92292 0.0013953 0.99591 0.6203 0.0018799 0.43153 1.9407 1.9403 15.9977 144.9977 0.00015454 -85.6668 0.95021
1.0542 0.98803 5.5191e-05 3.8182 0.012036 1.3878e-05 0.0011541 0.14519 0.00065819 0.14584 0.1328 0 0.037312 0.0389 0 0.89302 0.24807 0.066388 0.009283 4.2294 0.057983 6.9602e-05 0.83209 0.0052469 0.0059841 0.0013828 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13164 0.96197 0.92295 0.0013953 0.99592 0.62043 0.0018798 0.43154 1.941 1.9406 15.9977 144.9977 0.00015449 -85.6668 0.95121
1.0552 0.98803 5.5191e-05 3.8182 0.012036 1.3891e-05 0.0011541 0.14526 0.00065819 0.14591 0.13287 0 0.037308 0.0389 0 0.89309 0.2481 0.0664 0.0092844 4.2298 0.057992 6.9612e-05 0.83208 0.0052473 0.0059844 0.0013828 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13164 0.96203 0.92298 0.0013953 0.99593 0.62056 0.0018798 0.43155 1.9413 1.9409 15.9976 144.9977 0.00015444 -85.6668 0.95221
1.0562 0.98803 5.5191e-05 3.8182 0.012036 1.3904e-05 0.0011541 0.14533 0.00065819 0.14598 0.13293 0 0.037303 0.0389 0 0.89316 0.24814 0.066412 0.0092859 4.2301 0.058001 6.9621e-05 0.83207 0.0052476 0.0059848 0.0013828 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13164 0.9621 0.92301 0.0013953 0.99593 0.62069 0.0018798 0.43156 1.9416 1.9412 15.9976 144.9978 0.00015439 -85.6668 0.95321
1.0572 0.98803 5.5191e-05 3.8182 0.012036 1.3918e-05 0.0011541 0.1454 0.00065819 0.14606 0.133 0 0.037298 0.0389 0 0.89324 0.24817 0.066424 0.0092873 4.2304 0.05801 6.9638e-05 0.83206 0.0052479 0.0059851 0.0013828 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13164 0.96217 0.92304 0.0013953 0.99594 0.62083 0.0018798 0.43157 1.942 1.9415 15.9976 144.9978 0.00015434 -85.6669 0.95421
1.0582 0.98803 5.5191e-05 3.8182 0.012036 1.3931e-05 0.0011541 0.14548 0.00065819 0.14613 0.13307 0 0.037293 0.0389 0 0.89331 0.2482 0.066436 0.0092888 4.2307 0.058019 6.9646e-05 0.83205 0.0052483 0.0059855 0.0013828 0.98699 0.99173 2.9813e-06 1.1925e-05 0.13165 0.96223 0.92307 0.0013953 0.99595 0.62096 0.0018798 0.43159 1.9423 1.9418 15.9975 144.9978 0.00015429 -85.6669 0.95521
1.0592 0.98803 5.5191e-05 3.8182 0.012036 1.3944e-05 0.0011541 0.14555 0.00065819 0.1462 0.13314 0 0.037289 0.0389 0 0.89339 0.24824 0.066448 0.0092903 4.231 0.058028 6.9654e-05 0.83204 0.0052486 0.0059858 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13165 0.9623 0.9231 0.0013953 0.99596 0.62109 0.0018798 0.4316 1.9426 1.9421 15.9975 144.9978 0.00015425 -85.6669 0.95621
1.0602 0.98803 5.519e-05 3.8182 0.012036 1.3957e-05 0.0011541 0.14562 0.00065819 0.14627 0.1332 0 0.037284 0.0389 0 0.89346 0.24827 0.06646 0.0092917 4.2313 0.058037 6.9671e-05 0.83203 0.0052489 0.0059861 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13165 0.96237 0.92313 0.0013952 0.99597 0.62122 0.0018798 0.43161 1.9429 1.9424 15.9975 144.9978 0.0001542 -85.6669 0.95721
1.0612 0.98803 5.519e-05 3.8182 0.012036 1.397e-05 0.0011541 0.14569 0.0006582 0.14635 0.13327 0 0.037279 0.0389 0 0.89354 0.2483 0.066471 0.0092932 4.2316 0.058046 6.9682e-05 0.83202 0.0052493 0.0059865 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13166 0.96243 0.92317 0.0013952 0.99597 0.62135 0.0018798 0.43162 1.9432 1.9427 15.9974 144.9979 0.00015415 -85.667 0.95821
1.0622 0.98803 5.519e-05 3.8182 0.012036 1.3983e-05 0.0011541 0.14576 0.0006582 0.14642 0.13334 0 0.037275 0.0389 0 0.89361 0.24833 0.066483 0.0092946 4.2319 0.058055 6.9689e-05 0.83202 0.0052496 0.0059868 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13166 0.9625 0.9232 0.0013952 0.99598 0.62149 0.0018798 0.43163 1.9435 1.943 15.9974 144.9979 0.0001541 -85.667 0.95921
1.0632 0.98803 5.519e-05 3.8182 0.012036 1.3996e-05 0.0011541 0.14584 0.0006582 0.14649 0.13341 0 0.03727 0.0389 0 0.89368 0.24837 0.066495 0.0092961 4.2322 0.058063 6.9704e-05 0.83201 0.0052499 0.0059871 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13166 0.96257 0.92323 0.0013952 0.99599 0.62162 0.0018798 0.43164 1.9438 1.9433 15.9974 144.9979 0.00015406 -85.667 0.96021
1.0642 0.98803 5.519e-05 3.8182 0.012036 1.401e-05 0.0011541 0.14591 0.0006582 0.14656 0.13347 0 0.037265 0.0389 0 0.89376 0.2484 0.066507 0.0092976 4.2325 0.058072 6.9715e-05 0.832 0.0052503 0.0059875 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13166 0.96263 0.92325 0.0013952 0.996 0.62175 0.0018798 0.43165 1.9441 1.9436 15.9973 144.9979 0.00015401 -85.667 0.96121
1.0652 0.98803 5.519e-05 3.8182 0.012036 1.4023e-05 0.0011541 0.14598 0.0006582 0.14663 0.13354 0 0.037261 0.0389 0 0.89383 0.24843 0.066519 0.009299 4.2329 0.058081 6.9726e-05 0.83199 0.0052506 0.0059878 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13167 0.9627 0.92328 0.0013952 0.99601 0.62188 0.0018798 0.43167 1.9444 1.9439 15.9973 144.998 0.00015396 -85.6671 0.96221
1.0662 0.98803 5.519e-05 3.8182 0.012036 1.4036e-05 0.0011541 0.14605 0.0006582 0.14671 0.13361 0 0.037256 0.0389 0 0.89391 0.24847 0.066531 0.0093005 4.2332 0.05809 6.9738e-05 0.83198 0.0052509 0.0059881 0.0013828 0.98699 0.99173 2.9812e-06 1.1925e-05 0.13167 0.96276 0.92331 0.0013952 0.99601 0.62201 0.0018798 0.43168 1.9447 1.9442 15.9973 144.998 0.00015392 -85.6671 0.96321
1.0672 0.98803 5.519e-05 3.8182 0.012036 1.4049e-05 0.0011541 0.14612 0.0006582 0.14678 0.13367 0 0.037251 0.0389 0 0.89398 0.2485 0.066543 0.009302 4.2335 0.058099 6.975e-05 0.83197 0.0052513 0.0059885 0.0013828 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13167 0.96283 0.92334 0.0013952 0.99602 0.62214 0.0018798 0.43169 1.945 1.9445 15.9972 144.998 0.00015387 -85.6671 0.96421
1.0682 0.98803 5.519e-05 3.8182 0.012036 1.4062e-05 0.0011541 0.1462 0.00065821 0.14685 0.13374 0 0.037246 0.0389 0 0.89406 0.24853 0.066555 0.0093034 4.2338 0.058108 6.9761e-05 0.83196 0.0052516 0.0059888 0.0013828 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13167 0.96289 0.92337 0.0013952 0.99603 0.62227 0.0018798 0.4317 1.9453 1.9448 15.9972 144.998 0.00015382 -85.6671 0.96521
1.0692 0.98803 5.519e-05 3.8182 0.012036 1.4075e-05 0.0011541 0.14627 0.00065821 0.14692 0.13381 0 0.037242 0.0389 0 0.89413 0.24857 0.066567 0.0093049 4.2341 0.058117 6.9773e-05 0.83195 0.0052519 0.0059892 0.0013828 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13168 0.96296 0.9234 0.0013952 0.99604 0.62241 0.0018798 0.43171 1.9455 1.9451 15.9972 144.998 0.00015378 -85.6671 0.96621
1.0702 0.98803 5.519e-05 3.8182 0.012036 1.4088e-05 0.0011541 0.14634 0.00065821 0.14699 0.13388 0 0.037237 0.0389 0 0.89421 0.2486 0.066579 0.0093064 4.2344 0.058126 6.9784e-05 0.83194 0.0052523 0.0059895 0.0013828 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13168 0.96302 0.92343 0.0013952 0.99604 0.62254 0.0018798 0.43172 1.9458 1.9454 15.9971 144.9981 0.00015373 -85.6672 0.96721
1.0712 0.98803 5.519e-05 3.8182 0.012036 1.4102e-05 0.0011541 0.14641 0.00065821 0.14706 0.13394 0 0.037232 0.0389 0 0.89428 0.24863 0.066591 0.0093078 4.2347 0.058135 6.9796e-05 0.83193 0.0052526 0.0059898 0.0013827 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13168 0.96308 0.92346 0.0013952 0.99605 0.62267 0.0018798 0.43173 1.9461 1.9457 15.9971 144.9981 0.00015369 -85.6672 0.96821
1.0722 0.98803 5.519e-05 3.8182 0.012036 1.4115e-05 0.0011541 0.14648 0.00065821 0.14713 0.13401 0 0.037228 0.0389 0 0.89435 0.24867 0.066603 0.0093093 4.2351 0.058144 6.9807e-05 0.83193 0.0052529 0.0059902 0.0013827 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13169 0.96315 0.92349 0.0013952 0.99606 0.6228 0.0018798 0.43174 1.9464 1.946 15.9971 144.9981 0.00015364 -85.6672 0.96921
1.0732 0.98803 5.519e-05 3.8182 0.012036 1.4128e-05 0.0011541 0.14655 0.00065821 0.14721 0.13408 0 0.037223 0.0389 0 0.89443 0.2487 0.066615 0.0093108 4.2354 0.058153 6.9819e-05 0.83192 0.0052533 0.0059905 0.0013827 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13169 0.96321 0.92352 0.0013952 0.99606 0.62293 0.0018798 0.43176 1.9467 1.9463 15.997 144.9981 0.00015359 -85.6672 0.97021
1.0742 0.98803 5.519e-05 3.8182 0.012036 1.4141e-05 0.0011541 0.14662 0.00065821 0.14728 0.13414 0 0.037219 0.0389 0 0.8945 0.24873 0.066627 0.0093122 4.2357 0.058162 6.983e-05 0.83191 0.0052536 0.0059909 0.0013827 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13169 0.96328 0.92355 0.0013952 0.99607 0.62306 0.0018798 0.43177 1.947 1.9466 15.997 144.9981 0.00015355 -85.6673 0.97121
1.0752 0.98803 5.519e-05 3.8182 0.012036 1.4154e-05 0.0011541 0.1467 0.00065822 0.14735 0.13421 0 0.037214 0.0389 0 0.89458 0.24876 0.066639 0.0093137 4.236 0.058171 6.9842e-05 0.8319 0.005254 0.0059912 0.0013827 0.98699 0.99173 2.9811e-06 1.1924e-05 0.13169 0.96334 0.92358 0.0013952 0.99608 0.62319 0.0018798 0.43178 1.9473 1.9469 15.997 144.9982 0.0001535 -85.6673 0.97221
1.0762 0.98803 5.5189e-05 3.8182 0.012036 1.4167e-05 0.0011541 0.14677 0.00065822 0.14742 0.13428 0 0.037209 0.0389 0 0.89465 0.2488 0.06665 0.0093152 4.2363 0.05818 6.9853e-05 0.83189 0.0052543 0.0059915 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.1317 0.9634 0.92361 0.0013952 0.99609 0.62332 0.0018798 0.43179 1.9476 1.9472 15.9969 144.9982 0.00015346 -85.6673 0.97321
1.0772 0.98803 5.5189e-05 3.8182 0.012036 1.418e-05 0.0011541 0.14684 0.00065822 0.14749 0.13434 0 0.037205 0.0389 0 0.89473 0.24883 0.066662 0.0093166 4.2366 0.058189 6.9865e-05 0.83188 0.0052546 0.0059919 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.1317 0.96346 0.92363 0.0013952 0.99609 0.62346 0.0018798 0.4318 1.9479 1.9475 15.9969 144.9982 0.00015341 -85.6673 0.97421
1.0782 0.98803 5.5189e-05 3.8182 0.012036 1.4194e-05 0.0011541 0.14691 0.00065822 0.14756 0.13441 0 0.0372 0.0389 0 0.8948 0.24886 0.066674 0.0093181 4.237 0.058198 6.9876e-05 0.83187 0.005255 0.0059922 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.1317 0.96353 0.92366 0.0013952 0.9961 0.62359 0.0018798 0.43181 1.9482 1.9478 15.9969 144.9982 0.00015337 -85.6673 0.97521
1.0792 0.98803 5.5189e-05 3.8182 0.012036 1.4207e-05 0.0011541 0.14698 0.00065822 0.14763 0.13448 0 0.037195 0.0389 0 0.89488 0.2489 0.066686 0.0093196 4.2373 0.058207 6.9888e-05 0.83186 0.0052553 0.0059926 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13171 0.96359 0.92369 0.0013952 0.99611 0.62372 0.0018798 0.43182 1.9485 1.9481 15.9968 144.9982 0.00015332 -85.6674 0.97621
1.0802 0.98803 5.5189e-05 3.8182 0.012036 1.422e-05 0.0011541 0.14705 0.00065822 0.1477 0.13454 0 0.037191 0.0389 0 0.89495 0.24893 0.066698 0.0093211 4.2376 0.058216 6.9899e-05 0.83185 0.0052557 0.0059929 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13171 0.96365 0.92372 0.0013952 0.99611 0.62385 0.0018798 0.43184 1.9488 1.9484 15.9968 144.9983 0.00015328 -85.6674 0.97721
1.0812 0.98803 5.5189e-05 3.8182 0.012036 1.4233e-05 0.0011541 0.14712 0.00065822 0.14778 0.13461 0 0.037186 0.0389 0 0.89503 0.24896 0.06671 0.0093225 4.2379 0.058225 6.9911e-05 0.83184 0.005256 0.0059932 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13171 0.96371 0.92375 0.0013952 0.99612 0.62398 0.0018797 0.43185 1.9491 1.9486 15.9967 144.9983 0.00015323 -85.6674 0.97821
1.0822 0.98803 5.5189e-05 3.8182 0.012036 1.4246e-05 0.0011541 0.14719 0.00065823 0.14785 0.13467 0 0.037182 0.0389 0 0.8951 0.249 0.066722 0.009324 4.2382 0.058234 6.9923e-05 0.83184 0.0052563 0.0059936 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13171 0.96378 0.92378 0.0013952 0.99613 0.62411 0.0018797 0.43186 1.9494 1.9489 15.9967 144.9983 0.00015319 -85.6674 0.97921
1.0832 0.98803 5.5189e-05 3.8182 0.012036 1.4259e-05 0.0011541 0.14726 0.00065823 0.14792 0.13474 0 0.037177 0.0389 0 0.89518 0.24903 0.066734 0.0093255 4.2386 0.058243 6.9934e-05 0.83183 0.0052567 0.0059939 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13172 0.96384 0.9238 0.0013952 0.99613 0.62424 0.0018797 0.43187 1.9497 1.9492 15.9967 144.9983 0.00015315 -85.6674 0.98021
1.0842 0.98803 5.5189e-05 3.8182 0.012036 1.4272e-05 0.0011541 0.14733 0.00065823 0.14799 0.13481 0 0.037172 0.0389 0 0.89525 0.24906 0.066746 0.0093269 4.2389 0.058252 6.9946e-05 0.83182 0.005257 0.0059943 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13172 0.9639 0.92383 0.0013952 0.99614 0.62437 0.0018797 0.43188 1.95 1.9495 15.9966 144.9983 0.0001531 -85.6675 0.98121
1.0852 0.98803 5.5189e-05 3.8182 0.012036 1.4286e-05 0.0011541 0.14741 0.00065823 0.14806 0.13487 0 0.037168 0.0389 0 0.89533 0.2491 0.066758 0.0093284 4.2392 0.058261 6.9958e-05 0.83181 0.0052574 0.0059946 0.0013827 0.98699 0.99173 2.981e-06 1.1924e-05 0.13172 0.96396 0.92386 0.0013952 0.99615 0.6245 0.0018797 0.43189 1.9502 1.9498 15.9966 144.9984 0.00015306 -85.6675 0.98221
1.0862 0.98803 5.5189e-05 3.8182 0.012036 1.4299e-05 0.0011541 0.14748 0.00065823 0.14813 0.13494 0 0.037163 0.0389 0 0.8954 0.24913 0.066771 0.0093299 4.2395 0.05827 6.9969e-05 0.8318 0.0052577 0.005995 0.0013827 0.98699 0.99173 2.9809e-06 1.1924e-05 0.13173 0.96402 0.92389 0.0013952 0.99615 0.62463 0.0018797 0.4319 1.9505 1.9501 15.9966 144.9984 0.00015301 -85.6675 0.98321
1.0872 0.98803 5.5189e-05 3.8182 0.012036 1.4312e-05 0.0011541 0.14755 0.00065823 0.1482 0.13501 0 0.037159 0.0389 0 0.89548 0.24916 0.066783 0.0093314 4.2398 0.058279 6.998e-05 0.83179 0.0052581 0.0059953 0.0013827 0.98699 0.99173 2.9809e-06 1.1924e-05 0.13173 0.96408 0.92392 0.0013952 0.99616 0.62476 0.0018797 0.43191 1.9508 1.9504 15.9965 144.9984 0.00015297 -85.6675 0.98421
1.0882 0.98803 5.5189e-05 3.8182 0.012036 1.4325e-05 0.0011541 0.14762 0.00065823 0.14827 0.13507 0 0.037154 0.0389 0 0.89555 0.2492 0.066795 0.0093329 4.2402 0.058288 6.9992e-05 0.83178 0.0052584 0.0059957 0.0013827 0.98699 0.99173 2.9809e-06 1.1924e-05 0.13173 0.96414 0.92394 0.0013952 0.99617 0.62489 0.0018797 0.43193 1.9511 1.9507 15.9965 144.9984 0.00015293 -85.6675 0.98521
1.0892 0.98803 5.5189e-05 3.8182 0.012036 1.4338e-05 0.0011542 0.14769 0.00065824 0.14834 0.13514 0 0.037149 0.0389 0 0.89563 0.24923 0.066807 0.0093343 4.2405 0.058297 7.0005e-05 0.83177 0.0052587 0.005996 0.0013827 0.98699 0.99173 2.9809e-06 1.1924e-05 0.13173 0.9642 0.92397 0.0013952 0.99617 0.62503 0.0018797 0.43194 1.9514 1.951 15.9965 144.9984 0.00015288 -85.6676 0.98621
1.0902 0.98803 5.5189e-05 3.8182 0.012035 1.4351e-05 0.0011542 0.14776 0.00065824 0.14841 0.1352 0 0.037145 0.0389 0 0.8957 0.24926 0.066819 0.0093358 4.2408 0.058306 7.0015e-05 0.83176 0.0052591 0.0059964 0.0013827 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13174 0.96427 0.924 0.0013952 0.99618 0.62516 0.0018797 0.43195 1.9517 1.9513 15.9964 144.9985 0.00015284 -85.6676 0.98721
1.0912 0.98803 5.5189e-05 3.8182 0.012035 1.4364e-05 0.0011542 0.14783 0.00065824 0.14848 0.13527 0 0.03714 0.0389 0 0.89578 0.2493 0.066831 0.0093373 4.2411 0.058315 7.0026e-05 0.83175 0.0052594 0.0059967 0.0013827 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13174 0.96433 0.92403 0.0013952 0.99619 0.62529 0.0018797 0.43196 1.952 1.9516 15.9964 144.9985 0.0001528 -85.6676 0.98821
1.0922 0.98803 5.5188e-05 3.8182 0.012035 1.4378e-05 0.0011542 0.1479 0.00065824 0.14855 0.13533 0 0.037136 0.0389 0 0.89585 0.24933 0.066843 0.0093388 4.2415 0.058324 7.004e-05 0.83175 0.0052598 0.0059971 0.0013827 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13174 0.96439 0.92405 0.0013952 0.99619 0.62542 0.0018797 0.43197 1.9523 1.9518 15.9964 144.9985 0.00015275 -85.6676 0.98921
1.0932 0.98803 5.5188e-05 3.8182 0.012035 1.4391e-05 0.0011542 0.14797 0.00065824 0.14862 0.1354 0 0.037131 0.0389 0 0.89593 0.24936 0.066855 0.0093402 4.2418 0.058334 7.0052e-05 0.83174 0.0052601 0.0059974 0.0013826 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13175 0.96445 0.92408 0.0013952 0.9962 0.62555 0.0018797 0.43198 1.9526 1.9521 15.9963 144.9985 0.00015271 -85.6676 0.99021
1.0942 0.98803 5.5188e-05 3.8182 0.012035 1.4404e-05 0.0011542 0.14804 0.00065824 0.14869 0.13547 0 0.037127 0.0389 0 0.89601 0.2494 0.066867 0.0093417 4.2421 0.058343 7.0062e-05 0.83173 0.0052605 0.0059977 0.0013826 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13175 0.9645 0.92411 0.0013952 0.99621 0.62568 0.0018797 0.43199 1.9528 1.9524 15.9963 144.9985 0.00015267 -85.6676 0.99121
1.0952 0.98803 5.5188e-05 3.8182 0.012035 1.4417e-05 0.0011542 0.14811 0.00065824 0.14876 0.13553 0 0.037122 0.0389 0 0.89608 0.24943 0.066879 0.0093432 4.2424 0.058352 7.0077e-05 0.83172 0.0052608 0.0059981 0.0013826 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13175 0.96456 0.92413 0.0013952 0.99621 0.62581 0.0018797 0.43201 1.9531 1.9527 15.9963 144.9986 0.00015263 -85.6677 0.99221
1.0962 0.98803 5.5188e-05 3.8182 0.012035 1.443e-05 0.0011542 0.14818 0.00065825 0.14883 0.1356 0 0.037117 0.0389 0 0.89616 0.24946 0.066891 0.0093447 4.2428 0.058361 7.0088e-05 0.83171 0.0052612 0.0059984 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13175 0.96462 0.92416 0.0013952 0.99622 0.62594 0.0018797 0.43202 1.9534 1.953 15.9962 144.9986 0.00015258 -85.6677 0.99321
1.0972 0.98803 5.5188e-05 3.8182 0.012035 1.4443e-05 0.0011542 0.14825 0.00065825 0.1489 0.13566 0 0.037113 0.0389 0 0.89623 0.2495 0.066903 0.0093462 4.2431 0.05837 7.0097e-05 0.8317 0.0052615 0.0059988 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96468 0.92419 0.0013952 0.99623 0.62607 0.0018797 0.43203 1.9537 1.9533 15.9962 144.9986 0.00015254 -85.6677 0.99421
1.0982 0.98803 5.5188e-05 3.8182 0.012035 1.4456e-05 0.0011542 0.14832 0.00065825 0.14897 0.13573 0 0.037108 0.0389 0 0.89631 0.24953 0.066915 0.0093477 4.2434 0.058379 7.0109e-05 0.83169 0.0052619 0.0059991 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96474 0.92421 0.0013952 0.99623 0.6262 0.0018797 0.43204 1.954 1.9536 15.9962 144.9986 0.0001525 -85.6677 0.99521
1.0992 0.98803 5.5188e-05 3.8182 0.012035 1.447e-05 0.0011542 0.14839 0.00065825 0.14904 0.13579 0 0.037104 0.0389 0 0.89638 0.24957 0.066927 0.0093491 4.2437 0.058388 7.0121e-05 0.83168 0.0052622 0.0059995 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.9648 0.92424 0.0013952 0.99624 0.62633 0.0018797 0.43205 1.9543 1.9538 15.9961 144.9986 0.00015246 -85.6677 0.99621
1.0995 0.98803 5.5188e-05 3.8182 0.012035 1.4473e-05 0.0011542 0.14841 0.00065825 0.14906 0.13581 0 0.037103 0.0389 0 0.8964 0.24957 0.06693 0.0093495 4.2438 0.05839 7.0123e-05 0.83168 0.0052623 0.0059996 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96482 0.92425 0.0013952 0.99624 0.62636 0.0018797 0.43205 1.9543 1.9539 15.9961 144.9987 0.00015245 -85.6677 0.99646
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.4479e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066936 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96484 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99696
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.4479e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066936 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96484 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99697
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.4479e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96484 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99697
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013951 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6677 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.667 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6663 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013826 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.665 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013827 0.98699 0.99173 2.9808e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6623 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013829 0.98699 0.99173 2.9809e-06 1.1923e-05 0.13176 0.96485 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.657 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013837 0.98699 0.99173 2.9813e-06 1.1924e-05 0.13176 0.96485 0.92426 0.0013952 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6464 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013863 0.98699 0.99173 2.9827e-06 1.1927e-05 0.13177 0.96485 0.92426 0.0013953 0.99624 0.62643 0.0018797 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.6251 0.99698
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-05 0.83168 0.0052625 0.0059998 0.0013935 0.98699 0.99173 2.9877e-06 1.1938e-05 0.13177 0.96485 0.92426 0.0013958 0.99624 0.62643 0.0018798 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.5826 0.99699
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.013e-05 0.83168 0.0052625 0.0059998 0.001402 0.98699 0.99173 2.9948e-06 1.1954e-05 0.13177 0.96485 0.92426 0.0013965 0.99624 0.62643 0.0018799 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.5401 0.99699
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.013e-05 0.83167 0.0052625 0.0059998 0.0014208 0.98699 0.99173 3.0156e-06 1.2003e-05 0.13177 0.96485 0.92426 0.0013987 0.99624 0.62643 0.0018802 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.4552 0.997
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14845 0.00065825 0.1491 0.13585 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.013e-05 0.83167 0.0052625 0.0059998 0.0014406 0.98699 0.99173 3.0416e-06 1.2068e-05 0.13177 0.96485 0.92426 0.0014016 0.99624 0.62643 0.0018807 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015243 -85.3705 0.99701
1.1 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14845 0.00065825 0.1491 0.13585 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.013e-05 0.83167 0.0052625 0.0059998 0.0014815 0.98698 0.99173 3.1079e-06 1.2247e-05 0.13177 0.96485 0.92426 0.0014098 0.99624 0.62643 0.001882 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -85.2013 0.99703
1.1001 0.98803 5.5188e-05 3.8182 0.012035 1.448e-05 0.0011542 0.14845 0.00065825 0.1491 0.13585 0 0.0371 0.0389 0 0.89645 0.24959 0.066937 0.0093504 4.244 0.058396 7.013e-05 0.83167 0.0052625 0.0059998 0.0015193 0.98697 0.99173 3.176e-06 1.2443e-05 0.13177 0.96485 0.92426 0.0014188 0.99624 0.62644 0.0018837 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -85.0493 0.99704
1.1001 0.98803 5.5188e-05 3.8182 0.012035 1.4481e-05 0.0011542 0.14845 0.00065825 0.1491 0.13585 0 0.0371 0.0389 0 0.89645 0.24959 0.066938 0.0093504 4.244 0.058396 7.013e-05 0.83167 0.0052625 0.0059998 0.001558 0.98696 0.99173 3.2506e-06 1.2668e-05 0.13177 0.96485 0.92426 0.0014293 0.99624 0.62644 0.0018857 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -84.8976 0.99706
1.1001 0.98803 5.5188e-05 3.8182 0.012035 1.4481e-05 0.0011542 0.14845 0.00065825 0.1491 0.13585 0 0.0371 0.0389 0 0.89645 0.24959 0.066938 0.0093504 4.244 0.058396 7.013e-05 0.83167 0.0052625 0.0059998 0.0015975 0.98695 0.99173 3.3301e-06 1.2918e-05 0.13177 0.96485 0.92426 0.0014409 0.99624 0.62644 0.001888 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -84.7462 0.99707
1.1001 0.98803 5.5188e-05 3.8182 0.012035 1.4481e-05 0.0011542 0.14845 0.00065825 0.14911 0.13585 0 0.0371 0.0389 0 0.89645 0.24959 0.066938 0.0093505 4.244 0.058396 7.0131e-05 0.83167 0.0052625 0.0059998 0.0016794 0.98692 0.99172 3.4989e-06 1.3465e-05 0.13177 0.96485 0.92426 0.0014664 0.99624 0.62644 0.0018935 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -84.4441 0.9971
1.1002 0.98803 5.5188e-05 3.8182 0.012035 1.4482e-05 0.0011542 0.14845 0.00065825 0.14911 0.13585 0 0.0371 0.0389 0 0.89645 0.2496 0.066938 0.0093505 4.244 0.058396 7.0131e-05 0.83167 0.0052625 0.0059998 0.0017652 0.98688 0.99172 3.6813e-06 1.4081e-05 0.13177 0.96485 0.92427 0.0014951 0.99624 0.62645 0.0019002 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -84.143 0.99713
1.1002 0.98803 5.5188e-05 3.8182 0.012035 1.4482e-05 0.0011542 0.14846 0.00065825 0.14911 0.13586 0 0.0371 0.0389 0 0.89645 0.2496 0.066939 0.0093505 4.2441 0.058397 7.0132e-05 0.83167 0.0052625 0.0059998 0.001855 0.98684 0.99171 3.8757e-06 1.476e-05 0.13177 0.96485 0.92427 0.0015265 0.99624 0.62645 0.001908 0.43206 1.9545 1.9541 15.9961 144.9987 0.00015242 -83.8429 0.99716
1.1002 0.98803 5.5188e-05 3.8182 0.012035 1.4483e-05 0.0011542 0.14846 0.00065825 0.14911 0.13586 0 0.037099 0.0389 0 0.89646 0.2496 0.06694 0.0093506 4.2441 0.058397 7.0132e-05 0.83167 0.0052626 0.0059999 0.0020471 0.98673 0.9917 4.2963e-06 1.6267e-05 0.13177 0.96486 0.92427 0.0015948 0.99624 0.62646 0.001927 0.43206 1.9546 1.9541 15.9961 144.9987 0.00015242 -83.2459 0.99723
1.1003 0.98803 5.5188e-05 3.8182 0.012035 1.4484e-05 0.0011542 0.14846 0.00065825 0.14912 0.13586 0 0.037099 0.0389 0 0.89646 0.2496 0.06694 0.0093507 4.2441 0.058398 7.0133e-05 0.83167 0.0052626 0.0059999 0.0022571 0.98659 0.99167 4.7607e-06 1.7964e-05 0.13177 0.96486 0.92427 0.0016692 0.99624 0.62647 0.00195 0.43206 1.9546 1.9542 15.9961 144.9987 0.00015241 -82.6529 0.99729
1.1004 0.98803 5.5188e-05 3.8182 0.012035 1.4484e-05 0.0011542 0.14847 0.00065825 0.14912 0.13587 0 0.037099 0.0389 0 0.89647 0.2496 0.066941 0.0093508 4.2441 0.058398 7.0134e-05 0.83167 0.0052626 0.0059999 0.0024865 0.98643 0.99165 5.2712e-06 1.9841e-05 0.13177 0.96486 0.92427 0.0017484 0.99624 0.62647 0.0019767 0.43206 1.9546 1.9542 15.9961 144.9987 0.00015241 -82.0637 0.99735
1.1004 0.98803 5.5188e-05 3.8182 0.012035 1.4485e-05 0.0011542 0.14847 0.00065825 0.14913 0.13587 0 0.037098 0.0389 0 0.89647 0.24961 0.066942 0.0093509 4.2441 0.058399 7.0134e-05 0.83167 0.0052626 0.0059999 0.002737 0.98624 0.99162 5.8319e-06 2.1906e-05 0.13177 0.96486 0.92427 0.0018314 0.99624 0.62648 0.0020065 0.43205 1.9546 1.9542 15.9961 144.9987 0.00015241 -81.478 0.99741
1.1006 0.98803 5.5188e-05 3.8182 0.012035 1.4487e-05 0.0011542 0.14848 0.00065825 0.14914 0.13588 0 0.037098 0.0389 0 0.89648 0.24961 0.066943 0.0093511 4.2442 0.0584 7.0136e-05 0.83167 0.0052627 0.006 0.0033093 0.98578 0.99153 7.1241e-06 2.6648e-05 0.13177 0.96486 0.92428 0.0020083 0.99624 0.62649 0.0020749 0.43205 1.9546 1.9542 15.9961 144.9987 0.00015241 -80.3164 0.99753
1.1007 0.98803 5.5188e-05 3.8182 0.012035 1.4488e-05 0.0011542 0.14849 0.00065825 0.14914 0.13589 0 0.037097 0.0389 0 0.89649 0.24961 0.066945 0.0093513 4.2442 0.058401 7.0137e-05 0.83167 0.0052627 0.006 0.0039896 0.98522 0.99143 8.6803e-06 3.232e-05 0.13177 0.96486 0.92428 0.0021985 0.99624 0.62651 0.0021528 0.43204 1.9547 1.9543 15.9961 144.9987 0.0001524 -79.1667 0.99765
1.1008 0.98803 5.5188e-05 3.8182 0.012035 1.449e-05 0.0011542 0.1485 0.00065825 0.14915 0.1359 0 0.037097 0.0389 0 0.8965 0.24962 0.066946 0.0093515 4.2443 0.058402 7.0139e-05 0.83167 0.0052628 0.006 0.0047963 0.98456 0.99129 1.0552e-05 3.9094e-05 0.13177 0.96486 0.92428 0.0024023 0.99624 0.62652 0.0022387 0.43203 1.9547 1.9543 15.9961 144.9987 0.0001524 -78.0273 0.99778
1.1009 0.98803 5.5188e-05 3.8182 0.012035 1.4492e-05 0.0011542 0.14851 0.00065825 0.14916 0.1359 0 0.037096 0.0389 0 0.89651 0.24962 0.066948 0.0093516 4.2443 0.058403 7.014e-05 0.83167 0.0052628 0.0060001 0.005752 0.9838 0.99113 1.2801e-05 4.7182e-05 0.13177 0.96486 0.92429 0.0026207 0.99624 0.62653 0.0023311 0.43202 1.9547 1.9543 15.9961 144.9987 0.0001524 -76.8967 0.9979
1.101 0.98803 5.5188e-05 3.8182 0.012035 1.4493e-05 0.0011542 0.14852 0.00065825 0.14917 0.13591 0 0.037096 0.0389 0 0.89652 0.24963 0.066949 0.0093518 4.2443 0.058404 7.0142e-05 0.83167 0.0052628 0.0060001 0.0068837 0.98293 0.99093 1.5501e-05 5.6833e-05 0.13177 0.96485 0.92429 0.0028551 0.99623 0.62654 0.0024294 0.43201 1.9548 1.9544 15.9961 144.9987 0.00015239 -75.7737 0.99802
1.1012 0.98803 5.5188e-05 3.8182 0.012035 1.4495e-05 0.0011542 0.14852 0.00065825 0.14918 0.13592 0 0.037095 0.0389 0 0.89653 0.24963 0.066951 0.009352 4.2444 0.058406 7.0143e-05 0.83166 0.0052629 0.0060002 0.008223 0.98194 0.99069 1.8744e-05 6.8337e-05 0.13177 0.96484 0.92429 0.0031061 0.99623 0.62656 0.0025328 0.432 1.9548 1.9544 15.9961 144.9987 0.00015239 -74.6571 0.99815
1.1013 0.98803 5.5188e-05 3.8182 0.012035 1.4497e-05 0.0011542 0.14853 0.00065825 0.14919 0.13593 0 0.037095 0.0389 0 0.89654 0.24963 0.066952 0.0093522 4.2444 0.058407 7.0144e-05 0.83166 0.0052629 0.0060002 0.0098038 0.98084 0.99042 2.2633e-05 8.2019e-05 0.13177 0.96482 0.9243 0.0033739 0.99623 0.62657 0.0026409 0.43199 1.9549 1.9544 15.996 144.9986 0.00015239 -73.546 0.99827
1.1014 0.98803 5.5188e-05 3.8182 0.012035 1.4498e-05 0.0011542 0.14854 0.00065825 0.1492 0.13594 0 0.037094 0.0389 0 0.89655 0.24964 0.066954 0.0093524 4.2445 0.058408 7.0146e-05 0.83166 0.005263 0.0060003 0.011661 0.97962 0.99009 2.7284e-05 9.8255e-05 0.13177 0.96481 0.9243 0.0036589 0.99622 0.62658 0.002753 0.43198 1.9549 1.9545 15.996 144.9986 0.00015239 -72.4393 0.99839
1.1015 0.98803 5.5188e-05 3.8182 0.012035 1.45e-05 0.0011542 0.14855 0.00065825 0.1492 0.13594 0 0.037093 0.0389 0 0.89656 0.24964 0.066955 0.0093526 4.2445 0.058409 7.0147e-05 0.83166 0.005263 0.0060003 0.013842 0.97827 0.98972 3.2845e-05 0.00011751 0.13177 0.96478 0.9243 0.0039623 0.99622 0.62659 0.0028687 0.43196 1.9549 1.9545 15.996 144.9986 0.00015239 -71.3361 0.99851
1.1017 0.98803 5.5188e-05 3.8182 0.012035 1.4501e-05 0.0011542 0.14856 0.00065825 0.14921 0.13595 0 0.037093 0.0389 0 0.89657 0.24965 0.066957 0.0093527 4.2445 0.05841 7.0149e-05 0.83166 0.0052631 0.0060003 0.016405 0.97677 0.98928 3.9492e-05 0.00014033 0.13177 0.96475 0.9243 0.0042852 0.99621 0.6266 0.0029874 0.43195 1.955 1.9545 15.996 144.9986 0.00015239 -70.2355 0.99864
1.1018 0.98803 5.5188e-05 3.8182 0.012035 1.4503e-05 0.0011542 0.14857 0.00065825 0.14922 0.13596 0 0.037092 0.0389 0 0.89657 0.24965 0.066958 0.0093529 4.2446 0.058411 7.015e-05 0.83166 0.0052631 0.0060004 0.019415 0.97513 0.98878 4.7437e-05 0.00016734 0.13177 0.96472 0.92431 0.0046279 0.9962 0.62662 0.0031089 0.43193 1.955 1.9546 15.996 144.9986 0.00015238 -69.1368 0.99876
1.1019 0.98803 5.5188e-05 3.8182 0.012035 1.4505e-05 0.0011542 0.14858 0.00065825 0.14923 0.13597 0 0.037092 0.0389 0 0.89658 0.24965 0.06696 0.0093531 4.2446 0.058412 7.0152e-05 0.83166 0.0052631 0.0060004 0.022932 0.97332 0.98821 5.692e-05 0.00019928 0.13177 0.96468 0.92431 0.0049906 0.99619 0.62663 0.003233 0.43191 1.955 1.9546 15.996 144.9986 0.00015238 -68.0392 0.99888
1.102 0.98803 5.5188e-05 3.8182 0.012035 1.4506e-05 0.0011542 0.14858 0.00065825 0.14924 0.13598 0 0.037091 0.0389 0 0.89659 0.24966 0.066961 0.0093533 4.2447 0.058413 7.0153e-05 0.83166 0.0052632 0.0060005 0.027037 0.97134 0.98754 6.8241e-05 0.00023702 0.13177 0.96463 0.92431 0.0053741 0.99618 0.62664 0.0033594 0.43189 1.9551 1.9546 15.996 144.9986 0.00015238 -66.9421 0.999
1.1021 0.98803 5.5188e-05 3.8182 0.012035 1.4508e-05 0.0011542 0.14859 0.00065825 0.14925 0.13598 0 0.037091 0.0389 0 0.8966 0.24966 0.066962 0.0093534 4.2447 0.058414 7.0154e-05 0.83166 0.0052632 0.0060005 0.031309 0.96939 0.98686 8.0283e-05 0.00027676 0.13177 0.96458 0.92432 0.0057375 0.99617 0.62665 0.0034749 0.43188 1.9551 1.9547 15.996 144.9986 0.00015238 -65.9542 0.99911
1.1022 0.98803 5.5188e-05 3.8182 0.012035 1.4509e-05 0.0011542 0.1486 0.00065825 0.14925 0.13599 0 0.03709 0.0389 0 0.89661 0.24967 0.066964 0.0093536 4.2447 0.058415 7.0156e-05 0.83165 0.0052633 0.0060006 0.036206 0.96728 0.98609 9.4385e-05 0.00032286 0.13177 0.96452 0.92432 0.0061188 0.99615 0.62666 0.0035919 0.43186 1.9551 1.9547 15.996 144.9986 0.00015238 -64.9652 0.99922
1.1024 0.98803 5.5188e-05 3.8182 0.012035 1.4511e-05 0.0011542 0.14861 0.00065825 0.14926 0.136 0 0.03709 0.0389 0 0.89662 0.24967 0.066965 0.0093538 4.2448 0.058416 7.0157e-05 0.83165 0.0052633 0.0060006 0.041808 0.965 0.98522 0.0001109 0.00037631 0.13177 0.96446 0.92432 0.0065182 0.99614 0.62667 0.0037102 0.43184 1.9552 1.9547 15.996 144.9986 0.00015238 -63.974 0.99933
1.1025 0.98803 5.5188e-05 3.8182 0.012035 1.4512e-05 0.0011542 0.14862 0.00065825 0.14927 0.136 0 0.037089 0.0389 0 0.89663 0.24967 0.066966 0.0093539 4.2448 0.058417 7.0158e-05 0.83165 0.0052633 0.0060006 0.048211 0.96253 0.98424 0.00013024 0.00043826 0.13177 0.96438 0.92433 0.0069362 0.99612 0.62668 0.0038297 0.43182 1.9552 1.9548 15.9959 144.9986 0.00015239 -62.9795 0.99944
1.1026 0.98803 5.5188e-05 3.8182 0.012035 1.4513e-05 0.0011542 0.14862 0.00065825 0.14928 0.13601 0 0.037089 0.0389 0 0.89664 0.24968 0.066968 0.0093541 4.2448 0.058418 7.0159e-05 0.83165 0.0052634 0.0060007 0.055521 0.95985 0.98313 0.0001529 0.00051006 0.13177 0.9643 0.92433 0.0073732 0.99609 0.62669 0.0039504 0.43181 1.9552 1.9548 15.9959 144.9986 0.00015239 -61.98 0.99955
1.1027 0.98803 5.5188e-05 3.8182 0.012035 1.4515e-05 0.0011542 0.14863 0.00065825 0.14928 0.13602 0 0.037088 0.0389 0 0.89664 0.24968 0.066969 0.0093543 4.2449 0.058419 7.0161e-05 0.83165 0.0052634 0.0060007 0.063867 0.95694 0.98187 0.00017948 0.00059328 0.13177 0.96421 0.92433 0.0078296 0.99606 0.62669 0.004072 0.43179 1.9552 1.9548 15.9959 144.9986 0.00015239 -60.973 0.99966
1.1028 0.98803 5.5188e-05 3.8182 0.012035 1.4516e-05 0.0011542 0.14864 0.00065825 0.14929 0.13603 0 0.037088 0.0389 0 0.89665 0.24968 0.06697 0.0093544 4.2449 0.05842 7.0162e-05 0.83165 0.0052635 0.0060007 0.073394 0.9538 0.98046 0.00021072 0.00068986 0.13177 0.9641 0.92433 0.0083062 0.99602 0.6267 0.0041946 0.43177 1.9553 1.9549 15.9959 144.9986 0.00015239 -59.955 0.99978
1.1029 0.98803 5.5188e-05 3.8182 0.012035 1.4518e-05 0.0011542 0.14865 0.00065825 0.1493 0.13603 0 0.037087 0.0389 0 0.89666 0.24969 0.066972 0.0093546 4.245 0.058421 7.0163e-05 0.83165 0.0052635 0.0060008 0.084275 0.95039 0.97886 0.00024751 0.00080214 0.13177 0.96399 0.92434 0.0088036 0.99597 0.62671 0.004318 0.43175 1.9553 1.9549 15.9959 144.9986 0.00015239 -58.9208 0.99989
1.103 0.98803 5.5188e-05 3.8182 0.012035 1.4519e-05 0.0011542 0.14865 0.00065825 0.14931 0.13604 0 0.037087 0.0389 0 0.89667 0.24969 0.066973 0.0093547 4.245 0.058422 7.0164e-05 0.83165 0.0052635 0.0060008 0.093316 0.94768 0.97755 0.00027892 0.00089679 0.13177 0.9639 0.92434 0.0091847 0.99593 0.62672 0.0044097 0.43173 1.9553 1.9549 15.9959 144.9986 0.00015239 -58.1426 0.99997
1.1031 0.98803 5.5188e-05 3.8182 0.012035 1.452e-05 0.0011542 0.14866 0.00065826 0.14931 0.13604 0 0.037087 0.0389 0 0.89667 0.24969 0.066974 0.0093548 4.245 0.058423 7.0165e-05 0.83165 0.0052635 0.0060008 0.10335 0.9448 0.97612 0.00031461 0.0010031 0.13177 0.9638 0.92434 0.0095783 0.99587 0.62672 0.0045017 0.43172 1.9554 1.9549 15.9959 144.9986 0.0001524 -57.3473 1
1.1031 0.98803 5.5188e-05 3.8182 0.012035 1.4521e-05 0.0011542 0.14866 0.00065826 0.14932 0.13605 0 0.037086 0.0389 0 0.89668 0.2497 0.066975 0.009355 4.245 0.058424 7.0166e-05 0.83165 0.0052636 0.0060009 0.11453 0.94172 0.97455 0.00035533 0.0011228 0.13177 0.96369 0.92434 0.009985 0.99581 0.62673 0.0045942 0.4317 1.9554 1.955 15.9959 144.9986 0.0001524 -56.529 1.0001
1.1032 0.98803 5.5188e-05 3.8182 0.012035 1.4522e-05 0.0011542 0.14867 0.00065826 0.14932 0.13605 0 0.037086 0.0389 0 0.89668 0.2497 0.066976 0.0093551 4.2451 0.058424 7.0167e-05 0.83165 0.0052636 0.0060009 0.12704 0.93843 0.97282 0.00040207 0.0012583 0.13177 0.96357 0.92434 0.010406 0.99574 0.62674 0.0046872 0.43169 1.9554 1.955 15.9959 144.9986 0.0001524 -55.6795 1.0002
1.1033 0.98803 5.5188e-05 3.8182 0.012035 1.4523e-05 0.0011542 0.14867 0.00065826 0.14933 0.13606 0 0.037085 0.0389 0 0.89669 0.2497 0.066977 0.0093552 4.2451 0.058425 7.0168e-05 0.83165 0.0052636 0.0060009 0.13968 0.93526 0.97112 0.00045035 0.0013962 0.13177 0.96346 0.92435 0.010798 0.99566 0.62674 0.0047712 0.43168 1.9554 1.955 15.9959 144.9986 0.0001524 -54.8792 1.0003
1.1034 0.98803 5.5188e-05 3.8182 0.012035 1.4524e-05 0.0011542 0.14868 0.00065826 0.14933 0.13606 0 0.037085 0.0389 0 0.8967 0.2497 0.066977 0.0093553 4.2451 0.058426 7.0169e-05 0.83164 0.0052637 0.006001 0.15239 0.93222 0.96945 0.00049994 0.0015357 0.13177 0.96336 0.92435 0.011162 0.99557 0.62674 0.0048472 0.43166 1.9554 1.955 15.9959 144.9986 0.0001524 -54.1204 1.0004
1.1034 0.98803 5.5188e-05 3.8182 0.012035 1.4525e-05 0.0011542 0.14868 0.00065826 0.14934 0.13607 0 0.037085 0.0389 0 0.8967 0.24971 0.066978 0.0093554 4.2451 0.058426 7.017e-05 0.83164 0.0052637 0.006001 0.16664 0.92897 0.96764 0.00055662 0.0016926 0.13177 0.96324 0.92435 0.011538 0.99547 0.62675 0.0049236 0.43165 1.9555 1.955 15.9959 144.9986 0.00015241 -53.3133 1.0004
1.1035 0.98803 5.5188e-05 3.8182 0.012035 1.4526e-05 0.0011542 0.14869 0.00065826 0.14934 0.13607 0 0.037085 0.0389 0 0.8967 0.24971 0.066979 0.0093555 4.2451 0.058427 7.017e-05 0.83164 0.0052637 0.006001 0.18108 0.92583 0.96586 0.00061511 0.0018517 0.13178 0.96314 0.92435 0.011888 0.99536 0.62675 0.0049927 0.43164 1.9555 1.9551 15.9959 144.9986 0.00015241 -52.5328 1.0005
1.1035 0.98803 5.5188e-05 3.8182 0.012035 1.4526e-05 0.0011542 0.14869 0.00065826 0.14934 0.13608 0 0.037084 0.0389 0 0.89671 0.24971 0.06698 0.0093555 4.2452 0.058427 7.0171e-05 0.83164 0.0052637 0.006001 0.19569 0.9228 0.96413 0.00067525 0.0020126 0.13178 0.96304 0.92435 0.012213 0.99524 0.62675 0.0050553 0.43163 1.9555 1.9551 15.9959 144.9986 0.00015241 -51.7729 1.0005
1.1036 0.98803 5.5188e-05 3.8182 0.012035 1.4527e-05 0.0011542 0.14869 0.00065826 0.14935 0.13608 0 0.037084 0.0389 0 0.89671 0.24971 0.06698 0.0093556 4.2452 0.058428 7.0171e-05 0.83164 0.0052637 0.006001 0.21043 0.91988 0.96245 0.00073689 0.0021747 0.13178 0.96294 0.92435 0.012515 0.99511 0.62675 0.0051119 0.43162 1.9555 1.9551 15.996 144.9986 0.00015241 -51.029 1.0006
1.1036 0.98803 5.5188e-05 3.8182 0.012035 1.4527e-05 0.0011542 0.1487 0.00065826 0.14935 0.13608 0 0.037084 0.0389 0 0.89672 0.24971 0.066981 0.0093557 4.2452 0.058428 7.0172e-05 0.83164 0.0052637 0.006001 0.22528 0.91705 0.96082 0.0007999 0.0023376 0.13178 0.96285 0.92435 0.012796 0.99498 0.62675 0.0051631 0.43161 1.9555 1.9551 15.996 144.9986 0.00015241 -50.2973 1.0006
1.1037 0.98803 5.5188e-05 3.8182 0.012035 1.4528e-05 0.0011542 0.1487 0.00065826 0.14935 0.13608 0 0.037084 0.0389 0 0.89672 0.24971 0.066981 0.0093557 4.2452 0.058429 7.0172e-05 0.83164 0.0052638 0.0060011 0.24197 0.914 0.95906 0.00087178 0.0025202 0.13178 0.96276 0.92435 0.013086 0.99482 0.62676 0.0052147 0.4316 1.9555 1.9551 15.996 144.9986 0.00015242 -49.4906 1.0007
1.1037 0.98803 5.5188e-05 3.8182 0.012035 1.4529e-05 0.0011542 0.1487 0.00065826 0.14936 0.13609 0 0.037084 0.0389 0 0.89672 0.24972 0.066982 0.0093558 4.2452 0.058429 7.0173e-05 0.83164 0.0052638 0.0060011 0.2589 0.91101 0.95735 0.00094591 0.0027052 0.13178 0.96267 0.92435 0.013356 0.99466 0.62676 0.0052615 0.4316 1.9555 1.9551 15.996 144.9986 0.00015242 -48.6831 1.0007
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.4529e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89672 0.24972 0.066982 0.0093559 4.2452 0.058429 7.0173e-05 0.83164 0.0052638 0.0060011 0.27602 0.90805 0.95569 0.0010222 0.0028923 0.13178 0.96258 0.92436 0.013607 0.99448 0.62676 0.005304 0.43159 1.9556 1.9551 15.9961 144.9986 0.00015242 -47.8729 1.0007
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.4529e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2452 0.058429 7.0174e-05 0.83164 0.0052638 0.0060011 0.29327 0.90512 0.95409 0.0011006 0.0030812 0.13178 0.9625 0.92436 0.013842 0.9943 0.62675 0.0053426 0.43158 1.9556 1.9551 15.9961 144.9986 0.00015242 -47.0588 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.4529e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2452 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.29743 0.90441 0.95371 0.0011197 0.0031269 0.13178 0.96249 0.92436 0.013895 0.99426 0.62675 0.0053513 0.43158 1.9556 1.9551 15.9961 144.9986 0.00015242 -46.8626 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2452 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30607 0.90295 0.95294 0.0011597 0.003222 0.13178 0.96245 0.92436 0.014004 0.99416 0.62675 0.0053688 0.43158 1.9556 1.9551 15.9961 144.9986 0.00015242 -46.454 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30663 0.90286 0.95289 0.0011623 0.0032281 0.13178 0.96245 0.92436 0.014011 0.99415 0.62675 0.0053699 0.43158 1.9556 1.9551 15.9961 144.9986 0.00015242 -46.4277 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30775 0.90267 0.95279 0.0011676 0.0032405 0.13178 0.96244 0.92436 0.014025 0.99414 0.62675 0.0053721 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3749 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30789 0.90264 0.95277 0.0011682 0.0032421 0.13178 0.96244 0.92436 0.014027 0.99414 0.62675 0.0053724 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.368 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30818 0.90259 0.95275 0.0011696 0.0032453 0.13178 0.96244 0.92436 0.01403 0.99414 0.62675 0.005373 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3543 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30822 0.90259 0.95275 0.0011698 0.0032457 0.13178 0.96244 0.92436 0.014031 0.99414 0.62675 0.0053731 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3526 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30825 0.90258 0.95274 0.0011699 0.0032461 0.13178 0.96244 0.92436 0.014031 0.99414 0.62675 0.0053731 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3508 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30828 0.90257 0.95274 0.0011701 0.0032464 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053732 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3495 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30828 0.90257 0.95274 0.0011701 0.0032464 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053732 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3493 1.0008
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30829 0.90257 0.95274 0.0011701 0.0032465 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053732 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.349 1.0007
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.3083 0.90257 0.95274 0.0011701 0.0032465 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053732 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3488 1.0006
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.3083 0.90257 0.95274 0.0011701 0.0032466 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053732 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3487 1.0006
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.3083 0.90257 0.95274 0.0011702 0.0032466 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053732 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3484 1.0005
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30832 0.90257 0.95274 0.0011702 0.0032468 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053733 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3478 1.0003
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30834 0.90256 0.95273 0.0011703 0.0032471 0.13178 0.96244 0.92436 0.014032 0.99414 0.62675 0.0053733 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3466 0.99987
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30839 0.90256 0.95273 0.0011706 0.0032476 0.13178 0.96244 0.92436 0.014033 0.99413 0.62675 0.0053734 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3443 0.99909
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30849 0.90254 0.95272 0.001171 0.0032487 0.13178 0.96244 0.92436 0.014034 0.99413 0.62675 0.0053736 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3395 0.99752
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30869 0.90251 0.9527 0.001172 0.0032509 0.13178 0.96244 0.92436 0.014037 0.99413 0.62675 0.005374 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3301 0.99439
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30889 0.90247 0.95269 0.0011729 0.0032531 0.13178 0.96244 0.92436 0.014039 0.99413 0.62675 0.0053744 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3206 0.99127
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30909 0.90244 0.95267 0.0011739 0.0032553 0.13178 0.96244 0.92436 0.014041 0.99413 0.62675 0.0053748 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.3111 0.98816
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.30949 0.90237 0.95263 0.0011757 0.0032598 0.13178 0.96244 0.92436 0.014046 0.99412 0.62675 0.0053756 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.2921 0.98197
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.3099 0.9023 0.9526 0.0011776 0.0032642 0.13178 0.96243 0.92436 0.014051 0.99412 0.62675 0.0053763 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.2731 0.97581
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.3103 0.90223 0.95256 0.0011795 0.0032687 0.13178 0.96243 0.92436 0.014056 0.99411 0.62675 0.0053771 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.254 0.96969
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.0093559 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.31111 0.90209 0.95249 0.0011833 0.0032776 0.13178 0.96243 0.92436 0.014066 0.9941 0.62675 0.0053787 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.2156 0.95756
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.31274 0.90182 0.95235 0.001191 0.0032956 0.13178 0.96242 0.92436 0.014086 0.99409 0.62675 0.0053818 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.1384 0.93376
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.31422 0.90156 0.95222 0.0011979 0.003312 0.13178 0.96242 0.92436 0.014104 0.99407 0.62675 0.0053846 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -46.0682 0.91285
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.31571 0.90131 0.95209 0.001205 0.0033285 0.13178 0.96241 0.92436 0.014121 0.99405 0.62675 0.0053875 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -45.9973 0.8924
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.31722 0.90105 0.95196 0.0012121 0.0033452 0.13178 0.9624 0.92436 0.014139 0.99403 0.62675 0.0053903 0.43158 1.9556 1.9552 15.9961 144.9986 0.00015242 -45.9257 0.87241
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.31874 0.90079 0.95182 0.0012193 0.0033621 0.13178 0.9624 0.92436 0.014157 0.99402 0.62675 0.0053931 0.43158 1.9556 1.9552 15.9962 144.9986 0.00015242 -45.8535 0.85287
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.32183 0.90026 0.95156 0.001234 0.0033963 0.13178 0.96239 0.92436 0.014193 0.99398 0.62675 0.0053988 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015242 -45.707 0.81509
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.32496 0.89972 0.95129 0.001249 0.0034313 0.13178 0.96237 0.92436 0.01423 0.99395 0.62675 0.0054045 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015242 -45.5576 0.77899
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14936 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.32816 0.89917 0.95102 0.0012643 0.0034669 0.13178 0.96236 0.92436 0.014266 0.99391 0.62675 0.0054102 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015242 -45.4052 0.7445
1.1038 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14937 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.33199 0.8985 0.95069 0.0012828 0.0035097 0.13178 0.96235 0.92436 0.014309 0.99386 0.62675 0.0054169 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015242 -45.2223 0.7059
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14937 0.13609 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0174e-05 0.83164 0.0052638 0.0060011 0.33591 0.89782 0.95036 0.0013018 0.0035536 0.13178 0.96233 0.92436 0.014353 0.99382 0.62675 0.0054236 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015243 -45.0349 0.66931
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0175e-05 0.83164 0.0052638 0.0060011 0.33991 0.89711 0.95003 0.0013213 0.0035986 0.13178 0.96232 0.92436 0.014397 0.99377 0.62675 0.0054304 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015243 -44.8429 0.63461
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0175e-05 0.83164 0.0052638 0.0060011 0.344 0.89638 0.94969 0.0013414 0.0036447 0.13178 0.9623 0.92436 0.014441 0.99372 0.62675 0.0054372 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015243 -44.6461 0.60172
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.453e-05 0.0011542 0.14871 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89673 0.24972 0.066983 0.009356 4.2453 0.05843 7.0175e-05 0.83164 0.0052638 0.0060011 0.34819 0.89563 0.94934 0.0013621 0.0036921 0.13178 0.96229 0.92436 0.014486 0.99367 0.62675 0.005444 0.43157 1.9556 1.9552 15.9962 144.9986 0.00015243 -44.4444 0.57052
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14871 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89673 0.24972 0.066984 0.009356 4.2453 0.05843 7.0175e-05 0.83164 0.0052638 0.0060011 0.35685 0.89404 0.94863 0.0014054 0.0037907 0.13178 0.96225 0.92436 0.014577 0.99356 0.62675 0.0054577 0.43157 1.9556 1.9552 15.9963 144.9986 0.00015243 -44.0251 0.51291
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14871 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89673 0.24972 0.066984 0.0093561 4.2453 0.05843 7.0175e-05 0.83164 0.0052638 0.0060011 0.36591 0.89233 0.9479 0.0014515 0.003895 0.13178 0.96222 0.92436 0.014669 0.99345 0.62675 0.0054715 0.43156 1.9556 1.9552 15.9963 144.9986 0.00015243 -43.5831 0.46111
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066984 0.0093561 4.2453 0.05843 7.0175e-05 0.83164 0.0052638 0.0060011 0.37541 0.89047 0.94715 0.0015007 0.0040055 0.13178 0.96219 0.92436 0.014763 0.99333 0.62675 0.0054854 0.43156 1.9556 1.9552 15.9963 144.9986 0.00015243 -43.1164 0.41454
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066984 0.0093561 4.2453 0.058431 7.0175e-05 0.83164 0.0052638 0.0060011 0.38537 0.88844 0.94637 0.0015532 0.0041228 0.13178 0.96216 0.92436 0.014859 0.9932 0.62675 0.0054994 0.43156 1.9556 1.9552 15.9963 144.9986 0.00015243 -42.6228 0.37268
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066984 0.0093561 4.2453 0.058431 7.0175e-05 0.83164 0.0052638 0.0060011 0.39583 0.88619 0.94556 0.0016096 0.0042478 0.13178 0.96212 0.92436 0.014957 0.99307 0.62674 0.0055137 0.43156 1.9556 1.9552 15.9964 144.9986 0.00015243 -42.0999 0.33504
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066984 0.0093561 4.2453 0.058431 7.0175e-05 0.83164 0.0052638 0.0060012 0.4068 0.88367 0.94472 0.0016701 0.0043813 0.13178 0.96209 0.92436 0.015058 0.99292 0.62674 0.0055281 0.43155 1.9556 1.9552 15.9964 144.9986 0.00015243 -41.545 0.30121
1.1039 0.98803 5.5188e-05 3.8182 0.012035 1.4531e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066984 0.0093561 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.41832 0.88082 0.94385 0.0017355 0.0045245 0.13178 0.96206 0.92436 0.015161 0.99277 0.62674 0.0055427 0.43155 1.9556 1.9552 15.9964 144.9986 0.00015243 -40.9553 0.27079
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43044 0.87755 0.94295 0.0018063 0.0046784 0.13178 0.96202 0.92436 0.015267 0.9926 0.62674 0.0055576 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -40.3275 0.24345
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43239 0.87699 0.94281 0.0018179 0.0047036 0.13178 0.96201 0.92436 0.015284 0.99258 0.62674 0.0055599 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -40.2254 0.23942
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43634 0.87583 0.94252 0.0018416 0.0047549 0.13178 0.962 0.92436 0.015318 0.99252 0.62674 0.0055647 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -40.0182 0.23157
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43663 0.87574 0.9425 0.0018434 0.0047588 0.13178 0.962 0.92436 0.015321 0.99252 0.62674 0.005565 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -40.0028 0.231
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43687 0.87565 0.94248 0.0018448 0.0047619 0.13178 0.962 0.92436 0.015323 0.99251 0.62674 0.0055653 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.9902 0.23054
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43708 0.87557 0.94246 0.0018461 0.0047646 0.13178 0.962 0.92436 0.015325 0.99251 0.62674 0.0055656 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.9792 0.23014
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037083 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.4375 0.87541 0.94243 0.0018486 0.0047701 0.13178 0.962 0.92436 0.015328 0.99251 0.62674 0.0055661 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.9571 0.22934
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43792 0.87526 0.9424 0.0018512 0.0047756 0.13178 0.962 0.92436 0.015332 0.9925 0.62674 0.0055666 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.935 0.22854
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43834 0.8751 0.94237 0.0018537 0.0047811 0.13178 0.962 0.92436 0.015335 0.99249 0.62674 0.0055671 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.9129 0.22774
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.43919 0.87478 0.94231 0.0018589 0.0047922 0.13178 0.96199 0.92436 0.015343 0.99248 0.62674 0.005568 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.8684 0.22615
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.44003 0.87447 0.94225 0.001864 0.0048033 0.13178 0.96199 0.92436 0.01535 0.99247 0.62674 0.0055691 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.8238 0.22458
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.44088 0.87415 0.94219 0.0018692 0.0048145 0.13178 0.96199 0.92436 0.015357 0.99246 0.62674 0.0055701 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.779 0.22301
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.44259 0.87351 0.94206 0.0018797 0.004837 0.13178 0.96198 0.92436 0.015372 0.99244 0.62674 0.0055721 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.6888 0.21991
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.44603 0.87222 0.94181 0.0019009 0.0048828 0.13178 0.96197 0.92436 0.015401 0.99239 0.62674 0.0055761 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.5061 0.21384
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.44952 0.87091 0.94155 0.0019227 0.0049296 0.13178 0.96196 0.92436 0.015431 0.99234 0.62673 0.0055802 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.3203 0.20794
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.45306 0.86958 0.94129 0.001945 0.0049774 0.13178 0.96195 0.92436 0.015461 0.99229 0.62673 0.0055842 0.43155 1.9556 1.9552 15.9965 144.9986 0.00015243 -39.1313 0.2022
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.45664 0.86823 0.94103 0.0019678 0.0050262 0.13178 0.96194 0.92436 0.015491 0.99224 0.62673 0.0055883 0.43155 1.9556 1.9552 15.9966 144.9986 0.00015243 -38.939 0.19662
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.46395 0.86548 0.9405 0.0020151 0.0051273 0.13178 0.96192 0.92436 0.015552 0.99214 0.62673 0.0055966 0.43155 1.9556 1.9552 15.9966 144.9986 0.00015243 -38.5444 0.18591
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14937 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.47145 0.86264 0.93995 0.0020648 0.0052332 0.13178 0.9619 0.92436 0.015615 0.99204 0.62673 0.0056051 0.43154 1.9556 1.9552 15.9966 144.9986 0.00015243 -38.1357 0.1758
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14938 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.47914 0.85971 0.93939 0.002117 0.0053441 0.13178 0.96188 0.92436 0.015679 0.99193 0.62673 0.0056136 0.43154 1.9556 1.9552 15.9966 144.9986 0.00015243 -37.7124 0.16623
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14938 0.1361 0 0.037082 0.0389 0 0.89674 0.24973 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.48703 0.85668 0.93881 0.002172 0.0054605 0.13178 0.96186 0.92436 0.015744 0.99182 0.62673 0.0056223 0.43154 1.9556 1.9552 15.9967 144.9986 0.00015244 -37.2738 0.15718
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14938 0.1361 0 0.037082 0.0389 0 0.89674 0.24973 0.066985 0.0093562 4.2453 0.058431 7.0176e-05 0.83164 0.0052639 0.0060012 0.49512 0.85356 0.93822 0.0022301 0.005583 0.13178 0.96184 0.92436 0.015811 0.99171 0.62672 0.0056311 0.43154 1.9556 1.9552 15.9967 144.9986 0.00015244 -36.8193 0.14863
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4532e-05 0.0011542 0.14872 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89674 0.24973 0.066985 0.0093562 4.2453 0.058432 7.0176e-05 0.83164 0.0052639 0.0060012 0.51192 0.84696 0.93698 0.0023562 0.0058478 0.13178 0.96179 0.92436 0.015951 0.99147 0.62672 0.0056493 0.43154 1.9556 1.9552 15.9968 144.9986 0.00015244 -35.8594 0.13289
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14872 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89674 0.24973 0.066985 0.0093563 4.2453 0.058432 7.0176e-05 0.83164 0.0052639 0.0060012 0.52753 0.8407 0.93582 0.002481 0.0061083 0.13178 0.96175 0.92436 0.016081 0.99126 0.62672 0.0056662 0.43154 1.9556 1.9552 15.9968 144.9986 0.00015244 -34.9476 0.12033
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14872 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093563 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.54379 0.83399 0.9346 0.0026199 0.0063969 0.13178 0.96171 0.92436 0.01622 0.99103 0.62671 0.0056838 0.43153 1.9556 1.9552 15.9969 144.9986 0.00015244 -33.9749 0.10895
1.104 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093563 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.56071 0.82677 0.93331 0.0027754 0.0067185 0.13178 0.96166 0.92436 0.016367 0.9908 0.62671 0.0057024 0.43153 1.9556 1.9552 15.997 144.9986 0.00015244 -32.9373 0.098659
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093563 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.57827 0.81899 0.93195 0.0029506 0.007079 0.13178 0.96161 0.92436 0.016525 0.99056 0.6267 0.005722 0.43153 1.9556 1.9552 15.997 144.9986 0.00015244 -31.831 0.089338
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093563 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.59646 0.81056 0.93051 0.0031491 0.0074857 0.13178 0.96156 0.92436 0.016697 0.99032 0.62669 0.0057431 0.43153 1.9556 1.9552 15.9971 144.9986 0.00015244 -30.6525 0.080898
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093563 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.61523 0.8014 0.92898 0.0033754 0.0079476 0.13178 0.96151 0.92436 0.016884 0.99007 0.62668 0.0057657 0.43153 1.9556 1.9552 15.9972 144.9986 0.00015244 -29.3989 0.073256
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093563 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.63453 0.79142 0.92738 0.0036352 0.0084759 0.13178 0.96145 0.92436 0.01709 0.98981 0.62668 0.0057904 0.43152 1.9556 1.9552 15.9973 144.9986 0.00015244 -28.0679 0.066336
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4533e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093564 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.6543 0.78051 0.92568 0.0039355 0.0090844 0.13178 0.96139 0.92436 0.017319 0.98955 0.62667 0.0058176 0.43152 1.9556 1.9552 15.9974 144.9986 0.00015244 -26.6583 0.060072
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093564 4.2453 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.67444 0.76855 0.9239 0.0042849 0.0097903 0.13178 0.96132 0.92436 0.017576 0.98929 0.62665 0.0058477 0.43152 1.9557 1.9552 15.9975 144.9986 0.00015245 -25.1702 0.0544
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066986 0.0093564 4.2454 0.058432 7.0177e-05 0.83164 0.0052639 0.0060012 0.69484 0.75545 0.92202 0.0046943 0.010615 0.13178 0.96125 0.92436 0.017868 0.98902 0.62664 0.0058815 0.43152 1.9557 1.9552 15.9976 144.9986 0.00015245 -23.6054 0.049264
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14938 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066987 0.0093564 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.7154 0.74109 0.92006 0.0051772 0.011585 0.13178 0.96116 0.92436 0.018202 0.98875 0.62662 0.0059196 0.43152 1.9557 1.9552 15.9977 144.9986 0.00015245 -21.9674 0.044615
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14939 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066987 0.0093564 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.73595 0.72537 0.91801 0.0057502 0.012734 0.13178 0.96107 0.92436 0.018586 0.98848 0.6266 0.0059631 0.43151 1.9557 1.9552 15.9978 144.9986 0.00015245 -20.262 0.040404
1.1041 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14939 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066987 0.0093564 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.75637 0.70822 0.91588 0.0064341 0.014102 0.13178 0.96097 0.92436 0.019032 0.9882 0.62658 0.0060129 0.43151 1.9557 1.9552 15.998 144.9986 0.00015245 -18.497 0.036593
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14939 0.13611 0 0.037082 0.0389 0 0.89675 0.24973 0.066987 0.0093564 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.77648 0.68959 0.91368 0.0072539 0.015738 0.13178 0.96086 0.92436 0.01955 0.98793 0.62655 0.0060702 0.43151 1.9557 1.9552 15.9981 144.9986 0.00015245 -16.6825 0.033141
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14939 0.13612 0 0.037082 0.0389 0 0.89676 0.24973 0.066987 0.0093565 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.79613 0.66948 0.91141 0.0082404 0.017703 0.13178 0.96073 0.92436 0.020153 0.98765 0.62651 0.0061364 0.43151 1.9557 1.9553 15.9982 144.9986 0.00015245 -14.8307 0.030016
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4534e-05 0.0011542 0.14873 0.00065826 0.14939 0.13612 0 0.037082 0.0389 0 0.89676 0.24973 0.066987 0.0093565 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.81515 0.64795 0.90907 0.0094303 0.020069 0.13178 0.96059 0.92436 0.020855 0.98737 0.62647 0.0062127 0.43151 1.9557 1.9553 15.9984 144.9986 0.00015246 -12.9552 0.027187
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14873 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066987 0.0093565 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.83341 0.62511 0.90669 0.010867 0.022919 0.13178 0.96043 0.92436 0.021671 0.98709 0.62642 0.0063006 0.4315 1.9557 1.9553 15.9985 144.9986 0.00015246 -11.0711 0.024625
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066987 0.0093565 4.2454 0.058433 7.0178e-05 0.83164 0.0052639 0.0060012 0.85075 0.60112 0.90426 0.0126 0.02635 0.13178 0.96025 0.92436 0.022612 0.98682 0.62636 0.0064014 0.4315 1.9557 1.9553 15.9986 144.9986 0.00015246 -9.1937 0.022305
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093565 4.2454 0.058433 7.0179e-05 0.83164 0.0052639 0.0060012 0.86709 0.57621 0.9018 0.014687 0.030472 0.13178 0.96005 0.92436 0.023693 0.98654 0.62629 0.0065164 0.4315 1.9557 1.9553 15.9988 144.9986 0.00015246 -7.3382 0.020205
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093565 4.2454 0.058433 7.0179e-05 0.83164 0.0052639 0.0060012 0.88231 0.55063 0.89931 0.017192 0.035405 0.13178 0.95983 0.92436 0.024925 0.98626 0.62621 0.0066468 0.4315 1.9557 1.9553 15.9989 144.9986 0.00015246 -5.5191 0.018304
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058433 7.0179e-05 0.83164 0.005264 0.0060013 0.89638 0.52464 0.8968 0.020183 0.041277 0.13178 0.95959 0.92436 0.026315 0.98598 0.62612 0.0067933 0.4315 1.9557 1.9553 15.999 144.9986 0.00015246 -3.7493 0.016582
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.90926 0.49852 0.89427 0.023731 0.04822 0.13178 0.95933 0.92436 0.027873 0.9857 0.62602 0.0069569 0.43149 1.9557 1.9553 15.9991 144.9986 0.00015247 -2.0397 0.015023
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.91787 0.47961 0.89242 0.026702 0.054012 0.13178 0.95913 0.92436 0.029111 0.9855 0.62593 0.0070867 0.43149 1.9557 1.9553 15.9992 144.9986 0.00015247 -0.84053 0.013984
1.1042 0.98803 5.5188e-05 3.8182 0.012035 1.4535e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.92586 0.46085 0.89057 0.030035 0.060488 0.13178 0.95891 0.92436 0.030441 0.98529 0.62585 0.0072259 0.43149 1.9557 1.9553 15.9993 144.9986 0.00015247 0.31947 0.013017
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.93253 0.44417 0.88889 0.033366 0.066938 0.13178 0.95871 0.92436 0.031715 0.98511 0.62576 0.0073591 0.43149 1.9557 1.9553 15.9994 144.9986 0.00015247 1.3282 0.012204
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.93871 0.42773 0.88722 0.037032 0.07401 0.13178 0.95851 0.92436 0.033064 0.98493 0.62568 0.0075001 0.43149 1.9557 1.9553 15.9995 144.9986 0.00015247 2.3024 0.011443
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.94443 0.41157 0.88554 0.041051 0.08173 0.13178 0.9583 0.92436 0.034486 0.98475 0.62559 0.0076486 0.43149 1.9557 1.9552 15.9995 144.9986 0.00015248 3.2413 0.01073
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.14939 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.9497 0.39575 0.88387 0.045438 0.090121 0.13178 0.95808 0.92436 0.03598 0.98456 0.6255 0.0078048 0.43149 1.9557 1.9552 15.9996 144.9986 0.00015248 4.1445 0.010061
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.1494 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066988 0.0093566 4.2454 0.058434 7.0179e-05 0.83164 0.005264 0.0060013 0.95455 0.38028 0.88219 0.050209 0.099202 0.13178 0.95786 0.92435 0.037545 0.98438 0.6254 0.0079684 0.43148 1.9557 1.9552 15.9996 144.9986 0.00015248 5.012 0.0094343
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.1494 0.13612 0 0.037081 0.0389 0 0.89676 0.24973 0.066989 0.0093566 4.2454 0.058434 7.018e-05 0.83164 0.005264 0.0060013 0.95899 0.36519 0.88051 0.055376 0.10899 0.13178 0.95763 0.92435 0.039181 0.9842 0.6253 0.0081394 0.43148 1.9557 1.9552 15.9997 144.9986 0.00015248 5.8438 0.0088472
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.1494 0.13612 0 0.037081 0.0389 0 0.89677 0.24973 0.066989 0.0093567 4.2454 0.058434 7.018e-05 0.83164 0.005264 0.0060013 0.96305 0.35051 0.87883 0.06095 0.11948 0.13178 0.95739 0.92435 0.040884 0.98402 0.6252 0.0083176 0.43148 1.9557 1.9551 15.9998 144.9986 0.00015249 6.6404 0.0082969
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.1494 0.13612 0 0.037081 0.0389 0 0.89677 0.24974 0.066989 0.0093567 4.2454 0.058434 7.018e-05 0.83164 0.005264 0.0060013 0.96675 0.33625 0.87716 0.066939 0.13068 0.13178 0.95716 0.92435 0.042654 0.98383 0.6251 0.0085029 0.43148 1.9557 1.9551 15.9998 144.9986 0.00015249 7.4023 0.0077813
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.1494 0.13612 0 0.037081 0.0389 0 0.89677 0.24974 0.066989 0.0093567 4.2454 0.058434 7.018e-05 0.83164 0.005264 0.0060013 0.97317 0.30904 0.8738 0.080181 0.1552 0.13178 0.95667 0.92435 0.046386 0.98347 0.6249 0.0088943 0.43148 1.9557 1.9549 15.9999 144.9986 0.00015251 8.8252 0.0068453
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4536e-05 0.0011542 0.14874 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.066989 0.0093567 4.2454 0.058434 7.018e-05 0.83164 0.005264 0.0060013 0.97843 0.28358 0.87046 0.095119 0.18244 0.13178 0.95617 0.92435 0.05036 0.9831 0.62468 0.0093121 0.43147 1.9557 1.9545 16 144.9986 0.00015253 10.1198 0.0060234
1.1043 0.98803 5.5188e-05 3.8182 0.012035 1.4537e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.066989 0.0093567 4.2454 0.058434 7.018e-05 0.83164 0.005264 0.0060013 0.98272 0.25989 0.86712 0.11172 0.21219 0.13178 0.95567 0.92434 0.054557 0.98274 0.62447 0.0097547 0.43147 1.9557 1.9541 16.0001 144.9986 0.00015255 11.2946 0.0053017
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4537e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.066989 0.0093567 4.2454 0.058435 7.018e-05 0.83164 0.005264 0.0060013 0.98617 0.23793 0.86379 0.12993 0.24418 0.13178 0.95515 0.92434 0.058961 0.98237 0.62425 0.010221 0.43147 1.9557 1.9534 16.0001 144.9986 0.00015259 12.3588 0.0046678
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4537e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.06699 0.0093568 4.2454 0.058435 7.018e-05 0.83164 0.005264 0.0060013 0.98895 0.21762 0.86046 0.14965 0.27807 0.13178 0.95463 0.92433 0.063552 0.98201 0.62403 0.010708 0.43147 1.9557 1.9524 16.0002 144.9986 0.00015264 13.3216 0.0041112
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4537e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.06699 0.0093568 4.2454 0.058435 7.0181e-05 0.83164 0.005264 0.0060013 0.99117 0.19889 0.85715 0.17074 0.31346 0.13178 0.9541 0.92433 0.068314 0.98164 0.62381 0.011216 0.43146 1.9557 1.9511 16.0003 144.9986 0.00015271 14.1921 0.0036225
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4537e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.06699 0.0093568 4.2454 0.058435 7.0181e-05 0.83164 0.005264 0.0060013 0.99293 0.18166 0.85385 0.19306 0.34993 0.13178 0.95357 0.92433 0.073228 0.98128 0.62358 0.011743 0.43146 1.9557 1.9495 16.0003 144.9986 0.00015279 14.9787 0.0031933
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4537e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.037081 0.0389 0 0.89677 0.24974 0.06699 0.0093568 4.2454 0.058435 7.0181e-05 0.83164 0.005264 0.0060013 0.99433 0.16582 0.85055 0.21643 0.38708 0.13178 0.95304 0.92432 0.07828 0.98092 0.62336 0.012287 0.43146 1.9557 1.9474 16.0004 144.9986 0.0001529 15.6894 0.0028163
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14875 0.00065826 0.1494 0.13613 0 0.03708 0.0389 0 0.89677 0.24974 0.06699 0.0093568 4.2455 0.058435 7.0181e-05 0.83163 0.005264 0.0060013 0.99543 0.1513 0.84727 0.24069 0.42447 0.13178 0.9525 0.92431 0.083454 0.98055 0.62314 0.012847 0.43146 1.9557 1.9449 16.0004 144.9986 0.00015303 16.3318 0.0024854
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14875 0.00065826 0.14941 0.13613 0 0.03708 0.0389 0 0.89678 0.24974 0.06699 0.0093569 4.2455 0.058435 7.0181e-05 0.83163 0.005264 0.0060013 0.99629 0.13799 0.844 0.26566 0.46171 0.13178 0.95196 0.92431 0.088735 0.98019 0.62291 0.013421 0.43145 1.9557 1.942 16.0004 144.9986 0.00015318 16.9126 0.0021947
1.1044 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14875 0.00065826 0.14941 0.13613 0 0.03708 0.0389 0 0.89678 0.24974 0.06699 0.0093569 4.2455 0.058435 7.0181e-05 0.83163 0.005264 0.0060013 0.99697 0.12581 0.84074 0.29115 0.49845 0.13178 0.95142 0.9243 0.09411 0.97982 0.62268 0.014009 0.43145 1.9556 1.9385 16.0005 144.9986 0.00015336 17.4379 0.0019395
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14875 0.00065826 0.14941 0.13613 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0181e-05 0.83163 0.005264 0.0060013 0.99751 0.11467 0.83749 0.31699 0.53437 0.13178 0.95088 0.92429 0.099568 0.97946 0.62246 0.014609 0.43145 1.9556 1.9344 16.0005 144.9986 0.00015357 17.9132 0.0017153
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14875 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.99793 0.10448 0.83425 0.34301 0.56921 0.13178 0.95034 0.92429 0.1051 0.9791 0.62223 0.01522 0.43145 1.9555 1.9296 16.0005 144.9986 0.00015381 18.3437 0.0015185
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14875 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.99799 0.10273 0.83367 0.34774 0.57539 0.13178 0.95024 0.92428 0.10611 0.97903 0.62219 0.015332 0.43144 1.9555 1.9287 16.0005 144.9986 0.00015386 18.4174 0.0014854
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.99811 0.099315 0.8325 0.3572 0.58762 0.13178 0.95005 0.92428 0.10813 0.9789 0.62211 0.015557 0.43144 1.9555 1.9268 16.0005 144.9986 0.00015396 18.5608 0.001451
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4538e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.99823 0.09601 0.83133 0.36665 0.59967 0.13178 0.94985 0.92428 0.11016 0.97877 0.62203 0.015783 0.43144 1.9555 1.9247 16.0005 144.9986 0.00015406 18.6993 0.0014539
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.99833 0.092812 0.83016 0.3761 0.61153 0.13178 0.94965 0.92427 0.1122 0.97864 0.62194 0.016011 0.43144 1.9555 1.9227 16.0005 144.9986 0.00015417 18.8329 0.0014676
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.0093569 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.99842 0.089718 0.82899 0.38552 0.62318 0.13178 0.94945 0.92427 0.11425 0.9785 0.62186 0.016239 0.43144 1.9554 1.9205 16.0005 144.9986 0.00015428 18.962 0.0014738
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060013 0.9985 0.087019 0.82795 0.39397 0.63349 0.13178 0.94928 0.92427 0.11609 0.97838 0.62179 0.016446 0.43144 1.9554 1.9186 16.0006 144.9986 0.00015439 19.0743 0.001475
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060014 0.99857 0.084401 0.8269 0.40241 0.64362 0.13178 0.9491 0.92426 0.11794 0.97827 0.62171 0.016654 0.43144 1.9554 1.9165 16.0006 144.9986 0.00015449 19.1831 0.0014771
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.005264 0.0060014 0.99864 0.081859 0.82585 0.41081 0.65358 0.13178 0.94892 0.92426 0.1198 0.97815 0.62164 0.016862 0.43144 1.9554 1.9144 16.0006 144.9986 0.0001546 19.2886 0.0014811
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.0052641 0.0060014 0.9987 0.079393 0.82481 0.41918 0.66336 0.13178 0.94875 0.92426 0.12166 0.97803 0.62156 0.017072 0.43144 1.9553 1.9122 16.0006 144.9986 0.00015472 19.3909 0.0014859
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.0052641 0.0060014 0.99876 0.077 0.82376 0.42752 0.67296 0.13178 0.94857 0.92425 0.12352 0.97791 0.62149 0.017282 0.43144 1.9553 1.9099 16.0006 144.9986 0.00015484 19.49 0.0014905
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.0052641 0.0060014 0.99881 0.074677 0.82272 0.43582 0.68238 0.13178 0.94839 0.92425 0.12539 0.97779 0.62141 0.017493 0.43144 1.9553 1.9076 16.0006 144.9986 0.00015496 19.5862 0.0014948
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.0052641 0.0060014 0.99886 0.072424 0.82168 0.44407 0.69161 0.13178 0.94821 0.92424 0.12725 0.97767 0.62134 0.017705 0.43143 1.9552 1.9051 16.0006 144.9986 0.00015509 19.6794 0.0014989
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066991 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.0052641 0.0060014 0.99895 0.068115 0.8196 0.46043 0.70951 0.13178 0.94786 0.92424 0.131 0.97744 0.62119 0.018131 0.43143 1.9552 1.8999 16.0006 144.9986 0.00015536 19.8576 0.0015068
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066992 0.009357 4.2455 0.058436 7.0182e-05 0.83163 0.0052641 0.0060014 0.99902 0.06406 0.81753 0.47658 0.72665 0.13178 0.9475 0.92423 0.13476 0.9772 0.62104 0.01856 0.43143 1.9551 1.8942 16.0006 144.9986 0.00015567 20.0254 0.0015149
1.1045 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89678 0.24974 0.066992 0.009357 4.2455 0.058436 7.0183e-05 0.83163 0.0052641 0.0060014 0.99909 0.060242 0.81546 0.49251 0.74304 0.13178 0.94715 0.92422 0.13852 0.97696 0.62089 0.018992 0.43143 1.955 1.888 16.0006 144.9986 0.000156 20.1836 0.0015233
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.4539e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89679 0.24974 0.066992 0.009357 4.2455 0.058436 7.0183e-05 0.83163 0.0052641 0.0060014 0.99914 0.056649 0.8134 0.50818 0.75867 0.13178 0.94679 0.9242 0.14229 0.97673 0.62075 0.019426 0.43143 1.9549 1.8811 16.0006 144.9986 0.00015637 20.3328 0.0015319
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14941 0.13614 0 0.03708 0.0389 0 0.89679 0.24974 0.066992 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99919 0.053268 0.81134 0.52358 0.77356 0.13178 0.94644 0.92419 0.14607 0.97649 0.6206 0.019862 0.43143 1.9548 1.8734 16.0006 144.9986 0.00015678 20.4737 0.0015405
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24974 0.066992 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99923 0.050087 0.80929 0.5387 0.78771 0.13178 0.94608 0.92418 0.14985 0.97625 0.62045 0.020301 0.43142 1.9547 1.8648 16.0006 144.9986 0.00015724 20.6069 0.0015489
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24974 0.066992 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99926 0.047094 0.80724 0.55353 0.80115 0.13178 0.94573 0.92417 0.15363 0.97602 0.6203 0.020742 0.43142 1.9546 1.8553 16.0006 144.9986 0.00015775 20.733 0.0015574
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24974 0.066992 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99929 0.044278 0.8052 0.56806 0.81388 0.13178 0.94537 0.92415 0.15742 0.97578 0.62015 0.021185 0.43142 1.9544 1.8446 16.0006 144.9986 0.00015833 20.8525 0.0015659
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24975 0.066992 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99932 0.041629 0.80316 0.58227 0.82593 0.13178 0.94502 0.92414 0.1612 0.97554 0.62 0.021629 0.43142 1.9543 1.8326 16.0006 144.9986 0.00015898 20.9659 0.0015744
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24975 0.066992 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99934 0.039137 0.80113 0.59616 0.83733 0.13178 0.94466 0.92412 0.16499 0.97531 0.61985 0.022076 0.43142 1.9541 1.8193 16.0006 144.9985 0.00015971 21.0737 0.0015829
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14876 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24975 0.066993 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99936 0.036793 0.79911 0.60973 0.84808 0.13178 0.94431 0.9241 0.16877 0.97507 0.6197 0.022524 0.43142 1.9539 1.8045 16.0006 144.9985 0.00016053 21.1763 0.0015914
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14877 0.00065826 0.14942 0.13614 0 0.03708 0.0389 0 0.89679 0.24975 0.066993 0.0093571 4.2455 0.058437 7.0183e-05 0.83163 0.0052641 0.0060014 0.99938 0.034588 0.79708 0.62297 0.85822 0.13178 0.94395 0.92408 0.17255 0.97483 0.61956 0.022974 0.43141 1.9537 1.788 16.0006 144.9985 0.00016144 21.2742 0.0015999
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.454e-05 0.0011542 0.14877 0.00065826 0.14942 0.13615 0 0.037079 0.0389 0 0.89679 0.24975 0.066993 0.0093572 4.2455 0.058437 7.0184e-05 0.83163 0.0052641 0.0060014 0.9994 0.032515 0.79507 0.63589 0.86776 0.13178 0.9436 0.92406 0.17632 0.9746 0.61941 0.023426 0.43141 1.9534 1.77 16.0006 144.9985 0.00016246 21.3676 0.0016084
1.1046 0.98803 5.5188e-05 3.8182 0.012035 1.4541e-05 0.0011542 0.14877 0.00065826 0.14942 0.13615 0 0.037079 0.0389 0 0.89679 0.24975 0.066993 0.0093572 4.2455 0.058437 7.0184e-05 0.83163 0.0052641 0.0060014 0.99942 0.028731 0.79105 0.66071 0.88518 0.13178 0.94289 0.92402 0.18386 0.97412 0.61911 0.024333 0.43141 1.9529 1.7292 16.0006 144.9985 0.0001648 21.5426 0.0016254
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4541e-05 0.0011542 0.14877 0.00065826 0.14942 0.13615 0 0.037079 0.0389 0 0.89679 0.24975 0.066993 0.0093572 4.2455 0.058437 7.0184e-05 0.83163 0.0052641 0.0060014 0.99944 0.025804 0.78757 0.68119 0.89862 0.13178 0.94227 0.92397 0.19039 0.97371 0.61885 0.025124 0.43141 1.9523 1.689 16.0006 144.9985 0.00016717 21.6834 0.0016401
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4541e-05 0.0011542 0.14877 0.00065826 0.14942 0.13615 0 0.037079 0.0389 0 0.89679 0.24975 0.066993 0.0093572 4.2455 0.058438 7.0184e-05 0.83163 0.0052641 0.0060014 0.99946 0.023424 0.78446 0.69878 0.9095 0.13178 0.94172 0.92393 0.19624 0.97335 0.61862 0.02584 0.4314 1.9517 1.6501 16.0006 144.9985 0.00016954 21.8024 0.0016534
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4541e-05 0.0011542 0.14877 0.00065826 0.14942 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066993 0.0093572 4.2455 0.058438 7.0184e-05 0.83163 0.0052641 0.0060014 0.99947 0.021469 0.78167 0.71393 0.91837 0.13178 0.94122 0.92389 0.2015 0.97301 0.61841 0.026487 0.4314 1.9511 1.6136 16.0006 144.9985 0.00017182 21.9042 0.0016653
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4541e-05 0.0011542 0.14877 0.00065826 0.14942 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093573 4.2455 0.058438 7.0184e-05 0.83163 0.0052641 0.0060014 0.99948 0.019677 0.77889 0.72846 0.92645 0.13178 0.94072 0.92384 0.20674 0.97268 0.6182 0.027135 0.4314 1.9504 1.5764 16.0006 144.9985 0.00017423 22.0015 0.0016772
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14877 0.00065826 0.14943 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093573 4.2455 0.058438 7.0184e-05 0.83163 0.0052641 0.0060014 0.99949 0.018034 0.77612 0.74238 0.93379 0.13178 0.94022 0.92379 0.21196 0.97235 0.61799 0.027786 0.4314 1.9496 1.5391 16.0006 144.9985 0.00017671 22.0949 0.0016892
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14877 0.00065826 0.14943 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093573 4.2456 0.058438 7.0185e-05 0.83163 0.0052641 0.0060014 0.99949 0.016527 0.77336 0.75569 0.94045 0.13178 0.93973 0.92374 0.21717 0.97202 0.61778 0.028439 0.43139 1.9488 1.5023 16.0006 144.9985 0.00017925 22.1849 0.0017011
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14877 0.00065826 0.14943 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093573 4.2456 0.058438 7.0185e-05 0.83163 0.0052641 0.0060014 0.9995 0.015146 0.77061 0.76843 0.94648 0.13178 0.93923 0.92368 0.22236 0.97169 0.61758 0.029093 0.43139 1.9479 1.4665 16.0006 144.9985 0.00018181 22.2718 0.001713
1.1047 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14877 0.00065826 0.14943 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093573 4.2456 0.058438 7.0185e-05 0.83163 0.0052641 0.0060014 0.99951 0.01388 0.76787 0.7806 0.95195 0.13178 0.93873 0.92362 0.22753 0.97136 0.61737 0.02975 0.43139 1.9469 1.4317 16.0006 144.9985 0.00018438 22.356 0.001725
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14877 0.00065826 0.14943 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093573 4.2456 0.058438 7.0185e-05 0.83163 0.0052641 0.0060014 0.99951 0.012719 0.76513 0.79222 0.95689 0.13178 0.93824 0.92355 0.23268 0.97103 0.61716 0.030408 0.43139 1.9458 1.3984 16.0006 144.9985 0.00018693 22.4379 0.0017369
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14878 0.00065826 0.14943 0.13615 0 0.037079 0.0389 0 0.8968 0.24975 0.066994 0.0093574 4.2456 0.058438 7.0185e-05 0.83163 0.0052641 0.0060014 0.99952 0.011655 0.76241 0.8033 0.96135 0.13178 0.93774 0.92348 0.23782 0.97069 0.61695 0.031068 0.43138 1.9447 1.3664 16.0006 144.9985 0.00018946 22.5177 0.0017488
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4542e-05 0.0011542 0.14878 0.00065826 0.14943 0.13616 0 0.037079 0.0389 0 0.8968 0.24975 0.066995 0.0093574 4.2456 0.058439 7.0185e-05 0.83163 0.0052641 0.0060015 0.99952 0.010679 0.7597 0.81387 0.96538 0.13178 0.93724 0.92341 0.24293 0.97036 0.61674 0.031729 0.43138 1.9436 1.3359 16.0006 144.9984 0.00019197 22.5957 0.0017608
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4543e-05 0.0011542 0.14878 0.00065826 0.14943 0.13616 0 0.037079 0.0389 0 0.8968 0.24975 0.066995 0.0093574 4.2456 0.058439 7.0185e-05 0.83163 0.0052642 0.0060015 0.99953 0.0097851 0.757 0.82395 0.96901 0.13178 0.93675 0.92334 0.24802 0.97003 0.61653 0.032392 0.43138 1.9424 1.3069 16.0006 144.9984 0.00019444 22.6721 0.0017727
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4543e-05 0.0011542 0.14878 0.00065826 0.14943 0.13616 0 0.037079 0.0389 0 0.89681 0.24975 0.066995 0.0093574 4.2456 0.058439 7.0186e-05 0.83163 0.0052642 0.0060015 0.99954 0.0082146 0.75162 0.84268 0.97522 0.13178 0.93576 0.92317 0.25814 0.96937 0.61611 0.033722 0.43137 1.9398 1.2529 16.0006 144.9984 0.00019926 22.8207 0.0017966
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4543e-05 0.0011542 0.14878 0.00065826 0.14943 0.13616 0 0.037079 0.0389 0 0.89681 0.24975 0.066995 0.0093575 4.2456 0.058439 7.0186e-05 0.83163 0.0052642 0.0060015 0.99954 0.0074048 0.74845 0.85294 0.97833 0.13178 0.93517 0.92306 0.2641 0.96898 0.61587 0.034514 0.43137 1.9382 1.2233 16.0006 144.9984 0.00020205 22.9065 0.0018107
1.1048 0.98803 5.5188e-05 3.8182 0.012035 1.4543e-05 0.0011542 0.14878 0.00065826 0.14943 0.13616 0 0.037079 0.0389 0 0.89681 0.24975 0.066995 0.0093575 4.2456 0.058439 7.0186e-05 0.83163 0.0052642 0.0060015 0.99955 0.0066746 0.74529 0.8626 0.98106 0.13178 0.93458 0.92295 0.27003 0.96859 0.61562 0.035308 0.43137 1.9365 1.1954 16.0006 144.9984 0.00020478 22.9907 0.0018249
1.1049 0.98803 5.5188e-05 3.8182 0.012035 1.4543e-05 0.0011542 0.14878 0.00065826 0.14944 0.13616 0 0.037078 0.0389 0 0.89681 0.24975 0.066996 0.0093575 4.2456 0.058439 7.0186e-05 0.83163 0.0052642 0.0060015 0.99955 0.0060162 0.74215 0.8717 0.98346 0.13178 0.934 0.92284 0.27593 0.9682 0.61537 0.036104 0.43136 1.9347 1.1691 16.0006 144.9984 0.00020746 23.0736 0.001839
1.1049 0.98803 5.5188e-05 3.8182 0.012035 1.4544e-05 0.0011542 0.14878 0.00065826 0.14944 0.13616 0 0.037078 0.0389 0 0.89681 0.24975 0.066996 0.0093575 4.2456 0.058439 7.0186e-05 0.83163 0.0052642 0.0060015 0.99955 0.0054225 0.73902 0.88026 0.98557 0.13178 0.93341 0.92271 0.2818 0.96781 0.61513 0.036901 0.43136 1.9329 1.1442 16.0006 144.9984 0.00021008 23.1552 0.0018532
1.1049 0.98803 5.5188e-05 3.8182 0.012035 1.4544e-05 0.0011542 0.14878 0.00065826 0.14944 0.13616 0 0.037078 0.0389 0 0.89681 0.24975 0.066996 0.0093575 4.2456 0.058439 7.0187e-05 0.83163 0.0052642 0.0060015 0.99956 0.0048873 0.7359 0.8883 0.98741 0.13178 0.93282 0.92258 0.28764 0.96741 0.61488 0.037701 0.43136 1.9311 1.1207 16.0006 144.9984 0.00021265 23.2355 0.0018673
1.1049 0.98803 5.5188e-05 3.8182 0.012035 1.4544e-05 0.0011542 0.14879 0.00065826 0.14944 0.13616 0 0.037078 0.0389 0 0.89681 0.24976 0.066996 0.0093576 4.2456 0.05844 7.0187e-05 0.83163 0.0052642 0.0060015 0.99956 0.0044047 0.73279 0.89586 0.98903 0.13178 0.93224 0.92245 0.29344 0.96702 0.61463 0.038502 0.43136 1.9292 1.0984 16.0006 144.9984 0.00021518 23.3146 0.0018815
1.1049 0.98803 5.5188e-05 3.8182 0.012035 1.4544e-05 0.0011542 0.14879 0.00065826 0.14944 0.13616 0 0.037078 0.0389 0 0.89681 0.24976 0.066996 0.0093576 4.2456 0.05844 7.0187e-05 0.83163 0.0052642 0.0060015 0.99957 0.0039696 0.7297 0.90295 0.99044 0.13178 0.93165 0.92231 0.29922 0.96663 0.61439 0.039306 0.43135 1.9272 1.0773 16.0006 144.9983 0.00021765 23.3924 0.0018956
1.1049 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14944 0.13617 0 0.037078 0.0389 0 0.89681 0.24976 0.066997 0.0093576 4.2456 0.05844 7.0187e-05 0.83163 0.0052642 0.0060015 0.99957 0.0032238 0.72356 0.91584 0.99276 0.13178 0.93048 0.92202 0.31067 0.96585 0.61389 0.040917 0.43135 1.9232 1.0382 16.0006 144.9983 0.00022247 23.5444 0.0019239
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14944 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99958 0.0026728 0.71807 0.92609 0.99436 0.13178 0.92943 0.92174 0.32086 0.96515 0.61345 0.042374 0.43134 1.9194 1.0063 16.0006 144.9983 0.00022667 23.6768 0.0019494
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0022157 0.71262 0.93518 0.99561 0.13178 0.92838 0.92145 0.33095 0.96445 0.613 0.043836 0.43134 1.9156 0.97704 16.0006 144.9983 0.00023073 23.8046 0.0019748
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021898 0.71228 0.93572 0.99568 0.13178 0.92832 0.92143 0.33157 0.9644 0.61298 0.043927 0.43134 1.9153 0.97529 16.0006 144.9983 0.00023098 23.8124 0.0019764
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021879 0.71226 0.93576 0.99568 0.13178 0.92831 0.92142 0.33162 0.9644 0.61298 0.043934 0.43134 1.9153 0.97516 16.0006 144.9983 0.000231 23.813 0.0019766
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021841 0.71221 0.93584 0.99569 0.13178 0.9283 0.92142 0.33171 0.96439 0.61297 0.043948 0.43134 1.9153 0.9749 16.0006 144.9983 0.00023104 23.8142 0.0019768
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021836 0.7122 0.93585 0.99569 0.13178 0.9283 0.92142 0.33173 0.96439 0.61297 0.043949 0.43134 1.9153 0.97487 16.0006 144.9983 0.00023105 23.8143 0.0019768
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021826 0.71219 0.93587 0.99569 0.13178 0.9283 0.92142 0.33175 0.96439 0.61297 0.043953 0.43134 1.9152 0.9748 16.0006 144.9983 0.00023105 23.8146 0.0019769
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021821 0.71218 0.93588 0.9957 0.13178 0.9283 0.92142 0.33176 0.96439 0.61297 0.043955 0.43134 1.9152 0.97477 16.0006 144.9983 0.00023106 23.8144 0.0019769
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021816 0.71218 0.93589 0.9957 0.13178 0.92829 0.92142 0.33177 0.96439 0.61297 0.043956 0.43134 1.9152 0.97474 16.0006 144.9983 0.00023106 23.8143 0.0019769
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021807 0.71216 0.9359 0.9957 0.13178 0.92829 0.92142 0.3318 0.96439 0.61297 0.04396 0.43134 1.9152 0.97468 16.0006 144.9983 0.00023107 23.814 0.001977
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.002179 0.71214 0.93594 0.9957 0.13178 0.92829 0.92142 0.33184 0.96438 0.61297 0.043966 0.43134 1.9152 0.97455 16.0006 144.9983 0.00023109 23.8134 0.0019771
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021754 0.71209 0.93602 0.99571 0.13178 0.92828 0.92142 0.33193 0.96438 0.61296 0.043979 0.43134 1.9152 0.97431 16.0006 144.9983 0.00023113 23.8123 0.0019773
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021683 0.712 0.93616 0.99573 0.13178 0.92826 0.92141 0.3321 0.96437 0.61295 0.044004 0.43134 1.9151 0.97383 16.0006 144.9983 0.0002312 23.81 0.0019778
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021541 0.71181 0.93646 0.99577 0.13178 0.92822 0.9214 0.33245 0.96434 0.61294 0.044056 0.43134 1.915 0.97286 16.0006 144.9983 0.00023134 23.8055 0.0019787
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021401 0.71162 0.93675 0.99581 0.13178 0.92819 0.92139 0.3328 0.96432 0.61292 0.044107 0.43134 1.9148 0.97189 16.0006 144.9983 0.00023147 23.801 0.0019796
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0021262 0.71143 0.93704 0.99584 0.13178 0.92815 0.92138 0.33315 0.96429 0.61291 0.044158 0.43134 1.9147 0.97093 16.0006 144.9983 0.00023161 23.7964 0.0019805
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0020985 0.71105 0.93762 0.99591 0.13178 0.92808 0.92136 0.33385 0.96424 0.61288 0.04426 0.43134 1.9144 0.96901 16.0006 144.9983 0.00023189 23.7873 0.0019822
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0020711 0.71067 0.93819 0.99598 0.13178 0.928 0.92134 0.33455 0.96419 0.61285 0.044363 0.43134 1.9141 0.9671 16.0006 144.9983 0.00023217 23.7783 0.001984
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0020175 0.70992 0.93931 0.99612 0.13178 0.92786 0.92129 0.33594 0.9641 0.61278 0.044567 0.43133 1.9136 0.96332 16.0006 144.9983 0.00023272 23.7601 0.0019876
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4545e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0019652 0.70916 0.94042 0.99625 0.13178 0.92771 0.92125 0.33733 0.964 0.61272 0.044771 0.43133 1.913 0.95958 16.0006 144.9983 0.00023328 23.7419 0.0019911
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0018647 0.70765 0.94256 0.9965 0.13178 0.92742 0.92116 0.34009 0.9638 0.6126 0.045179 0.43133 1.9119 0.95223 16.0006 144.9982 0.00023437 23.7055 0.0019983
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066998 0.0093577 4.2457 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0017694 0.70614 0.94461 0.99672 0.13178 0.92712 0.92107 0.34284 0.9636 0.61247 0.045586 0.43133 1.9108 0.94504 16.0006 144.9982 0.00023546 23.669 0.0020054
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066998 0.0093578 4.2457 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.0016789 0.70464 0.94658 0.99693 0.13178 0.92683 0.92098 0.34557 0.96341 0.61235 0.045993 0.43133 1.9097 0.93802 16.0006 144.9982 0.00023654 23.6324 0.0020125
1.105 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066998 0.0093578 4.2457 0.058441 7.0188e-05 0.83163 0.0052642 0.0060015 0.99959 0.001593 0.70314 0.94847 0.99713 0.13178 0.92654 0.92089 0.34828 0.96321 0.61223 0.046399 0.43133 1.9085 0.93115 16.0005 144.9982 0.00023761 23.5957 0.0020197
1.1051 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.1488 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066998 0.0093578 4.2457 0.058441 7.0189e-05 0.83163 0.0052642 0.0060015 0.99959 0.0014344 0.70015 0.95203 0.99748 0.13178 0.92595 0.92071 0.35366 0.96282 0.61198 0.047207 0.43132 1.9062 0.91787 16.0005 144.9982 0.00023973 23.5221 0.0020339
1.1051 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.1488 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066998 0.0093578 4.2457 0.058441 7.0189e-05 0.83163 0.0052642 0.0060016 0.99959 0.0012917 0.69718 0.95531 0.99777 0.13178 0.92536 0.92052 0.35897 0.96243 0.61173 0.048013 0.43132 1.9039 0.90516 16.0005 144.9982 0.00024182 23.4481 0.0020482
1.1051 0.98803 5.5188e-05 3.8182 0.012035 1.4546e-05 0.0011542 0.1488 0.00065826 0.14945 0.13618 0 0.037077 0.0389 0 0.89683 0.24976 0.066998 0.0093578 4.2457 0.058441 7.0189e-05 0.83163 0.0052643 0.0060016 0.99958 0.0011632 0.69421 0.95834 0.99802 0.13178 0.92478 0.92032 0.36422 0.96204 0.61148 0.048816 0.43132 1.9016 0.89299 16.0005 144.9982 0.00024388 23.3736 0.0020624
1.1051 0.98803 5.5188e-05 3.8182 0.012035 1.4547e-05 0.0011542 0.1488 0.00065826 0.14945 0.13618 0 0.037077 0.0389 0 0.89683 0.24976 0.066998 0.0093579 4.2457 0.058441 7.0189e-05 0.83163 0.0052643 0.0060016 0.99958 0.0010475 0.69126 0.96113 0.99824 0.13178 0.9242 0.92013 0.36941 0.96164 0.61124 0.049615 0.43132 1.8992 0.88132 16.0005 144.9982 0.0002459 23.2986 0.0020767
1.1051 0.98803 5.5188e-05 3.8182 0.012035 1.4547e-05 0.0011542 0.1488 0.00065826 0.14945 0.13618 0 0.037077 0.0389 0 0.89683 0.24976 0.066999 0.0093579 4.2457 0.058442 7.0189e-05 0.83163 0.0052643 0.0060016 0.99958 0.00094323 0.68832 0.96371 0.99843 0.13178 0.92361 0.91993 0.37453 0.96125 0.61099 0.050412 0.43131 1.8968 0.87013 16.0005 144.9982 0.0002479 23.2231 0.0020909
1.1051 0.98803 5.5188e-05 3.8182 0.012035 1.4547e-05 0.0011542 0.1488 0.00065826 0.14946 0.13618 0 0.037077 0.0389 0 0.89683 0.24976 0.066999 0.0093579 4.2457 0.058442 7.019e-05 0.83163 0.0052643 0.0060016 0.99957 0.00076483 0.68248 0.9683 0.99873 0.13178 0.92244 0.91952 0.3846 0.96047 0.61049 0.051995 0.43131 1.892 0.84908 16.0005 144.9981 0.00025182 23.0703 0.0021195
1.1052 0.98803 5.5188e-05 3.8182 0.012035 1.4547e-05 0.0011542 0.1488 0.00065826 0.14946 0.13618 0 0.037077 0.0389 0 0.89683 0.24976 0.066999 0.009358 4.2457 0.058442 7.019e-05 0.83163 0.0052643 0.0060016 0.99957 0.00063729 0.67744 0.97175 0.99892 0.13178 0.92143 0.91915 0.39317 0.95979 0.61006 0.053364 0.4313 1.8877 0.83208 16.0005 144.9981 0.00025515 22.9351 0.0021443
1.1052 0.98803 5.5188e-05 3.8182 0.012035 1.4548e-05 0.0011542 0.14881 0.00065826 0.14946 0.13618 0 0.037077 0.0389 0 0.89683 0.24977 0.067 0.009358 4.2457 0.058442 7.019e-05 0.83163 0.0052643 0.0060016 0.99956 0.00053111 0.67243 0.97476 0.99907 0.13178 0.92042 0.91878 0.40156 0.95911 0.60963 0.054724 0.4313 1.8834 0.8162 16.0005 144.9981 0.00025841 22.7978 0.0021691
1.1052 0.98803 5.5188e-05 3.8182 0.012035 1.4548e-05 0.0011542 0.14881 0.00065826 0.14946 0.13618 0 0.037077 0.0389 0 0.89684 0.24977 0.067 0.009358 4.2457 0.058442 7.019e-05 0.83163 0.0052643 0.0060016 0.99956 0.0004427 0.66746 0.9774 0.99918 0.13178 0.9194 0.9184 0.40978 0.95843 0.60921 0.056073 0.43129 1.879 0.80134 16.0005 144.998 0.0002616 22.6584 0.0021939
1.1053 0.98803 5.5188e-05 3.8182 0.012035 1.4549e-05 0.0011542 0.14881 0.00065826 0.14946 0.13619 0 0.037077 0.0389 0 0.89684 0.24977 0.067 0.0093581 4.2457 0.058443 7.0191e-05 0.83163 0.0052643 0.0060016 0.99954 0.00030753 0.65763 0.98172 0.99933 0.13178 0.91738 0.91761 0.42569 0.95707 0.60835 0.058743 0.43128 1.8702 0.77437 16.0005 144.998 0.00026778 22.3729 0.0022436
1.1053 0.98803 5.5188e-05 3.8182 0.012035 1.4549e-05 0.0011542 0.14881 0.00065826 0.14947 0.13619 0 0.037076 0.0389 0 0.89684 0.24977 0.067001 0.0093582 4.2457 0.058443 7.0191e-05 0.83163 0.0052643 0.0060016 0.99953 0.00022584 0.64942 0.9846 0.99941 0.13178 0.91568 0.91692 0.43865 0.95592 0.60762 0.060974 0.43127 1.8626 0.75403 16.0004 144.9979 0.00027282 22.1242 0.0022857
1.1054 0.98803 5.5188e-05 3.8182 0.012035 1.455e-05 0.0011542 0.14882 0.00065826 0.14947 0.13619 0 0.037076 0.0389 0 0.89685 0.24977 0.067001 0.0093582 4.2458 0.058444 7.0192e-05 0.83163 0.0052643 0.0060017 0.99952 0.0001658 0.64132 0.98691 0.99946 0.13178 0.91397 0.91621 0.45114 0.95477 0.6069 0.063176 0.43126 1.8549 0.73568 16.0004 144.9979 0.00027771 21.869 0.0023277
1.1054 0.98803 5.5188e-05 3.8182 0.012035 1.455e-05 0.0011542 0.14882 0.00065826 0.14947 0.13619 0 0.037076 0.0389 0 0.89685 0.24977 0.067002 0.0093583 4.2458 0.058444 7.0192e-05 0.83163 0.0052644 0.0060017 0.99951 0.00012563 0.63411 0.9886 0.99948 0.13178 0.91244 0.91555 0.462 0.95374 0.60625 0.065134 0.43126 1.8479 0.72067 16.0004 144.9978 0.00028198 21.6341 0.0023656
1.1054 0.98803 5.5188e-05 3.8182 0.012035 1.4551e-05 0.0011542 0.14882 0.00065826 0.14948 0.1362 0 0.037076 0.0389 0 0.89685 0.24977 0.067002 0.0093583 4.2458 0.058444 7.0193e-05 0.83163 0.0052644 0.0060017 0.99949 9.5223e-05 0.62699 0.99 0.99949 0.13178 0.91092 0.91489 0.47251 0.95271 0.6056 0.067069 0.43125 1.8409 0.70694 16.0004 144.9978 0.00028615 21.3945 0.0024034
1.1055 0.98803 5.5188e-05 3.8182 0.012035 1.4551e-05 0.0011542 0.14882 0.00065826 0.14948 0.1362 0 0.037076 0.0389 0 0.89685 0.24977 0.067003 0.0093584 4.2458 0.058445 7.0193e-05 0.83163 0.0052644 0.0060017 0.99948 7.2216e-05 0.61994 0.99114 0.99949 0.13178 0.90939 0.91421 0.48268 0.95168 0.60495 0.06898 0.43124 1.8339 0.69435 16.0004 144.9977 0.00029021 21.1505 0.0024413
1.1055 0.98803 5.5188e-05 3.8182 0.012035 1.4552e-05 0.0011542 0.14883 0.00065826 0.14948 0.1362 0 0.037076 0.0389 0 0.89686 0.24978 0.067003 0.0093585 4.2458 0.058445 7.0194e-05 0.83163 0.0052644 0.0060017 0.99947 5.212e-05 0.61173 0.99225 0.99948 0.13178 0.9076 0.91339 0.49426 0.95047 0.60419 0.071205 0.43123 1.8255 0.68081 16.0004 144.9977 0.00029487 20.8574 0.0024859
1.1056 0.98803 5.5188e-05 3.8182 0.012035 1.4553e-05 0.0011542 0.14883 0.00065826 0.14948 0.13621 0 0.037075 0.0389 0 0.89686 0.24978 0.067004 0.0093585 4.2458 0.058446 7.0194e-05 0.83162 0.0052644 0.0060017 0.99945 3.7619e-05 0.60363 0.99312 0.99947 0.13178 0.90581 0.91256 0.50539 0.94925 0.60343 0.073399 0.43122 1.8172 0.66855 16.0004 144.9976 0.00029941 20.5591 0.0025306
1.1056 0.98803 5.5188e-05 3.8182 0.012035 1.4553e-05 0.0011542 0.14883 0.00065826 0.14949 0.13621 0 0.037075 0.0389 0 0.89686 0.24978 0.067004 0.0093586 4.2458 0.058446 7.0195e-05 0.83162 0.0052644 0.0060017 0.99943 2.7155e-05 0.59563 0.99382 0.99945 0.13178 0.90403 0.91172 0.51609 0.94804 0.60267 0.075559 0.43121 1.8088 0.65743 16.0003 144.9976 0.00030383 20.2565 0.0025753
1.1056 0.98803 5.5188e-05 3.8182 0.012035 1.4554e-05 0.0011542 0.14884 0.00065826 0.14949 0.13621 0 0.037075 0.0389 0 0.89687 0.24978 0.067005 0.0093587 4.2459 0.058446 7.0195e-05 0.83162 0.0052644 0.0060018 0.99941 1.9607e-05 0.58775 0.99438 0.99943 0.13178 0.90225 0.91086 0.52637 0.94683 0.60191 0.077687 0.4312 1.8003 0.64733 16.0003 144.9975 0.00030814 19.9502 0.00262
1.1057 0.98803 5.5188e-05 3.8182 0.012035 1.4554e-05 0.0011542 0.14884 0.00065826 0.14949 0.13621 0 0.037075 0.0389 0 0.89687 0.24978 0.067006 0.0093587 4.2459 0.058447 7.0196e-05 0.83162 0.0052645 0.0060018 0.99939 1.4167e-05 0.57997 0.99482 0.9994 0.13178 0.90048 0.90999 0.53626 0.94563 0.60115 0.079783 0.4312 1.7919 0.63816 16.0003 144.9974 0.00031235 19.6408 0.0026646
1.1057 0.98803 5.5188e-05 3.8182 0.012035 1.4555e-05 0.0011542 0.14884 0.00065826 0.1495 0.13622 0 0.037075 0.0389 0 0.89687 0.24978 0.067006 0.0093588 4.2459 0.058447 7.0196e-05 0.83162 0.0052645 0.0060018 0.99937 1.0243e-05 0.57229 0.99516 0.99938 0.13178 0.89871 0.90911 0.54576 0.94442 0.6004 0.081846 0.43119 1.7835 0.62983 16.0003 144.9974 0.00031646 19.329 0.0027093
1.1058 0.98803 5.5188e-05 3.8182 0.012035 1.4556e-05 0.0011542 0.14885 0.00065826 0.1495 0.13622 0 0.037074 0.0389 0 0.89688 0.24978 0.067007 0.0093589 4.2459 0.058448 7.0197e-05 0.83162 0.0052645 0.0060018 0.99935 7.4177e-06 0.56472 0.99542 0.99935 0.13178 0.89695 0.90822 0.55489 0.94322 0.59964 0.083878 0.43118 1.7751 0.62226 16.0003 144.9973 0.00032048 19.0154 0.002754
1.1058 0.98803 5.5188e-05 3.8182 0.012035 1.4556e-05 0.0011542 0.14885 0.00065826 0.1495 0.13622 0 0.037074 0.0389 0 0.89688 0.24979 0.067007 0.0093589 4.2459 0.058448 7.0197e-05 0.83162 0.0052645 0.0060018 0.99933 5.3816e-06 0.55724 0.99562 0.99932 0.13178 0.89519 0.90732 0.56367 0.94201 0.59889 0.085878 0.43117 1.7667 0.61538 16.0002 144.9972 0.00032441 18.7007 0.0027987
1.1059 0.98803 5.5188e-05 3.8182 0.012035 1.4557e-05 0.0011542 0.14886 0.00065826 0.14951 0.13623 0 0.037074 0.0389 0 0.89689 0.24979 0.067008 0.0093591 4.2459 0.058449 7.0199e-05 0.83162 0.0052645 0.0060018 0.99929 2.8794e-06 0.5426 0.99586 0.99924 0.13178 0.8917 0.90548 0.5802 0.93961 0.59739 0.089785 0.43115 1.7499 0.60345 16.0002 144.9971 0.00033202 18.0703 0.002888
1.106 0.98803 5.5188e-05 3.8182 0.012035 1.4558e-05 0.0011542 0.14886 0.00065826 0.14951 0.13623 0 0.037073 0.0389 0 0.89689 0.24979 0.067009 0.0093592 4.246 0.05845 7.0199e-05 0.83162 0.0052646 0.0060019 0.99924 1.7015e-06 0.53015 0.99593 0.99918 0.13178 0.88867 0.90384 0.59358 0.93752 0.59609 0.093092 0.43113 1.7353 0.5948 16.0002 144.997 0.00033841 17.5222 0.0029659
1.1061 0.98803 5.5188e-05 3.8182 0.012035 1.4559e-05 0.0011542 0.14887 0.00065826 0.14952 0.13624 0 0.037073 0.0389 0 0.8969 0.24979 0.06701 0.0093593 4.246 0.05845 7.02e-05 0.83162 0.0052646 0.0060019 0.9992 9.6018e-07 0.518 0.99592 0.9991 0.13178 0.88566 0.90218 0.60606 0.93544 0.59479 0.09631 0.43112 1.7209 0.58755 16.0002 144.9969 0.00034459 16.9783 0.0030438
1.1061 0.98803 5.5188e-05 3.8182 0.012035 1.456e-05 0.0011542 0.14887 0.00065826 0.14952 0.13624 0 0.037073 0.0389 0 0.89691 0.2498 0.067011 0.0093594 4.246 0.058451 7.0201e-05 0.83162 0.0052646 0.0060019 0.99915 4.7678e-07 0.50612 0.99584 0.99902 0.13178 0.88267 0.90049 0.6177 0.93336 0.5935 0.09944 0.4311 1.7065 0.58152 16.0001 144.9967 0.00035058 16.4407 0.0031217
1.1062 0.98803 5.5188e-05 3.8182 0.012035 1.4561e-05 0.0011542 0.14888 0.00065826 0.14953 0.13625 0 0.037072 0.0389 0 0.89691 0.2498 0.067012 0.0093595 4.246 0.058452 7.0202e-05 0.83162 0.0052647 0.006002 0.9991 2.482e-07 0.49453 0.99569 0.99893 0.13178 0.8797 0.89877 0.62857 0.93129 0.59222 0.10249 0.43109 1.6923 0.57657 16.0001 144.9966 0.00035639 15.9113 0.0031995
1.1063 0.98803 5.5188e-05 3.8182 0.012035 1.4562e-05 0.0011542 0.14888 0.00065826 0.14954 0.13625 0 0.037072 0.0389 0 0.89692 0.2498 0.067013 0.0093596 4.2461 0.058452 7.0203e-05 0.83162 0.0052647 0.006002 0.99905 2.0022e-07 0.4832 0.99549 0.99884 0.13178 0.87676 0.89704 0.63871 0.92922 0.59094 0.10545 0.43107 1.6782 0.57256 16.0001 144.9965 0.00036203 15.3917 0.0032774
1.1064 0.98803 5.5188e-05 3.8182 0.012035 1.4563e-05 0.0011542 0.14889 0.00065826 0.14954 0.13626 0 0.037072 0.0389 0 0.89692 0.24981 0.067014 0.0093598 4.2461 0.058453 7.0204e-05 0.83162 0.0052647 0.006002 0.999 1.4231e-07 0.47214 0.99525 0.99874 0.13178 0.87383 0.89528 0.64817 0.92715 0.58967 0.10834 0.43105 1.6642 0.56939 16 144.9964 0.00036751 14.8831 0.0033553
1.1065 0.98803 5.5188e-05 3.8182 0.012035 1.4564e-05 0.0011542 0.14889 0.00065826 0.14955 0.13626 0 0.037071 0.0389 0 0.89693 0.24981 0.067015 0.0093599 4.2461 0.058454 7.0205e-05 0.83162 0.0052647 0.006002 0.99894 4.1074e-09 0.46134 0.99498 0.99863 0.13178 0.87093 0.8935 0.657 0.92509 0.58841 0.11115 0.43104 1.6504 0.56696 16 144.9963 0.00037284 14.3866 0.0034332
1.1065 0.98803 5.5188e-05 3.8182 0.012035 1.4565e-05 0.0011542 0.1489 0.00065826 0.14955 0.13627 0 0.037071 0.0389 0 0.89693 0.24981 0.067016 0.00936 4.2461 0.058454 7.0206e-05 0.83162 0.0052648 0.0060021 0.99888 -6.3536e-08 0.45078 0.99467 0.99851 0.13178 0.86805 0.8917 0.66525 0.92303 0.58715 0.1139 0.43102 1.6367 0.56521 16 144.9961 0.00037804 13.9029 0.0035111
1.1066 0.98803 5.5188e-05 3.8182 0.012035 1.4566e-05 0.0011542 0.1489 0.00065826 0.14956 0.13627 0 0.037071 0.0389 0 0.89694 0.24981 0.067017 0.0093601 4.2462 0.058455 7.0207e-05 0.83162 0.0052648 0.0060021 0.99883 3.5708e-08 0.44048 0.99433 0.99839 0.13178 0.86519 0.88988 0.67295 0.92098 0.5859 0.11657 0.43101 1.6232 0.56405 16 144.996 0.0003831 13.4327 0.003589
1.1067 0.98803 5.5188e-05 3.8182 0.012035 1.4568e-05 0.0011542 0.14891 0.00065826 0.14956 0.13628 0 0.03707 0.0389 0 0.89695 0.24982 0.067018 0.0093602 4.2462 0.058456 7.0208e-05 0.83161 0.0052648 0.0060021 0.99877 1.2333e-07 0.43041 0.99396 0.99826 0.13178 0.86235 0.88804 0.68014 0.91894 0.58466 0.11918 0.43099 1.6098 0.56345 15.9999 144.9959 0.00038804 12.9763 0.0036669
1.1068 0.98803 5.5188e-05 3.8182 0.012035 1.4569e-05 0.0011542 0.14891 0.00065826 0.14957 0.13628 0 0.03707 0.0389 0 0.89695 0.24982 0.067019 0.0093603 4.2462 0.058457 7.0209e-05 0.83161 0.0052648 0.0060022 0.99871 7.823e-08 0.42058 0.99356 0.99813 0.13178 0.85954 0.88619 0.68685 0.91689 0.58342 0.12172 0.43097 1.5966 0.56333 15.9999 144.9957 0.00039286 12.5337 0.0037448
1.1068 0.98803 5.5188e-05 3.8182 0.012035 1.457e-05 0.0011542 0.14892 0.00065826 0.14957 0.13629 0 0.03707 0.0389 0 0.89696 0.24982 0.06702 0.0093604 4.2463 0.058457 7.0209e-05 0.83161 0.0052649 0.0060022 0.99864 -2.2228e-09 0.41098 0.99314 0.99799 0.13178 0.85676 0.88432 0.69312 0.91486 0.5822 0.12421 0.43096 1.5836 0.56365 15.9999 144.9956 0.00039756 12.1052 0.0038226
1.1069 0.98803 5.5188e-05 3.8182 0.012035 1.4571e-05 0.0011542 0.14893 0.00065826 0.14958 0.13629 0 0.037069 0.0389 0 0.89696 0.24982 0.067021 0.0093606 4.2463 0.058458 7.021e-05 0.83161 0.0052649 0.0060022 0.99858 5.3607e-09 0.40161 0.9927 0.99784 0.13179 0.85399 0.88243 0.69897 0.91282 0.58098 0.12664 0.43094 1.5708 0.56438 15.9999 144.9955 0.00040215 11.6908 0.0039005
1.107 0.98803 5.5188e-05 3.8182 0.012035 1.4572e-05 0.0011542 0.14893 0.00065826 0.14958 0.1363 0 0.037069 0.0389 0 0.89697 0.24983 0.067021 0.0093607 4.2463 0.058459 7.0211e-05 0.83161 0.0052649 0.0060022 0.99852 7.477e-08 0.39245 0.99223 0.99769 0.13179 0.85125 0.88053 0.70444 0.91079 0.57977 0.12901 0.43093 1.5581 0.56548 15.9998 144.9954 0.00040664 11.2902 0.0039784
1.1071 0.98803 5.5188e-05 3.8182 0.012035 1.4573e-05 0.0011542 0.14894 0.00065826 0.14959 0.1363 0 0.037068 0.0389 0 0.89698 0.24983 0.067022 0.0093608 4.2463 0.058459 7.0212e-05 0.83161 0.005265 0.0060023 0.99845 8.8029e-08 0.3835 0.99175 0.99753 0.13179 0.84854 0.87862 0.70954 0.90877 0.57856 0.13133 0.43091 1.5457 0.56691 15.9998 144.9952 0.00041102 10.9032 0.0040563
1.1072 0.98803 5.5188e-05 3.8182 0.012035 1.4574e-05 0.0011542 0.14894 0.00065826 0.1496 0.13631 0 0.037068 0.0389 0 0.89698 0.24983 0.067023 0.0093609 4.2464 0.05846 7.0213e-05 0.83161 0.005265 0.0060023 0.99839 1.498e-08 0.37477 0.99124 0.99737 0.13179 0.84585 0.8767 0.71431 0.90675 0.57737 0.13361 0.43089 1.5334 0.56865 15.9998 144.9951 0.00041531 10.5295 0.0041342
1.1072 0.98803 5.5188e-05 3.8182 0.012035 1.4575e-05 0.0011542 0.14895 0.00065826 0.1496 0.13631 0 0.037068 0.0389 0 0.89699 0.24983 0.067024 0.009361 4.2464 0.058461 7.0214e-05 0.83161 0.005265 0.0060023 0.99832 -4.8564e-08 0.36623 0.99071 0.9972 0.13179 0.84318 0.87476 0.71875 0.90474 0.57618 0.13583 0.43088 1.5212 0.57067 15.9998 144.995 0.0004195 10.1686 0.0042121
1.1073 0.98803 5.5188e-05 3.8182 0.012035 1.4576e-05 0.0011542 0.14895 0.00065826 0.14961 0.13632 0 0.037067 0.0389 0 0.89699 0.24984 0.067025 0.0093611 4.2464 0.058462 7.0215e-05 0.83161 0.005265 0.0060023 0.99826 -5.9055e-08 0.3579 0.99017 0.99702 0.13179 0.84054 0.87281 0.7229 0.90273 0.57501 0.13801 0.43086 1.5093 0.57295 15.9997 144.9949 0.00042361 9.8204 0.00429
1.1074 0.98803 5.5188e-05 3.8182 0.012035 1.4577e-05 0.0011542 0.14896 0.00065826 0.14961 0.13632 0 0.037067 0.0389 0 0.897 0.24984 0.067026 0.0093613 4.2464 0.058462 7.0216e-05 0.83161 0.0052651 0.0060024 0.99819 -4.2228e-08 0.34976 0.9896 0.99684 0.13179 0.83792 0.87085 0.72677 0.90072 0.57383 0.14015 0.43085 1.4976 0.57546 15.9997 144.9947 0.00042762 9.4842 0.0043679
1.1075 0.98803 5.5188e-05 3.8182 0.012035 1.4578e-05 0.0011542 0.14896 0.00065826 0.14962 0.13633 0 0.037067 0.0389 0 0.89701 0.24984 0.067027 0.0093614 4.2465 0.058463 7.0217e-05 0.83161 0.0052651 0.0060024 0.99813 -2.3138e-08 0.34181 0.98902 0.99666 0.13179 0.83532 0.86888 0.73038 0.89872 0.57267 0.14225 0.43083 1.486 0.5782 15.9997 144.9946 0.00043154 9.1596 0.0044458
1.1075 0.98803 5.5188e-05 3.8182 0.012035 1.4579e-05 0.0011542 0.14897 0.00065826 0.14962 0.13634 0 0.037066 0.0389 0 0.89701 0.24984 0.067028 0.0093615 4.2465 0.058464 7.0218e-05 0.83161 0.0052651 0.0060024 0.99806 -1.1031e-08 0.33404 0.98843 0.99647 0.13179 0.83274 0.8669 0.73375 0.89672 0.57152 0.1443 0.43081 1.4746 0.58113 15.9997 144.9945 0.00043538 8.8462 0.0045236
1.1076 0.98803 5.5187e-05 3.8182 0.012035 1.458e-05 0.0011542 0.14897 0.00065826 0.14963 0.13634 0 0.037066 0.0389 0 0.89702 0.24985 0.067029 0.0093616 4.2465 0.058464 7.0219e-05 0.83161 0.0052651 0.0060025 0.99799 -5.3552e-09 0.32645 0.98781 0.99628 0.13179 0.83019 0.86492 0.73688 0.89473 0.57037 0.14632 0.4308 1.4635 0.58425 15.9996 144.9943 0.00043914 8.5435 0.0046015
1.1077 0.98803 5.5187e-05 3.8182 0.012035 1.4581e-05 0.0011542 0.14898 0.00065826 0.14963 0.13635 0 0.037066 0.0389 0 0.89702 0.24985 0.06703 0.0093617 4.2465 0.058465 7.022e-05 0.83161 0.0052652 0.0060025 0.99793 -3.3216e-09 0.31904 0.98719 0.99608 0.13179 0.82766 0.86292 0.73979 0.89274 0.56924 0.1483 0.43078 1.4524 0.58754 15.9996 144.9942 0.00044282 8.251 0.0046794
1.1078 0.98803 5.5187e-05 3.8182 0.012035 1.4582e-05 0.0011542 0.14898 0.00065826 0.14964 0.13635 0 0.037065 0.0389 0 0.89703 0.24985 0.067031 0.0093618 4.2466 0.058466 7.022e-05 0.8316 0.0052652 0.0060025 0.99786 -2.4498e-09 0.3118 0.98655 0.99588 0.13179 0.82515 0.86092 0.7425 0.89076 0.56811 0.15025 0.43077 1.4416 0.59099 15.9996 144.9941 0.00044642 7.9681 0.0047573
1.1079 0.98803 5.5187e-05 3.8182 0.012035 1.4584e-05 0.0011542 0.149 0.00065826 0.14965 0.13636 0 0.037065 0.0389 0 0.89704 0.24986 0.067033 0.0093621 4.2466 0.058467 7.0222e-05 0.8316 0.0052653 0.0060026 0.99773 -1.5375e-09 0.29783 0.98522 0.99546 0.13179 0.8202 0.85689 0.74736 0.8868 0.56588 0.15405 0.43073 1.4206 0.5983 15.9995 144.9938 0.0004534 7.4296 0.0049131
1.1081 0.98803 5.5187e-05 3.8182 0.012035 1.4586e-05 0.0011542 0.14901 0.00065826 0.14966 0.13637 0 0.037064 0.0389 0 0.89705 0.24986 0.067035 0.0093623 4.2467 0.058469 7.0224e-05 0.8316 0.0052653 0.0060026 0.99761 -3.9402e-10 0.28579 0.98398 0.99507 0.13179 0.81582 0.85325 0.75113 0.88326 0.56389 0.15736 0.43071 1.4022 0.6053 15.9995 144.9936 0.00045943 6.9734 0.0050533
1.1082 0.98803 5.5187e-05 3.8182 0.012035 1.4588e-05 0.0011542 0.14902 0.00065826 0.14967 0.13638 0 0.037063 0.0389 0 0.89706 0.24987 0.067036 0.0093625 4.2467 0.05847 7.0226e-05 0.8316 0.0052654 0.0060027 0.9975 3.4705e-10 0.27426 0.98271 0.99467 0.13179 0.8115 0.8496 0.75441 0.87973 0.56194 0.16058 0.43068 1.3845 0.61264 15.9994 144.9934 0.00046523 6.5417 0.0051935
1.1084 0.98803 5.5187e-05 3.8182 0.012035 1.4589e-05 0.0011542 0.14902 0.00065826 0.14968 0.13639 0 0.037063 0.0389 0 0.89707 0.24987 0.067038 0.0093627 4.2468 0.058471 7.0227e-05 0.8316 0.0052654 0.0060027 0.99738 4.0512e-10 0.26319 0.9814 0.99426 0.13179 0.80725 0.84593 0.75723 0.87622 0.56001 0.16371 0.43065 1.3673 0.62027 15.9994 144.9932 0.00047082 6.1319 0.0053337
1.1085 0.98803 5.5187e-05 3.8182 0.012035 1.4591e-05 0.0011542 0.14903 0.00065826 0.14969 0.1364 0 0.037062 0.0389 0 0.89708 0.24988 0.06704 0.0093629 4.2468 0.058472 7.0229e-05 0.8316 0.0052655 0.0060028 0.99726 1.5069e-10 0.25259 0.98005 0.99385 0.13179 0.80306 0.84225 0.75964 0.87272 0.5581 0.16675 0.43062 1.3507 0.62814 15.9994 144.9929 0.00047619 5.7421 0.0054739
1.1086 0.98803 5.5187e-05 3.8182 0.012035 1.4593e-05 0.0011542 0.14904 0.00065826 0.1497 0.13641 0 0.037061 0.0389 0 0.89709 0.24988 0.067041 0.0093631 4.2468 0.058474 7.023e-05 0.8316 0.0052655 0.0060028 0.99715 -2.2673e-11 0.24242 0.97868 0.99342 0.13179 0.79893 0.83856 0.76167 0.86923 0.55622 0.16972 0.43059 1.3346 0.63621 15.9993 144.9927 0.00048136 5.3701 0.0056141
1.1088 0.98803 5.5187e-05 3.8182 0.012035 1.4595e-05 0.0011542 0.14905 0.00065826 0.14971 0.13642 0 0.037061 0.0389 0 0.8971 0.24989 0.067043 0.0093633 4.2469 0.058475 7.0232e-05 0.8316 0.0052655 0.0060029 0.99703 -3.2497e-11 0.23266 0.97727 0.99298 0.13179 0.79486 0.83487 0.76336 0.86576 0.55437 0.17262 0.43056 1.3192 0.64445 15.9993 144.9925 0.00048633 5.0142 0.0057543
1.1089 0.98803 5.5187e-05 3.8182 0.012035 1.4597e-05 0.0011542 0.14906 0.00065826 0.14972 0.13642 0 0.03706 0.0389 0 0.89712 0.24989 0.067045 0.0093635 4.2469 0.058476 7.0234e-05 0.83159 0.0052656 0.0060029 0.99692 4.9388e-12 0.22331 0.97583 0.99254 0.13179 0.79085 0.83118 0.76473 0.8623 0.55254 0.17545 0.43053 1.3042 0.65282 15.9992 144.9923 0.00049111 4.6726 0.0058945
1.1091 0.98803 5.5187e-05 3.8182 0.012035 1.4599e-05 0.0011542 0.14907 0.00065826 0.14973 0.13643 0 0.03706 0.0389 0 0.89713 0.2499 0.067046 0.0093637 4.247 0.058477 7.0235e-05 0.83159 0.0052656 0.006003 0.99681 3.6243e-12 0.21434 0.97436 0.99208 0.13179 0.78689 0.82749 0.76582 0.85886 0.55073 0.17821 0.4305 1.2898 0.66129 15.9992 144.9921 0.00049571 4.3441 0.0060347
1.1092 0.98803 5.5187e-05 3.8182 0.012035 1.46e-05 0.0011542 0.14908 0.00065826 0.14974 0.13644 0 0.037059 0.0389 0 0.89714 0.2499 0.067048 0.009364 4.247 0.058479 7.0237e-05 0.83159 0.0052657 0.006003 0.99669 -2.0807e-11 0.20574 0.97287 0.99162 0.13179 0.78299 0.8238 0.76665 0.85543 0.54895 0.18091 0.43048 1.276 0.66983 15.9991 144.9918 0.00050014 4.0271 0.0061749
1.1093 0.98803 5.5187e-05 3.8182 0.012035 1.4602e-05 0.0011542 0.14909 0.00065826 0.14975 0.13645 0 0.037058 0.0389 0 0.89715 0.2499 0.06705 0.0093642 4.2471 0.05848 7.0239e-05 0.83159 0.0052657 0.0060031 0.99658 -2.4597e-11 0.19749 0.97134 0.99114 0.13179 0.77914 0.82011 0.76723 0.85201 0.54719 0.18355 0.43045 1.2626 0.67842 15.9991 144.9916 0.00050439 3.7204 0.0063151
1.1095 0.98803 5.5187e-05 3.8182 0.012035 1.4604e-05 0.0011542 0.1491 0.00065826 0.14976 0.13646 0 0.037058 0.0389 0 0.89716 0.24991 0.067052 0.0093644 4.2471 0.058481 7.024e-05 0.83159 0.0052658 0.0060031 0.99646 -6.206e-12 0.18958 0.96979 0.99066 0.13179 0.77535 0.81643 0.76759 0.84861 0.54545 0.18613 0.43042 1.2498 0.68704 15.9991 144.9914 0.00050848 3.4231 0.0064553
1.1096 0.98803 5.5187e-05 3.8182 0.012035 1.4606e-05 0.0011542 0.14911 0.00065826 0.14977 0.13647 0 0.037057 0.0389 0 0.89717 0.24991 0.067053 0.0093646 4.2472 0.058483 7.0242e-05 0.83159 0.0052658 0.0060032 0.99635 7.2136e-12 0.18199 0.96821 0.99017 0.13179 0.77161 0.81276 0.76774 0.84522 0.54374 0.18865 0.43039 1.2374 0.69566 15.999 144.9912 0.0005124 3.1341 0.0065954
1.1098 0.98803 5.5187e-05 3.8182 0.012035 1.4608e-05 0.0011542 0.14912 0.00065826 0.14978 0.13648 0 0.037056 0.0389 0 0.89718 0.24992 0.067055 0.0093648 4.2472 0.058484 7.0244e-05 0.83159 0.0052659 0.0060032 0.99623 4.1609e-12 0.17471 0.9666 0.98967 0.13179 0.76791 0.8091 0.7677 0.84184 0.54205 0.19112 0.43036 1.2256 0.70426 15.999 144.991 0.00051618 2.8525 0.0067356
1.1099 0.98803 5.5187e-05 3.8182 0.012035 1.461e-05 0.0011542 0.14913 0.00065826 0.14979 0.13649 0 0.037056 0.0389 0 0.89719 0.24992 0.067057 0.009365 4.2473 0.058485 7.0245e-05 0.83159 0.0052659 0.0060033 0.99612 -3.3821e-12 0.16772 0.96497 0.98916 0.13179 0.76427 0.80545 0.76748 0.83848 0.54038 0.19354 0.43033 1.2142 0.71282 15.9989 144.9908 0.0005198 2.5775 0.0068758
1.1102 0.98803 5.5187e-05 3.8182 0.012035 1.4613e-05 0.0011542 0.14915 0.00065826 0.14981 0.13651 0 0.037055 0.0389 0 0.89721 0.24993 0.06706 0.0093654 4.2474 0.058488 7.0249e-05 0.83158 0.005266 0.0060034 0.99588 -2.0416e-11 0.1546 0.9616 0.9881 0.13179 0.75713 0.79819 0.76656 0.8318 0.53711 0.19823 0.43027 1.1927 0.72978 15.9989 144.9904 0.00052663 2.0446 0.0071562
1.1104 0.98803 5.5187e-05 3.8182 0.012035 1.4617e-05 0.0011542 0.14917 0.00065827 0.14982 0.13652 0 0.037053 0.0389 0 0.89723 0.24994 0.067063 0.0093658 4.2474 0.05849 7.0252e-05 0.83158 0.0052661 0.0060035 0.99566 -1.1911e-11 0.14368 0.95847 0.98712 0.1318 0.75086 0.79171 0.76523 0.82583 0.53424 0.2023 0.43022 1.1749 0.74476 15.9988 144.99 0.00053232 1.5811 0.0074086
1.1107 0.98803 5.5187e-05 3.8182 0.012035 1.462e-05 0.0011542 0.14919 0.00065827 0.14984 0.13654 0 0.037052 0.0389 0 0.89725 0.24995 0.067066 0.0093662 4.2475 0.058492 7.0254e-05 0.83158 0.0052662 0.0060035 0.99544 5.2587e-12 0.13356 0.95523 0.98609 0.1318 0.74474 0.78529 0.76348 0.8199 0.53144 0.20621 0.43017 1.1585 0.75939 15.9987 144.9896 0.0005376 1.1296 0.007661
1.1109 0.98803 5.5187e-05 3.8182 0.012035 1.4623e-05 0.0011542 0.1492 0.00065827 0.14986 0.13655 0 0.037051 0.0389 0 0.89727 0.24996 0.067069 0.0093665 4.2476 0.058495 7.0257e-05 0.83158 0.0052663 0.0060036 0.99521 -4.714e-12 0.12415 0.95188 0.98502 0.1318 0.73877 0.77893 0.76137 0.81402 0.52871 0.20999 0.43012 1.1433 0.77362 15.9986 144.9893 0.00054252 0.68757 0.0079133
1.1112 0.98803 5.5187e-05 3.8182 0.012035 1.4627e-05 0.0011542 0.14922 0.00065827 0.14987 0.13657 0 0.03705 0.0389 0 0.89729 0.24997 0.067072 0.0093669 4.2477 0.058497 7.026e-05 0.83157 0.0052664 0.0060037 0.99498 -1.842e-11 0.11543 0.94841 0.9839 0.1318 0.73293 0.77265 0.75891 0.80818 0.52604 0.21363 0.43007 1.1293 0.78738 15.9986 144.9889 0.00054709 0.2527 0.0081657
1.1114 0.98803 5.5187e-05 3.8182 0.012035 1.463e-05 0.0011542 0.14924 0.00065827 0.14989 0.13659 0 0.037049 0.0389 0 0.89731 0.24998 0.067075 0.0093673 4.2478 0.058499 7.0263e-05 0.83157 0.0052665 0.0060038 0.99473 5.7074e-12 0.10733 0.9448 0.98272 0.1318 0.72724 0.76645 0.75614 0.80239 0.52345 0.21715 0.43002 1.1164 0.80065 15.9985 144.9886 0.00055133 -0.17698 0.008418
1.1117 0.98803 5.5187e-05 3.8182 0.012035 1.4633e-05 0.0011542 0.14926 0.00065827 0.14991 0.1366 0 0.037048 0.0389 0 0.89733 0.24998 0.067078 0.0093677 4.2479 0.058502 7.0266e-05 0.83157 0.0052666 0.0060039 0.99448 2.712e-11 0.099811 0.94105 0.98149 0.1318 0.72168 0.76034 0.7531 0.79663 0.52092 0.22054 0.42996 1.1046 0.81339 15.9984 144.9883 0.00055528 -0.60327 0.0086704
1.1119 0.98803 5.5187e-05 3.8182 0.012035 1.4637e-05 0.0011542 0.14927 0.00065827 0.14993 0.13662 0 0.037047 0.0389 0 0.89735 0.24999 0.067082 0.009368 4.2479 0.058504 7.0269e-05 0.83157 0.0052667 0.006004 0.99421 1.1238e-11 0.09283 0.93715 0.98019 0.1318 0.71625 0.75431 0.74979 0.79092 0.51846 0.22381 0.42991 1.0938 0.82557 15.9984 144.9879 0.00055895 -1.0278 0.0089227
1.1122 0.98803 5.5187e-05 3.8182 0.012035 1.464e-05 0.0011542 0.14929 0.00065827 0.14994 0.13664 0 0.037046 0.0389 0 0.89736 0.25 0.067085 0.0093684 4.248 0.058506 7.0272e-05 0.83156 0.0052668 0.0060041 0.99393 -6.8208e-12 0.08635 0.93309 0.97882 0.1318 0.71096 0.74838 0.74625 0.78525 0.51607 0.22696 0.42986 1.0839 0.83717 15.9983 144.9876 0.00056236 -1.452 0.0091751
1.1125 0.98803 5.5187e-05 3.8182 0.012035 1.4643e-05 0.0011542 0.14931 0.00065827 0.14996 0.13665 0 0.037044 0.0389 0 0.89738 0.25001 0.067088 0.0093688 4.2481 0.058508 7.0275e-05 0.83156 0.0052668 0.0060042 0.99364 1.6717e-11 0.080333 0.92884 0.97738 0.1318 0.70579 0.74256 0.74247 0.77962 0.51374 0.23 0.42981 1.0749 0.8482 15.9982 144.9873 0.00056554 -1.8774 0.0094274
1.1127 0.98803 5.5187e-05 3.8182 0.012035 1.4647e-05 0.0011542 0.14933 0.00065827 0.14998 0.13667 0 0.037043 0.0389 0 0.8974 0.25002 0.067091 0.0093692 4.2482 0.058511 7.0278e-05 0.83156 0.0052669 0.0060043 0.99333 3.9469e-11 0.074746 0.9244 0.97585 0.1318 0.70076 0.73684 0.73848 0.77404 0.51148 0.23293 0.42976 1.0667 0.85864 15.9982 144.987 0.0005685 -2.3053 0.0096798
1.113 0.98803 5.5187e-05 3.8182 0.012035 1.465e-05 0.0011542 0.14934 0.00065827 0.15 0.13669 0 0.037042 0.0389 0 0.89742 0.25003 0.067094 0.0093696 4.2483 0.058513 7.0281e-05 0.83156 0.005267 0.0060043 0.99301 -3.6511e-12 0.069558 0.91976 0.97423 0.1318 0.69585 0.73122 0.73429 0.76849 0.50929 0.23574 0.42971 1.0592 0.86849 15.9981 144.9866 0.00057126 -2.737 0.0099322
1.1133 0.98803 5.5187e-05 3.8182 0.012035 1.4654e-05 0.0011542 0.14936 0.00065827 0.15002 0.1367 0 0.037041 0.0389 0 0.89744 0.25004 0.067097 0.00937 4.2484 0.058516 7.0285e-05 0.83155 0.0052671 0.0060045 0.9926 -3.3402e-11 0.063958 0.91403 0.9722 0.1318 0.69027 0.7248 0.72914 0.76205 0.50681 0.2389 0.42965 1.0514 0.8793 15.998 144.9863 0.00057426 -3.2486 0.010227
1.1135 0.98803 5.5187e-05 3.8182 0.012035 1.4658e-05 0.0011542 0.14938 0.00065827 0.15004 0.13672 0 0.03704 0.0389 0 0.89747 0.25005 0.067101 0.0093704 4.2485 0.058518 7.0288e-05 0.83155 0.0052672 0.0060046 0.99216 -1.5154e-11 0.058823 0.90796 0.97002 0.1318 0.68486 0.71855 0.72372 0.75567 0.50442 0.24191 0.42959 1.0444 0.88933 15.9979 144.9859 0.00057702 -3.7694 0.010522
1.1138 0.98803 5.5187e-05 3.8182 0.012035 1.4661e-05 0.0011542 0.1494 0.00065827 0.15006 0.13674 0 0.037038 0.0389 0 0.89749 0.25006 0.067105 0.0093709 4.2486 0.058521 7.0292e-05 0.83155 0.0052673 0.0060047 0.99168 6.1514e-12 0.054113 0.90152 0.96765 0.13181 0.67963 0.71246 0.71805 0.74935 0.50212 0.24477 0.42953 1.0382 0.89863 15.9979 144.9856 0.00057958 -4.3017 0.010818
1.1141 0.98803 5.5187e-05 3.8182 0.012035 1.4665e-05 0.0011542 0.14943 0.00065827 0.15008 0.13676 0 0.037037 0.0389 0 0.89751 0.25007 0.067108 0.0093713 4.2487 0.058524 7.0295e-05 0.83155 0.0052674 0.0060048 0.99116 7.4626e-12 0.049793 0.89466 0.9651 0.13181 0.67456 0.70654 0.71213 0.74308 0.49992 0.2475 0.42946 1.0328 0.90723 15.9978 144.9853 0.00058193 -4.8476 0.011113
1.1144 0.98803 5.5187e-05 3.8182 0.012035 1.4669e-05 0.0011542 0.14945 0.00065827 0.1501 0.13678 0 0.037036 0.0389 0 0.89753 0.25008 0.067112 0.0093718 4.2488 0.058527 7.0299e-05 0.83154 0.0052675 0.0060049 0.99059 -1.4676e-13 0.045832 0.88734 0.96231 0.13181 0.66967 0.70081 0.70596 0.73686 0.49781 0.25008 0.4294 1.028 0.91515 15.9977 144.9849 0.00058412 -5.4097 0.011408
1.1147 0.98803 5.5187e-05 3.8182 0.012035 1.4673e-05 0.0011542 0.14947 0.00065827 0.15012 0.1368 0 0.037034 0.0389 0 0.89756 0.25009 0.067115 0.0093722 4.2489 0.058529 7.0302e-05 0.83154 0.0052676 0.006005 0.98997 -3.122e-12 0.042199 0.87951 0.95928 0.13181 0.66495 0.69526 0.69954 0.7307 0.4958 0.25252 0.42934 1.0237 0.92243 15.9976 144.9846 0.00058613 -5.9907 0.011703
1.115 0.98803 5.5187e-05 3.8182 0.012035 1.4677e-05 0.0011542 0.14949 0.00065827 0.15014 0.13682 0 0.037033 0.0389 0 0.89758 0.2501 0.067119 0.0093726 4.249 0.058532 7.0305e-05 0.83154 0.0052678 0.0060051 0.98927 -1.989e-13 0.038866 0.87112 0.95596 0.13181 0.6604 0.6899 0.69286 0.72459 0.49389 0.25482 0.42928 1.0201 0.92912 15.9976 144.9843 0.000588 -6.5934 0.011998
1.1153 0.98803 5.5187e-05 3.8182 0.012035 1.4681e-05 0.0011542 0.14951 0.00065827 0.15016 0.13684 0 0.037032 0.0389 0 0.8976 0.25011 0.067123 0.0093731 4.2491 0.058535 7.0309e-05 0.83154 0.0052679 0.0060052 0.9885 1.5156e-12 0.035811 0.86211 0.95232 0.13181 0.65603 0.68474 0.68591 0.71854 0.49207 0.25698 0.42922 1.0169 0.93525 15.9975 144.984 0.00058973 -7.2209 0.012293
1.1156 0.98803 5.5187e-05 3.8182 0.012035 1.4685e-05 0.0011542 0.14953 0.00065827 0.15018 0.13686 0 0.03703 0.0389 0 0.89762 0.25012 0.067126 0.0093735 4.2492 0.058537 7.0312e-05 0.83153 0.005268 0.0060053 0.98763 -2.123e-13 0.033008 0.85239 0.9483 0.13181 0.65183 0.67979 0.6787 0.71254 0.49035 0.25901 0.42916 1.0141 0.94086 15.9974 144.9837 0.00059133 -7.8766 0.012589
1.1159 0.98803 5.5187e-05 3.8182 0.012035 1.4689e-05 0.0011542 0.14955 0.00065827 0.1502 0.13688 0 0.037029 0.0389 0 0.89765 0.25013 0.06713 0.009374 4.2493 0.05854 7.0316e-05 0.83153 0.0052681 0.0060054 0.98664 -1.2117e-12 0.030439 0.84191 0.94387 0.13181 0.64781 0.67505 0.67121 0.7066 0.48872 0.26089 0.4291 1.0117 0.946 15.9974 144.9834 0.0005928 -8.5645 0.012884
1.1165 0.98803 5.5187e-05 3.8182 0.012035 1.4696e-05 0.0011542 0.14959 0.00065827 0.15024 0.13691 0 0.037026 0.0389 0 0.89769 0.25015 0.067137 0.0093748 4.2495 0.058546 7.0323e-05 0.83152 0.0052683 0.0060056 0.98424 -3.6345e-12 0.025926 0.81823 0.93348 0.13181 0.64031 0.66622 0.65535 0.69487 0.48578 0.26423 0.42898 1.008 0.95499 15.9972 144.9829 0.00059539 -10.0534 0.013474
1.117 0.98803 5.5187e-05 3.8182 0.012035 1.4703e-05 0.0011542 0.14962 0.00065827 0.15028 0.13695 0 0.037024 0.0389 0 0.89773 0.25016 0.067143 0.0093756 4.2496 0.05855 7.0329e-05 0.83152 0.0052685 0.0060058 0.98145 -1.6262e-12 0.022553 0.79379 0.92221 0.13181 0.63432 0.65922 0.64034 0.68471 0.48352 0.26671 0.42888 1.0056 0.96167 15.9971 144.9824 0.00059732 -11.5167 0.013994
1.1174 0.98803 5.5187e-05 3.8182 0.012035 1.4709e-05 0.0011542 0.14965 0.00065827 0.15031 0.13697 0 0.037022 0.0389 0 0.89776 0.25018 0.067148 0.0093762 4.2498 0.058554 7.0334e-05 0.83152 0.0052686 0.0060059 0.97862 2.589e-12 0.020235 0.77159 0.91152 0.13182 0.62999 0.65421 0.62776 0.67681 0.48195 0.26835 0.42879 1.0043 0.96627 15.997 144.9821 0.00059861 -12.7948 0.014405
1.1178 0.98803 5.5187e-05 3.8182 0.012035 1.4714e-05 0.0011542 0.14968 0.00065827 0.15033 0.137 0 0.03702 0.0389 0 0.89779 0.25019 0.067153 0.0093768 4.2499 0.058558 7.0339e-05 0.83151 0.0052688 0.0060061 0.975 2.8116e-12 0.018188 0.74637 0.89886 0.13182 0.62603 0.64969 0.6145 0.66902 0.48058 0.26971 0.42871 1.0033 0.97033 15.9969 144.9818 0.00059969 -14.1986 0.014817
1.1183 0.98803 5.5187e-05 3.8182 0.012035 1.4719e-05 0.0011542 0.14971 0.00065828 0.15036 0.13703 0 0.037019 0.0389 0 0.89782 0.25021 0.067158 0.0093775 4.2501 0.058562 7.0343e-05 0.83151 0.0052689 0.0060062 0.9703 -1.6179e-12 0.016386 0.7176 0.88377 0.13182 0.62245 0.64568 0.60056 0.66135 0.4794 0.2708 0.42863 1.0026 0.97395 15.9969 144.9815 0.00060058 -15.7459 0.015228
1.1186 0.98803 5.5187e-05 3.8182 0.012035 1.4724e-05 0.0011542 0.14973 0.00065828 0.15039 0.13705 0 0.037017 0.0389 0 0.89785 0.25022 0.067163 0.009378 4.2502 0.058565 7.0348e-05 0.83151 0.005269 0.0060064 0.96479 -3.1542e-12 0.014952 0.68821 0.86764 0.13182 0.61954 0.6425 0.58741 0.65455 0.47849 0.27154 0.42855 1.0022 0.97689 15.9968 144.9812 0.00060119 -17.2758 0.015598
1.1189 0.98803 5.5187e-05 3.8182 0.012035 1.4728e-05 0.0011542 0.14975 0.00065828 0.15041 0.13707 0 0.037016 0.0389 0 0.89788 0.25023 0.067166 0.0093784 4.2503 0.058568 7.0351e-05 0.8315 0.0052691 0.0060065 0.95931 -1.1237e-12 0.013939 0.66246 0.85295 0.13182 0.61747 0.6403 0.57669 0.64928 0.47787 0.27197 0.42849 1.0021 0.97903 15.9967 144.981 0.00060155 -18.5773 0.015889
1.1192 0.98803 5.5187e-05 3.8182 0.012035 1.4732e-05 0.0011542 0.14977 0.00065828 0.15043 0.13709 0 0.037014 0.0389 0 0.8979 0.25024 0.06717 0.0093789 4.2504 0.05857 7.0355e-05 0.8315 0.0052692 0.0060066 0.9525 6.6139e-13 0.013021 0.63413 0.83619 0.13182 0.61557 0.63835 0.56563 0.6441 0.47733 0.27228 0.42843 1.002 0.98106 15.9967 144.9808 0.0006018 -19.9699 0.01618
1.1195 0.98803 5.5187e-05 3.8182 0.012035 1.4736e-05 0.0011542 0.14979 0.00065828 0.15045 0.13711 0 0.037013 0.0389 0 0.89792 0.25025 0.067174 0.0093793 4.2505 0.058573 7.0358e-05 0.8315 0.0052693 0.0060067 0.94399 2.2451e-13 0.01219 0.60302 0.81704 0.13182 0.61385 0.63665 0.55423 0.63899 0.47687 0.27246 0.42837 1.0021 0.98299 15.9966 144.9807 0.00060193 -21.455 0.016471
1.1198 0.98803 5.5187e-05 3.8182 0.012035 1.474e-05 0.0011542 0.14981 0.00065828 0.15047 0.13713 0 0.037012 0.0389 0 0.89794 0.25026 0.067177 0.0093798 4.2506 0.058576 7.0362e-05 0.83149 0.0052694 0.0060068 0.93333 -8.0189e-13 0.011441 0.56895 0.79517 0.13182 0.61229 0.63519 0.54251 0.63399 0.47648 0.27252 0.42831 1.0022 0.98484 15.9966 144.9805 0.00060195 -23.0307 0.016761
1.1201 0.98803 5.5187e-05 3.8182 0.012035 1.4743e-05 0.0011542 0.14983 0.00065828 0.15049 0.13714 0 0.03701 0.0389 0 0.89796 0.25027 0.067181 0.0093802 4.2507 0.058578 7.0365e-05 0.83149 0.0052695 0.0060069 0.91994 -2.7227e-13 0.01077 0.53181 0.77026 0.13182 0.61088 0.63395 0.53045 0.6291 0.47615 0.27247 0.42825 1.0024 0.98657 15.9965 144.9803 0.00060186 -24.6905 0.017052
1.1204 0.98803 5.5187e-05 3.8182 0.012035 1.4747e-05 0.0011542 0.14985 0.00065828 0.15051 0.13716 0 0.037009 0.0389 0 0.89799 0.25028 0.067184 0.0093806 4.2508 0.058581 7.0368e-05 0.83149 0.0052697 0.006007 0.90319 9.1361e-13 0.010171 0.49164 0.74196 0.13182 0.60961 0.63292 0.51805 0.62434 0.47587 0.27232 0.4282 1.0027 0.98818 15.9965 144.9802 0.00060169 -26.4229 0.017343
1.1207 0.98803 5.5187e-05 3.8182 0.012035 1.4751e-05 0.0011542 0.14987 0.00065828 0.15053 0.13718 0 0.037008 0.0389 0 0.89801 0.25029 0.067188 0.0093811 4.2509 0.058584 7.0372e-05 0.83149 0.0052698 0.0060071 0.88242 4.7279e-13 0.0096394 0.44861 0.71 0.13183 0.60846 0.63207 0.50528 0.61976 0.47565 0.27206 0.42814 1.003 0.98967 15.9964 144.9801 0.00060145 -28.2104 0.017634
1.1209 0.98803 5.5187e-05 3.8182 0.012035 1.4754e-05 0.0011542 0.14989 0.00065828 0.15055 0.1372 0 0.037007 0.0389 0 0.89803 0.2503 0.067191 0.0093814 4.251 0.058586 7.0375e-05 0.83148 0.0052698 0.0060072 0.85976 -6.7425e-13 0.0092147 0.4078 0.67795 0.13183 0.60753 0.63145 0.49341 0.6158 0.47548 0.27175 0.42808 1.0034 0.99091 15.9964 144.9799 0.00060117 -29.8476 0.017896
1.1212 0.98803 5.5187e-05 3.8182 0.012035 1.4758e-05 0.0011542 0.14991 0.00065828 0.15056 0.13721 0 0.037006 0.0389 0 0.89805 0.2503 0.067194 0.0093818 4.251 0.058588 7.0378e-05 0.83148 0.0052699 0.0060073 0.83588 -8.8022e-13 0.0088727 0.36981 0.64642 0.13183 0.60676 0.63097 0.4824 0.61241 0.47535 0.27141 0.42804 1.0037 0.99197 15.9964 144.9798 0.00060087 -31.3277 0.018131
1.1214 0.98803 5.5187e-05 3.8182 0.012035 1.4761e-05 0.0011542 0.14992 0.00065828 0.15058 0.13723 0 0.037005 0.0389 0 0.89806 0.25031 0.067197 0.0093822 4.2511 0.05859 7.038e-05 0.83148 0.00527 0.0060074 0.8086 -3.6171e-13 0.0085655 0.33115 0.61241 0.13183 0.60605 0.63056 0.471 0.60922 0.47525 0.27101 0.42799 1.0041 0.99296 15.9963 144.9797 0.00060055 -32.7987 0.018367
1.1216 0.98803 5.5187e-05 3.8182 0.012035 1.4764e-05 0.0011542 0.14994 0.00065828 0.15059 0.13724 0 0.037004 0.0389 0 0.89808 0.25032 0.0672 0.0093825 4.2512 0.058593 7.0383e-05 0.83148 0.0052701 0.0060075 0.77801 1.8879e-14 0.0082904 0.29244 0.5761 0.13183 0.60539 0.63021 0.45918 0.60624 0.47516 0.27054 0.42794 1.0045 0.99391 15.9963 144.9797 0.0006002 -34.2463 0.018603
1.1219 0.98803 5.5187e-05 3.8182 0.012035 1.4767e-05 0.0011542 0.14996 0.00065828 0.15061 0.13726 0 0.037003 0.0389 0 0.8981 0.25033 0.067202 0.0093829 4.2513 0.058595 7.0386e-05 0.83148 0.0052702 0.0060075 0.74441 -5.8673e-14 0.0080441 0.25438 0.5378 0.13183 0.60478 0.62991 0.44689 0.60351 0.47509 0.27001 0.42789 1.0049 0.99481 15.9963 144.9796 0.00059984 -35.658 0.018838
1.1221 0.98803 5.5187e-05 3.8182 0.012035 1.477e-05 0.0011542 0.14997 0.00065828 0.15063 0.13727 0 0.037002 0.0389 0 0.89812 0.25034 0.067205 0.0093832 4.2514 0.058597 7.0389e-05 0.83147 0.0052703 0.0060076 0.70831 -2.439e-13 0.0078237 0.21772 0.4979 0.13183 0.60421 0.62963 0.43407 0.60106 0.47503 0.26942 0.42785 1.0053 0.99567 15.9962 144.9795 0.00059946 -37.0242 0.019074
1.1223 0.98803 5.5187e-05 3.8182 0.012035 1.4773e-05 0.0011542 0.14999 0.00065828 0.15064 0.13729 0 0.037001 0.0389 0 0.89813 0.25034 0.067208 0.0093835 4.2514 0.058599 7.0391e-05 0.83147 0.0052703 0.0060077 0.6742 -2.2316e-13 0.007645 0.18651 0.46104 0.13183 0.60373 0.62941 0.42205 0.5991 0.47499 0.26882 0.4278 1.0057 0.99642 15.9962 144.9794 0.00059911 -38.2089 0.019286
1.1225 0.98803 5.5187e-05 3.8182 0.012035 1.4776e-05 0.0011542 0.15 0.00065828 0.15066 0.1373 0 0.037 0.0389 0 0.89815 0.25035 0.06721 0.0093838 4.2515 0.058601 7.0394e-05 0.83147 0.0052704 0.0060078 0.6391 -1.0357e-13 0.007483 0.15746 0.42372 0.13183 0.60328 0.62921 0.40956 0.5974 0.47496 0.26816 0.42776 1.0061 0.99714 15.9962 144.9794 0.00059876 -39.3482 0.019498
1.1227 0.98803 5.5187e-05 3.8182 0.012035 1.4778e-05 0.0011542 0.15002 0.00065828 0.15067 0.13732 0 0.036999 0.0389 0 0.89817 0.25036 0.067213 0.0093842 4.2516 0.058603 7.0396e-05 0.83147 0.0052705 0.0060078 0.60358 3.5738e-05 0.0073444 0.13096 0.3864 0.13183 0.60286 0.62902 0.39659 0.59594 0.47494 0.26744 0.42772 1.0065 0.99783 15.9962 144.9793 0.0005984 -40.4406 0.01971
1.1229 0.98803 5.5187e-05 3.8182 0.012035 1.478e-05 0.0011542 0.15003 0.00065828 0.15068 0.13733 0 0.036998 0.0389 0 0.89818 0.25036 0.067215 0.0093844 4.2516 0.058604 7.0398e-05 0.83147 0.0052705 0.0060079 0.57868 9.5469e-05 0.0072648 0.11403 0.36045 0.13183 0.60257 0.6289 0.3872 0.59506 0.47492 0.26689 0.42769 1.0068 0.99831 15.9962 144.9793 0.00059814 -41.1787 0.019859
1.123 0.98803 5.5187e-05 3.8182 0.012035 1.4782e-05 0.0011542 0.15004 0.00065828 0.15069 0.13733 0 0.036997 0.0389 0 0.89819 0.25037 0.067217 0.0093846 4.2517 0.058605 7.04e-05 0.83146 0.0052706 0.006008 0.55401 0.00016918 0.0071976 0.098532 0.33488 0.13183 0.6023 0.6288 0.37759 0.5943 0.47491 0.26631 0.42766 1.0071 0.99878 15.9962 144.9792 0.00059789 -41.8936 0.020008
1.1232 0.98803 5.5187e-05 3.8182 0.012035 1.4784e-05 0.0011542 0.15005 0.00065828 0.1507 0.13734 0 0.036997 0.0389 0 0.8982 0.25037 0.067219 0.0093848 4.2517 0.058607 7.0402e-05 0.83146 0.0052707 0.006008 0.5297 0.0002427 0.00714 0.084488 0.30985 0.13183 0.60204 0.6287 0.36775 0.59365 0.4749 0.26569 0.42763 1.0075 0.99924 15.9961 144.9792 0.00059763 -42.5857 0.020156
1.1233 0.98803 5.5187e-05 3.8182 0.012035 1.4786e-05 0.0011542 0.15006 0.00065828 0.15071 0.13735 0 0.036996 0.0389 0 0.89821 0.25038 0.06722 0.009385 4.2518 0.058608 7.0403e-05 0.83146 0.0052707 0.0060081 0.50826 0.00030928 0.0070958 0.073087 0.28788 0.13183 0.60181 0.62863 0.35872 0.59315 0.4749 0.2651 0.4276 1.0077 0.99965 15.9961 144.9792 0.0005974 -43.1894 0.02029
1.1234 0.98803 5.5187e-05 3.8182 0.012035 1.4788e-05 0.0011542 0.15007 0.00065828 0.15072 0.13736 0 0.036996 0.0389 0 0.89822 0.25038 0.067222 0.0093852 4.2518 0.058609 7.0405e-05 0.83146 0.0052708 0.0060081 0.48732 0.00038189 0.0070598 0.062836 0.26656 0.13183 0.6016 0.62857 0.34953 0.59273 0.4749 0.26449 0.42758 1.008 1 15.9961 144.9791 0.00059717 -43.7752 0.020424
1.1236 0.98803 5.5186e-05 3.8182 0.012035 1.4789e-05 0.0011542 0.15008 0.00065828 0.15073 0.13737 0 0.036995 0.0389 0 0.89823 0.25039 0.067223 0.0093854 4.2519 0.05861 7.0406e-05 0.83146 0.0052708 0.0060082 0.46695 0.00046351 0.0070324 0.053695 0.24595 0.13183 0.60139 0.62852 0.34019 0.59238 0.4749 0.26384 0.42755 1.0083 1.0004 15.9961 144.9791 0.00059694 -44.3435 0.020558
1.1237 0.98803 5.5186e-05 3.8182 0.012035 1.4791e-05 0.0011542 0.15008 0.00065828 0.15074 0.13738 0 0.036994 0.0389 0 0.89824 0.25039 0.067225 0.0093856 4.2519 0.058612 7.0408e-05 0.83146 0.0052708 0.0060082 0.44722 0.00055352 0.0070137 0.045613 0.22616 0.13183 0.60119 0.62848 0.33071 0.5921 0.4749 0.26316 0.42753 1.0086 1.0008 15.9961 144.9791 0.0005967 -44.8946 0.020692
1.1238 0.98803 5.5186e-05 3.8182 0.012035 1.4793e-05 0.0011542 0.15009 0.00065828 0.15075 0.13739 0 0.036994 0.0389 0 0.89825 0.25039 0.067227 0.0093858 4.2519 0.058613 7.041e-05 0.83146 0.0052709 0.0060083 0.42817 0.00065049 0.0070032 0.038526 0.20722 0.13183 0.60099 0.62846 0.32112 0.59187 0.4749 0.26244 0.4275 1.0089 1.0012 15.9961 144.979 0.00059647 -45.4289 0.020826
1.124 0.98803 5.5186e-05 3.8182 0.012035 1.4795e-05 0.0011542 0.1501 0.00065828 0.15076 0.1374 0 0.036993 0.0389 0 0.89826 0.2504 0.067228 0.009386 4.252 0.058614 7.0411e-05 0.83146 0.0052709 0.0060083 0.40983 0.00075428 0.0070007 0.032363 0.18921 0.13184 0.60081 0.62845 0.31144 0.5917 0.4749 0.2617 0.42747 1.0092 1.0016 15.9961 144.979 0.00059623 -45.9468 0.020959
1.1241 0.98803 5.5186e-05 3.8182 0.012035 1.4796e-05 0.0011542 0.15011 0.00065828 0.15077 0.1374 0 0.036993 0.0389 0 0.89827 0.2504 0.06723 0.0093862 4.252 0.058615 7.0413e-05 0.83146 0.005271 0.0060083 0.39224 0.00086589 0.0070061 0.027048 0.17216 0.13184 0.60063 0.62845 0.30167 0.59157 0.4749 0.26092 0.42745 1.0095 1.002 15.9961 144.979 0.00059599 -46.4486 0.021093
1.1243 0.98803 5.5186e-05 3.8182 0.012035 1.4798e-05 0.0011542 0.15012 0.00065828 0.15077 0.13741 0 0.036992 0.0389 0 0.89828 0.25041 0.067232 0.0093864 4.2521 0.058617 7.0414e-05 0.83145 0.005271 0.0060084 0.37541 0.00098633 0.0070196 0.0225 0.1561 0.13184 0.60046 0.62848 0.29184 0.59149 0.47491 0.2601 0.42742 1.0098 1.0023 15.9961 144.979 0.00059576 -46.9347 0.021227
1.1244 0.98803 5.5186e-05 3.8182 0.012035 1.48e-05 0.0011542 0.15013 0.00065828 0.15078 0.13742 0 0.036991 0.0389 0 0.89829 0.25041 0.067233 0.0093866 4.2521 0.058618 7.0416e-05 0.83145 0.0052711 0.0060084 0.35935 0.001116 0.0070412 0.018641 0.14106 0.13184 0.60029 0.62851 0.28197 0.59144 0.47491 0.25926 0.42739 1.0101 1.0027 15.9961 144.9789 0.00059552 -47.4056 0.021361
1.1245 0.98803 5.5186e-05 3.8182 0.012035 1.4802e-05 0.0011542 0.15014 0.00065828 0.15079 0.13743 0 0.036991 0.0389 0 0.8983 0.25042 0.067235 0.0093868 4.2522 0.058619 7.0417e-05 0.83145 0.0052711 0.0060085 0.34404 0.001255 0.0070707 0.015392 0.12703 0.13184 0.60014 0.62856 0.27209 0.59143 0.47492 0.25837 0.42737 1.0104 1.0031 15.9961 144.9789 0.00059528 -47.8615 0.021495
1.1247 0.98803 5.5186e-05 3.8182 0.012035 1.4803e-05 0.0011542 0.15015 0.00065828 0.1508 0.13744 0 0.03699 0.0389 0 0.89831 0.25042 0.067237 0.009387 4.2522 0.05862 7.0419e-05 0.83145 0.0052712 0.0060085 0.3295 0.0014033 0.0071081 0.012676 0.11401 0.13184 0.59999 0.62863 0.26221 0.59144 0.47493 0.25745 0.42734 1.0107 1.0034 15.996 144.9789 0.00059504 -48.3028 0.021629
1.1248 0.98803 5.5186e-05 3.8182 0.012035 1.4805e-05 0.0011542 0.15016 0.00065828 0.15081 0.13745 0 0.03699 0.0389 0 0.89832 0.25043 0.067238 0.0093872 4.2523 0.058622 7.0421e-05 0.83145 0.0052712 0.0060086 0.31569 0.0015615 0.0071533 0.010422 0.10199 0.13184 0.59984 0.62871 0.25236 0.59148 0.47494 0.2565 0.42732 1.011 1.0038 15.996 144.9789 0.0005948 -48.7301 0.021763
1.1249 0.98803 5.5186e-05 3.8182 0.012035 1.4807e-05 0.0011542 0.15017 0.00065828 0.15082 0.13746 0 0.036989 0.0389 0 0.89833 0.25043 0.06724 0.0093874 4.2523 0.058623 7.0422e-05 0.83145 0.0052713 0.0060086 0.3026 0.0017298 0.0072063 0.0085658 0.090948 0.13184 0.59971 0.62881 0.24257 0.59154 0.47495 0.25551 0.42729 1.0113 1.0042 15.996 144.9789 0.00059456 -49.1436 0.021897
1.1251 0.98803 5.5186e-05 3.8182 0.012035 1.4809e-05 0.0011542 0.15018 0.00065828 0.15083 0.13746 0 0.036988 0.0389 0 0.89834 0.25044 0.067241 0.0093876 4.2524 0.058624 7.0424e-05 0.83145 0.0052713 0.0060087 0.29021 0.0019087 0.007267 0.007046 0.08085 0.13184 0.59957 0.62892 0.23285 0.59162 0.47496 0.25449 0.42727 1.0116 1.0045 15.996 144.9788 0.00059432 -49.5438 0.02203
1.1252 0.98803 5.5186e-05 3.8182 0.012035 1.4811e-05 0.0011542 0.15019 0.00065828 0.15084 0.13747 0 0.036988 0.0389 0 0.89835 0.25044 0.067243 0.0093878 4.2524 0.058625 7.0425e-05 0.83145 0.0052714 0.0060087 0.27849 0.0020983 0.0073354 0.0058093 0.071659 0.13184 0.59945 0.62904 0.22324 0.59172 0.47497 0.25343 0.42724 1.0119 1.0049 15.996 144.9788 0.00059408 -49.9311 0.022164
1.1253 0.98803 5.5186e-05 3.8182 0.012035 1.4812e-05 0.0011542 0.15019 0.00065828 0.15085 0.13748 0 0.036987 0.0389 0 0.89836 0.25044 0.067245 0.009388 4.2524 0.058626 7.0427e-05 0.83144 0.0052714 0.0060088 0.26741 0.0022989 0.0074114 0.0048084 0.063333 0.13184 0.59933 0.62917 0.21374 0.59182 0.47498 0.25234 0.42721 1.0122 1.0052 15.996 144.9788 0.00059384 -50.3059 0.022298
1.1256 0.98803 5.5186e-05 3.8182 0.012035 1.4816e-05 0.0011542 0.15021 0.00065829 0.15087 0.1375 0 0.036986 0.0389 0 0.89838 0.25045 0.067248 0.0093884 4.2525 0.058629 7.043e-05 0.83144 0.0052715 0.0060089 0.24707 0.0027336 0.0075858 0.0033542 0.049083 0.13184 0.59911 0.62947 0.1952 0.59207 0.475 0.25006 0.42716 1.0128 1.0059 15.996 144.9788 0.00059336 -51.0196 0.022566
1.1259 0.98803 5.5186e-05 3.8182 0.012035 1.4819e-05 0.0011542 0.15023 0.00065829 0.15088 0.13752 0 0.036985 0.0389 0 0.89841 0.25046 0.067251 0.0093888 4.2526 0.058631 7.0433e-05 0.83144 0.0052716 0.006009 0.22893 0.0032148 0.0077899 0.0024211 0.037695 0.13184 0.59891 0.6298 0.17738 0.59235 0.47502 0.24764 0.42711 1.0134 1.0066 15.996 144.9787 0.00059287 -51.6884 0.022834
1.1261 0.98803 5.5186e-05 3.8182 0.012035 1.4823e-05 0.0011542 0.15025 0.00065829 0.1509 0.13753 0 0.036984 0.0389 0 0.89843 0.25047 0.067255 0.0093892 4.2527 0.058634 7.0436e-05 0.83144 0.0052717 0.0060091 0.21277 0.0037439 0.008023 0.0018242 0.028744 0.13184 0.59873 0.63017 0.16043 0.59265 0.47505 0.24508 0.42706 1.014 1.0073 15.996 144.9787 0.00059239 -52.3157 0.023101
1.1264 0.98803 5.5186e-05 3.8182 0.012035 1.4826e-05 0.0011542 0.15027 0.00065829 0.15092 0.13755 0 0.036983 0.0389 0 0.89845 0.25048 0.067258 0.0093896 4.2528 0.058636 7.044e-05 0.83143 0.0052718 0.0060092 0.19834 0.0043221 0.0082847 0.0014393 0.02182 0.13184 0.59857 0.63056 0.14445 0.59297 0.47508 0.24241 0.42701 1.0146 1.0079 15.996 144.9787 0.0005919 -52.9047 0.023369
1.1267 0.98803 5.5186e-05 3.8182 0.012035 1.483e-05 0.0011542 0.15029 0.00065829 0.15094 0.13757 0 0.036981 0.0389 0 0.89847 0.25049 0.067261 0.00939 4.2529 0.058639 7.0443e-05 0.83143 0.0052719 0.0060093 0.18543 0.0049504 0.0085744 0.0011854 0.016541 0.13184 0.59842 0.63096 0.12952 0.5933 0.4751 0.23961 0.42696 1.0153 1.0086 15.996 144.9787 0.00059141 -53.4588 0.023637
1.1269 0.98803 5.5186e-05 3.8182 0.012035 1.4833e-05 0.0011542 0.1503 0.00065829 0.15096 0.13758 0 0.03698 0.0389 0 0.89849 0.2505 0.067264 0.0093904 4.253 0.058641 7.0446e-05 0.83143 0.005272 0.0060094 0.17386 0.0056295 0.0088915 0.0010113 0.012569 0.13184 0.5983 0.63138 0.11569 0.59364 0.47513 0.2367 0.42691 1.0159 1.0093 15.996 144.9786 0.00059092 -53.9812 0.023905
1.1272 0.98803 5.5186e-05 3.8182 0.012035 1.4837e-05 0.0011542 0.15032 0.00065829 0.15098 0.1376 0 0.036979 0.0389 0 0.89851 0.25051 0.067268 0.0093909 4.2531 0.058644 7.0449e-05 0.83143 0.0052721 0.0060095 0.16344 0.0063602 0.0092356 0.00088608 0.0096141 0.13184 0.59818 0.63182 0.103 0.59397 0.47516 0.23368 0.42686 1.0165 1.0099 15.996 144.9786 0.00059043 -54.4749 0.024172
1.1275 0.98803 5.5186e-05 3.8182 0.012035 1.484e-05 0.0011542 0.15034 0.00065829 0.15099 0.13762 0 0.036978 0.0389 0 0.89853 0.25052 0.067271 0.0093913 4.2532 0.058646 7.0452e-05 0.83142 0.0052722 0.0060096 0.15403 0.0071432 0.0096062 0.00079123 0.0074372 0.13185 0.59809 0.63226 0.091447 0.59432 0.47519 0.23055 0.42681 1.0171 1.0106 15.9959 144.9786 0.00058993 -54.943 0.02444
1.1277 0.98803 5.5186e-05 3.8182 0.012035 1.4844e-05 0.0011542 0.15036 0.00065829 0.15101 0.13764 0 0.036977 0.0389 0 0.89855 0.25053 0.067274 0.0093917 4.2533 0.058649 7.0455e-05 0.83142 0.0052723 0.0060097 0.14549 0.0079793 0.010003 0.00071606 0.0058443 0.13185 0.59801 0.6327 0.081006 0.59466 0.47522 0.22733 0.42676 1.0178 1.0113 15.9959 144.9786 0.00058944 -55.3882 0.024708
1.128 0.98803 5.5186e-05 3.8182 0.012035 1.4847e-05 0.0011542 0.15038 0.00065829 0.15103 0.13765 0 0.036976 0.0389 0 0.89857 0.25054 0.067277 0.0093921 4.2534 0.058651 7.0459e-05 0.83142 0.0052724 0.0060098 0.13771 0.0088689 0.010426 0.00065426 0.0046831 0.13185 0.59794 0.63315 0.071644 0.595 0.47525 0.22401 0.42672 1.0184 1.0119 15.9959 144.9786 0.00058895 -55.8129 0.024976
1.1283 0.98803 5.5186e-05 3.8182 0.012035 1.4851e-05 0.0011542 0.1504 0.00065829 0.15105 0.13767 0 0.036974 0.0389 0 0.89859 0.25054 0.067281 0.0093925 4.2534 0.058654 7.0462e-05 0.83142 0.0052725 0.0060098 0.13058 0.0098129 0.010874 0.00060196 0.0038366 0.13185 0.59788 0.6336 0.063307 0.59534 0.47528 0.22061 0.42667 1.019 1.0126 15.9959 144.9786 0.00058845 -56.2196 0.025243
1.1285 0.98803 5.5186e-05 3.8182 0.012035 1.4855e-05 0.0011542 0.15041 0.00065829 0.15107 0.13769 0 0.036973 0.0389 0 0.89861 0.25055 0.067284 0.0093929 4.2535 0.058656 7.0465e-05 0.83141 0.0052726 0.0060099 0.12403 0.010812 0.011347 0.00055675 0.0032168 0.13185 0.59783 0.63405 0.055934 0.59568 0.47531 0.21713 0.42662 1.0196 1.0132 15.9959 144.9786 0.00058796 -56.6105 0.025511
1.1288 0.98803 5.5186e-05 3.8182 0.012035 1.4858e-05 0.0011542 0.15043 0.00065829 0.15109 0.1377 0 0.036972 0.0389 0 0.89863 0.25056 0.067287 0.0093933 4.2536 0.058658 7.0468e-05 0.83141 0.0052727 0.00601 0.11797 0.011867 0.011845 0.00051703 0.0027586 0.13185 0.5978 0.6345 0.049454 0.59601 0.47535 0.21358 0.42657 1.0203 1.0139 15.9959 144.9786 0.00058746 -56.9875 0.025779
1.129 0.98803 5.5186e-05 3.8182 0.012035 1.4861e-05 0.0011542 0.15045 0.00065829 0.1511 0.13772 0 0.036971 0.0389 0 0.89865 0.25057 0.06729 0.0093936 4.2537 0.05866 7.047e-05 0.83141 0.0052727 0.0060101 0.11384 0.012671 0.012224 0.00049094 0.0024991 0.13185 0.59778 0.63483 0.045255 0.59625 0.47537 0.21095 0.42653 1.0207 1.0143 15.9959 144.9785 0.0005871 -57.2542 0.025974
1.1292 0.98803 5.5186e-05 3.8182 0.012035 1.4863e-05 0.0011542 0.15046 0.00065829 0.15111 0.13773 0 0.03697 0.0389 0 0.89866 0.25058 0.067292 0.0093938 4.2538 0.058662 7.0473e-05 0.83141 0.0052728 0.0060102 0.10992 0.013506 0.012616 0.00046689 0.0022862 0.13185 0.59777 0.63516 0.041461 0.5965 0.47539 0.20828 0.4265 1.0212 1.0148 15.9959 144.9785 0.00058674 -57.5151 0.026169
1.1294 0.98803 5.5186e-05 3.8182 0.012035 1.4866e-05 0.0011542 0.15047 0.00065829 0.15113 0.13774 0 0.036969 0.0389 0 0.89867 0.25058 0.067294 0.0093941 4.2538 0.058664 7.0475e-05 0.83141 0.0052729 0.0060103 0.1062 0.014371 0.013021 0.00044468 0.0021095 0.13185 0.59776 0.63549 0.038041 0.59673 0.47542 0.20559 0.42647 1.0216 1.0153 15.9959 144.9785 0.00058638 -57.7707 0.026364
1.1296 0.98803 5.5186e-05 3.8182 0.012035 1.4868e-05 0.0011542 0.15049 0.00065829 0.15114 0.13775 0 0.036969 0.0389 0 0.89869 0.25059 0.067297 0.0093944 4.2539 0.058666 7.0477e-05 0.8314 0.005273 0.0060103 0.10264 0.015268 0.01344 0.00042407 0.001961 0.13185 0.59776 0.63582 0.034968 0.59697 0.47544 0.20286 0.42643 1.0221 1.0157 15.9959 144.9785 0.00058601 -58.0216 0.026558
1.1298 0.98803 5.5186e-05 3.8182 0.012035 1.4871e-05 0.0011542 0.1505 0.00065829 0.15115 0.13777 0 0.036968 0.0389 0 0.8987 0.2506 0.067299 0.0093947 4.254 0.058667 7.048e-05 0.8314 0.005273 0.0060104 0.099254 0.016198 0.013871 0.00040486 0.0018342 0.13185 0.59777 0.63614 0.032211 0.59721 0.47546 0.2001 0.4264 1.0226 1.0162 15.9959 144.9785 0.00058565 -58.2681 0.026753
1.13 0.98803 5.5186e-05 3.8182 0.012035 1.4873e-05 0.0011542 0.15051 0.00065829 0.15117 0.13778 0 0.036967 0.0389 0 0.89872 0.2506 0.067302 0.009395 4.254 0.058669 7.0482e-05 0.8314 0.0052731 0.0060105 0.096014 0.01716 0.014317 0.00038688 0.0017246 0.13185 0.59777 0.63647 0.029744 0.59744 0.47549 0.19731 0.42636 1.023 1.0167 15.9959 144.9785 0.00058529 -58.5108 0.026948
1.1302 0.98803 5.5186e-05 3.8182 0.012035 1.4876e-05 0.0011542 0.15053 0.00065829 0.15118 0.13779 0 0.036966 0.0389 0 0.89873 0.25061 0.067304 0.0093953 4.2541 0.058671 7.0484e-05 0.8314 0.0052732 0.0060105 0.092912 0.018156 0.014776 0.00037002 0.0016285 0.13185 0.59779 0.6368 0.027541 0.59767 0.47551 0.1945 0.42633 1.0235 1.0171 15.9959 144.9785 0.00058493 -58.7499 0.027143
1.1304 0.98803 5.5186e-05 3.8182 0.012035 1.4879e-05 0.0011542 0.15054 0.00065829 0.15119 0.1378 0 0.036965 0.0389 0 0.89875 0.25062 0.067306 0.0093956 4.2542 0.058673 7.0487e-05 0.8314 0.0052732 0.0060106 0.089939 0.019185 0.015248 0.00035416 0.0015432 0.13185 0.59781 0.63713 0.025576 0.5979 0.47554 0.19167 0.42629 1.0239 1.0176 15.9959 144.9785 0.00058456 -58.9859 0.027338
1.1306 0.98803 5.5186e-05 3.8182 0.012035 1.4881e-05 0.0011542 0.15055 0.00065829 0.15121 0.13782 0 0.036964 0.0389 0 0.89876 0.25062 0.067309 0.0093959 4.2542 0.058675 7.0489e-05 0.8314 0.0052733 0.0060107 0.087083 0.020249 0.015735 0.0003392 0.0014664 0.13185 0.59783 0.63745 0.023826 0.59813 0.47556 0.18881 0.42626 1.0244 1.0181 15.9959 144.9785 0.0005842 -59.219 0.027533
1.1308 0.98803 5.5186e-05 3.8182 0.012035 1.4884e-05 0.0011542 0.15057 0.00065829 0.15122 0.13783 0 0.036963 0.0389 0 0.89878 0.25063 0.067311 0.0093962 4.2543 0.058676 7.0491e-05 0.83139 0.0052734 0.0060107 0.08434 0.021349 0.016235 0.00032508 0.0013964 0.13186 0.59786 0.63778 0.02227 0.59836 0.47558 0.18593 0.42623 1.0249 1.0185 15.9959 144.9785 0.00058384 -59.4495 0.027728
1.1309 0.98803 5.5186e-05 3.8182 0.012035 1.4886e-05 0.0011542 0.15058 0.00065829 0.15123 0.13784 0 0.036963 0.0389 0 0.89879 0.25064 0.067314 0.0093965 4.2544 0.058678 7.0493e-05 0.83139 0.0052734 0.0060108 0.081698 0.022485 0.016749 0.00031172 0.0013322 0.13186 0.59789 0.63811 0.020885 0.59859 0.47561 0.18304 0.42619 1.0253 1.019 15.9959 144.9785 0.00058347 -59.6777 0.027923
1.1311 0.98803 5.5186e-05 3.8182 0.012035 1.4889e-05 0.0011542 0.15059 0.00065829 0.15125 0.13785 0 0.036962 0.0389 0 0.89881 0.25064 0.067316 0.0093968 4.2544 0.05868 7.0496e-05 0.83139 0.0052735 0.0060109 0.079152 0.023658 0.017278 0.00029906 0.0012728 0.13186 0.59792 0.63843 0.019655 0.59881 0.47563 0.18012 0.42616 1.0258 1.0195 15.9959 144.9785 0.00058311 -59.9037 0.028118
1.1313 0.98803 5.5186e-05 3.8182 0.012035 1.4891e-05 0.0011542 0.1506 0.00065829 0.15126 0.13786 0 0.036961 0.0389 0 0.89882 0.25065 0.067318 0.009397 4.2545 0.058682 7.0498e-05 0.83139 0.0052736 0.006011 0.076942 0.024746 0.017765 0.00028821 0.0012229 0.13186 0.59796 0.63873 0.018665 0.59901 0.47566 0.17748 0.42613 1.0262 1.0199 15.9959 144.9785 0.00058278 -60.1053 0.028293
1.1315 0.98803 5.5186e-05 3.8182 0.012035 1.4893e-05 0.0011542 0.15062 0.00065829 0.15127 0.13788 0 0.03696 0.0389 0 0.89884 0.25065 0.06732 0.0093973 4.2545 0.058683 7.05e-05 0.83139 0.0052736 0.006011 0.074803 0.025866 0.018265 0.00027785 0.0011758 0.13186 0.598 0.63902 0.017774 0.59921 0.47568 0.17484 0.4261 1.0266 1.0203 15.9959 144.9785 0.00058246 -60.3055 0.028469
1.1317 0.98803 5.5186e-05 3.8182 0.012035 1.4896e-05 0.0011542 0.15063 0.00065829 0.15128 0.13789 0 0.036959 0.0389 0 0.89885 0.25066 0.067322 0.0093976 4.2546 0.058685 7.0502e-05 0.83139 0.0052737 0.0060111 0.072731 0.027018 0.018777 0.00026794 0.0011314 0.13186 0.59804 0.63931 0.016971 0.5994 0.4757 0.17218 0.42607 1.027 1.0207 15.9959 144.9785 0.00058213 -60.5044 0.028644
1.1319 0.98803 5.5186e-05 3.8182 0.012035 1.4899e-05 0.0011542 0.15064 0.00065829 0.1513 0.1379 0 0.036958 0.0389 0 0.89887 0.25067 0.067325 0.0093979 4.2547 0.058687 7.0505e-05 0.83138 0.0052738 0.0060112 0.070071 0.028601 0.019476 0.00025541 0.0010758 0.13186 0.5981 0.6397 0.016024 0.59966 0.47573 0.16862 0.42603 1.0276 1.0213 15.9959 144.9785 0.00058169 -60.767 0.028878
1.1321 0.98803 5.5186e-05 3.8182 0.012035 1.4902e-05 0.0011542 0.15066 0.00065829 0.15131 0.13792 0 0.036957 0.0389 0 0.89889 0.25068 0.067328 0.0093983 4.2548 0.058689 7.0508e-05 0.83138 0.0052739 0.0060113 0.06752 0.030244 0.020197 0.00024359 0.0010237 0.13186 0.59817 0.64009 0.015197 0.59992 0.47576 0.16506 0.42599 1.0281 1.0219 15.9959 144.9785 0.00058126 -61.0276 0.029111
1.1324 0.98803 5.5186e-05 3.8182 0.012035 1.4905e-05 0.0011542 0.15068 0.00065829 0.15133 0.13793 0 0.036956 0.0389 0 0.8989 0.25068 0.067331 0.0093986 4.2548 0.058691 7.051e-05 0.83138 0.005274 0.0060113 0.06507 0.031949 0.020941 0.0002324 0.00097488 0.13186 0.59824 0.64047 0.014471 0.60018 0.47579 0.16148 0.42595 1.0287 1.0224 15.9959 144.9785 0.00058082 -61.2862 0.029345
1.1326 0.98803 5.5186e-05 3.8182 0.012035 1.4908e-05 0.0011542 0.15069 0.00065829 0.15134 0.13795 0 0.036955 0.0389 0 0.89892 0.25069 0.067334 0.009399 4.2549 0.058693 7.0513e-05 0.83138 0.005274 0.0060114 0.062717 0.033717 0.021706 0.00022181 0.0009289 0.13186 0.59832 0.64086 0.01383 0.60043 0.47582 0.15789 0.42591 1.0292 1.023 15.9959 144.9785 0.00058038 -61.5431 0.029578
1.1328 0.98803 5.5186e-05 3.8182 0.012035 1.4911e-05 0.0011542 0.15071 0.00065829 0.15136 0.13796 0 0.036954 0.0389 0 0.89894 0.2507 0.067337 0.0093993 4.255 0.058696 7.0516e-05 0.83137 0.0052741 0.0060115 0.060455 0.03555 0.022495 0.00021178 0.00088554 0.13186 0.5984 0.64124 0.013263 0.60068 0.47585 0.15429 0.42587 1.0298 1.0235 15.9959 144.9784 0.00057995 -61.7983 0.029812
1.1331 0.98803 5.5186e-05 3.8182 0.012035 1.4914e-05 0.0011542 0.15072 0.00065829 0.15138 0.13798 0 0.036953 0.0389 0 0.89896 0.25071 0.06734 0.0093997 4.2551 0.058698 7.0519e-05 0.83137 0.0052742 0.0060116 0.058281 0.03745 0.023307 0.00020227 0.00084458 0.13186 0.59849 0.64163 0.012756 0.60093 0.47588 0.15069 0.42583 1.0303 1.0241 15.9959 144.9784 0.00057951 -62.0519 0.030045
1.1333 0.98803 5.5186e-05 3.8182 0.012035 1.4917e-05 0.0011542 0.15074 0.0006583 0.15139 0.13799 0 0.036952 0.0389 0 0.89897 0.25072 0.067343 0.0094 4.2552 0.0587 7.0521e-05 0.83137 0.0052743 0.0060117 0.05619 0.039418 0.024142 0.00019325 0.00080584 0.13186 0.59858 0.64201 0.0123 0.60118 0.47591 0.1471 0.42579 1.0309 1.0246 15.9959 144.9784 0.00057907 -62.304 0.030279
1.1335 0.98803 5.5186e-05 3.8182 0.012035 1.492e-05 0.0011542 0.15075 0.0006583 0.15141 0.13801 0 0.036951 0.0389 0 0.89899 0.25072 0.067345 0.0094004 4.2552 0.058702 7.0524e-05 0.83137 0.0052744 0.0060118 0.054179 0.041458 0.025002 0.00018469 0.00076917 0.13186 0.59868 0.64239 0.011888 0.60142 0.47594 0.1435 0.42576 1.0314 1.0252 15.9959 144.9784 0.00057863 -62.5547 0.030512
1.1338 0.98803 5.5186e-05 3.8182 0.012035 1.4923e-05 0.0011542 0.15077 0.0006583 0.15142 0.13802 0 0.03695 0.0389 0 0.89901 0.25073 0.067348 0.0094007 4.2553 0.058704 7.0527e-05 0.83137 0.0052745 0.0060118 0.052245 0.043571 0.025887 0.00017655 0.00073444 0.13186 0.59879 0.64278 0.011512 0.60167 0.47597 0.13991 0.42572 1.032 1.0257 15.9959 144.9784 0.0005782 -62.804 0.030746
1.1342 0.98803 5.5186e-05 3.8182 0.012035 1.4929e-05 0.0011542 0.1508 0.0006583 0.15146 0.13805 0 0.036948 0.0389 0 0.89905 0.25075 0.067354 0.0094014 4.2555 0.058709 7.0532e-05 0.83136 0.0052746 0.006012 0.048593 0.048023 0.027731 0.00016147 0.00067026 0.13187 0.59901 0.64354 0.010847 0.60215 0.47603 0.13275 0.42564 1.0331 1.0268 15.9959 144.9784 0.00057732 -63.2986 0.031212
1.1347 0.98803 5.5186e-05 3.8182 0.012035 1.4935e-05 0.0011542 0.15083 0.0006583 0.15148 0.13808 0 0.036946 0.0389 0 0.89908 0.25076 0.067359 0.0094021 4.2556 0.058712 7.0537e-05 0.83136 0.0052748 0.0060122 0.045538 0.052301 0.02948 0.00014913 0.00061795 0.13187 0.59922 0.64422 0.010325 0.60258 0.47608 0.12635 0.42557 1.0341 1.0278 15.9959 144.9784 0.00057653 -63.7393 0.031633
1.1351 0.98803 5.5186e-05 3.8182 0.012035 1.494e-05 0.0011542 0.15086 0.0006583 0.15151 0.1381 0 0.036945 0.0389 0 0.89911 0.25078 0.067364 0.0094027 4.2558 0.058716 7.0542e-05 0.83135 0.0052749 0.0060123 0.042686 0.056848 0.031317 0.00013784 0.00057024 0.13187 0.59945 0.6449 0.0098565 0.603 0.47613 0.12001 0.42551 1.035 1.0288 15.9959 144.9784 0.00057575 -64.1761 0.032053
1.1355 0.98803 5.5186e-05 3.8182 0.012035 1.4946e-05 0.0011542 0.15089 0.0006583 0.15154 0.13813 0 0.036943 0.0389 0 0.89914 0.25079 0.067369 0.0094033 4.2559 0.05872 7.0547e-05 0.83135 0.0052751 0.0060125 0.040024 0.061677 0.033244 0.00012751 0.00052668 0.13187 0.59969 0.64558 0.0094298 0.60342 0.47619 0.11374 0.42544 1.036 1.0298 15.9959 144.9784 0.00057496 -64.6089 0.032473
1.1359 0.98803 5.5186e-05 3.8182 0.012035 1.4951e-05 0.0011542 0.15092 0.0006583 0.15157 0.13816 0 0.036941 0.0389 0 0.89918 0.2508 0.067375 0.0094039 4.2561 0.058724 7.0552e-05 0.83135 0.0052752 0.0060126 0.037539 0.066802 0.035265 0.00011804 0.00048686 0.13187 0.59994 0.64626 0.0090358 0.60383 0.47624 0.10757 0.42538 1.037 1.0308 15.996 144.9784 0.00057417 -65.0379 0.032894
1.1363 0.98803 5.5186e-05 3.8182 0.012035 1.4957e-05 0.0011542 0.15095 0.0006583 0.1516 0.13818 0 0.036939 0.0389 0 0.89921 0.25082 0.06738 0.0094046 4.2562 0.058728 7.0557e-05 0.83134 0.0052754 0.0060128 0.035216 0.072235 0.037384 0.00010936 0.00045042 0.13187 0.6002 0.64693 0.0086685 0.60425 0.4763 0.1015 0.42531 1.038 1.0318 15.996 144.9784 0.00057338 -65.463 0.033314
1.1368 0.98803 5.5186e-05 3.8182 0.012035 1.4963e-05 0.0011542 0.15097 0.0006583 0.15163 0.13821 0 0.036937 0.0389 0 0.89924 0.25083 0.067385 0.0094052 4.2564 0.058732 7.0562e-05 0.83134 0.0052755 0.0060129 0.03306 0.077991 0.039603 0.00010138 0.00041705 0.13187 0.60048 0.64761 0.0083239 0.60465 0.47635 0.095557 0.42525 1.039 1.0328 15.996 144.9783 0.00057259 -65.8843 0.033734
1.137 0.98803 5.5186e-05 3.8182 0.012035 1.4966e-05 0.0011542 0.15099 0.0006583 0.15165 0.13823 0 0.036936 0.0389 0 0.89926 0.25084 0.067388 0.0094056 4.2564 0.058734 7.0566e-05 0.83134 0.0052756 0.006013 0.031725 0.081909 0.0411 9.6556e-05 0.00039688 0.13187 0.60066 0.64804 0.0081108 0.60492 0.47639 0.091769 0.42521 1.0396 1.0335 15.996 144.9783 0.00057207 -66.1559 0.034007
1.1373 0.98803 5.5186e-05 3.8182 0.012035 1.497e-05 0.0011542 0.15101 0.0006583 0.15166 0.13825 0 0.036935 0.0389 0 0.89928 0.25085 0.067392 0.009406 4.2565 0.058737 7.0569e-05 0.83133 0.0052757 0.0060131 0.030449 0.085972 0.042642 9.1988e-05 0.00037781 0.13188 0.60085 0.64847 0.0079055 0.60518 0.47642 0.088043 0.42517 1.0403 1.0341 15.996 144.9783 0.00057156 -66.4259 0.03428
1.1375 0.98803 5.5186e-05 3.8182 0.012035 1.4973e-05 0.0011542 0.15103 0.0006583 0.15168 0.13826 0 0.036934 0.0389 0 0.8993 0.25086 0.067395 0.0094064 4.2566 0.058739 7.0572e-05 0.83133 0.0052758 0.0060132 0.029352 0.089755 0.04407 8.8086e-05 0.00036154 0.13188 0.60103 0.64886 0.007727 0.60541 0.47645 0.084747 0.42513 1.0408 1.0347 15.996 144.9783 0.0005711 -66.6675 0.034526
1.1378 0.98803 5.5186e-05 3.8182 0.012035 1.4976e-05 0.0011542 0.15104 0.0006583 0.1517 0.13828 0 0.036933 0.0389 0 0.89932 0.25087 0.067398 0.0094068 4.2567 0.058741 7.0575e-05 0.83133 0.0052759 0.0060133 0.028298 0.093662 0.045536 8.437e-05 0.00034606 0.13188 0.6012 0.64925 0.0075541 0.60565 0.47649 0.081506 0.42509 1.0414 1.0353 15.996 144.9783 0.00057064 -66.9078 0.034772
1.138 0.98803 5.5186e-05 3.8182 0.012035 1.4979e-05 0.0011542 0.15106 0.0006583 0.15171 0.13829 0 0.036932 0.0389 0 0.89934 0.25088 0.067401 0.0094071 4.2568 0.058744 7.0578e-05 0.83133 0.005276 0.0060134 0.027285 0.097694 0.047041 8.0831e-05 0.00033133 0.13188 0.60139 0.64964 0.0073864 0.60588 0.47652 0.078325 0.42506 1.042 1.0359 15.996 144.9783 0.00057017 -67.1467 0.035017
1.1383 0.98803 5.5186e-05 3.8182 0.012035 1.4983e-05 0.0011542 0.15108 0.0006583 0.15173 0.13831 0 0.036931 0.0389 0 0.89936 0.25089 0.067404 0.0094075 4.2569 0.058746 7.0581e-05 0.83132 0.0052761 0.0060135 0.026311 0.10185 0.048585 7.746e-05 0.00031732 0.13188 0.60157 0.65003 0.0072237 0.60611 0.47655 0.075204 0.42502 1.0426 1.0364 15.996 144.9783 0.00056971 -67.3843 0.035263
1.1385 0.98803 5.5186e-05 3.8182 0.012035 1.4986e-05 0.0011542 0.15109 0.0006583 0.15175 0.13832 0 0.036929 0.0389 0 0.89938 0.25089 0.067407 0.0094079 4.257 0.058748 7.0583e-05 0.83132 0.0052762 0.0060136 0.025376 0.10615 0.050171 7.4248e-05 0.00030398 0.13188 0.60176 0.65042 0.0070659 0.60635 0.47658 0.072148 0.42499 1.0431 1.037 15.996 144.9783 0.00056925 -67.6205 0.035509
1.1388 0.98803 5.5186e-05 3.8182 0.012035 1.4989e-05 0.0011542 0.15111 0.0006583 0.15176 0.13834 0 0.036928 0.0389 0 0.89939 0.2509 0.06741 0.0094083 4.257 0.05875 7.0586e-05 0.83132 0.0052763 0.0060137 0.024478 0.11057 0.051798 7.1188e-05 0.00029128 0.13188 0.60195 0.6508 0.0069128 0.60658 0.47661 0.069157 0.42495 1.0437 1.0376 15.996 144.9783 0.00056879 -67.8554 0.035754
1.139 0.98803 5.5186e-05 3.8182 0.012035 1.4992e-05 0.0011542 0.15113 0.0006583 0.15178 0.13835 0 0.036927 0.0389 0 0.89941 0.25091 0.067413 0.0094086 4.2571 0.058753 7.0589e-05 0.83132 0.0052764 0.0060138 0.023615 0.11513 0.053468 6.8272e-05 0.00027919 0.13188 0.60214 0.65119 0.0067642 0.60681 0.47665 0.066234 0.42492 1.0443 1.0382 15.996 144.9783 0.00056832 -68.0889 0.036
1.1393 0.98803 5.5186e-05 3.8182 0.012035 1.4996e-05 0.0011542 0.15114 0.0006583 0.1518 0.13837 0 0.036926 0.0389 0 0.89943 0.25092 0.067416 0.009409 4.2572 0.058755 7.0592e-05 0.83132 0.0052765 0.0060139 0.022785 0.11983 0.055181 6.5492e-05 0.00026767 0.13188 0.60234 0.65157 0.0066198 0.60704 0.47668 0.06338 0.42489 1.0449 1.0388 15.9961 144.9783 0.00056786 -68.321 0.036246
1.1398 0.98803 5.5185e-05 3.8182 0.012035 1.5002e-05 0.0011542 0.15118 0.0006583 0.15183 0.1384 0 0.036924 0.0389 0 0.89947 0.25094 0.067422 0.0094097 4.2574 0.05876 7.0598e-05 0.83131 0.0052766 0.006014 0.021223 0.12964 0.058741 6.0314e-05 0.00024625 0.13188 0.60274 0.65234 0.0063436 0.60751 0.47674 0.057889 0.42482 1.046 1.0399 15.9961 144.9783 0.00056694 -68.7809 0.036737
1.1402 0.98803 5.5185e-05 3.8182 0.012035 1.5008e-05 0.0011542 0.15121 0.0006583 0.15186 0.13843 0 0.036922 0.0389 0 0.8995 0.25095 0.067427 0.0094104 4.2575 0.058764 7.0603e-05 0.83131 0.0052768 0.0060142 0.01992 0.13896 0.062105 5.6056e-05 0.00022866 0.13188 0.60311 0.65302 0.0061083 0.60792 0.4768 0.053201 0.42476 1.0471 1.041 15.9961 144.9782 0.0005661 -69.1899 0.03718
1.1406 0.98803 5.5185e-05 3.8182 0.012035 1.5014e-05 0.0011542 0.15124 0.0006583 0.15189 0.13846 0 0.03692 0.0389 0 0.89954 0.25097 0.067433 0.0094111 4.2577 0.058768 7.0609e-05 0.8313 0.005277 0.0060144 0.018707 0.14877 0.065625 5.2145e-05 0.00021252 0.13189 0.60348 0.65371 0.0058849 0.60834 0.47686 0.048761 0.4247 1.0481 1.042 15.9961 144.9782 0.00056527 -69.5942 0.037622
1.1411 0.98803 5.5185e-05 3.8182 0.012035 1.5019e-05 0.0011542 0.15127 0.00065831 0.15192 0.13849 0 0.036918 0.0389 0 0.89957 0.25098 0.067438 0.0094117 4.2578 0.058772 7.0614e-05 0.8313 0.0052771 0.0060145 0.017578 0.15905 0.069309 4.855e-05 0.00019771 0.13189 0.60387 0.65439 0.0056728 0.60876 0.47692 0.044572 0.42464 1.0491 1.043 15.9961 144.9782 0.00056444 -69.9936 0.038064
1.142 0.98803 5.5185e-05 3.8182 0.012035 1.5031e-05 0.0011542 0.15133 0.00065831 0.15198 0.13854 0 0.036915 0.0389 0 0.89964 0.25101 0.067449 0.0094131 4.2582 0.05878 7.0624e-05 0.83129 0.0052774 0.0060148 0.01555 0.18112 0.077192 4.2203e-05 0.00017159 0.13189 0.60466 0.65574 0.0052797 0.6096 0.47704 0.03696 0.42453 1.0512 1.0451 15.9962 144.9782 0.00056277 -70.7772 0.038949
1.1429 0.98803 5.5185e-05 3.8182 0.012035 1.5043e-05 0.0011542 0.15139 0.00065831 0.15204 0.1386 0 0.036911 0.0389 0 0.89971 0.25104 0.06746 0.0094144 4.2585 0.058788 7.0635e-05 0.83128 0.0052778 0.0060152 0.013793 0.20519 0.085809 3.6827e-05 0.00014952 0.13189 0.60547 0.65709 0.0049246 0.61045 0.47716 0.030363 0.42442 1.0532 1.0472 15.9962 144.9782 0.00056111 -71.5399 0.039833
1.1437 0.98803 5.5185e-05 3.8182 0.012035 1.5054e-05 0.0011542 0.15145 0.00065831 0.1521 0.13865 0 0.036907 0.0389 0 0.89978 0.25107 0.067471 0.0094157 4.2588 0.058796 7.0645e-05 0.83127 0.0052781 0.0060155 0.01227 0.23128 0.09522 3.2264e-05 0.00013083 0.13189 0.60631 0.65842 0.0046037 0.61131 0.47728 0.024749 0.42432 1.0553 1.0493 15.9963 144.9781 0.00055944 -72.2805 0.040718
1.1446 0.98803 5.5185e-05 3.8182 0.012035 1.5066e-05 0.0011542 0.15151 0.00065831 0.15216 0.13871 0 0.036903 0.0389 0 0.89984 0.2511 0.067482 0.0094171 4.2591 0.058805 7.0656e-05 0.83127 0.0052784 0.0060158 0.010951 0.25934 0.10548 2.8386e-05 0.00011497 0.1319 0.60716 0.65975 0.0043137 0.61218 0.4774 0.020061 0.42422 1.0574 1.0513 15.9963 144.9781 0.00055778 -72.9978 0.041603
1.1455 0.98803 5.5185e-05 3.8182 0.012035 1.5078e-05 0.0011542 0.15157 0.00065831 0.15222 0.13876 0 0.036899 0.0389 0 0.89991 0.25113 0.067493 0.0094184 4.2594 0.058813 7.0667e-05 0.83126 0.0052787 0.0060162 0.0098056 0.2893 0.11665 2.5084e-05 0.00010148 0.1319 0.60804 0.66106 0.0040515 0.61307 0.47752 0.016219 0.42413 1.0594 1.0534 15.9964 144.9781 0.00055612 -73.6908 0.042487
1.1464 0.98803 5.5185e-05 3.8182 0.012035 1.5089e-05 0.0011542 0.15162 0.00065831 0.15228 0.13882 0 0.036895 0.0389 0 0.89998 0.25116 0.067504 0.0094197 4.2597 0.058821 7.0677e-05 0.83125 0.0052791 0.0060165 0.008819 0.321 0.12878 2.2269e-05 9.0003e-05 0.1319 0.60892 0.66237 0.0038145 0.61398 0.47764 0.013128 0.42404 1.0615 1.0555 15.9964 144.9781 0.00055446 -74.3582 0.043372
1.1472 0.98803 5.5185e-05 3.8182 0.012035 1.51e-05 0.0011542 0.15168 0.00065831 0.15233 0.13887 0 0.036892 0.0389 0 0.90004 0.25119 0.067513 0.0094209 4.26 0.058828 7.0687e-05 0.83124 0.0052793 0.0060168 0.0080358 0.35089 0.14055 2.0089e-05 8.1123e-05 0.13191 0.60973 0.66354 0.0036209 0.61482 0.47775 0.010903 0.42396 1.0633 1.0573 15.9965 144.978 0.00055296 -74.9363 0.044168
1.1479 0.98803 5.5185e-05 3.8182 0.012035 1.5109e-05 0.0011542 0.15173 0.00065831 0.15238 0.13892 0 0.036889 0.0389 0 0.9001 0.25121 0.067522 0.009422 4.2602 0.058835 7.0695e-05 0.83124 0.0052796 0.006017 0.0074123 0.37872 0.15185 1.8371e-05 7.4135e-05 0.13191 0.61047 0.66458 0.0034612 0.61559 0.47785 0.0092862 0.4239 1.065 1.059 15.9965 144.978 0.00055162 -75.4377 0.044884
1.1486 0.98803 5.5185e-05 3.8182 0.012035 1.5117e-05 0.0011542 0.15177 0.00065831 0.15242 0.13896 0 0.036886 0.0389 0 0.90015 0.25124 0.06753 0.009423 4.2604 0.058841 7.0703e-05 0.83123 0.0052798 0.0060173 0.0069103 0.40441 0.1626 1.6999e-05 6.8557e-05 0.13191 0.61114 0.66551 0.0033283 0.6163 0.47794 0.0080979 0.42384 1.0665 1.0605 15.9966 144.978 0.00055041 -75.8732 0.045529
1.1492 0.98803 5.5185e-05 3.8182 0.012035 1.5126e-05 0.0011542 0.15181 0.00065832 0.15247 0.139 0 0.036883 0.0389 0 0.9002 0.25126 0.067538 0.009424 4.2607 0.058847 7.0711e-05 0.83122 0.0052801 0.0060175 0.0064585 0.43057 0.17391 1.5771e-05 6.3571e-05 0.13191 0.61181 0.66644 0.003205 0.61702 0.47803 0.0071244 0.42379 1.0679 1.062 15.9966 144.978 0.00054921 -76.2937 0.046174
1.1498 0.98803 5.5185e-05 3.8182 0.012035 1.5134e-05 0.0011542 0.15186 0.00065832 0.15251 0.13904 0 0.036881 0.0389 0 0.90025 0.25128 0.067546 0.009425 4.2609 0.058853 7.0718e-05 0.83122 0.0052803 0.0060178 0.0060488 0.45708 0.18575 1.4673e-05 5.9113e-05 0.13191 0.61249 0.66737 0.0030906 0.61776 0.47813 0.0063314 0.42374 1.0694 1.0635 15.9967 144.978 0.000548 -76.699 0.046819
1.1505 0.98803 5.5185e-05 3.8182 0.012035 1.5143e-05 0.0011542 0.1519 0.00065832 0.15255 0.13908 0 0.036878 0.0389 0 0.9003 0.2513 0.067554 0.0094259 4.2611 0.058859 7.0726e-05 0.83121 0.0052806 0.006018 0.0056776 0.4838 0.19812 1.3689e-05 5.512e-05 0.13192 0.61317 0.66828 0.0029845 0.61852 0.47822 0.0056881 0.42369 1.0709 1.065 15.9967 144.978 0.0005468 -77.0888 0.047464
1.1511 0.98803 5.5185e-05 3.8182 0.012035 1.5151e-05 0.0011542 0.15194 0.00065832 0.1526 0.13912 0 0.036875 0.0389 0 0.90035 0.25132 0.067562 0.0094269 4.2613 0.058865 7.0734e-05 0.83121 0.0052808 0.0060182 0.0053441 0.51058 0.21099 1.2805e-05 5.154e-05 0.13192 0.61386 0.6692 0.0028862 0.61928 0.47831 0.0051674 0.42364 1.0724 1.0665 15.9968 144.9779 0.0005456 -77.4632 0.048109
1.1518 0.98803 5.5185e-05 3.8182 0.012035 1.516e-05 0.0011542 0.15199 0.00065832 0.15264 0.13916 0 0.036872 0.0389 0 0.9004 0.25135 0.06757 0.0094279 4.2616 0.058871 7.0741e-05 0.8312 0.005281 0.0060185 0.0050408 0.53728 0.22435 1.2012e-05 4.8328e-05 0.13192 0.61454 0.67011 0.002795 0.62007 0.47841 0.0047462 0.4236 1.0739 1.068 15.9968 144.9779 0.0005444 -77.8222 0.048754
1.1524 0.98803 5.5185e-05 3.8182 0.012035 1.5168e-05 0.0011542 0.15203 0.00065832 0.15268 0.1392 0 0.036869 0.0389 0 0.90045 0.25137 0.067578 0.0094289 4.2618 0.058877 7.0749e-05 0.83119 0.0052813 0.0060187 0.0047666 0.56375 0.23815 1.13e-05 4.5442e-05 0.13192 0.61523 0.67101 0.0027104 0.62087 0.4785 0.0044049 0.42355 1.0754 1.0695 15.9969 144.9779 0.00054321 -78.1658 0.049399
1.1531 0.98803 5.5185e-05 3.8182 0.012035 1.5177e-05 0.0011542 0.15207 0.00065832 0.15273 0.13924 0 0.036867 0.0389 0 0.90049 0.25139 0.067586 0.0094298 4.262 0.058883 7.0757e-05 0.83119 0.0052815 0.006019 0.0045184 0.58985 0.25237 1.0658e-05 4.2845e-05 0.13192 0.61593 0.67191 0.0026321 0.62169 0.4786 0.004127 0.42351 1.0769 1.071 15.9969 144.9779 0.00054201 -78.4942 0.050043
1.1537 0.98803 5.5185e-05 3.8182 0.012035 1.5185e-05 0.0011542 0.15212 0.00065832 0.15277 0.13928 0 0.036864 0.0389 0 0.90054 0.25141 0.067594 0.0094308 4.2623 0.058889 7.0764e-05 0.83118 0.0052817 0.0060192 0.0042934 0.61544 0.26696 1.008e-05 4.0506e-05 0.13192 0.61662 0.67281 0.0025595 0.62252 0.47869 0.0038991 0.42347 1.0783 1.0725 15.997 144.9779 0.00054082 -78.8076 0.050688
1.1544 0.98803 5.5185e-05 3.8182 0.012035 1.5194e-05 0.0011542 0.15216 0.00065832 0.15281 0.13932 0 0.036861 0.0389 0 0.90059 0.25144 0.067602 0.0094318 4.2625 0.058895 7.0772e-05 0.83118 0.005282 0.0060194 0.0040889 0.6404 0.28188 9.5579e-06 3.8397e-05 0.13193 0.61732 0.6737 0.0024922 0.62337 0.47879 0.0037106 0.42344 1.0798 1.074 15.997 144.9779 0.00053963 -79.1061 0.051333
1.155 0.98803 5.5185e-05 3.8182 0.012035 1.5202e-05 0.0011542 0.1522 0.00065832 0.15286 0.13936 0 0.036858 0.0389 0 0.90064 0.25146 0.06761 0.0094328 4.2627 0.058901 7.078e-05 0.83117 0.0052822 0.0060197 0.0039035 0.66462 0.29709 9.0868e-06 3.6493e-05 0.13193 0.61802 0.67458 0.0024299 0.62424 0.47889 0.0035529 0.4234 1.0813 1.0755 15.9971 144.9779 0.00053844 -79.3901 0.051978
1.1556 0.98803 5.5184e-05 3.8182 0.012035 1.5211e-05 0.0011542 0.15225 0.00065832 0.1529 0.1394 0 0.036856 0.0389 0 0.90069 0.25148 0.067618 0.0094337 4.2629 0.058907 7.0788e-05 0.83116 0.0052825 0.0060199 0.0037343 0.688 0.31253 8.6606e-06 3.4772e-05 0.13193 0.61871 0.67546 0.0023722 0.62513 0.47899 0.0034195 0.42337 1.0828 1.077 15.9971 144.9779 0.00053725 -79.66 0.052623
1.1563 0.98803 5.5184e-05 3.8182 0.012035 1.5219e-05 0.0011542 0.15229 0.00065832 0.15294 0.13944 0 0.036853 0.0389 0 0.90074 0.2515 0.067626 0.0094347 4.2632 0.058913 7.0795e-05 0.83116 0.0052827 0.0060202 0.0035822 0.71043 0.32815 8.2751e-06 3.3215e-05 0.13193 0.61941 0.67634 0.0023187 0.62603 0.47909 0.0033052 0.42334 1.0842 1.0785 15.9972 144.9778 0.00053607 -79.916 0.053268
1.1569 0.98803 5.5184e-05 3.8182 0.012035 1.5228e-05 0.0011542 0.15233 0.00065833 0.15299 0.13948 0 0.03685 0.0389 0 0.90079 0.25152 0.067634 0.0094357 4.2634 0.058919 7.0803e-05 0.83115 0.0052829 0.0060204 0.0034393 0.73186 0.34392 7.9251e-06 3.1803e-05 0.13193 0.62011 0.67721 0.0022692 0.62694 0.47918 0.003206 0.42331 1.0857 1.0799 15.9972 144.9778 0.00053489 -80.1587 0.053913
1.1576 0.98803 5.5184e-05 3.8182 0.012035 1.5236e-05 0.0011542 0.15237 0.00065833 0.15303 0.13952 0 0.036847 0.0389 0 0.90084 0.25155 0.067642 0.0094367 4.2636 0.058925 7.0811e-05 0.83115 0.0052832 0.0060206 0.0033148 0.75223 0.35978 7.608e-06 3.0523e-05 0.13194 0.62082 0.67808 0.0022232 0.62787 0.47928 0.0031192 0.42328 1.0872 1.0814 15.9973 144.9778 0.00053371 -80.3884 0.054558
1.1582 0.98803 5.5184e-05 3.8182 0.012035 1.5244e-05 0.0011542 0.15241 0.00065833 0.15307 0.13956 0 0.036845 0.0389 0 0.90089 0.25157 0.067649 0.0094375 4.2638 0.05893 7.0818e-05 0.83114 0.0052834 0.0060209 0.003209 0.76963 0.3741 7.3473e-06 2.9472e-05 0.13194 0.62145 0.67885 0.0021848 0.62872 0.47937 0.0030496 0.42326 1.0885 1.0828 15.9973 144.9778 0.00053266 -80.5844 0.055138
1.1587 0.98803 5.5184e-05 3.8182 0.012035 1.5251e-05 0.0011542 0.15245 0.00065833 0.1531 0.13959 0 0.036843 0.0389 0 0.90093 0.25158 0.067656 0.0094383 4.264 0.058935 7.0824e-05 0.83114 0.0052836 0.006021 0.0031213 0.7845 0.387 7.131e-06 2.8599e-05 0.13194 0.62202 0.67955 0.0021524 0.6295 0.47946 0.0029927 0.42323 1.0897 1.084 15.9974 144.9778 0.00053171 -80.7524 0.05566
1.1592 0.98803 5.5184e-05 3.8182 0.012035 1.5257e-05 0.0011542 0.15248 0.00065833 0.15314 0.13962 0 0.036841 0.0389 0 0.90097 0.2516 0.067662 0.0094391 4.2642 0.05894 7.083e-05 0.83113 0.0052838 0.0060212 0.0030401 0.79863 0.39988 6.9305e-06 2.7791e-05 0.13194 0.62258 0.68024 0.002122 0.63028 0.47954 0.0029405 0.42321 1.0909 1.0852 15.9974 144.9778 0.00053076 -80.9127 0.056183
1.1597 0.98803 5.5184e-05 3.8182 0.012035 1.5264e-05 0.0011542 0.15252 0.00065833 0.15317 0.13966 0 0.036838 0.0389 0 0.90101 0.25162 0.067669 0.0094399 4.2644 0.058945 7.0837e-05 0.83113 0.005284 0.0060214 0.0029651 0.81201 0.41273 6.7445e-06 2.7041e-05 0.13194 0.62315 0.68093 0.0020933 0.63107 0.47962 0.0028924 0.4232 1.0921 1.0864 15.9975 144.9778 0.00052982 -81.0657 0.056705
1.1603 0.98803 5.5184e-05 3.8182 0.012035 1.5271e-05 0.0011542 0.15255 0.00065833 0.15321 0.13969 0 0.036836 0.0389 0 0.90105 0.25164 0.067675 0.0094407 4.2646 0.05895 7.0843e-05 0.83112 0.0052842 0.0060216 0.0028944 0.82465 0.42553 6.572e-06 2.6346e-05 0.13195 0.62372 0.68162 0.0020664 0.63188 0.4797 0.0028479 0.42318 1.0933 1.0876 15.9975 144.9778 0.00052887 -81.2115 0.057227
1.1608 0.98803 5.5184e-05 3.8182 0.012035 1.5278e-05 0.0011542 0.15259 0.00065833 0.15324 0.13972 0 0.036834 0.0389 0 0.90109 0.25166 0.067682 0.0094415 4.2647 0.058955 7.0849e-05 0.83112 0.0052844 0.0060218 0.0028304 0.83655 0.43825 6.4114e-06 2.5699e-05 0.13195 0.62429 0.68231 0.002041 0.63269 0.47979 0.0028067 0.42316 1.0945 1.0888 15.9976 144.9778 0.00052793 -81.3504 0.05775
1.1613 0.98803 5.5184e-05 3.8182 0.012035 1.5285e-05 0.0011542 0.15262 0.00065833 0.15328 0.13975 0 0.036832 0.0389 0 0.90113 0.25167 0.067688 0.0094423 4.2649 0.05896 7.0855e-05 0.83111 0.0052845 0.006022 0.0027691 0.84774 0.45088 6.2623e-06 2.5099e-05 0.13195 0.62486 0.68299 0.0020172 0.6335 0.47987 0.0027684 0.42314 1.0956 1.09 15.9976 144.9778 0.00052699 -81.4827 0.058272
1.1618 0.98803 5.5184e-05 3.8182 0.012035 1.5292e-05 0.0011542 0.15266 0.00065833 0.15331 0.13979 0 0.036829 0.0389 0 0.90117 0.25169 0.067695 0.0094431 4.2651 0.058964 7.0862e-05 0.83111 0.0052847 0.0060222 0.0027109 0.85822 0.46342 6.1238e-06 2.454e-05 0.13195 0.62543 0.68367 0.0019948 0.63433 0.47995 0.0027328 0.42313 1.0968 1.0912 15.9977 144.9778 0.00052605 -81.6086 0.058794
1.1623 0.98803 5.5184e-05 3.8182 0.012035 1.5299e-05 0.0011542 0.15269 0.00065833 0.15335 0.13982 0 0.036827 0.0389 0 0.90121 0.25171 0.067701 0.0094439 4.2653 0.058969 7.0868e-05 0.8311 0.0052849 0.0060224 0.0026592 0.86802 0.47583 5.9947e-06 2.402e-05 0.13195 0.62599 0.68434 0.0019737 0.63516 0.48004 0.0026995 0.42311 1.098 1.0923 15.9977 144.9778 0.00052512 -81.7284 0.059317
1.1629 0.98803 5.5184e-05 3.8182 0.012035 1.5305e-05 0.0011542 0.15273 0.00065833 0.15338 0.13985 0 0.036825 0.0389 0 0.90125 0.25173 0.067708 0.0094447 4.2655 0.058974 7.0874e-05 0.8311 0.0052851 0.0060226 0.0026099 0.87716 0.48811 5.8744e-06 2.3536e-05 0.13195 0.62656 0.68502 0.0019538 0.636 0.48012 0.0026685 0.4231 1.0992 1.0935 15.9977 144.9778 0.00052419 -81.8424 0.059839
1.1634 0.98803 5.5184e-05 3.8182 0.012035 1.5312e-05 0.0011542 0.15276 0.00065833 0.15341 0.13988 0 0.036823 0.0389 0 0.90129 0.25175 0.067714 0.0094455 4.2657 0.058979 7.088e-05 0.83109 0.0052853 0.0060228 0.0025616 0.88567 0.50025 5.7624e-06 2.3085e-05 0.13195 0.62713 0.68569 0.0019351 0.63684 0.4802 0.0026394 0.42308 1.1004 1.0947 15.9978 144.9778 0.00052326 -81.9507 0.060361
1.1639 0.98803 5.5184e-05 3.8182 0.012035 1.5319e-05 0.0011542 0.1528 0.00065833 0.15345 0.13992 0 0.036821 0.0389 0 0.90133 0.25176 0.067721 0.0094463 4.2659 0.058984 7.0887e-05 0.83109 0.0052855 0.006023 0.0025203 0.89357 0.51223 5.6578e-06 2.2664e-05 0.13196 0.6277 0.68636 0.0019175 0.6377 0.48029 0.0026123 0.42307 1.1016 1.0959 15.9978 144.9778 0.00052233 -82.0538 0.060884
1.1644 0.98803 5.5184e-05 3.8182 0.012034 1.5326e-05 0.0011542 0.15283 0.00065833 0.15348 0.13995 0 0.036818 0.0389 0 0.90137 0.25178 0.067727 0.0094471 4.266 0.058989 7.0893e-05 0.83108 0.0052857 0.0060232 0.0024785 0.90089 0.52405 5.5602e-06 2.2271e-05 0.13196 0.62826 0.68702 0.001901 0.63855 0.48037 0.0025868 0.42306 1.1027 1.0971 15.9979 144.9778 0.0005214 -82.1517 0.061406
1.165 0.98803 5.5184e-05 3.8182 0.012034 1.5333e-05 0.0011542 0.15286 0.00065833 0.15352 0.13998 0 0.036816 0.0389 0 0.90141 0.2518 0.067734 0.0094479 4.2662 0.058994 7.0899e-05 0.83108 0.0052859 0.0060234 0.002442 0.90767 0.5357 5.469e-06 2.1904e-05 0.13196 0.62883 0.68768 0.0018854 0.63942 0.48046 0.002563 0.42305 1.1039 1.0983 15.9979 144.9778 0.00052048 -82.2447 0.061928
1.1654 0.98803 5.5184e-05 3.8182 0.012034 1.5339e-05 0.0011542 0.1529 0.00065834 0.15355 0.14001 0 0.036814 0.0389 0 0.90145 0.25182 0.067739 0.0094486 4.2664 0.058998 7.0905e-05 0.83107 0.0052861 0.0060236 0.0024089 0.91333 0.54603 5.3921e-06 2.1595e-05 0.13196 0.62934 0.68828 0.0018721 0.6402 0.48053 0.0025428 0.42304 1.105 1.0994 15.998 144.9778 0.00051965 -82.3244 0.062399
1.1659 0.98803 5.5184e-05 3.8182 0.012034 1.5345e-05 0.0011542 0.15293 0.00065834 0.15358 0.14004 0 0.036812 0.0389 0 0.90149 0.25183 0.067745 0.0094493 4.2666 0.059002 7.0911e-05 0.83107 0.0052863 0.0060238 0.0023795 0.91858 0.55621 5.3196e-06 2.1303e-05 0.13196 0.62985 0.68887 0.0018595 0.64098 0.48061 0.0025237 0.42303 1.106 1.1004 15.998 144.9778 0.00051882 -82.4005 0.062869
1.1664 0.98803 5.5184e-05 3.8182 0.012034 1.5351e-05 0.0011542 0.15296 0.00065834 0.15361 0.14007 0 0.03681 0.0389 0 0.90152 0.25185 0.067751 0.00945 4.2667 0.059007 7.0916e-05 0.83106 0.0052864 0.0060239 0.0023517 0.92346 0.56623 5.2513e-06 2.1028e-05 0.13196 0.63036 0.68946 0.0018476 0.64177 0.48069 0.0025056 0.42302 1.1071 1.1015 15.9981 144.9778 0.000518 -82.4732 0.063339
1.1668 0.98803 5.5184e-05 3.8182 0.012034 1.5358e-05 0.0011542 0.15299 0.00065834 0.15364 0.1401 0 0.036808 0.0389 0 0.90156 0.25186 0.067757 0.0094507 4.2669 0.059011 7.0922e-05 0.83106 0.0052866 0.0060241 0.0023241 0.92799 0.5761 5.187e-06 2.077e-05 0.13197 0.63086 0.69005 0.0018362 0.64257 0.48076 0.0024886 0.42301 1.1082 1.1026 15.9981 144.9778 0.00051717 -82.5426 0.063809
1.1675 0.98803 5.5184e-05 3.8182 0.012034 1.5366e-05 0.0011542 0.15303 0.00065834 0.15369 0.14014 0 0.036805 0.0389 0 0.90161 0.25189 0.067765 0.0094517 4.2671 0.059017 7.093e-05 0.83105 0.0052869 0.0060244 0.0022885 0.93379 0.58969 5.1027e-06 2.043e-05 0.13197 0.63158 0.69087 0.0018213 0.64368 0.48087 0.0024662 0.42299 1.1096 1.1041 15.9982 144.9778 0.00051602 -82.6348 0.06447
1.1682 0.98803 5.5184e-05 3.8182 0.012034 1.5375e-05 0.0011542 0.15308 0.00065834 0.15373 0.14018 0 0.036803 0.0389 0 0.90166 0.25191 0.067773 0.0094527 4.2674 0.059024 7.0938e-05 0.83105 0.0052871 0.0060246 0.0022569 0.93899 0.60297 5.025e-06 2.0118e-05 0.13197 0.63229 0.69169 0.0018074 0.64481 0.48098 0.0024454 0.42298 1.1111 1.1056 15.9982 144.9778 0.00051487 -82.7211 0.06513
1.1688 0.98803 5.5184e-05 3.8182 0.012034 1.5384e-05 0.0011542 0.15312 0.00065834 0.15377 0.14022 0 0.0368 0.0389 0 0.90171 0.25193 0.067782 0.0094537 4.2676 0.05903 7.0946e-05 0.83104 0.0052874 0.0060249 0.0022268 0.94363 0.61591 4.9532e-06 1.983e-05 0.13197 0.633 0.6925 0.0017945 0.64594 0.48109 0.0024262 0.42297 1.1126 1.1071 15.9983 144.9778 0.00051372 -82.802 0.065791
1.1695 0.98803 5.5184e-05 3.8182 0.012034 1.5392e-05 0.0011542 0.15316 0.00065834 0.15382 0.14026 0 0.036797 0.0389 0 0.90177 0.25196 0.06779 0.0094547 4.2679 0.059036 7.0954e-05 0.83104 0.0052876 0.0060251 0.002198 0.94778 0.62852 4.887e-06 1.9563e-05 0.13197 0.63371 0.69331 0.0017825 0.64708 0.4812 0.0024084 0.42296 1.1141 1.1086 15.9983 144.9778 0.00051258 -82.8778 0.066452
1.1701 0.98803 5.5184e-05 3.8182 0.012034 1.5401e-05 0.0011542 0.15321 0.00065834 0.15386 0.1403 0 0.036794 0.0389 0 0.90182 0.25198 0.067798 0.0094557 4.2681 0.059042 7.0962e-05 0.83103 0.0052878 0.0060254 0.0021724 0.95148 0.64079 4.8258e-06 1.9317e-05 0.13198 0.63442 0.69412 0.0017714 0.64822 0.48131 0.0023919 0.42295 1.1156 1.11 15.9984 144.9778 0.00051144 -82.9488 0.067112
1.1708 0.98803 5.5184e-05 3.8182 0.012034 1.541e-05 0.0011542 0.15325 0.00065834 0.15391 0.14034 0 0.036791 0.0389 0 0.90187 0.252 0.067806 0.0094568 4.2683 0.059048 7.097e-05 0.83102 0.0052881 0.0060256 0.0021492 0.95477 0.65273 4.769e-06 1.9089e-05 0.13198 0.63513 0.69492 0.001761 0.64936 0.48142 0.0023765 0.42294 1.117 1.1115 15.9985 144.9778 0.0005103 -83.0153 0.067773
1.1715 0.98803 5.5183e-05 3.8182 0.012034 1.5418e-05 0.0011542 0.15329 0.00065834 0.15395 0.14038 0 0.036789 0.0389 0 0.90192 0.25202 0.067814 0.0094578 4.2686 0.059054 7.0978e-05 0.83102 0.0052883 0.0060259 0.0021264 0.95769 0.66434 4.7165e-06 1.8878e-05 0.13198 0.63584 0.69572 0.0017513 0.65051 0.48153 0.0023623 0.42293 1.1185 1.113 15.9985 144.9778 0.00050917 -83.0777 0.068434
1.1721 0.98803 5.5183e-05 3.8182 0.012034 1.5427e-05 0.0011542 0.15334 0.00065834 0.15399 0.14042 0 0.036786 0.0389 0 0.90197 0.25205 0.067823 0.0094588 4.2688 0.059061 7.0985e-05 0.83101 0.0052886 0.0060261 0.0021054 0.96029 0.67561 4.6678e-06 1.8682e-05 0.13198 0.63654 0.69651 0.0017422 0.65166 0.48164 0.002349 0.42292 1.12 1.1145 15.9986 144.9778 0.00050804 -83.1362 0.069094
1.1728 0.98803 5.5183e-05 3.8182 0.012034 1.5436e-05 0.0011542 0.15338 0.00065834 0.15404 0.14047 0 0.036783 0.0389 0 0.90202 0.25207 0.067831 0.0094598 4.269 0.059067 7.0993e-05 0.831 0.0052888 0.0060264 0.0020878 0.96259 0.68655 4.6224e-06 1.85e-05 0.13198 0.63725 0.6973 0.0017338 0.65281 0.48175 0.0023367 0.42291 1.1215 1.116 15.9986 144.9778 0.00050692 -83.1911 0.069755
1.1734 0.98803 5.5183e-05 3.8182 0.012034 1.5444e-05 0.0011542 0.15343 0.00065835 0.15408 0.14051 0 0.03678 0.0389 0 0.90207 0.25209 0.067839 0.0094608 4.2693 0.059073 7.1001e-05 0.831 0.0052891 0.0060266 0.0020708 0.96463 0.69717 4.5803e-06 1.8331e-05 0.13199 0.63795 0.69809 0.0017259 0.65396 0.48186 0.0023252 0.42291 1.1229 1.1175 15.9987 144.9778 0.0005058 -83.2426 0.070416
1.1741 0.98803 5.5183e-05 3.8182 0.012034 1.5453e-05 0.0011542 0.15347 0.00065835 0.15412 0.14055 0 0.036778 0.0389 0 0.90213 0.25212 0.067847 0.0094618 4.2695 0.059079 7.1009e-05 0.83099 0.0052893 0.0060269 0.0020519 0.96644 0.70747 4.5412e-06 1.8173e-05 0.13199 0.63865 0.69887 0.0017186 0.65512 0.48197 0.0023144 0.4229 1.1244 1.119 15.9988 144.9778 0.00050468 -83.291 0.071076
1.1748 0.98803 5.5183e-05 3.8182 0.012034 1.5462e-05 0.0011542 0.15351 0.00065835 0.15417 0.14059 0 0.036775 0.0389 0 0.90218 0.25214 0.067856 0.0094628 4.2698 0.059085 7.1017e-05 0.83099 0.0052896 0.0060271 0.0020374 0.96804 0.71744 4.5047e-06 1.8027e-05 0.13199 0.63935 0.69965 0.0017117 0.65628 0.48208 0.0023044 0.42289 1.1259 1.1204 15.9988 144.9778 0.00050357 -83.3364 0.071737
1.1754 0.98803 5.5183e-05 3.8182 0.012034 1.547e-05 0.0011542 0.15356 0.00065835 0.15421 0.14063 0 0.036772 0.0389 0 0.90223 0.25216 0.067864 0.0094638 4.27 0.059092 7.1025e-05 0.83098 0.0052898 0.0060274 0.0020244 0.96946 0.72711 4.4706e-06 1.789e-05 0.13199 0.64005 0.70043 0.0017052 0.65744 0.48219 0.0022951 0.42288 1.1273 1.1219 15.9989 144.9778 0.00050246 -83.3791 0.072398
1.1761 0.98803 5.5183e-05 3.8182 0.012034 1.5479e-05 0.0011542 0.1536 0.00065835 0.15425 0.14067 0 0.036769 0.0389 0 0.90228 0.25218 0.067872 0.0094648 4.2702 0.059098 7.1033e-05 0.83097 0.0052901 0.0060276 0.0020098 0.97072 0.73647 4.4388e-06 1.7762e-05 0.13199 0.64075 0.7012 0.0016992 0.6586 0.4823 0.0022864 0.42288 1.1288 1.1234 15.9989 144.9778 0.00050136 -83.4193 0.073059
1.1767 0.98803 5.5183e-05 3.8182 0.012034 1.5488e-05 0.0011542 0.15364 0.00065835 0.1543 0.14071 0 0.036767 0.0389 0 0.90233 0.25221 0.06788 0.0094658 4.2705 0.059104 7.1041e-05 0.83097 0.0052903 0.0060279 0.0019964 0.97183 0.74553 4.4091e-06 1.7643e-05 0.132 0.64145 0.70197 0.0016935 0.65976 0.48241 0.0022782 0.42287 1.1303 1.1249 15.999 144.9778 0.00050026 -83.4572 0.073719
1.1774 0.98803 5.5183e-05 3.8182 0.012034 1.5496e-05 0.0011542 0.15369 0.00065835 0.15434 0.14075 0 0.036764 0.0389 0 0.90238 0.25223 0.067889 0.0094668 4.2707 0.05911 7.1049e-05 0.83096 0.0052906 0.0060281 0.0019856 0.97281 0.75429 4.3812e-06 1.7531e-05 0.132 0.64215 0.70273 0.0016882 0.66092 0.48252 0.0022705 0.42286 1.1317 1.1264 15.9991 144.9778 0.00049916 -83.4929 0.07438
1.1781 0.98803 5.5183e-05 3.8182 0.012034 1.5505e-05 0.0011542 0.15373 0.00065835 0.15438 0.14079 0 0.036761 0.0389 0 0.90243 0.25225 0.067897 0.0094678 4.2709 0.059116 7.1057e-05 0.83095 0.0052908 0.0060284 0.0019748 0.97369 0.76277 4.3551e-06 1.7426e-05 0.132 0.64284 0.70349 0.0016832 0.66208 0.48263 0.0022634 0.42286 1.1332 1.1278 15.9991 144.9778 0.00049807 -83.5265 0.075041
1.1787 0.98803 5.5183e-05 3.8182 0.012034 1.5514e-05 0.0011542 0.15377 0.00065835 0.15443 0.14083 0 0.036758 0.0389 0 0.90249 0.25228 0.067905 0.0094688 4.2712 0.059123 7.1065e-05 0.83095 0.0052911 0.0060286 0.0019638 0.97446 0.77097 4.3307e-06 1.7328e-05 0.132 0.64354 0.70424 0.0016785 0.66324 0.48274 0.0022566 0.42285 1.1347 1.1293 15.9992 144.9778 0.00049698 -83.5583 0.075701
1.1794 0.98803 5.5183e-05 3.8182 0.012034 1.5523e-05 0.0011542 0.15382 0.00065835 0.15447 0.14087 0 0.036755 0.0389 0 0.90254 0.2523 0.067913 0.0094699 4.2714 0.059129 7.1073e-05 0.83094 0.0052913 0.0060289 0.0019542 0.97515 0.77889 4.3076e-06 1.7235e-05 0.132 0.64423 0.705 0.001674 0.6644 0.48286 0.0022503 0.42285 1.1361 1.1308 15.9992 144.9778 0.0004959 -83.5883 0.076362
1.1804 0.98803 5.5183e-05 3.8182 0.012034 1.5536e-05 0.0011542 0.15388 0.00065835 0.15454 0.14093 0 0.036751 0.0389 0 0.90262 0.25233 0.067926 0.0094714 4.2718 0.059138 7.1085e-05 0.83093 0.0052917 0.0060293 0.0019405 0.97605 0.79038 4.2753e-06 1.7106e-05 0.13201 0.64528 0.70613 0.0016678 0.66615 0.48302 0.0022414 0.42284 1.1383 1.133 15.9993 144.9778 0.00049426 -83.6307 0.077362
1.1814 0.98803 5.5183e-05 3.8182 0.012034 1.5549e-05 0.0011542 0.15395 0.00065835 0.1546 0.14099 0 0.036747 0.0389 0 0.90269 0.25237 0.067938 0.0094729 4.2722 0.059148 7.1097e-05 0.83092 0.0052921 0.0060296 0.0019279 0.9768 0.80128 4.2458e-06 1.6987e-05 0.13201 0.64632 0.70725 0.001662 0.6679 0.48319 0.0022332 0.42283 1.1405 1.1352 15.9994 144.9778 0.00049264 -83.6698 0.078362
1.1824 0.98803 5.5183e-05 3.8182 0.012034 1.5562e-05 0.0011542 0.15401 0.00065836 0.15467 0.14106 0 0.036743 0.0389 0 0.90277 0.2524 0.067951 0.0094744 4.2725 0.059157 7.1109e-05 0.83091 0.0052925 0.00603 0.0019164 0.97743 0.81162 4.2187e-06 1.6878e-05 0.13201 0.64736 0.70837 0.0016567 0.66965 0.48336 0.0022258 0.42283 1.1427 1.1374 15.9995 144.9778 0.00049102 -83.7059 0.079362
1.1834 0.98803 5.5183e-05 3.8182 0.012034 1.5575e-05 0.0011542 0.15408 0.00065836 0.15473 0.14112 0 0.036739 0.0389 0 0.90285 0.25244 0.067963 0.009476 4.2729 0.059166 7.1122e-05 0.8309 0.0052928 0.0060304 0.0019058 0.97796 0.82142 4.1937e-06 1.6778e-05 0.13202 0.6484 0.70948 0.0016519 0.6714 0.48353 0.0022189 0.42282 1.1449 1.1396 15.9996 144.9778 0.00048941 -83.7394 0.080362
1.1844 0.98803 5.5183e-05 3.8182 0.012034 1.5588e-05 0.0011542 0.15414 0.00065836 0.1548 0.14118 0 0.036735 0.0389 0 0.90293 0.25247 0.067976 0.0094775 4.2733 0.059176 7.1134e-05 0.8309 0.0052932 0.0060308 0.0018961 0.97842 0.8307 4.1706e-06 1.6686e-05 0.13202 0.64943 0.71058 0.0016473 0.67314 0.4837 0.0022126 0.42281 1.1471 1.1418 15.9997 144.9778 0.00048781 -83.7705 0.081362
1.1854 0.98803 5.5183e-05 3.8182 0.012034 1.5601e-05 0.0011542 0.15421 0.00065836 0.15486 0.14124 0 0.036731 0.0389 0 0.90301 0.25251 0.067989 0.009479 4.2736 0.059185 7.1146e-05 0.83089 0.0052936 0.0060312 0.0018868 0.9788 0.8395 4.1492e-06 1.66e-05 0.13202 0.65046 0.71167 0.0016431 0.67488 0.48387 0.0022067 0.42281 1.1493 1.144 15.9997 144.9778 0.00048622 -83.7995 0.082362
1.1864 0.98803 5.5183e-05 3.8182 0.012034 1.5614e-05 0.0011542 0.15427 0.00065836 0.15493 0.1413 0 0.036726 0.0389 0 0.90308 0.25254 0.068001 0.0094806 4.274 0.059195 7.1158e-05 0.83088 0.005294 0.0060316 0.0018784 0.97914 0.84783 4.1293e-06 1.652e-05 0.13203 0.65149 0.71275 0.0016392 0.67661 0.48404 0.0022013 0.4228 1.1514 1.1462 15.9998 144.9778 0.00048464 -83.8266 0.083362
1.1874 0.98803 5.5182e-05 3.8182 0.012034 1.5628e-05 0.0011542 0.15434 0.00065836 0.15499 0.14136 0 0.036722 0.0389 0 0.90316 0.25258 0.068014 0.0094821 4.2743 0.059204 7.117e-05 0.83087 0.0052944 0.0060319 0.0018704 0.97942 0.85571 4.1107e-06 1.6445e-05 0.13203 0.65252 0.71383 0.0016355 0.67834 0.48421 0.0021962 0.4228 1.1536 1.1484 15.9999 144.9779 0.00048306 -83.852 0.084362
1.1884 0.98803 5.5182e-05 3.8182 0.012034 1.5641e-05 0.0011542 0.1544 0.00065836 0.15506 0.14142 0 0.036718 0.0389 0 0.90324 0.25261 0.068026 0.0094836 4.2747 0.059213 7.1182e-05 0.83086 0.0052948 0.0060323 0.0018632 0.97967 0.86317 4.0933e-06 1.6376e-05 0.13203 0.65354 0.7149 0.0016321 0.68007 0.48438 0.0021914 0.42279 1.1558 1.1506 16 144.9779 0.0004815 -83.876 0.085362
1.1894 0.98803 5.5182e-05 3.8182 0.012034 1.5654e-05 0.0011542 0.15447 0.00065836 0.15512 0.14148 0 0.036714 0.0389 0 0.90332 0.25265 0.068039 0.0094852 4.2751 0.059223 7.1194e-05 0.83085 0.0052951 0.0060327 0.001856 0.97989 0.87022 4.077e-06 1.631e-05 0.13204 0.65456 0.71596 0.0016289 0.68178 0.48455 0.002187 0.42279 1.158 1.1528 16.0001 144.9779 0.00047994 -83.8985 0.086362
1.1904 0.98803 5.5182e-05 3.8182 0.012034 1.5667e-05 0.0011542 0.15453 0.00065837 0.15519 0.14154 0 0.03671 0.0389 0 0.9034 0.25268 0.068051 0.0094867 4.2755 0.059232 7.1206e-05 0.83084 0.0052955 0.0060331 0.0018498 0.98008 0.8769 4.0615e-06 1.6248e-05 0.13204 0.65558 0.71701 0.0016258 0.6835 0.48472 0.0021828 0.42278 1.1601 1.155 16.0002 144.9779 0.0004784 -83.9199 0.087362
1.1914 0.98803 5.5182e-05 3.8182 0.012034 1.568e-05 0.0011542 0.1546 0.00065837 0.15525 0.1416 0 0.036706 0.0389 0 0.90348 0.25272 0.068064 0.0094882 4.2758 0.059242 7.1219e-05 0.83083 0.0052959 0.0060335 0.001843 0.98025 0.88321 4.047e-06 1.619e-05 0.13204 0.65659 0.71806 0.0016229 0.6852 0.48489 0.0021788 0.42278 1.1623 1.1572 16.0003 144.9779 0.00047686 -83.9402 0.088362
1.1924 0.98803 5.5182e-05 3.8182 0.012034 1.5693e-05 0.0011542 0.15466 0.00065837 0.15532 0.14167 0 0.036702 0.0389 0 0.90355 0.25275 0.068076 0.0094898 4.2762 0.059251 7.1231e-05 0.83082 0.0052963 0.0060339 0.0018373 0.9804 0.88917 4.0331e-06 1.6134e-05 0.13205 0.6576 0.7191 0.0016202 0.68691 0.48505 0.002175 0.42278 1.1644 1.1593 16.0003 144.9779 0.00047532 -83.9595 0.089362
1.1934 0.98803 5.5182e-05 3.8182 0.012034 1.5706e-05 0.0011542 0.15473 0.00065837 0.15538 0.14173 0 0.036697 0.0389 0 0.90363 0.25278 0.068089 0.0094913 4.2766 0.059261 7.1243e-05 0.83081 0.0052967 0.0060343 0.0018314 0.98053 0.89481 4.02e-06 1.6082e-05 0.13205 0.65861 0.72013 0.0016175 0.6886 0.48522 0.0021715 0.42277 1.1666 1.1615 16.0004 144.9779 0.0004738 -83.978 0.090362
1.1944 0.98803 5.5182e-05 3.8182 0.012034 1.572e-05 0.0011542 0.15479 0.00065837 0.15545 0.14179 0 0.036693 0.0389 0 0.90371 0.25282 0.068102 0.0094928 4.2769 0.05927 7.1255e-05 0.8308 0.005297 0.0060346 0.0018269 0.98065 0.90014 4.0074e-06 1.6031e-05 0.13205 0.65961 0.72116 0.001615 0.69029 0.48539 0.0021681 0.42277 1.1687 1.1637 16.0005 144.9779 0.00047229 -83.9956 0.091362
1.1954 0.98803 5.5182e-05 3.8182 0.012034 1.5733e-05 0.0011542 0.15486 0.00065837 0.15551 0.14185 0 0.036689 0.0389 0 0.90379 0.25285 0.068114 0.0094944 4.2773 0.05928 7.1267e-05 0.83079 0.0052974 0.006035 0.0018206 0.98077 0.90517 3.9954e-06 1.5983e-05 0.13206 0.66061 0.72218 0.0016126 0.69197 0.48556 0.0021648 0.42277 1.1709 1.1658 16.0006 144.9779 0.00047078 -84.0126 0.092362
1.1964 0.98803 5.5182e-05 3.8182 0.012034 1.5746e-05 0.0011542 0.15492 0.00065837 0.15558 0.14191 0 0.036685 0.0389 0 0.90387 0.25289 0.068127 0.0094959 4.2777 0.059289 7.1279e-05 0.83078 0.0052978 0.0060354 0.0018175 0.98087 0.90993 3.9838e-06 1.5937e-05 0.13206 0.66161 0.72319 0.0016103 0.69365 0.48573 0.0021617 0.42276 1.173 1.168 16.0007 144.9779 0.00046928 -84.0289 0.093362
1.1974 0.98803 5.5182e-05 3.8182 0.012034 1.5759e-05 0.0011542 0.15499 0.00065837 0.15564 0.14197 0 0.036681 0.0389 0 0.90395 0.25292 0.068139 0.0094974 4.278 0.059298 7.1292e-05 0.83077 0.0052982 0.0060358 0.0018119 0.98096 0.91442 3.9727e-06 1.5892e-05 0.13206 0.66261 0.72419 0.0016081 0.69532 0.4859 0.0021587 0.42276 1.1752 1.1702 16.0007 144.9779 0.00046779 -84.0447 0.094362
1.1984 0.98803 5.5182e-05 3.8182 0.012034 1.5772e-05 0.0011542 0.15505 0.00065837 0.15571 0.14203 0 0.036677 0.0389 0 0.90402 0.25296 0.068152 0.009499 4.2784 0.059308 7.1304e-05 0.83076 0.0052986 0.0060362 0.0018068 0.98105 0.91867 3.962e-06 1.5849e-05 0.13206 0.6636 0.72519 0.0016059 0.69698 0.48607 0.0021558 0.42276 1.1773 1.1723 16.0008 144.9779 0.00046631 -84.06 0.095362
1.1994 0.98803 5.5182e-05 3.8182 0.012034 1.5785e-05 0.0011542 0.15512 0.00065838 0.15577 0.14209 0 0.036673 0.0389 0 0.9041 0.25299 0.068164 0.0095005 4.2788 0.059317 7.1316e-05 0.83075 0.005299 0.0060366 0.0018027 0.98114 0.92268 3.9516e-06 1.5808e-05 0.13207 0.66459 0.72618 0.0016039 0.69864 0.48624 0.0021531 0.42275 1.1794 1.1744 16.0009 144.9779 0.00046484 -84.0748 0.096362
1.2004 0.98803 5.5182e-05 3.8182 0.012034 1.5798e-05 0.0011542 0.15518 0.00065838 0.15584 0.14215 0 0.036669 0.0389 0 0.90418 0.25303 0.068177 0.009502 4.2792 0.059327 7.1328e-05 0.83074 0.0052994 0.006037 0.0017979 0.98121 0.92646 3.9416e-06 1.5767e-05 0.13207 0.66557 0.72716 0.0016018 0.70029 0.48641 0.0021504 0.42275 1.1816 1.1766 16.001 144.978 0.00046337 -84.0891 0.097362
1.2014 0.98803 5.5182e-05 3.8182 0.012034 1.5812e-05 0.0011542 0.15525 0.00065838 0.1559 0.14221 0 0.036665 0.0389 0 0.90426 0.25306 0.06819 0.0095036 4.2795 0.059336 7.134e-05 0.83074 0.0052997 0.0060374 0.0017946 0.98129 0.93004 3.9318e-06 1.5728e-05 0.13207 0.66656 0.72814 0.0015999 0.70193 0.48658 0.0021477 0.42275 1.1837 1.1787 16.001 144.978 0.00046191 -84.1031 0.098362
1.2024 0.98803 5.5182e-05 3.8182 0.012034 1.5825e-05 0.0011542 0.15531 0.00065838 0.15596 0.14227 0 0.036661 0.0389 0 0.90434 0.2531 0.068202 0.0095051 4.2799 0.059346 7.1353e-05 0.83073 0.0053001 0.0060378 0.0017902 0.98136 0.93341 3.9223e-06 1.5691e-05 0.13208 0.66754 0.72911 0.001598 0.70357 0.48675 0.0021452 0.42275 1.1858 1.1809 16.0011 144.978 0.00046046 -84.1167 0.099362
1.2034 0.98803 5.5181e-05 3.8182 0.012034 1.5838e-05 0.0011542 0.15537 0.00065838 0.15603 0.14233 0 0.036657 0.0389 0 0.90442 0.25313 0.068215 0.0095067 4.2803 0.059355 7.1365e-05 0.83072 0.0053005 0.0060382 0.0017868 0.98142 0.93659 3.9131e-06 1.5654e-05 0.13208 0.66851 0.73007 0.0015961 0.7052 0.48692 0.0021427 0.42275 1.1879 1.183 16.0012 144.978 0.00045902 -84.13 0.10036
1.2044 0.98803 5.5181e-05 3.8182 0.012034 1.5851e-05 0.0011542 0.15544 0.00065838 0.15609 0.14239 0 0.036653 0.0389 0 0.9045 0.25317 0.068227 0.0095082 4.2806 0.059365 7.1377e-05 0.83071 0.0053009 0.0060385 0.0017815 0.98149 0.9396 3.9041e-06 1.5618e-05 0.13208 0.66949 0.73103 0.0015943 0.70682 0.48709 0.0021403 0.42274 1.19 1.1851 16.0013 144.978 0.00045759 -84.143 0.10136
1.2054 0.98803 5.5181e-05 3.8182 0.012034 1.5864e-05 0.0011542 0.1555 0.00065838 0.15616 0.14245 0 0.036648 0.0389 0 0.90457 0.2532 0.06824 0.0095097 4.281 0.059374 7.1389e-05 0.8307 0.0053013 0.0060389 0.0017797 0.98155 0.94243 3.8953e-06 1.5582e-05 0.13209 0.67046 0.73198 0.0015925 0.70844 0.48726 0.002138 0.42274 1.1921 1.1872 16.0014 144.978 0.00045616 -84.1558 0.10236
1.2064 0.98803 5.5181e-05 3.8182 0.012034 1.5877e-05 0.0011542 0.15557 0.00065838 0.15622 0.14251 0 0.036644 0.0389 0 0.90465 0.25324 0.068253 0.0095113 4.2814 0.059384 7.1401e-05 0.83069 0.0053017 0.0060393 0.0017752 0.98161 0.94511 3.8867e-06 1.5548e-05 0.13209 0.67143 0.73293 0.0015908 0.71005 0.48743 0.0021357 0.42274 1.1942 1.1894 16.0014 144.978 0.00045474 -84.1683 0.10336
1.2074 0.98803 5.5181e-05 3.8182 0.012034 1.589e-05 0.0011542 0.15563 0.00065839 0.15629 0.14257 0 0.03664 0.0389 0 0.90473 0.25327 0.068265 0.0095128 4.2818 0.059393 7.1414e-05 0.83068 0.0053021 0.0060397 0.0017709 0.98167 0.94764 3.8783e-06 1.5514e-05 0.13209 0.67239 0.73386 0.0015891 0.71165 0.4876 0.0021334 0.42274 1.1963 1.1915 16.0015 144.978 0.00045333 -84.1805 0.10436
1.2084 0.98803 5.5181e-05 3.8182 0.012034 1.5903e-05 0.0011542 0.1557 0.00065839 0.15635 0.14263 0 0.036636 0.0389 0 0.90481 0.25331 0.068278 0.0095144 4.2821 0.059403 7.1426e-05 0.83067 0.0053025 0.0060401 0.0017679 0.98172 0.95002 3.87e-06 1.5481e-05 0.1321 0.67336 0.7348 0.0015874 0.71324 0.48777 0.0021312 0.42274 1.1984 1.1936 16.0016 144.978 0.00045193 -84.1926 0.10536
1.2094 0.98803 5.5181e-05 3.8182 0.012034 1.5917e-05 0.0011542 0.15576 0.00065839 0.15641 0.14269 0 0.036632 0.0389 0 0.90489 0.25334 0.068291 0.0095159 4.2825 0.059412 7.1438e-05 0.83066 0.0053028 0.0060405 0.0017636 0.98177 0.95227 3.8619e-06 1.5449e-05 0.1321 0.67432 0.73572 0.0015857 0.71483 0.48794 0.002129 0.42274 1.2005 1.1957 16.0017 144.978 0.00045053 -84.2044 0.10636
1.2104 0.98803 5.5181e-05 3.8182 0.012034 1.593e-05 0.0011542 0.15582 0.00065839 0.15648 0.14275 0 0.036628 0.0389 0 0.90497 0.25338 0.068303 0.0095175 4.2829 0.059422 7.145e-05 0.83065 0.0053032 0.0060409 0.0017615 0.98183 0.9544 3.8539e-06 1.5417e-05 0.1321 0.67527 0.73664 0.0015841 0.71641 0.48811 0.0021269 0.42274 1.2026 1.1978 16.0017 144.978 0.00044914 -84.2161 0.10736
1.2114 0.98803 5.5181e-05 3.8182 0.012034 1.5943e-05 0.0011542 0.15589 0.00065839 0.15654 0.14281 0 0.036624 0.0389 0 0.90505 0.25341 0.068316 0.009519 4.2833 0.059431 7.1462e-05 0.83064 0.0053036 0.0060413 0.0017561 0.98188 0.9564 3.8461e-06 1.5385e-05 0.13211 0.67623 0.73756 0.0015825 0.71799 0.48828 0.0021248 0.42274 1.2047 1.1999 16.0018 144.9781 0.00044776 -84.2276 0.10836
1.2124 0.98803 5.5181e-05 3.8182 0.012034 1.5956e-05 0.0011542 0.15595 0.00065839 0.1566 0.14287 0 0.03662 0.0389 0 0.90513 0.25345 0.068329 0.0095205 4.2837 0.059441 7.1475e-05 0.83063 0.005304 0.0060417 0.0017535 0.98193 0.95829 3.8384e-06 1.5354e-05 0.13211 0.67718 0.73847 0.001581 0.71955 0.48845 0.0021227 0.42273 1.2068 1.202 16.0019 144.9781 0.00044638 -84.2389 0.10936
1.2134 0.98803 5.5181e-05 3.8182 0.012034 1.5969e-05 0.0011542 0.15601 0.00065839 0.15667 0.14293 0 0.036616 0.0389 0 0.90521 0.25348 0.068341 0.0095221 4.284 0.05945 7.1487e-05 0.83062 0.0053044 0.0060421 0.00175 0.98198 0.96007 3.8308e-06 1.5324e-05 0.13211 0.67813 0.73937 0.0015794 0.72111 0.48862 0.0021207 0.42273 1.2088 1.2041 16.0019 144.9781 0.00044502 -84.2501 0.11036
1.2144 0.98803 5.5181e-05 3.8182 0.012034 1.5982e-05 0.0011542 0.15608 0.00065839 0.15673 0.14299 0 0.036612 0.0389 0 0.90528 0.25352 0.068354 0.0095236 4.2844 0.05946 7.1499e-05 0.83061 0.0053048 0.0060425 0.0017482 0.98202 0.96175 3.8233e-06 1.5294e-05 0.13212 0.67907 0.74026 0.0015779 0.72267 0.48879 0.0021187 0.42273 1.2109 1.2062 16.002 144.9781 0.00044366 -84.2612 0.11136
1.2154 0.98803 5.5181e-05 3.8182 0.012034 1.5995e-05 0.0011542 0.15614 0.00065839 0.1568 0.14305 0 0.036608 0.0389 0 0.90536 0.25355 0.068367 0.0095252 4.2848 0.059469 7.1511e-05 0.8306 0.0053052 0.0060429 0.0017434 0.98207 0.96334 3.816e-06 1.5265e-05 0.13212 0.68002 0.74116 0.0015764 0.72421 0.48896 0.0021167 0.42273 1.213 1.2082 16.0021 144.9781 0.00044231 -84.2721 0.11236
1.2164 0.98803 5.5181e-05 3.8182 0.012034 1.6009e-05 0.0011542 0.15621 0.0006584 0.15686 0.14311 0 0.036604 0.0389 0 0.90544 0.25359 0.068379 0.0095267 4.2852 0.059479 7.1524e-05 0.83059 0.0053056 0.0060433 0.0017408 0.98212 0.96484 3.8087e-06 1.5236e-05 0.13212 0.68096 0.74204 0.0015749 0.72575 0.48913 0.0021148 0.42273 1.215 1.2103 16.0022 144.9781 0.00044096 -84.2828 0.11336
1.2174 0.98803 5.5181e-05 3.8182 0.012034 1.6022e-05 0.0011542 0.15627 0.0006584 0.15692 0.14317 0 0.0366 0.0389 0 0.90552 0.25362 0.068392 0.0095283 4.2856 0.059488 7.1536e-05 0.83058 0.005306 0.0060437 0.0017376 0.98216 0.96625 3.8015e-06 1.5207e-05 0.13213 0.68189 0.74292 0.0015734 0.72728 0.4893 0.0021128 0.42273 1.2171 1.2124 16.0022 144.9781 0.00043962 -84.2935 0.11436
1.2184 0.98803 5.5181e-05 3.8182 0.012034 1.6035e-05 0.0011542 0.15633 0.0006584 0.15699 0.14323 0 0.036596 0.0389 0 0.9056 0.25366 0.068405 0.0095298 4.2859 0.059498 7.1548e-05 0.83057 0.0053064 0.0060441 0.0017356 0.98221 0.96758 3.7944e-06 1.5179e-05 0.13213 0.68283 0.74379 0.001572 0.72881 0.48947 0.0021109 0.42273 1.2191 1.2145 16.0023 144.9781 0.00043829 -84.304 0.11536
1.2194 0.98803 5.518e-05 3.8182 0.012034 1.6048e-05 0.0011542 0.1564 0.0006584 0.15705 0.14329 0 0.036592 0.0389 0 0.90568 0.25369 0.068417 0.0095314 4.2863 0.059507 7.1561e-05 0.83056 0.0053068 0.0060445 0.0017314 0.98225 0.96884 3.7874e-06 1.5151e-05 0.13213 0.68376 0.74466 0.0015705 0.73033 0.48964 0.0021091 0.42273 1.2212 1.2165 16.0024 144.9781 0.00043697 -84.3144 0.11636
1.2204 0.98803 5.518e-05 3.8182 0.012034 1.6061e-05 0.0011542 0.15646 0.0006584 0.15711 0.14335 0 0.036588 0.0389 0 0.90576 0.25373 0.06843 0.0095329 4.2867 0.059517 7.1573e-05 0.83055 0.0053071 0.0060449 0.0017288 0.98229 0.97002 3.7805e-06 1.5123e-05 0.13214 0.68469 0.74552 0.0015691 0.73184 0.48981 0.0021072 0.42273 1.2232 1.2186 16.0024 144.9781 0.00043565 -84.3247 0.11736
1.2214 0.98803 5.518e-05 3.8182 0.012034 1.6074e-05 0.0011542 0.15652 0.0006584 0.15718 0.14341 0 0.036584 0.0389 0 0.90584 0.25377 0.068443 0.0095345 4.2871 0.059526 7.1585e-05 0.83055 0.0053075 0.0060453 0.0017258 0.98233 0.97114 3.7737e-06 1.5096e-05 0.13214 0.68561 0.74638 0.0015677 0.73334 0.48998 0.0021054 0.42273 1.2253 1.2207 16.0025 144.9782 0.00043434 -84.3349 0.11836
1.2224 0.98803 5.518e-05 3.8182 0.012034 1.6087e-05 0.0011542 0.15659 0.0006584 0.15724 0.14347 0 0.03658 0.0389 0 0.90592 0.2538 0.068455 0.009536 4.2875 0.059536 7.1597e-05 0.83054 0.0053079 0.0060457 0.0017237 0.98238 0.9722 3.767e-06 1.5069e-05 0.13214 0.68653 0.74723 0.0015663 0.73484 0.49015 0.0021036 0.42274 1.2273 1.2227 16.0026 144.9782 0.00043304 -84.345 0.11936
1.2234 0.98803 5.518e-05 3.8182 0.012034 1.61e-05 0.0011542 0.15665 0.0006584 0.1573 0.14353 0 0.036576 0.0389 0 0.906 0.25384 0.068468 0.0095376 4.2878 0.059545 7.161e-05 0.83053 0.0053083 0.0060461 0.0017199 0.98242 0.97319 3.7603e-06 1.5042e-05 0.13215 0.68745 0.74808 0.001565 0.73633 0.49032 0.0021018 0.42274 1.2293 1.2248 16.0026 144.9782 0.00043175 -84.355 0.12036
1.2244 0.98803 5.518e-05 3.8182 0.012034 1.6114e-05 0.0011542 0.15671 0.0006584 0.15737 0.14359 0 0.036572 0.0389 0 0.90608 0.25387 0.068481 0.0095391 4.2882 0.059555 7.1622e-05 0.83052 0.0053087 0.0060465 0.0017187 0.98246 0.97413 3.7537e-06 1.5016e-05 0.13215 0.68837 0.74892 0.0015636 0.73781 0.49049 0.0021 0.42274 1.2314 1.2268 16.0027 144.9782 0.00043046 -84.3649 0.12136
1.2254 0.98803 5.518e-05 3.8182 0.012034 1.6127e-05 0.0011542 0.15678 0.00065841 0.15743 0.14364 0 0.036568 0.0389 0 0.90616 0.25391 0.068494 0.0095407 4.2886 0.059564 7.1634e-05 0.83051 0.0053091 0.0060469 0.0017154 0.9825 0.97501 3.7472e-06 1.499e-05 0.13215 0.68928 0.74976 0.0015623 0.73929 0.49066 0.0020982 0.42274 1.2334 1.2288 16.0028 144.9782 0.00042918 -84.3748 0.12236
1.2264 0.98803 5.518e-05 3.8182 0.012034 1.614e-05 0.0011542 0.15684 0.00065841 0.15749 0.1437 0 0.036564 0.0389 0 0.90623 0.25394 0.068506 0.0095422 4.289 0.059574 7.1647e-05 0.8305 0.0053095 0.0060473 0.0017128 0.98254 0.97585 3.7408e-06 1.4964e-05 0.13216 0.6902 0.75059 0.0015609 0.74076 0.49083 0.0020965 0.42274 1.2354 1.2309 16.0028 144.9782 0.0004279 -84.3845 0.12336
1.2274 0.98803 5.518e-05 3.8182 0.012034 1.6153e-05 0.0011542 0.1569 0.00065841 0.15756 0.14376 0 0.03656 0.0389 0 0.90631 0.25398 0.068519 0.0095438 4.2894 0.059584 7.1659e-05 0.83049 0.0053099 0.0060477 0.001709 0.98258 0.97664 3.7344e-06 1.4938e-05 0.13216 0.6911 0.75141 0.0015596 0.74222 0.491 0.0020948 0.42274 1.2374 1.2329 16.0029 144.9782 0.00042663 -84.3941 0.12436
1.2284 0.98803 5.518e-05 3.8182 0.012034 1.6166e-05 0.0011542 0.15697 0.00065841 0.15762 0.14382 0 0.036556 0.0389 0 0.90639 0.25401 0.068532 0.0095453 4.2898 0.059593 7.1671e-05 0.83048 0.0053103 0.0060481 0.0017076 0.98262 0.97738 3.7281e-06 1.4913e-05 0.13216 0.69201 0.75223 0.0015583 0.74368 0.49117 0.0020931 0.42274 1.2394 1.2349 16.003 144.9782 0.00042537 -84.4037 0.12536
1.2294 0.98803 5.518e-05 3.8182 0.012034 1.6179e-05 0.0011542 0.15703 0.00065841 0.15768 0.14388 0 0.036552 0.0389 0 0.90647 0.25405 0.068544 0.0095469 4.2901 0.059603 7.1684e-05 0.83047 0.0053107 0.0060485 0.0017045 0.98265 0.97808 3.7219e-06 1.4888e-05 0.13217 0.69291 0.75305 0.001557 0.74512 0.49134 0.0020914 0.42274 1.2414 1.237 16.003 144.9782 0.00042412 -84.4131 0.12636
1.2304 0.98803 5.518e-05 3.8182 0.012034 1.6192e-05 0.0011542 0.15709 0.00065841 0.15775 0.14394 0 0.036548 0.0389 0 0.90655 0.25408 0.068557 0.0095484 4.2905 0.059612 7.1696e-05 0.83046 0.0053111 0.0060489 0.0017019 0.98269 0.97874 3.7157e-06 1.4863e-05 0.13217 0.69381 0.75386 0.0015558 0.74657 0.49151 0.0020897 0.42274 1.2434 1.239 16.0031 144.9783 0.00042287 -84.4225 0.12736
1.2314 0.98803 5.518e-05 3.8182 0.012034 1.6206e-05 0.0011542 0.15715 0.00065841 0.15781 0.144 0 0.036544 0.0389 0 0.90663 0.25412 0.06857 0.00955 4.2909 0.059622 7.1708e-05 0.83045 0.0053115 0.0060493 0.0016984 0.98273 0.97936 3.7096e-06 1.4839e-05 0.13217 0.69471 0.75466 0.0015545 0.748 0.49168 0.0020881 0.42275 1.2454 1.241 16.0032 144.9783 0.00042162 -84.4318 0.12836
1.2324 0.98803 5.518e-05 3.8182 0.012034 1.6219e-05 0.0011542 0.15722 0.00065841 0.15787 0.14406 0 0.03654 0.0389 0 0.90671 0.25415 0.068583 0.0095515 4.2913 0.059631 7.1721e-05 0.83044 0.0053119 0.0060497 0.0016968 0.98277 0.97995 3.7035e-06 1.4815e-05 0.13218 0.69561 0.75546 0.0015532 0.74943 0.49185 0.0020864 0.42275 1.2474 1.243 16.0032 144.9783 0.00042039 -84.441 0.12936
1.2334 0.98803 5.518e-05 3.8182 0.012034 1.6232e-05 0.0011542 0.15728 0.00065841 0.15793 0.14412 0 0.036536 0.0389 0 0.90679 0.25419 0.068595 0.0095531 4.2917 0.059641 7.1733e-05 0.83043 0.0053123 0.0060501 0.0016924 0.9828 0.98051 3.6975e-06 1.4791e-05 0.13218 0.6965 0.75626 0.001552 0.75085 0.49202 0.0020848 0.42275 1.2494 1.245 16.0033 144.9783 0.00041916 -84.4502 0.13036
1.2344 0.98803 5.518e-05 3.8182 0.012034 1.6245e-05 0.0011542 0.15734 0.00065842 0.158 0.14418 0 0.036532 0.0389 0 0.90687 0.25422 0.068608 0.0095546 4.2921 0.059651 7.1745e-05 0.83042 0.0053127 0.0060505 0.0016904 0.98284 0.98103 3.6916e-06 1.4767e-05 0.13218 0.69739 0.75705 0.0015508 0.75226 0.49219 0.0020832 0.42275 1.2514 1.247 16.0034 144.9783 0.00041794 -84.4592 0.13136
1.2354 0.98803 5.5179e-05 3.8182 0.012034 1.6258e-05 0.0011542 0.15741 0.00065842 0.15806 0.14423 0 0.036528 0.0389 0 0.90695 0.25426 0.068621 0.0095562 4.2925 0.05966 7.1758e-05 0.83041 0.0053131 0.0060509 0.0016878 0.98287 0.98153 3.6857e-06 1.4744e-05 0.13219 0.69827 0.75783 0.0015495 0.75367 0.49236 0.0020816 0.42275 1.2534 1.249 16.0034 144.9783 0.00041672 -84.4682 0.13236
1.2364 0.98803 5.5179e-05 3.8182 0.012034 1.6271e-05 0.0011542 0.15747 0.00065842 0.15812 0.14429 0 0.036524 0.0389 0 0.90703 0.25429 0.068634 0.0095577 4.2929 0.05967 7.177e-05 0.8304 0.0053135 0.0060513 0.0016864 0.98291 0.98199 3.6799e-06 1.472e-05 0.13219 0.69916 0.75861 0.0015483 0.75507 0.49253 0.00208 0.42275 1.2554 1.251 16.0035 144.9783 0.00041551 -84.4771 0.13336
1.2374 0.98803 5.5179e-05 3.8182 0.012034 1.6284e-05 0.0011542 0.15753 0.00065842 0.15818 0.14435 0 0.036521 0.0389 0 0.90711 0.25433 0.068647 0.0095593 4.2932 0.059679 7.1782e-05 0.83039 0.0053139 0.0060517 0.0016826 0.98294 0.98243 3.6742e-06 1.4697e-05 0.13219 0.70004 0.75939 0.0015471 0.75647 0.4927 0.0020784 0.42276 1.2574 1.253 16.0035 144.9783 0.00041431 -84.486 0.13436
1.2384 0.98803 5.5179e-05 3.8182 0.012033 1.6297e-05 0.0011542 0.15759 0.00065842 0.15825 0.14441 0 0.036517 0.0389 0 0.90719 0.25437 0.068659 0.0095609 4.2936 0.059689 7.1795e-05 0.83038 0.0053143 0.0060521 0.0016805 0.98298 0.98285 3.6685e-06 1.4675e-05 0.1322 0.70092 0.76016 0.001546 0.75785 0.49287 0.0020769 0.42276 1.2593 1.255 16.0036 144.9783 0.00041311 -84.4947 0.13536
1.2394 0.98803 5.5179e-05 3.8182 0.012033 1.6311e-05 0.0011542 0.15766 0.00065842 0.15831 0.14447 0 0.036513 0.0389 0 0.90727 0.2544 0.068672 0.0095624 4.294 0.059698 7.1807e-05 0.83037 0.0053147 0.0060525 0.0016781 0.98301 0.98324 3.6628e-06 1.4652e-05 0.1322 0.70179 0.76093 0.0015448 0.75923 0.49304 0.0020753 0.42276 1.2613 1.257 16.0037 144.9784 0.00041192 -84.5034 0.13636
1.2404 0.98803 5.5179e-05 3.8182 0.012033 1.6324e-05 0.0011542 0.15772 0.00065842 0.15837 0.14453 0 0.036509 0.0389 0 0.90735 0.25444 0.068685 0.009564 4.2944 0.059708 7.1819e-05 0.83036 0.0053151 0.0060529 0.0016765 0.98305 0.98361 3.6573e-06 1.463e-05 0.1322 0.70267 0.76169 0.0015436 0.76061 0.49321 0.0020738 0.42276 1.2633 1.2589 16.0037 144.9784 0.00041074 -84.5121 0.13736
1.2414 0.98803 5.5179e-05 3.8182 0.012033 1.6337e-05 0.0011542 0.15778 0.00065842 0.15843 0.14459 0 0.036505 0.0389 0 0.90743 0.25447 0.068698 0.0095655 4.2948 0.059718 7.1832e-05 0.83035 0.0053155 0.0060533 0.0016731 0.98308 0.98396 3.6517e-06 1.4608e-05 0.13221 0.70354 0.76245 0.0015425 0.76197 0.49338 0.0020723 0.42277 1.2652 1.2609 16.0038 144.9784 0.00040956 -84.5206 0.13836
1.2424 0.98803 5.5179e-05 3.8182 0.012033 1.635e-05 0.0011542 0.15784 0.00065842 0.1585 0.14464 0 0.036501 0.0389 0 0.90751 0.25451 0.06871 0.0095671 4.2952 0.059727 7.1844e-05 0.83034 0.0053159 0.0060537 0.0016711 0.98311 0.98429 3.6462e-06 1.4586e-05 0.13221 0.70441 0.7632 0.0015413 0.76333 0.49355 0.0020708 0.42277 1.2672 1.2629 16.0038 144.9784 0.00040838 -84.5291 0.13936
1.2434 0.98803 5.5179e-05 3.8182 0.012033 1.6363e-05 0.0011542 0.15791 0.00065843 0.15856 0.1447 0 0.036497 0.0389 0 0.90759 0.25454 0.068723 0.0095686 4.2956 0.059737 7.1857e-05 0.83033 0.0053163 0.0060541 0.0016687 0.98315 0.9846 3.6408e-06 1.4564e-05 0.13221 0.70527 0.76395 0.0015402 0.76469 0.49372 0.0020693 0.42277 1.2691 1.2648 16.0039 144.9784 0.00040722 -84.5375 0.14036
1.2444 0.98803 5.5179e-05 3.8182 0.012033 1.6376e-05 0.0011542 0.15797 0.00065843 0.15862 0.14476 0 0.036493 0.0389 0 0.90767 0.25458 0.068736 0.0095702 4.296 0.059746 7.1869e-05 0.83033 0.0053167 0.0060545 0.001667 0.98318 0.98489 3.6354e-06 1.4542e-05 0.13222 0.70613 0.7647 0.001539 0.76603 0.49389 0.0020679 0.42277 1.2711 1.2668 16.004 144.9784 0.00040606 -84.5459 0.14136
1.2454 0.98803 5.5179e-05 3.8182 0.012033 1.6389e-05 0.0011542 0.15803 0.00065843 0.15868 0.14482 0 0.036489 0.0389 0 0.90775 0.25461 0.068749 0.0095718 4.2964 0.059756 7.1881e-05 0.83032 0.0053171 0.0060549 0.001664 0.98321 0.98517 3.6301e-06 1.4521e-05 0.13222 0.70699 0.76544 0.0015379 0.76737 0.49406 0.0020664 0.42278 1.273 1.2688 16.004 144.9784 0.0004049 -84.5542 0.14236
1.2464 0.98803 5.5179e-05 3.8182 0.012033 1.6403e-05 0.0011542 0.15809 0.00065843 0.15875 0.14488 0 0.036485 0.0389 0 0.90783 0.25465 0.068762 0.0095733 4.2968 0.059766 7.1894e-05 0.83031 0.0053175 0.0060553 0.0016631 0.98324 0.98544 3.6248e-06 1.45e-05 0.13222 0.70785 0.76617 0.0015368 0.76871 0.49423 0.002065 0.42278 1.2749 1.2707 16.0041 144.9784 0.00040375 -84.5624 0.14336
1.2474 0.98803 5.5179e-05 3.8182 0.012033 1.6416e-05 0.0011542 0.15815 0.00065843 0.15881 0.14494 0 0.036481 0.0389 0 0.90791 0.25468 0.068774 0.0095749 4.2972 0.059775 7.1906e-05 0.8303 0.0053179 0.0060557 0.0016605 0.98327 0.98568 3.6196e-06 1.4479e-05 0.13223 0.7087 0.7669 0.0015357 0.77003 0.4944 0.0020635 0.42278 1.2769 1.2727 16.0041 144.9784 0.00040261 -84.5705 0.14436
1.2484 0.98803 5.5179e-05 3.8182 0.012033 1.6429e-05 0.0011542 0.15822 0.00065843 0.15887 0.14499 0 0.036477 0.0389 0 0.90799 0.25472 0.068787 0.0095764 4.2976 0.059785 7.1919e-05 0.83029 0.0053183 0.0060562 0.0016583 0.9833 0.98592 3.6144e-06 1.4458e-05 0.13223 0.70956 0.76763 0.0015346 0.77135 0.49457 0.0020621 0.42279 1.2788 1.2746 16.0042 144.9785 0.00040148 -84.5786 0.14536
1.2494 0.98803 5.5179e-05 3.8182 0.012033 1.6442e-05 0.0011542 0.15828 0.00065843 0.15893 0.14505 0 0.036474 0.0389 0 0.90807 0.25476 0.0688 0.009578 4.298 0.059795 7.1931e-05 0.83028 0.0053187 0.0060566 0.0016552 0.98333 0.98614 3.6093e-06 1.4438e-05 0.13223 0.71041 0.76835 0.0015336 0.77267 0.49474 0.0020607 0.42279 1.2807 1.2765 16.0042 144.9785 0.00040034 -84.5867 0.14636
1.2504 0.98803 5.5179e-05 3.8182 0.012033 1.6455e-05 0.0011542 0.15834 0.00065843 0.15899 0.14511 0 0.03647 0.0389 0 0.90815 0.25479 0.068813 0.0095796 4.2983 0.059804 7.1943e-05 0.83027 0.0053191 0.006057 0.001654 0.98337 0.98635 3.6042e-06 1.4417e-05 0.13224 0.71125 0.76907 0.0015325 0.77398 0.49491 0.0020593 0.42279 1.2826 1.2785 16.0043 144.9785 0.00039922 -84.5946 0.14736
1.2514 0.98803 5.5178e-05 3.8182 0.012033 1.6468e-05 0.0011542 0.1584 0.00065843 0.15906 0.14517 0 0.036466 0.0389 0 0.90823 0.25483 0.068826 0.0095811 4.2987 0.059814 7.1956e-05 0.83026 0.0053195 0.0060574 0.0016516 0.9834 0.98655 3.5992e-06 1.4397e-05 0.13224 0.7121 0.76979 0.0015314 0.77528 0.49508 0.0020579 0.4228 1.2846 1.2804 16.0044 144.9785 0.0003981 -84.6025 0.14836
1.2524 0.98803 5.5178e-05 3.8182 0.012033 1.6481e-05 0.0011542 0.15846 0.00065843 0.15912 0.14523 0 0.036462 0.0389 0 0.90831 0.25486 0.068839 0.0095827 4.2991 0.059823 7.1968e-05 0.83025 0.0053199 0.0060578 0.0016494 0.98343 0.98673 3.5942e-06 1.4377e-05 0.13224 0.71294 0.7705 0.0015304 0.77657 0.49525 0.0020565 0.4228 1.2865 1.2823 16.0044 144.9785 0.00039699 -84.6104 0.14936
1.2534 0.98803 5.5178e-05 3.8182 0.012033 1.6494e-05 0.0011542 0.15853 0.00065844 0.15918 0.14528 0 0.036458 0.0389 0 0.90839 0.2549 0.068851 0.0095843 4.2995 0.059833 7.1981e-05 0.83024 0.0053203 0.0060582 0.0016467 0.98346 0.98691 3.5892e-06 1.4358e-05 0.13225 0.71378 0.7712 0.0015293 0.77786 0.49542 0.0020552 0.4228 1.2884 1.2843 16.0045 144.9785 0.00039588 -84.6181 0.15036
1.2544 0.98803 5.5178e-05 3.8182 0.012033 1.6508e-05 0.0011542 0.15859 0.00065844 0.15924 0.14534 0 0.036454 0.0389 0 0.90847 0.25493 0.068864 0.0095858 4.2999 0.059843 7.1993e-05 0.83023 0.0053207 0.0060586 0.0016452 0.98348 0.98708 3.5844e-06 1.4338e-05 0.13225 0.71462 0.7719 0.0015283 0.77914 0.49559 0.0020538 0.42281 1.2903 1.2862 16.0045 144.9785 0.00039478 -84.6258 0.15136
1.2554 0.98803 5.5178e-05 3.8182 0.012033 1.6521e-05 0.0011542 0.15865 0.00065844 0.1593 0.1454 0 0.03645 0.0389 0 0.90855 0.25497 0.068877 0.0095874 4.3003 0.059852 7.2006e-05 0.83022 0.0053211 0.006059 0.0016419 0.98351 0.98724 3.5795e-06 1.4319e-05 0.13225 0.71545 0.7726 0.0015273 0.78041 0.49576 0.0020525 0.42281 1.2922 1.2881 16.0046 144.9785 0.00039368 -84.6335 0.15236
1.2564 0.98803 5.5178e-05 3.8182 0.012033 1.6534e-05 0.0011542 0.15871 0.00065844 0.15936 0.14546 0 0.036446 0.0389 0 0.90863 0.25501 0.06889 0.009589 4.3007 0.059862 7.2018e-05 0.83021 0.0053215 0.0060594 0.0016401 0.98354 0.98739 3.5747e-06 1.4299e-05 0.13226 0.71628 0.7733 0.0015263 0.78168 0.49593 0.0020512 0.42281 1.2941 1.29 16.0046 144.9786 0.00039259 -84.6411 0.15336
1.2574 0.98803 5.5178e-05 3.8182 0.012033 1.6547e-05 0.0011542 0.15877 0.00065844 0.15943 0.14552 0 0.036443 0.0389 0 0.90871 0.25504 0.068903 0.0095905 4.3011 0.059872 7.203e-05 0.8302 0.0053219 0.0060598 0.0016381 0.98357 0.98753 3.5699e-06 1.428e-05 0.13226 0.71711 0.77399 0.0015253 0.78294 0.4961 0.0020498 0.42282 1.296 1.2919 16.0047 144.9786 0.00039151 -84.6486 0.15436
1.2584 0.98803 5.5178e-05 3.8182 0.012033 1.656e-05 0.0011542 0.15883 0.00065844 0.15949 0.14557 0 0.036439 0.0389 0 0.90879 0.25508 0.068916 0.0095921 4.3015 0.059881 7.2043e-05 0.83019 0.0053224 0.0060603 0.0016368 0.9836 0.98766 3.5652e-06 1.4261e-05 0.13226 0.71794 0.77467 0.0015243 0.7842 0.49627 0.0020485 0.42282 1.2978 1.2938 16.0047 144.9786 0.00039043 -84.6561 0.15536
1.2594 0.98803 5.5178e-05 3.8182 0.012033 1.6573e-05 0.0011542 0.1589 0.00065844 0.15955 0.14563 0 0.036435 0.0389 0 0.90887 0.25511 0.068929 0.0095936 4.3019 0.059891 7.2055e-05 0.83018 0.0053228 0.0060607 0.0016339 0.98363 0.98779 3.5605e-06 1.4243e-05 0.13227 0.71876 0.77535 0.0015233 0.78545 0.49644 0.0020473 0.42283 1.2997 1.2957 16.0048 144.9786 0.00038935 -84.6635 0.15636
1.2604 0.98803 5.5178e-05 3.8182 0.012033 1.6586e-05 0.0011542 0.15896 0.00065844 0.15961 0.14569 0 0.036431 0.0389 0 0.90895 0.25515 0.068941 0.0095952 4.3023 0.059901 7.2068e-05 0.83017 0.0053232 0.0060611 0.0016321 0.98365 0.98791 3.5559e-06 1.4224e-05 0.13227 0.71958 0.77603 0.0015223 0.78669 0.49661 0.002046 0.42283 1.3016 1.2976 16.0048 144.9786 0.00038828 -84.6709 0.15736
1.2614 0.98803 5.5178e-05 3.8182 0.012033 1.66e-05 0.0011542 0.15902 0.00065844 0.15967 0.14575 0 0.036427 0.0389 0 0.90903 0.25518 0.068954 0.0095968 4.3027 0.05991 7.208e-05 0.83016 0.0053236 0.0060615 0.0016302 0.98368 0.98803 3.5513e-06 1.4206e-05 0.13227 0.7204 0.77671 0.0015213 0.78793 0.49678 0.0020447 0.42284 1.3035 1.2995 16.0049 144.9786 0.00038722 -84.6782 0.15836
1.2624 0.98803 5.5178e-05 3.8182 0.012033 1.6613e-05 0.0011542 0.15908 0.00065845 0.15973 0.1458 0 0.036423 0.0389 0 0.90911 0.25522 0.068967 0.0095983 4.3031 0.05992 7.2093e-05 0.83015 0.005324 0.0060619 0.0016287 0.98371 0.98814 3.5468e-06 1.4187e-05 0.13228 0.72122 0.77738 0.0015204 0.78916 0.49695 0.0020434 0.42284 1.3053 1.3014 16.0049 144.9786 0.00038616 -84.6854 0.15936
1.2634 0.98803 5.5178e-05 3.8182 0.012033 1.6626e-05 0.0011542 0.15914 0.00065845 0.15979 0.14586 0 0.03642 0.0389 0 0.90919 0.25525 0.06898 0.0095999 4.3035 0.05993 7.2105e-05 0.83014 0.0053244 0.0060623 0.0016262 0.98374 0.98824 3.5422e-06 1.4169e-05 0.13228 0.72203 0.77805 0.0015194 0.79038 0.49712 0.0020422 0.42284 1.3072 1.3032 16.005 144.9786 0.00038511 -84.6926 0.16036
1.2644 0.98803 5.5178e-05 3.8182 0.012033 1.6639e-05 0.0011542 0.1592 0.00065845 0.15986 0.14592 0 0.036416 0.0389 0 0.90927 0.25529 0.068993 0.0096015 4.3039 0.059939 7.2118e-05 0.83013 0.0053248 0.0060627 0.0016254 0.98376 0.98834 3.5378e-06 1.4152e-05 0.13228 0.72284 0.77871 0.0015185 0.7916 0.49729 0.0020409 0.42285 1.3091 1.3051 16.005 144.9787 0.00038406 -84.6997 0.16136
1.2654 0.98803 5.5178e-05 3.8182 0.012033 1.6652e-05 0.0011542 0.15926 0.00065845 0.15992 0.14598 0 0.036412 0.0389 0 0.90935 0.25533 0.069006 0.0096031 4.3043 0.059949 7.213e-05 0.83012 0.0053252 0.0060632 0.0016232 0.98379 0.98843 3.5333e-06 1.4134e-05 0.13229 0.72365 0.77937 0.0015175 0.79281 0.49746 0.0020397 0.42285 1.3109 1.307 16.0051 144.9787 0.00038302 -84.7068 0.16236
1.2664 0.98803 5.5177e-05 3.8182 0.012033 1.6665e-05 0.0011542 0.15932 0.00065845 0.15998 0.14603 0 0.036408 0.0389 0 0.90943 0.25536 0.069019 0.0096046 4.3047 0.059959 7.2143e-05 0.83011 0.0053256 0.0060636 0.0016213 0.98382 0.98852 3.529e-06 1.4116e-05 0.13229 0.72446 0.78002 0.0015166 0.79401 0.49762 0.0020385 0.42286 1.3128 1.3088 16.0051 144.9787 0.00038198 -84.7138 0.16336
1.2674 0.98803 5.5177e-05 3.8182 0.012033 1.6678e-05 0.0011542 0.15939 0.00065845 0.16004 0.14609 0 0.036404 0.0389 0 0.90951 0.2554 0.069032 0.0096062 4.3051 0.059968 7.2155e-05 0.8301 0.005326 0.006064 0.0016188 0.98384 0.9886 3.5246e-06 1.4099e-05 0.13229 0.72526 0.78068 0.0015157 0.79521 0.49779 0.0020373 0.42286 1.3146 1.3107 16.0052 144.9787 0.00038095 -84.7208 0.16436
1.2684 0.98803 5.5177e-05 3.8182 0.012033 1.6691e-05 0.0011542 0.15945 0.00065845 0.1601 0.14615 0 0.0364 0.0389 0 0.90959 0.25543 0.069045 0.0096078 4.3055 0.059978 7.2168e-05 0.83009 0.0053264 0.0060644 0.0016177 0.98387 0.98868 3.5203e-06 1.4082e-05 0.1323 0.72606 0.78132 0.0015148 0.7964 0.49796 0.0020361 0.42287 1.3165 1.3126 16.0052 144.9787 0.00037993 -84.7277 0.16536
1.2694 0.98803 5.5177e-05 3.8182 0.012033 1.6705e-05 0.0011542 0.15951 0.00065845 0.16016 0.1462 0 0.036397 0.0389 0 0.90967 0.25547 0.069058 0.0096093 4.3059 0.059988 7.218e-05 0.83008 0.0053269 0.0060648 0.0016143 0.98389 0.98876 3.516e-06 1.4065e-05 0.1323 0.72686 0.78197 0.0015138 0.79759 0.49813 0.0020349 0.42287 1.3183 1.3144 16.0053 144.9787 0.00037891 -84.7346 0.16636
1.2704 0.98803 5.5177e-05 3.8182 0.012033 1.6718e-05 0.0011542 0.15957 0.00065845 0.16022 0.14626 0 0.036393 0.0389 0 0.90975 0.25551 0.06907 0.0096109 4.3063 0.059997 7.2193e-05 0.83007 0.0053273 0.0060652 0.0016128 0.98392 0.98883 3.5118e-06 1.4048e-05 0.1323 0.72766 0.78261 0.0015129 0.79877 0.4983 0.0020337 0.42288 1.3201 1.3163 16.0053 144.9787 0.00037789 -84.7414 0.16736
1.2714 0.98803 5.5177e-05 3.8182 0.012033 1.6731e-05 0.0011542 0.15963 0.00065845 0.16028 0.14632 0 0.036389 0.0389 0 0.90983 0.25554 0.069083 0.0096125 4.3067 0.060007 7.2205e-05 0.83007 0.0053277 0.0060656 0.0016111 0.98394 0.9889 3.5076e-06 1.4031e-05 0.13231 0.72845 0.78325 0.001512 0.79994 0.49847 0.0020326 0.42288 1.322 1.3181 16.0054 144.9788 0.00037688 -84.7482 0.16836
1.2724 0.98803 5.5177e-05 3.8182 0.012033 1.6744e-05 0.0011542 0.15969 0.00065846 0.16034 0.14638 0 0.036385 0.0389 0 0.90991 0.25558 0.069096 0.0096141 4.3071 0.060017 7.2218e-05 0.83006 0.0053281 0.0060661 0.0016101 0.98397 0.98896 3.5034e-06 1.4014e-05 0.13231 0.72924 0.78388 0.0015112 0.80111 0.49864 0.0020314 0.42289 1.3238 1.32 16.0054 144.9788 0.00037588 -84.7549 0.16936
1.2734 0.98803 5.5177e-05 3.8182 0.012033 1.6757e-05 0.0011542 0.15975 0.00065846 0.16041 0.14643 0 0.036381 0.0389 0 0.90999 0.25561 0.069109 0.0096156 4.3076 0.060027 7.223e-05 0.83005 0.0053285 0.0060665 0.0016074 0.98399 0.98903 3.4993e-06 1.3998e-05 0.13231 0.73003 0.78451 0.0015103 0.80227 0.49881 0.0020302 0.42289 1.3256 1.3218 16.0055 144.9788 0.00037487 -84.7615 0.17036
1.2744 0.98803 5.5177e-05 3.8182 0.012033 1.677e-05 0.0011542 0.15981 0.00065846 0.16047 0.14649 0 0.036378 0.0389 0 0.91007 0.25565 0.069122 0.0096172 4.308 0.060036 7.2243e-05 0.83004 0.0053289 0.0060669 0.0016058 0.98402 0.98909 3.4952e-06 1.3981e-05 0.13232 0.73082 0.78514 0.0015094 0.80343 0.49898 0.0020291 0.4229 1.3274 1.3236 16.0055 144.9788 0.00037388 -84.7681 0.17136
1.2754 0.98803 5.5177e-05 3.8182 0.012033 1.6783e-05 0.0011542 0.15987 0.00065846 0.16053 0.14655 0 0.036374 0.0389 0 0.91015 0.25568 0.069135 0.0096188 4.3084 0.060046 7.2255e-05 0.83003 0.0053293 0.0060673 0.0016042 0.98404 0.98914 3.4912e-06 1.3965e-05 0.13232 0.7316 0.78577 0.0015085 0.80458 0.49915 0.002028 0.4229 1.3292 1.3254 16.0056 144.9788 0.00037289 -84.7747 0.17236
1.2764 0.98803 5.5177e-05 3.8182 0.012033 1.6797e-05 0.0011542 0.15993 0.00065846 0.16059 0.1466 0 0.03637 0.0389 0 0.91023 0.25572 0.069148 0.0096203 4.3088 0.060056 7.2268e-05 0.83002 0.0053297 0.0060677 0.0016029 0.98406 0.9892 3.4872e-06 1.3949e-05 0.13232 0.73238 0.78639 0.0015077 0.80572 0.49932 0.0020269 0.42291 1.3311 1.3273 16.0056 144.9788 0.0003719 -84.7812 0.17336
1.2774 0.98803 5.5177e-05 3.8182 0.012033 1.681e-05 0.0011542 0.15999 0.00065846 0.16065 0.14666 0 0.036366 0.0389 0 0.91031 0.25576 0.069161 0.0096219 4.3092 0.060065 7.228e-05 0.83001 0.0053302 0.0060682 0.0016007 0.98409 0.98925 3.4832e-06 1.3933e-05 0.13233 0.73316 0.787 0.0015068 0.80686 0.49949 0.0020257 0.42291 1.3329 1.3291 16.0057 144.9788 0.00037092 -84.7876 0.17436
1.2784 0.98803 5.5177e-05 3.8182 0.012033 1.6823e-05 0.0011542 0.16005 0.00065846 0.16071 0.14672 0 0.036362 0.0389 0 0.9104 0.25579 0.069174 0.0096235 4.3096 0.060075 7.2293e-05 0.83 0.0053306 0.0060686 0.0016001 0.98411 0.9893 3.4792e-06 1.3917e-05 0.13233 0.73394 0.78762 0.001506 0.80799 0.49966 0.0020246 0.42292 1.3347 1.3309 16.0057 144.9788 0.00036995 -84.794 0.17536
1.2794 0.98803 5.5177e-05 3.8182 0.012033 1.6836e-05 0.0011542 0.16012 0.00065846 0.16077 0.14677 0 0.036359 0.0389 0 0.91048 0.25583 0.069187 0.0096251 4.31 0.060085 7.2305e-05 0.82999 0.005331 0.006069 0.0015981 0.98413 0.98935 3.4753e-06 1.3902e-05 0.13233 0.73472 0.78823 0.0015052 0.80912 0.49983 0.0020235 0.42293 1.3365 1.3327 16.0058 144.9789 0.00036898 -84.8004 0.17636
1.2804 0.98803 5.5177e-05 3.8182 0.012033 1.6849e-05 0.0011542 0.16018 0.00065846 0.16083 0.14683 0 0.036355 0.0389 0 0.91056 0.25586 0.0692 0.0096266 4.3104 0.060095 7.2318e-05 0.82998 0.0053314 0.0060694 0.0015964 0.98416 0.98939 3.4715e-06 1.3886e-05 0.13234 0.73549 0.78884 0.0015043 0.81023 0.5 0.0020225 0.42293 1.3383 1.3345 16.0058 144.9789 0.00036801 -84.8067 0.17736
1.2814 0.98803 5.5177e-05 3.8182 0.012033 1.6862e-05 0.0011542 0.16024 0.00065846 0.16089 0.14689 0 0.036351 0.0389 0 0.91064 0.2559 0.069213 0.0096282 4.3108 0.060104 7.233e-05 0.82997 0.0053318 0.0060698 0.0015942 0.98418 0.98943 3.4676e-06 1.3871e-05 0.13234 0.73626 0.78944 0.0015035 0.81135 0.50017 0.0020214 0.42294 1.34 1.3363 16.0059 144.9789 0.00036705 -84.8129 0.17836
1.2824 0.98803 5.5176e-05 3.8182 0.012033 1.6875e-05 0.0011542 0.1603 0.00065847 0.16095 0.14694 0 0.036347 0.0389 0 0.91072 0.25594 0.069226 0.0096298 4.3112 0.060114 7.2343e-05 0.82996 0.0053322 0.0060703 0.0015932 0.9842 0.98947 3.4638e-06 1.3856e-05 0.13234 0.73703 0.79004 0.0015027 0.81246 0.50034 0.0020203 0.42294 1.3418 1.3381 16.0059 144.9789 0.00036609 -84.8191 0.17936
1.2834 0.98803 5.5176e-05 3.8182 0.012033 1.6888e-05 0.0011542 0.16036 0.00065847 0.16101 0.147 0 0.036344 0.0389 0 0.9108 0.25597 0.069239 0.0096314 4.3116 0.060124 7.2356e-05 0.82995 0.0053326 0.0060707 0.0015902 0.98422 0.98951 3.46e-06 1.3841e-05 0.13235 0.73779 0.79064 0.0015019 0.81356 0.5005 0.0020193 0.42295 1.3436 1.3399 16.0059 144.9789 0.00036514 -84.8253 0.18036
1.2844 0.98803 5.5176e-05 3.8182 0.012033 1.6902e-05 0.0011542 0.16042 0.00065847 0.16107 0.14706 0 0.03634 0.0389 0 0.91088 0.25601 0.069252 0.009633 4.312 0.060133 7.2368e-05 0.82994 0.0053331 0.0060711 0.0015889 0.98425 0.98955 3.4563e-06 1.3826e-05 0.13235 0.73855 0.79123 0.0015011 0.81465 0.50067 0.0020182 0.42296 1.3454 1.3417 16.006 144.9789 0.0003642 -84.8314 0.18136
1.2854 0.98803 5.5176e-05 3.8182 0.012033 1.6915e-05 0.0011542 0.16048 0.00065847 0.16113 0.14711 0 0.036336 0.0389 0 0.91096 0.25604 0.069265 0.0096345 4.3124 0.060143 7.2381e-05 0.82993 0.0053335 0.0060715 0.0015874 0.98427 0.98959 3.4526e-06 1.3811e-05 0.13235 0.73932 0.79182 0.0015003 0.81574 0.50084 0.0020172 0.42296 1.3472 1.3435 16.006 144.9789 0.00036326 -84.8375 0.18236
1.2864 0.98803 5.5176e-05 3.8182 0.012033 1.6928e-05 0.0011542 0.16054 0.00065847 0.16119 0.14717 0 0.036332 0.0389 0 0.91104 0.25608 0.069278 0.0096361 4.3129 0.060153 7.2393e-05 0.82992 0.0053339 0.0060719 0.0015865 0.98429 0.98962 3.4489e-06 1.3796e-05 0.13236 0.74007 0.79241 0.0014995 0.81683 0.50101 0.0020161 0.42297 1.3489 1.3453 16.0061 144.979 0.00036232 -84.8435 0.18336
1.2874 0.98803 5.5176e-05 3.8182 0.012033 1.6941e-05 0.0011542 0.1606 0.00065847 0.16125 0.14723 0 0.036329 0.0389 0 0.91112 0.25612 0.069291 0.0096377 4.3133 0.060163 7.2406e-05 0.82991 0.0053343 0.0060724 0.0015841 0.98431 0.98966 3.4453e-06 1.3781e-05 0.13236 0.74083 0.793 0.0014987 0.81791 0.50118 0.0020151 0.42297 1.3507 1.347 16.0061 144.979 0.00036139 -84.8494 0.18436
1.2884 0.98803 5.5176e-05 3.8182 0.012033 1.6954e-05 0.0011542 0.16066 0.00065847 0.16131 0.14728 0 0.036325 0.0389 0 0.9112 0.25615 0.069304 0.0096393 4.3137 0.060172 7.2418e-05 0.8299 0.0053347 0.0060728 0.0015827 0.98433 0.98969 3.4417e-06 1.3767e-05 0.13236 0.74158 0.79358 0.0014979 0.81898 0.50135 0.0020141 0.42298 1.3524 1.3488 16.0062 144.979 0.00036046 -84.8554 0.18536
1.2894 0.98803 5.5176e-05 3.8182 0.012033 1.6967e-05 0.0011542 0.16072 0.00065847 0.16137 0.14734 0 0.036321 0.0389 0 0.91128 0.25619 0.069317 0.0096408 4.3141 0.060182 7.2431e-05 0.82989 0.0053351 0.0060732 0.0015813 0.98435 0.98972 3.4381e-06 1.3753e-05 0.13237 0.74233 0.79416 0.0014972 0.82005 0.50152 0.0020131 0.42299 1.3542 1.3506 16.0062 144.979 0.00035953 -84.8613 0.18636
1.2904 0.98803 5.5176e-05 3.8182 0.012033 1.698e-05 0.0011542 0.16078 0.00065847 0.16143 0.1474 0 0.036317 0.0389 0 0.91137 0.25622 0.06933 0.0096424 4.3145 0.060192 7.2444e-05 0.82988 0.0053356 0.0060736 0.0015801 0.98438 0.98975 3.4345e-06 1.3738e-05 0.13237 0.74308 0.79473 0.0014964 0.82111 0.50169 0.0020121 0.42299 1.3559 1.3523 16.0062 144.979 0.00035862 -84.8671 0.18736
1.2914 0.98803 5.5176e-05 3.8182 0.012033 1.6993e-05 0.0011542 0.16084 0.00065847 0.16149 0.14745 0 0.036314 0.0389 0 0.91145 0.25626 0.069343 0.009644 4.3149 0.060202 7.2456e-05 0.82987 0.005336 0.0060741 0.0015783 0.9844 0.98978 3.431e-06 1.3724e-05 0.13238 0.74383 0.7953 0.0014956 0.82216 0.50186 0.0020111 0.423 1.3577 1.3541 16.0063 144.979 0.0003577 -84.8729 0.18836
1.2924 0.98803 5.5176e-05 3.8182 0.012033 1.7007e-05 0.0011542 0.1609 0.00065848 0.16155 0.14751 0 0.03631 0.0389 0 0.91153 0.2563 0.069356 0.0096456 4.3153 0.060211 7.2469e-05 0.82986 0.0053364 0.0060745 0.0015775 0.98442 0.98981 3.4275e-06 1.371e-05 0.13238 0.74457 0.79587 0.0014949 0.82321 0.50203 0.0020101 0.42301 1.3594 1.3559 16.0063 144.979 0.00035679 -84.8786 0.18936
1.2934 0.98803 5.5176e-05 3.8182 0.012033 1.702e-05 0.0011542 0.16096 0.00065848 0.16161 0.14756 0 0.036306 0.0389 0 0.91161 0.25633 0.069369 0.0096472 4.3158 0.060221 7.2481e-05 0.82985 0.0053368 0.0060749 0.0015747 0.98444 0.98984 3.4241e-06 1.3697e-05 0.13238 0.74532 0.79644 0.0014941 0.82426 0.5022 0.0020091 0.42301 1.3612 1.3576 16.0064 144.9791 0.00035589 -84.8843 0.19036
1.2944 0.98803 5.5176e-05 3.8182 0.012033 1.7033e-05 0.0011542 0.16102 0.00065848 0.16167 0.14762 0 0.036303 0.0389 0 0.91169 0.25637 0.069382 0.0096488 4.3162 0.060231 7.2494e-05 0.82984 0.0053372 0.0060753 0.0015734 0.98446 0.98986 3.4206e-06 1.3683e-05 0.13239 0.74606 0.797 0.0014934 0.82529 0.50236 0.0020082 0.42302 1.3629 1.3594 16.0064 144.9791 0.00035499 -84.89 0.19136
1.2954 0.98803 5.5176e-05 3.8182 0.012033 1.7046e-05 0.0011542 0.16108 0.00065848 0.16173 0.14768 0 0.036299 0.0389 0 0.91177 0.2564 0.069395 0.0096503 4.3166 0.060241 7.2507e-05 0.82983 0.0053377 0.0060758 0.0015721 0.98448 0.98989 3.4172e-06 1.3669e-05 0.13239 0.74679 0.79757 0.0014927 0.82633 0.50253 0.0020072 0.42303 1.3646 1.3611 16.0064 144.9791 0.00035409 -84.8956 0.19236
1.2964 0.98803 5.5176e-05 3.8182 0.012033 1.7059e-05 0.0011542 0.16114 0.00065848 0.16179 0.14773 0 0.036295 0.0389 0 0.91185 0.25644 0.069408 0.0096519 4.317 0.060251 7.2519e-05 0.82982 0.0053381 0.0060762 0.0015712 0.9845 0.98991 3.4139e-06 1.3656e-05 0.13239 0.74753 0.79812 0.0014919 0.82735 0.5027 0.0020063 0.42303 1.3664 1.3628 16.0065 144.9791 0.0003532 -84.9012 0.19336
1.2974 0.98803 5.5176e-05 3.8182 0.012033 1.7072e-05 0.0011542 0.1612 0.00065848 0.16185 0.14779 0 0.036291 0.0389 0 0.91193 0.25648 0.069421 0.0096535 4.3174 0.06026 7.2532e-05 0.82981 0.0053385 0.0060766 0.0015692 0.98452 0.98993 3.4105e-06 1.3642e-05 0.1324 0.74826 0.79868 0.0014912 0.82837 0.50287 0.0020053 0.42304 1.3681 1.3646 16.0065 144.9791 0.00035231 -84.9067 0.19436
1.2984 0.98803 5.5175e-05 3.8182 0.012033 1.7085e-05 0.0011542 0.16126 0.00065848 0.16191 0.14784 0 0.036288 0.0389 0 0.91201 0.25651 0.069434 0.0096551 4.3178 0.06027 7.2544e-05 0.8298 0.0053389 0.006077 0.001569 0.98454 0.98996 3.4072e-06 1.3629e-05 0.1324 0.74899 0.79923 0.0014905 0.82939 0.50304 0.0020044 0.42305 1.3698 1.3663 16.0066 144.9791 0.00035143 -84.9122 0.19536
1.2994 0.98803 5.5175e-05 3.8182 0.012033 1.7099e-05 0.0011542 0.16132 0.00065848 0.16197 0.1479 0 0.036284 0.0389 0 0.9121 0.25655 0.069447 0.0096567 4.3182 0.06028 7.2557e-05 0.82979 0.0053393 0.0060775 0.0015674 0.98456 0.98998 3.4039e-06 1.3616e-05 0.1324 0.74972 0.79978 0.0014898 0.8304 0.50321 0.0020034 0.42305 1.3715 1.368 16.0066 144.9791 0.00035055 -84.9177 0.19636
1.3004 0.98803 5.5175e-05 3.8182 0.012033 1.7112e-05 0.0011542 0.16137 0.00065848 0.16203 0.14796 0 0.03628 0.0389 0 0.91218 0.25659 0.06946 0.0096583 4.3187 0.06029 7.257e-05 0.82978 0.0053398 0.0060779 0.0015658 0.98457 0.99 3.4007e-06 1.3603e-05 0.13241 0.75045 0.80033 0.0014891 0.83141 0.50338 0.0020025 0.42306 1.3732 1.3697 16.0066 144.9792 0.00034967 -84.9231 0.19736
1.3014 0.98803 5.5175e-05 3.8182 0.012033 1.7125e-05 0.0011542 0.16143 0.00065848 0.16209 0.14801 0 0.036277 0.0389 0 0.91226 0.25662 0.069473 0.0096598 4.3191 0.060299 7.2582e-05 0.82977 0.0053402 0.0060783 0.0015638 0.98459 0.99002 3.3975e-06 1.359e-05 0.13241 0.75117 0.80087 0.0014884 0.83241 0.50355 0.0020016 0.42307 1.3749 1.3715 16.0067 144.9792 0.0003488 -84.9284 0.19836
1.3024 0.98803 5.5175e-05 3.8182 0.012033 1.7138e-05 0.0011542 0.16149 0.00065849 0.16215 0.14807 0 0.036273 0.0389 0 0.91234 0.25666 0.069486 0.0096614 4.3195 0.060309 7.2595e-05 0.82976 0.0053406 0.0060788 0.0015631 0.98461 0.99004 3.3943e-06 1.3577e-05 0.13241 0.75189 0.80141 0.0014877 0.8334 0.50371 0.0020007 0.42307 1.3766 1.3732 16.0067 144.9792 0.00034794 -84.9338 0.19936
1.3034 0.98803 5.5175e-05 3.8182 0.012033 1.7151e-05 0.0011542 0.16155 0.00065849 0.16221 0.14812 0 0.036269 0.0389 0 0.91242 0.25669 0.069499 0.009663 4.3199 0.060319 7.2608e-05 0.82975 0.005341 0.0060792 0.0015603 0.98463 0.99006 3.3911e-06 1.3565e-05 0.13242 0.75261 0.80195 0.001487 0.83439 0.50388 0.0019998 0.42308 1.3783 1.3749 16.0068 144.9792 0.00034708 -84.9391 0.20036
1.3044 0.98803 5.5175e-05 3.8182 0.012033 1.7164e-05 0.0011542 0.16161 0.00065849 0.16227 0.14818 0 0.036266 0.0389 0 0.9125 0.25673 0.069512 0.0096646 4.3203 0.060329 7.262e-05 0.82974 0.0053414 0.0060796 0.0015592 0.98465 0.99008 3.3879e-06 1.3552e-05 0.13242 0.75333 0.80248 0.0014863 0.83537 0.50405 0.0019989 0.42309 1.38 1.3766 16.0068 144.9792 0.00034622 -84.9443 0.20136
1.3054 0.98803 5.5175e-05 3.8182 0.012033 1.7177e-05 0.0011542 0.16167 0.00065849 0.16233 0.14823 0 0.036262 0.0389 0 0.91258 0.25677 0.069525 0.0096662 4.3208 0.060339 7.2633e-05 0.82973 0.0053419 0.00608 0.001558 0.98467 0.9901 3.3848e-06 1.354e-05 0.13242 0.75405 0.80302 0.0014856 0.83635 0.50422 0.001998 0.4231 1.3817 1.3783 16.0068 144.9792 0.00034537 -84.9495 0.20236
1.3064 0.98803 5.5175e-05 3.8182 0.012033 1.719e-05 0.0011542 0.16173 0.00065849 0.16238 0.14829 0 0.036258 0.0389 0 0.91266 0.2568 0.069538 0.0096678 4.3212 0.060348 7.2646e-05 0.82972 0.0053423 0.0060805 0.0015573 0.98469 0.99012 3.3817e-06 1.3527e-05 0.13243 0.75476 0.80355 0.001485 0.83732 0.50439 0.0019972 0.4231 1.3834 1.38 16.0069 144.9793 0.00034452 -84.9547 0.20336
1.3074 0.98803 5.5175e-05 3.8182 0.012033 1.7204e-05 0.0011542 0.16179 0.00065849 0.16244 0.14834 0 0.036255 0.0389 0 0.91275 0.25684 0.069551 0.0096694 4.3216 0.060358 7.2658e-05 0.82971 0.0053427 0.0060809 0.0015553 0.9847 0.99013 3.3787e-06 1.3515e-05 0.13243 0.75547 0.80407 0.0014843 0.83829 0.50456 0.0019963 0.42311 1.3851 1.3817 16.0069 144.9793 0.00034367 -84.9598 0.20436
1.3084 0.98803 5.5175e-05 3.8182 0.012033 1.7217e-05 0.0011542 0.16185 0.00065849 0.1625 0.1484 0 0.036251 0.0389 0 0.91283 0.25687 0.069564 0.0096709 4.322 0.060368 7.2671e-05 0.8297 0.0053431 0.0060813 0.0015541 0.98472 0.99015 3.3756e-06 1.3503e-05 0.13243 0.75618 0.8046 0.0014836 0.83925 0.50473 0.0019954 0.42312 1.3867 1.3834 16.0069 144.9793 0.00034283 -84.9649 0.20536
1.3094 0.98803 5.5175e-05 3.8182 0.012033 1.723e-05 0.0011542 0.16191 0.00065849 0.16256 0.14846 0 0.036247 0.0389 0 0.91291 0.25691 0.069578 0.0096725 4.3224 0.060378 7.2684e-05 0.82969 0.0053436 0.0060818 0.001553 0.98474 0.99017 3.3726e-06 1.3491e-05 0.13244 0.75688 0.80512 0.001483 0.84021 0.50489 0.0019946 0.42312 1.3884 1.385 16.007 144.9793 0.000342 -84.9699 0.20636
1.3104 0.98803 5.5175e-05 3.8182 0.012033 1.7243e-05 0.0011542 0.16197 0.00065849 0.16262 0.14851 0 0.036244 0.0389 0 0.91299 0.25695 0.069591 0.0096741 4.3229 0.060388 7.2696e-05 0.82969 0.005344 0.0060822 0.0015519 0.98476 0.99019 3.3696e-06 1.3479e-05 0.13244 0.75759 0.80564 0.0014823 0.84116 0.50506 0.0019937 0.42313 1.3901 1.3867 16.007 144.9793 0.00034116 -84.975 0.20736
1.3114 0.98803 5.5175e-05 3.8182 0.012033 1.7256e-05 0.0011542 0.16203 0.00065849 0.16268 0.14857 0 0.03624 0.0389 0 0.91307 0.25698 0.069604 0.0096757 4.3233 0.060397 7.2709e-05 0.82968 0.0053444 0.0060826 0.0015505 0.98477 0.9902 3.3666e-06 1.3467e-05 0.13245 0.75829 0.80615 0.0014817 0.8421 0.50523 0.0019929 0.42314 1.3917 1.3884 16.0071 144.9793 0.00034033 -84.9799 0.20836
1.3124 0.98803 5.5175e-05 3.8182 0.012032 1.7269e-05 0.0011542 0.16209 0.0006585 0.16274 0.14862 0 0.036236 0.0389 0 0.91315 0.25702 0.069617 0.0096773 4.3237 0.060407 7.2722e-05 0.82967 0.0053448 0.0060831 0.0015496 0.98479 0.99022 3.3637e-06 1.3455e-05 0.13245 0.75899 0.80667 0.0014811 0.84304 0.5054 0.001992 0.42315 1.3934 1.3901 16.0071 144.9793 0.00033951 -84.9849 0.20936
1.3134 0.98803 5.5175e-05 3.8182 0.012032 1.7282e-05 0.0011542 0.16214 0.0006585 0.1628 0.14868 0 0.036233 0.0389 0 0.91324 0.25706 0.06963 0.0096789 4.3241 0.060417 7.2734e-05 0.82966 0.0053453 0.0060835 0.0015477 0.98481 0.99023 3.3608e-06 1.3443e-05 0.13245 0.75969 0.80718 0.0014804 0.84398 0.50557 0.0019912 0.42316 1.395 1.3917 16.0071 144.9794 0.00033869 -84.9898 0.21036
1.3144 0.98803 5.5174e-05 3.8182 0.012032 1.7295e-05 0.0011542 0.1622 0.0006585 0.16286 0.14873 0 0.036229 0.0389 0 0.91332 0.25709 0.069643 0.0096805 4.3246 0.060427 7.2747e-05 0.82965 0.0053457 0.0060839 0.0015477 0.98483 0.99025 3.3579e-06 1.3432e-05 0.13246 0.76038 0.80769 0.0014798 0.84491 0.50574 0.0019904 0.42316 1.3967 1.3934 16.0072 144.9794 0.00033787 -84.9946 0.21136
1.3154 0.98803 5.5174e-05 3.8182 0.012032 1.7309e-05 0.0011542 0.16226 0.0006585 0.16292 0.14879 0 0.036225 0.0389 0 0.9134 0.25713 0.069656 0.0096821 4.325 0.060437 7.276e-05 0.82964 0.0053461 0.0060844 0.0015462 0.98484 0.99026 3.355e-06 1.342e-05 0.13246 0.76108 0.80819 0.0014792 0.84583 0.50591 0.0019896 0.42317 1.3983 1.395 16.0072 144.9794 0.00033706 -84.9995 0.21236
1.3164 0.98803 5.5174e-05 3.8182 0.012032 1.7322e-05 0.0011542 0.16232 0.0006585 0.16297 0.14884 0 0.036222 0.0389 0 0.91348 0.25717 0.069669 0.0096837 4.3254 0.060447 7.2772e-05 0.82963 0.0053465 0.0060848 0.0015448 0.98486 0.99028 3.3522e-06 1.3409e-05 0.13246 0.76177 0.8087 0.0014785 0.84675 0.50607 0.0019887 0.42318 1.4 1.3967 16.0072 144.9794 0.00033625 -85.0042 0.21336
1.3174 0.98803 5.5174e-05 3.8182 0.012032 1.7335e-05 0.0011542 0.16238 0.0006585 0.16303 0.1489 0 0.036218 0.0389 0 0.91356 0.2572 0.069682 0.0096853 4.3258 0.060456 7.2785e-05 0.82962 0.005347 0.0060852 0.001543 0.98488 0.99029 3.3494e-06 1.3398e-05 0.13247 0.76246 0.8092 0.0014779 0.84767 0.50624 0.0019879 0.42319 1.4016 1.3983 16.0073 144.9794 0.00033545 -85.009 0.21436
1.3184 0.98803 5.5174e-05 3.8182 0.012032 1.7348e-05 0.0011542 0.16244 0.0006585 0.16309 0.14895 0 0.036214 0.0389 0 0.91364 0.25724 0.069695 0.0096868 4.3263 0.060466 7.2798e-05 0.82961 0.0053474 0.0060857 0.0015423 0.98489 0.9903 3.3466e-06 1.3387e-05 0.13247 0.76315 0.8097 0.0014773 0.84858 0.50641 0.0019871 0.42319 1.4033 1.4 16.0073 144.9794 0.00033465 -85.0137 0.21536
1.3194 0.98803 5.5174e-05 3.8182 0.012032 1.7361e-05 0.0011542 0.1625 0.0006585 0.16315 0.14901 0 0.036211 0.0389 0 0.91373 0.25727 0.069709 0.0096884 4.3267 0.060476 7.281e-05 0.8296 0.0053478 0.0060861 0.00154 0.98491 0.99032 3.3438e-06 1.3375e-05 0.13247 0.76383 0.81019 0.0014767 0.84948 0.50658 0.0019864 0.4232 1.4049 1.4016 16.0073 144.9794 0.00033385 -85.0184 0.21636
1.3204 0.98803 5.5174e-05 3.8182 0.012032 1.7374e-05 0.0011542 0.16255 0.0006585 0.16321 0.14906 0 0.036207 0.0389 0 0.91381 0.25731 0.069722 0.00969 4.3271 0.060486 7.2823e-05 0.82959 0.0053483 0.0060865 0.001539 0.98492 0.99033 3.341e-06 1.3364e-05 0.13248 0.76451 0.81069 0.0014761 0.85038 0.50675 0.0019856 0.42321 1.4065 1.4033 16.0074 144.9795 0.00033306 -85.0231 0.21736
1.3214 0.98803 5.5174e-05 3.8182 0.012032 1.7387e-05 0.0011542 0.16261 0.0006585 0.16327 0.14912 0 0.036204 0.0389 0 0.91389 0.25735 0.069735 0.0096916 4.3275 0.060496 7.2836e-05 0.82958 0.0053487 0.006087 0.001538 0.98494 0.99034 3.3383e-06 1.3353e-05 0.13248 0.76519 0.81118 0.0014755 0.85128 0.50691 0.0019848 0.42322 1.4081 1.4049 16.0074 144.9795 0.00033227 -85.0277 0.21836
1.3224 0.98803 5.5174e-05 3.8182 0.012032 1.7401e-05 0.0011542 0.16267 0.00065851 0.16333 0.14917 0 0.0362 0.0389 0 0.91397 0.25738 0.069748 0.0096932 4.328 0.060506 7.2849e-05 0.82957 0.0053491 0.0060874 0.0015373 0.98496 0.99036 3.3356e-06 1.3343e-05 0.13248 0.76587 0.81167 0.0014749 0.85216 0.50708 0.001984 0.42323 1.4097 1.4065 16.0074 144.9795 0.00033148 -85.0322 0.21936
1.3234 0.98803 5.5174e-05 3.8182 0.012032 1.7414e-05 0.0011542 0.16273 0.00065851 0.16338 0.14923 0 0.036196 0.0389 0 0.91405 0.25742 0.069761 0.0096948 4.3284 0.060515 7.2861e-05 0.82956 0.0053495 0.0060878 0.0015357 0.98497 0.99037 3.3329e-06 1.3332e-05 0.13249 0.76655 0.81215 0.0014743 0.85305 0.50725 0.0019832 0.42324 1.4114 1.4082 16.0075 144.9795 0.0003307 -85.0368 0.22036
1.3244 0.98803 5.5174e-05 3.8182 0.012032 1.7427e-05 0.0011542 0.16279 0.00065851 0.16344 0.14928 0 0.036193 0.0389 0 0.91413 0.25746 0.069774 0.0096964 4.3288 0.060525 7.2874e-05 0.82955 0.00535 0.0060883 0.0015355 0.98499 0.99038 3.3303e-06 1.3321e-05 0.13249 0.76722 0.81264 0.0014738 0.85393 0.50742 0.0019825 0.42324 1.413 1.4098 16.0075 144.9795 0.00032992 -85.0413 0.22136
1.3254 0.98803 5.5174e-05 3.8182 0.012032 1.744e-05 0.0011542 0.16285 0.00065851 0.1635 0.14934 0 0.036189 0.0389 0 0.91422 0.25749 0.069787 0.009698 4.3292 0.060535 7.2887e-05 0.82954 0.0053504 0.0060887 0.0015342 0.985 0.99039 3.3276e-06 1.3311e-05 0.13249 0.7679 0.81312 0.0014732 0.8548 0.50759 0.0019817 0.42325 1.4146 1.4114 16.0075 144.9795 0.00032915 -85.0458 0.22236
1.3264 0.98803 5.5174e-05 3.8182 0.012032 1.7453e-05 0.0011542 0.16291 0.00065851 0.16356 0.14939 0 0.036186 0.0389 0 0.9143 0.25753 0.069801 0.0096996 4.3297 0.060545 7.29e-05 0.82953 0.0053508 0.0060891 0.0015329 0.98502 0.99041 3.325e-06 1.33e-05 0.1325 0.76857 0.8136 0.0014726 0.85567 0.50776 0.001981 0.42326 1.4162 1.413 16.0075 144.9796 0.00032838 -85.0502 0.22336
1.3274 0.98803 5.5174e-05 3.8182 0.012032 1.7466e-05 0.0011543 0.16296 0.00065851 0.16362 0.14945 0 0.036182 0.0389 0 0.91438 0.25757 0.069814 0.0097012 4.3301 0.060555 7.2912e-05 0.82952 0.0053513 0.0060896 0.0015314 0.98503 0.99042 3.3224e-06 1.329e-05 0.1325 0.76923 0.81407 0.001472 0.85654 0.50792 0.0019802 0.42327 1.4178 1.4146 16.0076 144.9796 0.00032761 -85.0546 0.22436
1.3284 0.98803 5.5174e-05 3.8182 0.012032 1.7479e-05 0.0011543 0.16302 0.00065851 0.16368 0.1495 0 0.036178 0.0389 0 0.91446 0.2576 0.069827 0.0097028 4.3305 0.060565 7.2925e-05 0.82951 0.0053517 0.00609 0.0015306 0.98505 0.99043 3.3199e-06 1.328e-05 0.13251 0.7699 0.81455 0.0014715 0.8574 0.50809 0.0019795 0.42328 1.4194 1.4162 16.0076 144.9796 0.00032685 -85.059 0.22536
1.3294 0.98803 5.5174e-05 3.8182 0.012032 1.7492e-05 0.0011543 0.16308 0.00065851 0.16373 0.14955 0 0.036175 0.0389 0 0.91454 0.25764 0.06984 0.0097044 4.331 0.060575 7.2938e-05 0.8295 0.0053521 0.0060905 0.0015286 0.98506 0.99044 3.3173e-06 1.3269e-05 0.13251 0.77056 0.81502 0.0014709 0.85825 0.50826 0.0019788 0.42329 1.4209 1.4178 16.0076 144.9796 0.00032609 -85.0634 0.22636
1.3304 0.98803 5.5173e-05 3.8182 0.012032 1.7506e-05 0.0011543 0.16314 0.00065851 0.16379 0.14961 0 0.036171 0.0389 0 0.91463 0.25768 0.069853 0.009706 4.3314 0.060585 7.295e-05 0.82949 0.0053526 0.0060909 0.0015277 0.98508 0.99045 3.3148e-06 1.3259e-05 0.13251 0.77123 0.81549 0.0014704 0.8591 0.50843 0.001978 0.42329 1.4225 1.4194 16.0077 144.9796 0.00032533 -85.0677 0.22736
1.3314 0.98803 5.5173e-05 3.8182 0.012032 1.7519e-05 0.0011543 0.1632 0.00065851 0.16385 0.14966 0 0.036168 0.0389 0 0.91471 0.25771 0.069866 0.0097076 4.3318 0.060594 7.2963e-05 0.82948 0.005353 0.0060913 0.0015267 0.98509 0.99046 3.3123e-06 1.3249e-05 0.13252 0.77189 0.81596 0.0014698 0.85995 0.50859 0.0019773 0.4233 1.4241 1.421 16.0077 144.9796 0.00032458 -85.0719 0.22836
1.3324 0.98803 5.5173e-05 3.8182 0.012032 1.7532e-05 0.0011543 0.16325 0.00065851 0.16391 0.14972 0 0.036164 0.0389 0 0.91479 0.25775 0.06988 0.0097092 4.3323 0.060604 7.2976e-05 0.82947 0.0053534 0.0060918 0.001526 0.98511 0.99047 3.3098e-06 1.3239e-05 0.13252 0.77255 0.81642 0.0014693 0.86079 0.50876 0.0019766 0.42331 1.4257 1.4226 16.0077 144.9797 0.00032383 -85.0762 0.22936
1.3334 0.98803 5.5173e-05 3.8182 0.012032 1.7545e-05 0.0011543 0.16331 0.00065852 0.16397 0.14977 0 0.03616 0.0389 0 0.91487 0.25779 0.069893 0.0097108 4.3327 0.060614 7.2989e-05 0.82946 0.0053539 0.0060922 0.0015246 0.98512 0.99048 3.3073e-06 1.3229e-05 0.13252 0.7732 0.81689 0.0014687 0.86162 0.50893 0.0019759 0.42332 1.4273 1.4242 16.0078 144.9797 0.00032309 -85.0804 0.23036
1.3344 0.98803 5.5173e-05 3.8182 0.012032 1.7558e-05 0.0011543 0.16337 0.00065852 0.16402 0.14983 0 0.036157 0.0389 0 0.91495 0.25782 0.069906 0.0097124 4.3331 0.060624 7.3002e-05 0.82945 0.0053543 0.0060927 0.0015243 0.98514 0.99049 3.3049e-06 1.322e-05 0.13253 0.77386 0.81735 0.0014682 0.86245 0.5091 0.0019752 0.42333 1.4288 1.4258 16.0078 144.9797 0.00032235 -85.0846 0.23136
1.3354 0.98803 5.5173e-05 3.8182 0.012032 1.7571e-05 0.0011543 0.16343 0.00065852 0.16408 0.14988 0 0.036153 0.0389 0 0.91504 0.25786 0.069919 0.009714 4.3336 0.060634 7.3014e-05 0.82944 0.0053547 0.0060931 0.0015232 0.98515 0.99051 3.3024e-06 1.321e-05 0.13253 0.77451 0.81781 0.0014676 0.86328 0.50927 0.0019745 0.42334 1.4304 1.4273 16.0078 144.9797 0.00032161 -85.0887 0.23236
1.3364 0.98803 5.5173e-05 3.8182 0.012032 1.7584e-05 0.0011543 0.16349 0.00065852 0.16414 0.14994 0 0.03615 0.0389 0 0.91512 0.25789 0.069932 0.0097156 4.334 0.060644 7.3027e-05 0.82943 0.0053552 0.0060935 0.001522 0.98516 0.99052 3.3e-06 1.32e-05 0.13253 0.77516 0.81826 0.0014671 0.8641 0.50943 0.0019738 0.42335 1.432 1.4289 16.0078 144.9797 0.00032087 -85.0929 0.23336
1.3374 0.98803 5.5173e-05 3.8182 0.012032 1.7597e-05 0.0011543 0.16354 0.00065852 0.1642 0.14999 0 0.036146 0.0389 0 0.9152 0.25793 0.069946 0.0097172 4.3344 0.060654 7.304e-05 0.82942 0.0053556 0.006094 0.0015206 0.98518 0.99053 3.2976e-06 1.3191e-05 0.13254 0.77581 0.81872 0.0014666 0.86492 0.5096 0.0019731 0.42335 1.4335 1.4305 16.0079 144.9797 0.00032014 -85.097 0.23436
1.3384 0.98803 5.5173e-05 3.8182 0.012032 1.7611e-05 0.0011543 0.1636 0.00065852 0.16425 0.15004 0 0.036143 0.0389 0 0.91528 0.25797 0.069959 0.0097188 4.3349 0.060664 7.3053e-05 0.82941 0.005356 0.0060944 0.0015199 0.98519 0.99054 3.2953e-06 1.3181e-05 0.13254 0.77645 0.81917 0.0014661 0.86573 0.50977 0.0019724 0.42336 1.4351 1.432 16.0079 144.9797 0.00031941 -85.101 0.23536
1.3394 0.98803 5.5173e-05 3.8182 0.012032 1.7624e-05 0.0011543 0.16366 0.00065852 0.16431 0.1501 0 0.036139 0.0389 0 0.91536 0.258 0.069972 0.0097204 4.3353 0.060674 7.3065e-05 0.8294 0.0053565 0.0060949 0.0015182 0.98521 0.99055 3.2929e-06 1.3172e-05 0.13255 0.77709 0.81962 0.0014656 0.86654 0.50994 0.0019718 0.42337 1.4366 1.4336 16.0079 144.9798 0.00031869 -85.1051 0.23636
1.3404 0.98803 5.5173e-05 3.8182 0.012032 1.7637e-05 0.0011543 0.16372 0.00065852 0.16437 0.15015 0 0.036135 0.0389 0 0.91545 0.25804 0.069985 0.009722 4.3357 0.060683 7.3078e-05 0.82939 0.0053569 0.0060953 0.0015184 0.98522 0.99056 3.2906e-06 1.3162e-05 0.13255 0.77774 0.82007 0.001465 0.86734 0.5101 0.0019711 0.42338 1.4382 1.4351 16.008 144.9798 0.00031797 -85.1091 0.23736
1.3414 0.98803 5.5173e-05 3.8182 0.012032 1.765e-05 0.0011543 0.16377 0.00065852 0.16443 0.15021 0 0.036132 0.0389 0 0.91553 0.25808 0.069998 0.0097236 4.3362 0.060693 7.3091e-05 0.82938 0.0053573 0.0060957 0.0015172 0.98523 0.99056 3.2883e-06 1.3153e-05 0.13255 0.77838 0.82051 0.0014645 0.86814 0.51027 0.0019704 0.42339 1.4397 1.4367 16.008 144.9798 0.00031725 -85.113 0.23836
1.3424 0.98803 5.5173e-05 3.8182 0.012032 1.7663e-05 0.0011543 0.16383 0.00065852 0.16449 0.15026 0 0.036128 0.0389 0 0.91561 0.25811 0.070012 0.0097252 4.3366 0.060703 7.3104e-05 0.82937 0.0053578 0.0060962 0.001516 0.98525 0.99057 3.286e-06 1.3144e-05 0.13256 0.77901 0.82096 0.001464 0.86893 0.51044 0.0019698 0.4234 1.4412 1.4382 16.008 144.9798 0.00031654 -85.117 0.23936
1.3434 0.98803 5.5173e-05 3.8182 0.012032 1.7676e-05 0.0011543 0.16389 0.00065852 0.16454 0.15031 0 0.036125 0.0389 0 0.91569 0.25815 0.070025 0.0097268 4.337 0.060713 7.3117e-05 0.82936 0.0053582 0.0060966 0.0015147 0.98526 0.99058 3.2837e-06 1.3135e-05 0.13256 0.77965 0.8214 0.0014635 0.86972 0.51061 0.0019691 0.42341 1.4428 1.4398 16.008 144.9798 0.00031583 -85.1209 0.24036
1.3444 0.98803 5.5173e-05 3.8182 0.012032 1.7689e-05 0.0011543 0.16395 0.00065853 0.1646 0.15037 0 0.036121 0.0389 0 0.91578 0.25819 0.070038 0.0097284 4.3375 0.060723 7.3129e-05 0.82935 0.0053586 0.0060971 0.0015138 0.98527 0.99059 3.2814e-06 1.3126e-05 0.13256 0.78028 0.82184 0.001463 0.8705 0.51077 0.0019685 0.42342 1.4443 1.4413 16.0081 144.9798 0.00031512 -85.1248 0.24136
1.3454 0.98803 5.5172e-05 3.8182 0.012032 1.7702e-05 0.0011543 0.164 0.00065853 0.16466 0.15042 0 0.036118 0.0389 0 0.91586 0.25822 0.070051 0.00973 4.3379 0.060733 7.3142e-05 0.82934 0.0053591 0.0060975 0.0015128 0.98528 0.9906 3.2792e-06 1.3117e-05 0.13257 0.78092 0.82227 0.0014625 0.87128 0.51094 0.0019678 0.42343 1.4458 1.4429 16.0081 144.9799 0.00031442 -85.1286 0.24236
1.3464 0.98803 5.5172e-05 3.8182 0.012032 1.7716e-05 0.0011543 0.16406 0.00065853 0.16471 0.15048 0 0.036114 0.0389 0 0.91594 0.25826 0.070064 0.0097316 4.3384 0.060743 7.3155e-05 0.82933 0.0053595 0.006098 0.001512 0.9853 0.99061 3.277e-06 1.3108e-05 0.13257 0.78155 0.82271 0.001462 0.87206 0.51111 0.0019672 0.42344 1.4473 1.4444 16.0081 144.9799 0.00031372 -85.1325 0.24336
1.3474 0.98803 5.5172e-05 3.8182 0.012032 1.7729e-05 0.0011543 0.16412 0.00065853 0.16477 0.15053 0 0.036111 0.0389 0 0.91602 0.2583 0.070078 0.0097332 4.3388 0.060753 7.3168e-05 0.82932 0.00536 0.0060984 0.0015105 0.98531 0.99062 3.2748e-06 1.3099e-05 0.13257 0.78218 0.82314 0.0014616 0.87283 0.51128 0.0019665 0.42345 1.4489 1.4459 16.0081 144.9799 0.00031302 -85.1363 0.24436
1.3484 0.98803 5.5172e-05 3.8182 0.012032 1.7742e-05 0.0011543 0.16418 0.00065853 0.16483 0.15058 0 0.036107 0.0389 0 0.91611 0.25833 0.070091 0.0097348 4.3392 0.060763 7.3181e-05 0.82931 0.0053604 0.0060989 0.0015104 0.98532 0.99063 3.2726e-06 1.3091e-05 0.13258 0.7828 0.82357 0.0014611 0.8736 0.51144 0.0019659 0.42345 1.4504 1.4474 16.0082 144.9799 0.00031233 -85.14 0.24536
1.3494 0.98803 5.5172e-05 3.8182 0.012032 1.7755e-05 0.0011543 0.16423 0.00065853 0.16489 0.15064 0 0.036104 0.0389 0 0.91619 0.25837 0.070104 0.0097364 4.3397 0.060773 7.3194e-05 0.8293 0.0053608 0.0060993 0.0015093 0.98534 0.99064 3.2704e-06 1.3082e-05 0.13258 0.78343 0.824 0.0014606 0.87436 0.51161 0.0019653 0.42346 1.4519 1.449 16.0082 144.9799 0.00031164 -85.1438 0.24636
1.3504 0.98803 5.5172e-05 3.8182 0.012032 1.7768e-05 0.0011543 0.16429 0.00065853 0.16494 0.15069 0 0.0361 0.0389 0 0.91627 0.25841 0.070117 0.009738 4.3401 0.060783 7.3206e-05 0.82929 0.0053613 0.0060997 0.0015078 0.98535 0.99065 3.2683e-06 1.3073e-05 0.13258 0.78405 0.82443 0.0014601 0.87512 0.51178 0.0019647 0.42347 1.4534 1.4505 16.0082 144.9799 0.00031095 -85.1475 0.24736
1.3514 0.98803 5.5172e-05 3.8182 0.012032 1.7781e-05 0.0011543 0.16435 0.00065853 0.165 0.15074 0 0.036097 0.0389 0 0.91635 0.25844 0.070131 0.0097396 4.3406 0.060792 7.3219e-05 0.82928 0.0053617 0.0061002 0.0015074 0.98536 0.99066 3.2661e-06 1.3065e-05 0.13259 0.78467 0.82485 0.0014597 0.87587 0.51194 0.0019641 0.42348 1.4549 1.452 16.0082 144.98 0.00031026 -85.1512 0.24836
1.3524 0.98803 5.5172e-05 3.8182 0.012032 1.7794e-05 0.0011543 0.1644 0.00065853 0.16506 0.1508 0 0.036093 0.0389 0 0.91644 0.25848 0.070144 0.0097412 4.341 0.060802 7.3232e-05 0.82927 0.0053622 0.0061006 0.0015053 0.98537 0.99066 3.264e-06 1.3056e-05 0.13259 0.78529 0.82528 0.0014592 0.87662 0.51211 0.0019634 0.42349 1.4564 1.4535 16.0083 144.98 0.00030958 -85.1548 0.24936
1.3534 0.98803 5.5172e-05 3.8182 0.012032 1.7808e-05 0.0011543 0.16446 0.00065853 0.16511 0.15085 0 0.03609 0.0389 0 0.91652 0.25852 0.070157 0.0097428 4.3414 0.060812 7.3245e-05 0.82926 0.0053626 0.0061011 0.0015045 0.98539 0.99067 3.2619e-06 1.3048e-05 0.1326 0.7859 0.8257 0.0014587 0.87737 0.51228 0.0019628 0.4235 1.4579 1.455 16.0083 144.98 0.00030891 -85.1585 0.25036
1.3544 0.98803 5.5172e-05 3.8182 0.012032 1.7821e-05 0.0011543 0.16452 0.00065853 0.16517 0.1509 0 0.036086 0.0389 0 0.9166 0.25856 0.070171 0.0097444 4.3419 0.060822 7.3258e-05 0.82925 0.005363 0.0061015 0.0015039 0.9854 0.99068 3.2598e-06 1.304e-05 0.1326 0.78652 0.82611 0.0014583 0.87811 0.51245 0.0019622 0.42351 1.4594 1.4565 16.0083 144.98 0.00030823 -85.1621 0.25136
1.3554 0.98803 5.5172e-05 3.8182 0.012032 1.7834e-05 0.0011543 0.16457 0.00065854 0.16523 0.15096 0 0.036083 0.0389 0 0.91668 0.25859 0.070184 0.0097461 4.3423 0.060832 7.3271e-05 0.82924 0.0053635 0.006102 0.0015034 0.98541 0.99069 3.2578e-06 1.3031e-05 0.1326 0.78713 0.82653 0.0014578 0.87884 0.51261 0.0019616 0.42352 1.4608 1.458 16.0083 144.98 0.00030756 -85.1657 0.25236
1.3564 0.98803 5.5172e-05 3.8182 0.012032 1.7847e-05 0.0011543 0.16463 0.00065854 0.16529 0.15101 0 0.036079 0.0389 0 0.91677 0.25863 0.070197 0.0097477 4.3428 0.060842 7.3283e-05 0.82923 0.0053639 0.0061024 0.0015023 0.98542 0.9907 3.2557e-06 1.3023e-05 0.13261 0.78774 0.82695 0.0014574 0.87957 0.51278 0.001961 0.42353 1.4623 1.4595 16.0084 144.98 0.00030689 -85.1692 0.25336
1.3574 0.98803 5.5172e-05 3.8182 0.012032 1.786e-05 0.0011543 0.16469 0.00065854 0.16534 0.15106 0 0.036076 0.0389 0 0.91685 0.25867 0.07021 0.0097493 4.3432 0.060852 7.3296e-05 0.82922 0.0053644 0.0061029 0.0015021 0.98543 0.99071 3.2537e-06 1.3015e-05 0.13261 0.78835 0.82736 0.0014569 0.8803 0.51295 0.0019605 0.42354 1.4638 1.461 16.0084 144.9801 0.00030623 -85.1727 0.25436
1.3584 0.98803 5.5172e-05 3.8182 0.012032 1.7873e-05 0.0011543 0.16475 0.00065854 0.1654 0.15112 0 0.036072 0.0389 0 0.91693 0.2587 0.070224 0.0097509 4.3436 0.060862 7.3309e-05 0.82921 0.0053648 0.0061033 0.0014999 0.98544 0.99071 3.2517e-06 1.3007e-05 0.13261 0.78896 0.82777 0.0014565 0.88102 0.51311 0.0019599 0.42355 1.4653 1.4625 16.0084 144.9801 0.00030556 -85.1762 0.25536
1.3594 0.98803 5.5172e-05 3.8182 0.012032 1.7886e-05 0.0011543 0.1648 0.00065854 0.16546 0.15117 0 0.036069 0.0389 0 0.91701 0.25874 0.070237 0.0097525 4.3441 0.060872 7.3322e-05 0.8292 0.0053652 0.0061038 0.0014992 0.98546 0.99072 3.2497e-06 1.2999e-05 0.13262 0.78956 0.82818 0.001456 0.88174 0.51328 0.0019593 0.42356 1.4667 1.4639 16.0084 144.9801 0.00030491 -85.1797 0.25636
1.3604 0.98803 5.5172e-05 3.8182 0.012032 1.7899e-05 0.0011543 0.16486 0.00065854 0.16551 0.15122 0 0.036065 0.0389 0 0.9171 0.25878 0.07025 0.0097541 4.3445 0.060882 7.3335e-05 0.82919 0.0053657 0.0061042 0.0014986 0.98547 0.99073 3.2477e-06 1.2991e-05 0.13262 0.79017 0.82859 0.0014556 0.88246 0.51345 0.0019587 0.42357 1.4682 1.4654 16.0084 144.9801 0.00030425 -85.1832 0.25736
1.3614 0.98803 5.5171e-05 3.8182 0.012032 1.7913e-05 0.0011543 0.16492 0.00065854 0.16557 0.15128 0 0.036062 0.0389 0 0.91718 0.25881 0.070263 0.0097557 4.345 0.060892 7.3348e-05 0.82918 0.0053661 0.0061047 0.0014981 0.98548 0.99074 3.2457e-06 1.2983e-05 0.13263 0.79077 0.82899 0.0014551 0.88317 0.51361 0.0019581 0.42358 1.4697 1.4669 16.0085 144.9801 0.0003036 -85.1866 0.25836
1.3624 0.98803 5.5171e-05 3.8182 0.012032 1.7926e-05 0.0011543 0.16497 0.00065854 0.16563 0.15133 0 0.036058 0.0389 0 0.91726 0.25885 0.070277 0.0097573 4.3454 0.060902 7.3361e-05 0.82917 0.0053666 0.0061051 0.0014972 0.98549 0.99075 3.2438e-06 1.2975e-05 0.13263 0.79137 0.8294 0.0014547 0.88388 0.51378 0.0019576 0.42359 1.4711 1.4683 16.0085 144.9801 0.00030295 -85.19 0.25936
1.3634 0.98803 5.5171e-05 3.8182 0.012032 1.7939e-05 0.0011543 0.16503 0.00065854 0.16568 0.15138 0 0.036055 0.0389 0 0.91735 0.25889 0.07029 0.0097589 4.3459 0.060912 7.3374e-05 0.82916 0.005367 0.0061056 0.0014964 0.9855 0.99075 3.2418e-06 1.2968e-05 0.13263 0.79197 0.8298 0.0014543 0.88458 0.51395 0.001957 0.4236 1.4726 1.4698 16.0085 144.9802 0.0003023 -85.1934 0.26036
1.3644 0.98803 5.5171e-05 3.8182 0.012032 1.7952e-05 0.0011543 0.16509 0.00065854 0.16574 0.15144 0 0.036051 0.0389 0 0.91743 0.25892 0.070303 0.0097605 4.3463 0.060922 7.3386e-05 0.82915 0.0053675 0.006106 0.0014956 0.98551 0.99076 3.2399e-06 1.296e-05 0.13264 0.79256 0.8302 0.0014538 0.88528 0.51411 0.0019565 0.42361 1.474 1.4713 16.0085 144.9802 0.00030166 -85.1967 0.26136
1.3654 0.98803 5.5171e-05 3.8182 0.012032 1.7965e-05 0.0011543 0.16514 0.00065854 0.1658 0.15149 0 0.036048 0.0389 0 0.91751 0.25896 0.070317 0.0097621 4.3468 0.060932 7.3399e-05 0.82914 0.0053679 0.0061065 0.0014948 0.98552 0.99077 3.238e-06 1.2952e-05 0.13264 0.79316 0.8306 0.0014534 0.88597 0.51428 0.0019559 0.42362 1.4755 1.4727 16.0086 144.9802 0.00030102 -85.2 0.26236
1.3664 0.98803 5.5171e-05 3.8182 0.012032 1.7978e-05 0.0011543 0.1652 0.00065855 0.16585 0.15154 0 0.036044 0.0389 0 0.91759 0.259 0.07033 0.0097638 4.3472 0.060942 7.3412e-05 0.82913 0.0053683 0.0061069 0.0014938 0.98553 0.99078 3.2361e-06 1.2945e-05 0.13264 0.79375 0.83099 0.001453 0.88666 0.51445 0.0019554 0.42363 1.4769 1.4742 16.0086 144.9802 0.00030038 -85.2033 0.26336
1.3674 0.98803 5.5171e-05 3.8182 0.012032 1.7991e-05 0.0011543 0.16525 0.00065855 0.16591 0.1516 0 0.036041 0.0389 0 0.91768 0.25903 0.070343 0.0097654 4.3477 0.060952 7.3425e-05 0.82912 0.0053688 0.0061074 0.0014934 0.98555 0.99078 3.2343e-06 1.2937e-05 0.13265 0.79434 0.83139 0.0014526 0.88735 0.51461 0.0019548 0.42364 1.4784 1.4756 16.0086 144.9802 0.00029974 -85.2066 0.26436
1.3684 0.98803 5.5171e-05 3.8182 0.012032 1.8004e-05 0.0011543 0.16531 0.00065855 0.16596 0.15165 0 0.036037 0.0389 0 0.91776 0.25907 0.070357 0.009767 4.3481 0.060962 7.3438e-05 0.82911 0.0053692 0.0061078 0.0014926 0.98556 0.99079 3.2324e-06 1.293e-05 0.13265 0.79493 0.83178 0.0014522 0.88803 0.51478 0.0019543 0.42365 1.4798 1.4771 16.0086 144.9802 0.00029911 -85.2099 0.26536
1.3694 0.98803 5.5171e-05 3.8182 0.012032 1.8018e-05 0.0011543 0.16537 0.00065855 0.16602 0.1517 0 0.036034 0.0389 0 0.91784 0.25911 0.07037 0.0097686 4.3486 0.060972 7.3451e-05 0.8291 0.0053697 0.0061083 0.0014917 0.98557 0.9908 3.2306e-06 1.2922e-05 0.13265 0.79552 0.83217 0.0014518 0.88871 0.51495 0.0019537 0.42366 1.4812 1.4785 16.0086 144.9803 0.00029848 -85.2131 0.26636
1.3704 0.98803 5.5171e-05 3.8182 0.012032 1.8031e-05 0.0011543 0.16542 0.00065855 0.16608 0.15175 0 0.036031 0.0389 0 0.91793 0.25915 0.070383 0.0097702 4.349 0.060982 7.3464e-05 0.82909 0.0053701 0.0061087 0.0014907 0.98558 0.9908 3.2287e-06 1.2915e-05 0.13266 0.7961 0.83256 0.0014514 0.88938 0.51511 0.0019532 0.42367 1.4827 1.4799 16.0087 144.9803 0.00029786 -85.2163 0.26736
1.3714 0.98803 5.5171e-05 3.8182 0.012032 1.8044e-05 0.0011543 0.16548 0.00065855 0.16613 0.15181 0 0.036027 0.0389 0 0.91801 0.25918 0.070397 0.0097718 4.3495 0.060992 7.3477e-05 0.82908 0.0053706 0.0061092 0.00149 0.98559 0.99081 3.2269e-06 1.2908e-05 0.13266 0.79668 0.83294 0.001451 0.89005 0.51528 0.0019527 0.42368 1.4841 1.4814 16.0087 144.9803 0.00029723 -85.2195 0.26836
1.3724 0.98803 5.5171e-05 3.8182 0.012032 1.8057e-05 0.0011543 0.16554 0.00065855 0.16619 0.15186 0 0.036024 0.0389 0 0.91809 0.25922 0.07041 0.0097734 4.3499 0.061002 7.349e-05 0.82907 0.005371 0.0061096 0.001489 0.9856 0.99082 3.225e-06 1.29e-05 0.13267 0.79727 0.83333 0.0014506 0.89072 0.51545 0.0019521 0.42369 1.4855 1.4828 16.0087 144.9803 0.00029661 -85.2227 0.26936
1.3734 0.98803 5.5171e-05 3.8182 0.012032 1.807e-05 0.0011543 0.16559 0.00065855 0.16625 0.15191 0 0.03602 0.0389 0 0.91817 0.25926 0.070423 0.0097751 4.3504 0.061012 7.3503e-05 0.82906 0.0053715 0.0061101 0.0014886 0.98561 0.99083 3.2234e-06 1.2893e-05 0.13267 0.79785 0.83371 0.0014502 0.89138 0.51561 0.0019516 0.4237 1.4869 1.4842 16.0087 144.9803 0.000296 -85.2258 0.27036
1.3744 0.98803 5.5171e-05 3.8182 0.012032 1.8083e-05 0.0011543 0.16565 0.00065855 0.1663 0.15196 0 0.036017 0.0389 0 0.91826 0.25929 0.070437 0.0097767 4.3508 0.061022 7.3515e-05 0.82905 0.0053719 0.0061106 0.0014871 0.98562 0.99083 3.2214e-06 1.2886e-05 0.13267 0.79842 0.8341 0.0014498 0.89204 0.51578 0.0019511 0.42371 1.4883 1.4857 16.0087 144.9803 0.00029538 -85.2289 0.27136
1.3754 0.98803 5.5171e-05 3.8182 0.012032 1.8096e-05 0.0011543 0.1657 0.00065855 0.16636 0.15202 0 0.036013 0.0389 0 0.91834 0.25933 0.07045 0.0097783 4.3513 0.061032 7.3528e-05 0.82904 0.0053724 0.006111 0.0014864 0.98563 0.99084 3.2197e-06 1.2879e-05 0.13268 0.799 0.83448 0.0014494 0.89269 0.51594 0.0019506 0.42372 1.4897 1.4871 16.0088 144.9804 0.00029477 -85.232 0.27236
1.3764 0.98803 5.5171e-05 3.8182 0.012032 1.8109e-05 0.0011543 0.16576 0.00065855 0.16641 0.15207 0 0.03601 0.0389 0 0.91842 0.25937 0.070463 0.0097799 4.3517 0.061042 7.3541e-05 0.82903 0.0053728 0.0061115 0.0014859 0.98564 0.99085 3.2179e-06 1.2872e-05 0.13268 0.79957 0.83485 0.001449 0.89334 0.51611 0.0019501 0.42373 1.4911 1.4885 16.0088 144.9804 0.00029416 -85.2351 0.27336
1.3774 0.98803 5.517e-05 3.8182 0.012032 1.8123e-05 0.0011543 0.16582 0.00065856 0.16647 0.15212 0 0.036007 0.0389 0 0.91851 0.2594 0.070477 0.0097815 4.3522 0.061052 7.3554e-05 0.82902 0.0053732 0.0061119 0.0014853 0.98565 0.99085 3.2163e-06 1.2865e-05 0.13268 0.80015 0.83523 0.0014486 0.89399 0.51628 0.0019496 0.42374 1.4925 1.4899 16.0088 144.9804 0.00029355 -85.2381 0.27436
1.3784 0.98803 5.517e-05 3.8182 0.012032 1.8136e-05 0.0011543 0.16587 0.00065856 0.16653 0.15217 0 0.036003 0.0389 0 0.91859 0.25944 0.07049 0.0097831 4.3526 0.061062 7.3567e-05 0.82901 0.0053737 0.0061124 0.0014846 0.98566 0.99086 3.2145e-06 1.2858e-05 0.13269 0.80072 0.8356 0.0014482 0.89463 0.51644 0.0019491 0.42375 1.4939 1.4913 16.0088 144.9804 0.00029295 -85.2411 0.27536
1.3794 0.98803 5.517e-05 3.8182 0.012032 1.8149e-05 0.0011543 0.16593 0.00065856 0.16658 0.15223 0 0.036 0.0389 0 0.91867 0.25948 0.070503 0.0097847 4.3531 0.061072 7.358e-05 0.829 0.0053741 0.0061128 0.0014839 0.98567 0.99087 3.213e-06 1.2852e-05 0.13269 0.80129 0.83598 0.0014478 0.89527 0.51661 0.0019486 0.42376 1.4953 1.4927 16.0088 144.9804 0.00029235 -85.2441 0.27636
1.3804 0.98803 5.517e-05 3.8182 0.012032 1.8162e-05 0.0011543 0.16598 0.00065856 0.16664 0.15228 0 0.035996 0.0389 0 0.91876 0.25952 0.070517 0.0097864 4.3535 0.061082 7.3593e-05 0.82899 0.0053746 0.0061133 0.0014831 0.98568 0.99087 3.211e-06 1.2845e-05 0.1327 0.80185 0.83635 0.0014475 0.89591 0.51678 0.0019481 0.42377 1.4967 1.4941 16.0088 144.9805 0.00029175 -85.2471 0.27736
1.3814 0.98803 5.517e-05 3.8182 0.012032 1.8175e-05 0.0011543 0.16604 0.00065856 0.16669 0.15233 0 0.035993 0.0389 0 0.91884 0.25955 0.07053 0.009788 4.354 0.061092 7.3606e-05 0.82898 0.005375 0.0061137 0.0014825 0.98569 0.99088 3.2098e-06 1.2838e-05 0.1327 0.80242 0.83672 0.0014471 0.89654 0.51694 0.0019476 0.42378 1.4981 1.4955 16.0089 144.9805 0.00029116 -85.2501 0.27836
1.3824 0.98803 5.517e-05 3.8182 0.012032 1.8188e-05 0.0011543 0.16609 0.00065856 0.16675 0.15238 0 0.035989 0.0389 0 0.91892 0.25959 0.070544 0.0097896 4.3544 0.061102 7.3619e-05 0.82897 0.0053755 0.0061142 0.0014815 0.9857 0.99089 3.2073e-06 1.2831e-05 0.1327 0.80298 0.83709 0.0014467 0.89717 0.51711 0.0019471 0.42379 1.4995 1.4969 16.0089 144.9805 0.00029057 -85.253 0.27936
1.3834 0.98803 5.517e-05 3.8182 0.012032 1.8201e-05 0.0011543 0.16615 0.00065856 0.1668 0.15244 0 0.035986 0.0389 0 0.91901 0.25963 0.070557 0.0097912 4.3549 0.061112 7.3632e-05 0.82896 0.0053759 0.0061147 0.0014812 0.98571 0.99089 3.207e-06 1.2825e-05 0.13271 0.80354 0.83745 0.0014463 0.89779 0.51727 0.0019466 0.4238 1.5009 1.4983 16.0089 144.9805 0.00028998 -85.2559 0.28036
1.3844 0.98803 5.517e-05 3.8182 0.012032 1.8214e-05 0.0011543 0.16621 0.00065856 0.16686 0.15249 0 0.035983 0.0389 0 0.91909 0.25966 0.07057 0.0097928 4.3553 0.061122 7.3645e-05 0.82895 0.0053764 0.0061151 0.0014797 0.98572 0.9909 3.203e-06 1.2818e-05 0.13271 0.80411 0.83782 0.001446 0.89841 0.51744 0.0019462 0.42381 1.5022 1.4997 16.0089 144.9805 0.00028939 -85.2588 0.28136
1.3854 0.98803 5.517e-05 3.8182 0.012031 1.8228e-05 0.0011543 0.16626 0.00065856 0.16692 0.15254 0 0.035979 0.0389 0 0.91917 0.2597 0.070584 0.0097945 4.3558 0.061132 7.3658e-05 0.82894 0.0053768 0.0061156 0.0014791 0.98573 0.9909 3.2019e-06 1.2812e-05 0.13271 0.80466 0.83818 0.0014456 0.89903 0.5176 0.0019457 0.42382 1.5036 1.501 16.0089 144.9805 0.0002888 -85.2617 0.28236
1.3864 0.98803 5.517e-05 3.8182 0.012031 1.8241e-05 0.0011543 0.16632 0.00065856 0.16697 0.15259 0 0.035976 0.0389 0 0.91926 0.25974 0.070597 0.0097961 4.3563 0.061142 7.3671e-05 0.82893 0.0053773 0.006116 0.0014786 0.98574 0.99091 3.2004e-06 1.2805e-05 0.13272 0.80522 0.83854 0.0014452 0.89964 0.51777 0.0019452 0.42383 1.505 1.5024 16.0089 144.9806 0.00028822 -85.2645 0.28336
1.3874 0.98803 5.517e-05 3.8182 0.012031 1.8254e-05 0.0011543 0.16637 0.00065856 0.16703 0.15265 0 0.035972 0.0389 0 0.91934 0.25978 0.07061 0.0097977 4.3567 0.061152 7.3684e-05 0.82892 0.0053777 0.0061165 0.001478 0.98574 0.99092 3.2e-06 1.2799e-05 0.13272 0.80578 0.8389 0.0014449 0.90025 0.51794 0.0019447 0.42384 1.5063 1.5038 16.009 144.9806 0.00028764 -85.2674 0.28436
1.3884 0.98803 5.517e-05 3.8182 0.012031 1.8267e-05 0.0011543 0.16643 0.00065856 0.16708 0.1527 0 0.035969 0.0389 0 0.91942 0.25981 0.070624 0.0097993 4.3572 0.061162 7.3697e-05 0.82891 0.0053782 0.006117 0.0014774 0.98575 0.99092 3.1972e-06 1.2792e-05 0.13273 0.80633 0.83926 0.0014445 0.90086 0.5181 0.0019443 0.42385 1.5077 1.5052 16.009 144.9806 0.00028707 -85.2702 0.28536
1.3894 0.98803 5.517e-05 3.8182 0.012031 1.828e-05 0.0011543 0.16648 0.00065857 0.16714 0.15275 0 0.035966 0.0389 0 0.91951 0.25985 0.070637 0.0098009 4.3576 0.061172 7.371e-05 0.8289 0.0053786 0.0061174 0.0014767 0.98576 0.99093 3.1979e-06 1.2786e-05 0.13273 0.80688 0.83962 0.0014442 0.90146 0.51827 0.0019438 0.42386 1.5091 1.5065 16.009 144.9806 0.00028649 -85.273 0.28636
1.3904 0.98803 5.517e-05 3.8182 0.012031 1.8293e-05 0.0011543 0.16654 0.00065857 0.16719 0.1528 0 0.035962 0.0389 0 0.91959 0.25989 0.070651 0.0098026 4.3581 0.061182 7.3723e-05 0.82889 0.0053791 0.0061179 0.0014762 0.98577 0.99094 3.1926e-06 1.278e-05 0.13273 0.80743 0.83997 0.0014438 0.90206 0.51843 0.0019434 0.42387 1.5104 1.5079 16.009 144.9806 0.00028592 -85.2757 0.28736
1.3914 0.98803 5.517e-05 3.8182 0.012031 1.8306e-05 0.0011543 0.16659 0.00065857 0.16725 0.15285 0 0.035959 0.0389 0 0.91967 0.25992 0.070664 0.0098042 4.3585 0.061192 7.3736e-05 0.82888 0.0053796 0.0061183 0.0014751 0.98578 0.99094 3.1973e-06 1.2774e-05 0.13274 0.80798 0.84033 0.0014435 0.90265 0.5186 0.0019429 0.42389 1.5118 1.5093 16.009 144.9806 0.00028535 -85.2785 0.28836
1.3924 0.98803 5.517e-05 3.8182 0.012031 1.8319e-05 0.0011543 0.16665 0.00065857 0.1673 0.15291 0 0.035956 0.0389 0 0.91976 0.25996 0.070678 0.0098058 4.359 0.061202 7.3749e-05 0.82887 0.00538 0.0061188 0.0014752 0.98579 0.99095 3.1853e-06 1.2767e-05 0.13274 0.80853 0.84068 0.0014431 0.90325 0.51876 0.0019425 0.4239 1.5131 1.5106 16.009 144.9807 0.00028479 -85.2812 0.28936
1.3934 0.98803 5.5169e-05 3.8182 0.012031 1.8333e-05 0.0011543 0.1667 0.00065857 0.16736 0.15296 0 0.035952 0.0389 0 0.91984 0.26 0.070691 0.0098074 4.3595 0.061212 7.3762e-05 0.82886 0.0053805 0.0061193 0.0014744 0.9858 0.99095 3.1859e-06 1.2761e-05 0.13274 0.80907 0.84103 0.0014428 0.90383 0.51893 0.001942 0.42391 1.5145 1.512 16.0091 144.9807 0.00028422 -85.2839 0.29036
1.3944 0.98803 5.5169e-05 3.8182 0.012031 1.8346e-05 0.0011543 0.16676 0.00065857 0.16741 0.15301 0 0.035949 0.0389 0 0.91992 0.26004 0.070704 0.009809 4.3599 0.061222 7.3775e-05 0.82885 0.0053809 0.0061197 0.0014736 0.98581 0.99096 3.185e-06 1.2755e-05 0.13275 0.80961 0.84138 0.0014425 0.90442 0.5191 0.0019416 0.42392 1.5158 1.5133 16.0091 144.9807 0.00028366 -85.2866 0.29136
1.3954 0.98803 5.5169e-05 3.8182 0.012031 1.8359e-05 0.0011543 0.16682 0.00065857 0.16747 0.15306 0 0.035945 0.0389 0 0.92001 0.26007 0.070718 0.0098107 4.3604 0.061232 7.3788e-05 0.82884 0.0053814 0.0061202 0.0014728 0.98582 0.99096 3.1886e-06 1.2749e-05 0.13275 0.81015 0.84173 0.0014421 0.905 0.51926 0.0019411 0.42393 1.5171 1.5147 16.0091 144.9807 0.00028311 -85.2893 0.29236
1.3964 0.98803 5.5169e-05 3.8182 0.012031 1.8372e-05 0.0011543 0.16687 0.00065857 0.16752 0.15311 0 0.035942 0.0389 0 0.92009 0.26011 0.070731 0.0098123 4.3608 0.061242 7.3801e-05 0.82883 0.0053818 0.0061206 0.001472 0.98582 0.99097 3.1822e-06 1.2743e-05 0.13276 0.81069 0.84207 0.0014418 0.90558 0.51943 0.0019407 0.42394 1.5185 1.516 16.0091 144.9807 0.00028255 -85.2919 0.29336
1.3974 0.98803 5.5169e-05 3.8182 0.012031 1.8385e-05 0.0011543 0.16693 0.00065857 0.16758 0.15316 0 0.035939 0.0389 0 0.92017 0.26015 0.070745 0.0098139 4.3613 0.061252 7.3814e-05 0.82882 0.0053823 0.0061211 0.0014715 0.98583 0.99098 3.1904e-06 1.2737e-05 0.13276 0.81123 0.84242 0.0014415 0.90615 0.51959 0.0019403 0.42395 1.5198 1.5173 16.0091 144.9807 0.000282 -85.2946 0.29436
1.3984 0.98803 5.5169e-05 3.8182 0.012031 1.8398e-05 0.0011543 0.16698 0.00065857 0.16763 0.15322 0 0.035935 0.0389 0 0.92026 0.26018 0.070758 0.0098155 4.3618 0.061262 7.3827e-05 0.82881 0.0053827 0.0061216 0.0014706 0.98584 0.99098 3.1729e-06 1.2731e-05 0.13276 0.81177 0.84276 0.0014411 0.90672 0.51976 0.0019398 0.42396 1.5211 1.5187 16.0091 144.9808 0.00028145 -85.2972 0.29536
1.3994 0.98803 5.5169e-05 3.8182 0.012031 1.8411e-05 0.0011543 0.16704 0.00065857 0.16769 0.15327 0 0.035932 0.0389 0 0.92034 0.26022 0.070772 0.0098172 4.3622 0.061272 7.384e-05 0.8288 0.0053832 0.006122 0.0014706 0.98585 0.99099 3.1983e-06 1.2726e-05 0.13277 0.8123 0.8431 0.0014408 0.90729 0.51992 0.0019394 0.42397 1.5224 1.52 16.0091 144.9808 0.0002809 -85.2998 0.29636
1.4004 0.98803 5.5169e-05 3.8182 0.012031 1.8424e-05 0.0011543 0.16709 0.00065858 0.16774 0.15332 0 0.035929 0.0389 0 0.92042 0.26026 0.070785 0.0098188 4.3627 0.061282 7.3853e-05 0.82879 0.0053836 0.0061225 0.0014687 0.98586 0.99099 3.1515e-06 1.272e-05 0.13277 0.81284 0.84344 0.0014405 0.90785 0.52009 0.001939 0.42398 1.5237 1.5213 16.0092 144.9808 0.00028035 -85.3023 0.29736
1.4014 0.98803 5.5169e-05 3.8182 0.012031 1.8438e-05 0.0011543 0.16714 0.00065858 0.1678 0.15337 0 0.035925 0.0389 0 0.92051 0.2603 0.070798 0.0098204 4.3632 0.061292 7.3866e-05 0.82878 0.0053841 0.006123 0.0014681 0.98587 0.991 3.1591e-06 1.2714e-05 0.13277 0.81337 0.84378 0.0014402 0.90841 0.52025 0.0019385 0.42399 1.5251 1.5226 16.0092 144.9808 0.00027981 -85.3049 0.29836
1.4024 0.98803 5.5169e-05 3.8182 0.012031 1.8451e-05 0.0011543 0.1672 0.00065858 0.16785 0.15342 0 0.035922 0.0389 0 0.92059 0.26033 0.070812 0.009822 4.3636 0.061302 7.3879e-05 0.82877 0.0053846 0.0061234 0.0014683 0.98587 0.991 3.1764e-06 1.2708e-05 0.13278 0.8139 0.84411 0.0014398 0.90897 0.52042 0.0019381 0.424 1.5264 1.524 16.0092 144.9808 0.00027927 -85.3074 0.29936
1.4034 0.98803 5.5169e-05 3.8182 0.012031 1.8464e-05 0.0011543 0.16725 0.00065858 0.16791 0.15347 0 0.035919 0.0389 0 0.92067 0.26037 0.070825 0.0098237 4.3641 0.061313 7.3892e-05 0.82876 0.005385 0.0061239 0.0014677 0.98588 0.99101 3.1756e-06 1.2703e-05 0.13278 0.81443 0.84445 0.0014395 0.90952 0.52058 0.0019377 0.42402 1.5277 1.5253 16.0092 144.9809 0.00027873 -85.3099 0.30036
1.4044 0.98803 5.5169e-05 3.8182 0.012031 1.8477e-05 0.0011543 0.16731 0.00065858 0.16796 0.15352 0 0.035915 0.0389 0 0.92076 0.26041 0.070839 0.0098253 4.3646 0.061323 7.3905e-05 0.82875 0.0053855 0.0061244 0.001467 0.98589 0.99101 3.1742e-06 1.2697e-05 0.13279 0.81495 0.84478 0.0014392 0.91007 0.52075 0.0019373 0.42403 1.529 1.5266 16.0092 144.9809 0.0002782 -85.3124 0.30136
1.4054 0.98803 5.5169e-05 3.8182 0.012031 1.849e-05 0.0011543 0.16736 0.00065858 0.16802 0.15358 0 0.035912 0.0389 0 0.92084 0.26045 0.070852 0.0098269 4.365 0.061333 7.3918e-05 0.82874 0.0053859 0.0061248 0.0014664 0.9859 0.99102 3.1728e-06 1.2691e-05 0.13279 0.81548 0.84511 0.0014389 0.91062 0.52091 0.0019369 0.42404 1.5303 1.5279 16.0092 144.9809 0.00027766 -85.3149 0.30236
1.4064 0.98803 5.5169e-05 3.8182 0.012031 1.8503e-05 0.0011543 0.16742 0.00065858 0.16807 0.15363 0 0.035909 0.0389 0 0.92093 0.26048 0.070866 0.0098285 4.3655 0.061343 7.3931e-05 0.82873 0.0053864 0.0061253 0.0014658 0.98591 0.99103 3.1715e-06 1.2686e-05 0.13279 0.816 0.84544 0.0014386 0.91116 0.52108 0.0019365 0.42405 1.5316 1.5292 16.0092 144.9809 0.00027713 -85.3174 0.30336
1.4074 0.98803 5.5169e-05 3.8182 0.012031 1.8516e-05 0.0011543 0.16747 0.00065858 0.16813 0.15368 0 0.035905 0.0389 0 0.92101 0.26052 0.070879 0.0098302 4.3659 0.061353 7.3944e-05 0.82872 0.0053868 0.0061257 0.0014652 0.98591 0.99103 3.1701e-06 1.268e-05 0.1328 0.81652 0.84577 0.0014383 0.9117 0.52124 0.0019361 0.42406 1.5329 1.5305 16.0092 144.9809 0.0002766 -85.3198 0.30436
1.4084 0.98803 5.5168e-05 3.8182 0.012031 1.8529e-05 0.0011543 0.16753 0.00065858 0.16818 0.15373 0 0.035902 0.0389 0 0.92109 0.26056 0.070893 0.0098318 4.3664 0.061363 7.3957e-05 0.82871 0.0053873 0.0061262 0.0014646 0.98592 0.99104 3.1687e-06 1.2675e-05 0.1328 0.81704 0.8461 0.001438 0.91224 0.52141 0.0019357 0.42407 1.5342 1.5318 16.0093 144.9809 0.00027608 -85.3223 0.30536
1.4094 0.98803 5.5168e-05 3.8182 0.012031 1.8543e-05 0.0011543 0.16758 0.00065858 0.16824 0.15378 0 0.035899 0.0389 0 0.92118 0.2606 0.070906 0.0098334 4.3669 0.061373 7.397e-05 0.8287 0.0053878 0.0061267 0.0014641 0.98593 0.99104 3.1674e-06 1.267e-05 0.1328 0.81756 0.84643 0.0014377 0.91277 0.52157 0.0019353 0.42408 1.5354 1.5331 16.0093 144.981 0.00027555 -85.3247 0.30636
1.4104 0.98803 5.5168e-05 3.8182 0.012031 1.8556e-05 0.0011543 0.16764 0.00065858 0.16829 0.15383 0 0.035895 0.0389 0 0.92126 0.26063 0.07092 0.0098351 4.3673 0.061383 7.3983e-05 0.82869 0.0053882 0.0061271 0.0014635 0.98594 0.99105 3.166e-06 1.2664e-05 0.13281 0.81808 0.84675 0.0014374 0.9133 0.52174 0.0019349 0.42409 1.5367 1.5344 16.0093 144.981 0.00027503 -85.3271 0.30736
1.4114 0.98803 5.5168e-05 3.8182 0.012031 1.8569e-05 0.0011543 0.16769 0.00065858 0.16835 0.15388 0 0.035892 0.0389 0 0.92135 0.26067 0.070933 0.0098367 4.3678 0.061393 7.3996e-05 0.82868 0.0053887 0.0061276 0.0014629 0.98595 0.99105 3.1647e-06 1.2659e-05 0.13281 0.81859 0.84708 0.0014371 0.91383 0.5219 0.0019345 0.4241 1.538 1.5357 16.0093 144.981 0.00027451 -85.3295 0.30836
1.4124 0.98803 5.5168e-05 3.8182 0.012031 1.8582e-05 0.0011543 0.16775 0.00065859 0.1684 0.15393 0 0.035889 0.0389 0 0.92143 0.26071 0.070947 0.0098383 4.3683 0.061403 7.4009e-05 0.82867 0.0053891 0.0061281 0.0014623 0.98595 0.99106 3.1634e-06 1.2654e-05 0.13282 0.8191 0.8474 0.0014368 0.91435 0.52207 0.0019341 0.42411 1.5393 1.5369 16.0093 144.981 0.00027399 -85.3318 0.30936
1.4134 0.98803 5.5168e-05 3.8182 0.012031 1.8595e-05 0.0011543 0.1678 0.00065859 0.16845 0.15399 0 0.035885 0.0389 0 0.92151 0.26074 0.07096 0.0098399 4.3688 0.061413 7.4022e-05 0.82866 0.0053896 0.0061286 0.0014617 0.98596 0.99106 3.1621e-06 1.2648e-05 0.13282 0.81962 0.84772 0.0014365 0.91487 0.52223 0.0019337 0.42413 1.5405 1.5382 16.0093 144.981 0.00027348 -85.3342 0.31036
1.4144 0.98803 5.5168e-05 3.8182 0.012031 1.8608e-05 0.0011543 0.16785 0.00065859 0.16851 0.15404 0 0.035882 0.0389 0 0.9216 0.26078 0.070974 0.0098416 4.3692 0.061423 7.4035e-05 0.82865 0.0053901 0.006129 0.0014612 0.98597 0.99107 3.1608e-06 1.2643e-05 0.13282 0.82013 0.84804 0.0014362 0.91539 0.5224 0.0019333 0.42414 1.5418 1.5395 16.0093 144.981 0.00027297 -85.3365 0.31136
1.4154 0.98803 5.5168e-05 3.8182 0.012031 1.8621e-05 0.0011543 0.16791 0.00065859 0.16856 0.15409 0 0.035879 0.0389 0 0.92168 0.26082 0.070987 0.0098432 4.3697 0.061434 7.4048e-05 0.82864 0.0053905 0.0061295 0.0014606 0.98598 0.99107 3.1595e-06 1.2638e-05 0.13283 0.82064 0.84836 0.0014359 0.91591 0.52256 0.001933 0.42415 1.5431 1.5408 16.0093 144.9811 0.00027246 -85.3388 0.31236
1.4164 0.98803 5.5168e-05 3.8182 0.012031 1.8634e-05 0.0011543 0.16796 0.00065859 0.16862 0.15414 0 0.035876 0.0389 0 0.92176 0.26086 0.071001 0.0098448 4.3702 0.061444 7.4061e-05 0.82863 0.005391 0.00613 0.0014601 0.98598 0.99108 3.1582e-06 1.2633e-05 0.13283 0.82114 0.84867 0.0014356 0.91642 0.52272 0.0019326 0.42416 1.5443 1.542 16.0094 144.9811 0.00027195 -85.3411 0.31336
1.4174 0.98803 5.5168e-05 3.8182 0.012031 1.8648e-05 0.0011543 0.16802 0.00065859 0.16867 0.15419 0 0.035872 0.0389 0 0.92185 0.26089 0.071014 0.0098465 4.3706 0.061454 7.4075e-05 0.82862 0.0053914 0.0061304 0.0014595 0.98599 0.99108 3.1569e-06 1.2628e-05 0.13283 0.82165 0.84899 0.0014353 0.91693 0.52289 0.0019322 0.42417 1.5456 1.5433 16.0094 144.9811 0.00027144 -85.3434 0.31436
1.4184 0.98803 5.5168e-05 3.8182 0.012031 1.8661e-05 0.0011543 0.16807 0.00065859 0.16872 0.15424 0 0.035869 0.0389 0 0.92193 0.26093 0.071028 0.0098481 4.3711 0.061464 7.4088e-05 0.82861 0.0053919 0.0061309 0.0014589 0.986 0.99109 3.1557e-06 1.2623e-05 0.13284 0.82215 0.8493 0.001435 0.91743 0.52305 0.0019318 0.42418 1.5469 1.5446 16.0094 144.9811 0.00027094 -85.3456 0.31536
1.4194 0.98803 5.5168e-05 3.8182 0.012031 1.8674e-05 0.0011543 0.16812 0.00065859 0.16878 0.15429 0 0.035866 0.0389 0 0.92202 0.26097 0.071041 0.0098497 4.3716 0.061474 7.4101e-05 0.8286 0.0053924 0.0061314 0.0014584 0.986 0.99109 3.1544e-06 1.2618e-05 0.13284 0.82266 0.84961 0.0014347 0.91794 0.52322 0.0019315 0.42419 1.5481 1.5458 16.0094 144.9811 0.00027044 -85.3479 0.31636
1.4204 0.98803 5.5168e-05 3.8182 0.012031 1.8687e-05 0.0011543 0.16818 0.00065859 0.16883 0.15434 0 0.035862 0.0389 0 0.9221 0.26101 0.071055 0.0098514 4.372 0.061484 7.4114e-05 0.82859 0.0053928 0.0061318 0.0014579 0.98601 0.9911 3.1532e-06 1.2613e-05 0.13285 0.82316 0.84993 0.0014345 0.91844 0.52338 0.0019311 0.42421 1.5494 1.5471 16.0094 144.9812 0.00026994 -85.3501 0.31736
1.4214 0.98803 5.5168e-05 3.8182 0.012031 1.87e-05 0.0011543 0.16823 0.00065859 0.16889 0.15439 0 0.035859 0.0389 0 0.92219 0.26104 0.071068 0.009853 4.3725 0.061494 7.4127e-05 0.82858 0.0053933 0.0061323 0.0014573 0.98602 0.9911 3.1519e-06 1.2608e-05 0.13285 0.82366 0.85024 0.0014342 0.91893 0.52355 0.0019307 0.42422 1.5506 1.5483 16.0094 144.9812 0.00026944 -85.3523 0.31836
1.4224 0.98803 5.5168e-05 3.8182 0.012031 1.8713e-05 0.0011543 0.16829 0.00065859 0.16894 0.15444 0 0.035856 0.0389 0 0.92227 0.26108 0.071082 0.0098546 4.373 0.061504 7.414e-05 0.82857 0.0053937 0.0061328 0.0014568 0.98603 0.9911 3.1507e-06 1.2603e-05 0.13285 0.82416 0.85054 0.0014339 0.91943 0.52371 0.0019304 0.42423 1.5518 1.5496 16.0094 144.9812 0.00026895 -85.3545 0.31936
1.4234 0.98803 5.5168e-05 3.8182 0.012031 1.8726e-05 0.0011543 0.16834 0.00065859 0.16899 0.15449 0 0.035853 0.0389 0 0.92235 0.26112 0.071095 0.0098563 4.3735 0.061514 7.4153e-05 0.82856 0.0053942 0.0061333 0.0014563 0.98603 0.99111 3.1495e-06 1.2598e-05 0.13286 0.82465 0.85085 0.0014336 0.91992 0.52387 0.00193 0.42424 1.5531 1.5508 16.0094 144.9812 0.00026845 -85.3567 0.32036
1.4244 0.98803 5.5167e-05 3.8182 0.012031 1.8739e-05 0.0011543 0.16839 0.0006586 0.16905 0.15454 0 0.035849 0.0389 0 0.92244 0.26116 0.071109 0.0098579 4.3739 0.061525 7.4166e-05 0.82855 0.0053947 0.0061337 0.0014557 0.98604 0.99111 3.1483e-06 1.2593e-05 0.13286 0.82515 0.85116 0.0014334 0.9204 0.52404 0.0019297 0.42425 1.5543 1.5521 16.0094 144.9812 0.00026796 -85.3589 0.32136
1.4254 0.98803 5.5167e-05 3.8182 0.012031 1.8753e-05 0.0011543 0.16845 0.0006586 0.1691 0.15459 0 0.035846 0.0389 0 0.92252 0.26119 0.071122 0.0098595 4.3744 0.061535 7.4179e-05 0.82854 0.0053951 0.0061342 0.0014552 0.98605 0.99112 3.1471e-06 1.2588e-05 0.13287 0.82564 0.85146 0.0014331 0.92089 0.5242 0.0019293 0.42426 1.5555 1.5533 16.0094 144.9812 0.00026747 -85.361 0.32236
1.4264 0.98803 5.5167e-05 3.8182 0.012031 1.8766e-05 0.0011543 0.1685 0.0006586 0.16916 0.15464 0 0.035843 0.0389 0 0.92261 0.26123 0.071136 0.0098612 4.3749 0.061545 7.4192e-05 0.82853 0.0053956 0.0061347 0.0014547 0.98605 0.99112 3.1459e-06 1.2584e-05 0.13287 0.82613 0.85177 0.0014328 0.92137 0.52437 0.001929 0.42427 1.5568 1.5545 16.0094 144.9813 0.00026699 -85.3632 0.32336
1.4274 0.98803 5.5167e-05 3.8182 0.012031 1.8779e-05 0.0011543 0.16856 0.0006586 0.16921 0.1547 0 0.035839 0.0389 0 0.92269 0.26127 0.071149 0.0098628 4.3754 0.061555 7.4206e-05 0.82852 0.0053961 0.0061351 0.0014542 0.98606 0.99113 3.1447e-06 1.2579e-05 0.13287 0.82662 0.85207 0.0014326 0.92185 0.52453 0.0019286 0.42428 1.558 1.5558 16.0095 144.9813 0.0002665 -85.3653 0.32436
1.4284 0.98803 5.5167e-05 3.8182 0.012031 1.8792e-05 0.0011543 0.16861 0.0006586 0.16926 0.15475 0 0.035836 0.0389 0 0.92277 0.26131 0.071163 0.0098644 4.3758 0.061565 7.4219e-05 0.82851 0.0053965 0.0061356 0.0014537 0.98607 0.99113 3.1435e-06 1.2574e-05 0.13288 0.82711 0.85237 0.0014323 0.92232 0.52469 0.0019283 0.4243 1.5592 1.557 16.0095 144.9813 0.00026602 -85.3674 0.32536
1.4294 0.98803 5.5167e-05 3.8182 0.012031 1.8805e-05 0.0011543 0.16866 0.0006586 0.16932 0.1548 0 0.035833 0.0389 0 0.92286 0.26134 0.071176 0.0098661 4.3763 0.061575 7.4232e-05 0.8285 0.005397 0.0061361 0.0014532 0.98607 0.99114 3.1424e-06 1.257e-05 0.13288 0.8276 0.85267 0.001432 0.9228 0.52486 0.0019279 0.42431 1.5604 1.5582 16.0095 144.9813 0.00026554 -85.3695 0.32636
1.4304 0.98803 5.5167e-05 3.8182 0.012031 1.8818e-05 0.0011543 0.16872 0.0006586 0.16937 0.15485 0 0.03583 0.0389 0 0.92294 0.26138 0.07119 0.0098677 4.3768 0.061585 7.4245e-05 0.82849 0.0053975 0.0061366 0.0014527 0.98608 0.99114 3.1412e-06 1.2565e-05 0.13288 0.82808 0.85297 0.0014318 0.92327 0.52502 0.0019276 0.42432 1.5616 1.5595 16.0095 144.9813 0.00026507 -85.3716 0.32736
1.4314 0.98803 5.5167e-05 3.8182 0.012031 1.8831e-05 0.0011543 0.16877 0.0006586 0.16942 0.1549 0 0.035826 0.0389 0 0.92303 0.26142 0.071204 0.0098693 4.3773 0.061595 7.4258e-05 0.82848 0.0053979 0.006137 0.0014522 0.98609 0.99114 3.1401e-06 1.256e-05 0.13289 0.82857 0.85326 0.0014315 0.92373 0.52519 0.0019273 0.42433 1.5629 1.5607 16.0095 144.9814 0.00026459 -85.3736 0.32836
1.4324 0.98803 5.5167e-05 3.8182 0.012031 1.8844e-05 0.0011543 0.16882 0.0006586 0.16948 0.15495 0 0.035823 0.0389 0 0.92311 0.26146 0.071217 0.009871 4.3777 0.061606 7.4271e-05 0.82847 0.0053984 0.0061375 0.0014517 0.98609 0.99115 3.1389e-06 1.2556e-05 0.13289 0.82905 0.85356 0.0014313 0.9242 0.52535 0.0019269 0.42434 1.5641 1.5619 16.0095 144.9814 0.00026412 -85.3757 0.32936
1.4334 0.98803 5.5167e-05 3.8182 0.012031 1.8858e-05 0.0011543 0.16888 0.0006586 0.16953 0.155 0 0.03582 0.0389 0 0.9232 0.2615 0.071231 0.0098726 4.3782 0.061616 7.4284e-05 0.82846 0.0053989 0.006138 0.0014512 0.9861 0.99115 3.1378e-06 1.2551e-05 0.1329 0.82953 0.85385 0.001431 0.92466 0.52551 0.0019266 0.42435 1.5653 1.5631 16.0095 144.9814 0.00026364 -85.3777 0.33036
1.4344 0.98803 5.5167e-05 3.8182 0.012031 1.8871e-05 0.0011543 0.16893 0.0006586 0.16958 0.15505 0 0.035817 0.0389 0 0.92328 0.26153 0.071244 0.0098742 4.3787 0.061626 7.4297e-05 0.82845 0.0053993 0.0061385 0.0014507 0.98611 0.99116 3.1367e-06 1.2547e-05 0.1329 0.83001 0.85414 0.0014308 0.92512 0.52568 0.0019263 0.42437 1.5665 1.5643 16.0095 144.9814 0.00026318 -85.3797 0.33136
1.4354 0.98803 5.5167e-05 3.8182 0.012031 1.8884e-05 0.0011543 0.16898 0.0006586 0.16964 0.1551 0 0.035814 0.0389 0 0.92336 0.26157 0.071258 0.0098759 4.3792 0.061636 7.4311e-05 0.82844 0.0053998 0.0061389 0.0014502 0.98611 0.99116 3.1356e-06 1.2542e-05 0.1329 0.83049 0.85444 0.0014305 0.92557 0.52584 0.0019259 0.42438 1.5677 1.5655 16.0095 144.9814 0.00026271 -85.3817 0.33236
1.4364 0.98803 5.5167e-05 3.8182 0.012031 1.8897e-05 0.0011543 0.16904 0.0006586 0.16969 0.15515 0 0.03581 0.0389 0 0.92345 0.26161 0.071271 0.0098775 4.3797 0.061646 7.4324e-05 0.82843 0.0054003 0.0061394 0.0014497 0.98612 0.99117 3.1345e-06 1.2538e-05 0.13291 0.83097 0.85473 0.0014303 0.92603 0.52601 0.0019256 0.42439 1.5689 1.5667 16.0095 144.9814 0.00026224 -85.3837 0.33336
1.4374 0.98803 5.5167e-05 3.8182 0.012031 1.891e-05 0.0011543 0.16909 0.00065861 0.16974 0.1552 0 0.035807 0.0389 0 0.92353 0.26165 0.071285 0.0098792 4.3801 0.061656 7.4337e-05 0.82842 0.0054007 0.0061399 0.0014492 0.98613 0.99117 3.1334e-06 1.2534e-05 0.13291 0.83144 0.85502 0.00143 0.92648 0.52617 0.0019253 0.4244 1.5701 1.5679 16.0095 144.9815 0.00026178 -85.3857 0.33436
1.4384 0.98803 5.5167e-05 3.8182 0.012031 1.8923e-05 0.0011543 0.16914 0.00065861 0.1698 0.15525 0 0.035804 0.0389 0 0.92362 0.26168 0.071299 0.0098808 4.3806 0.061667 7.435e-05 0.82841 0.0054012 0.0061404 0.0014488 0.98613 0.99117 3.1323e-06 1.2529e-05 0.13292 0.83192 0.8553 0.0014298 0.92693 0.52633 0.001925 0.42441 1.5712 1.5691 16.0095 144.9815 0.00026132 -85.3876 0.33536
1.4394 0.98803 5.5167e-05 3.8182 0.012031 1.8936e-05 0.0011543 0.1692 0.00065861 0.16985 0.1553 0 0.035801 0.0389 0 0.9237 0.26172 0.071312 0.0098824 4.3811 0.061677 7.4363e-05 0.8284 0.0054017 0.0061408 0.0014483 0.98614 0.99118 3.1312e-06 1.2525e-05 0.13292 0.83239 0.85559 0.0014295 0.92737 0.5265 0.0019246 0.42442 1.5724 1.5703 16.0095 144.9815 0.00026086 -85.3896 0.33636
1.4404 0.98803 5.5166e-05 3.8182 0.012031 1.8949e-05 0.0011543 0.16925 0.00065861 0.1699 0.15535 0 0.035797 0.0389 0 0.92379 0.26176 0.071326 0.0098841 4.3816 0.061687 7.4376e-05 0.82839 0.0054021 0.0061413 0.0014478 0.98614 0.99118 3.1301e-06 1.2521e-05 0.13292 0.83286 0.85588 0.0014293 0.92781 0.52666 0.0019243 0.42444 1.5736 1.5715 16.0096 144.9815 0.0002604 -85.3915 0.33736
1.4414 0.98803 5.5166e-05 3.8182 0.012031 1.8963e-05 0.0011543 0.1693 0.00065861 0.16996 0.1554 0 0.035794 0.0389 0 0.92387 0.2618 0.071339 0.0098857 4.3821 0.061697 7.439e-05 0.82838 0.0054026 0.0061418 0.0014474 0.98615 0.99119 3.1291e-06 1.2516e-05 0.13293 0.83333 0.85616 0.001429 0.92825 0.52682 0.001924 0.42445 1.5748 1.5727 16.0096 144.9815 0.00025995 -85.3934 0.33836
1.4424 0.98803 5.5166e-05 3.8182 0.012031 1.8976e-05 0.0011543 0.16936 0.00065861 0.17001 0.15545 0 0.035791 0.0389 0 0.92396 0.26183 0.071353 0.0098873 4.3825 0.061707 7.4403e-05 0.82837 0.0054031 0.0061423 0.0014469 0.98616 0.99119 3.128e-06 1.2512e-05 0.13293 0.8338 0.85644 0.0014288 0.92869 0.52699 0.0019237 0.42446 1.576 1.5739 16.0096 144.9816 0.00025949 -85.3953 0.33936
1.4434 0.98803 5.5166e-05 3.8182 0.012031 1.8989e-05 0.0011543 0.16941 0.00065861 0.17006 0.1555 0 0.035788 0.0389 0 0.92404 0.26187 0.071367 0.009889 4.383 0.061717 7.4416e-05 0.82836 0.0054035 0.0061428 0.0014465 0.98616 0.99119 3.127e-06 1.2508e-05 0.13294 0.83426 0.85673 0.0014286 0.92912 0.52715 0.0019234 0.42447 1.5771 1.575 16.0096 144.9816 0.00025904 -85.3972 0.34036
1.4444 0.98803 5.5166e-05 3.8182 0.012031 1.9002e-05 0.0011543 0.16946 0.00065861 0.17012 0.15555 0 0.035785 0.0389 0 0.92413 0.26191 0.07138 0.0098906 4.3835 0.061727 7.4429e-05 0.82835 0.005404 0.0061432 0.001446 0.98617 0.9912 3.1259e-06 1.2504e-05 0.13294 0.83473 0.85701 0.0014283 0.92955 0.52731 0.0019231 0.42448 1.5783 1.5762 16.0096 144.9816 0.00025859 -85.3991 0.34136
1.4454 0.98803 5.5166e-05 3.8182 0.012031 1.9015e-05 0.0011543 0.16952 0.00065861 0.17017 0.1556 0 0.035781 0.0389 0 0.92421 0.26195 0.071394 0.0098923 4.384 0.061738 7.4442e-05 0.82834 0.0054045 0.0061437 0.0014455 0.98617 0.9912 3.1249e-06 1.25e-05 0.13294 0.83519 0.85729 0.0014281 0.92998 0.52748 0.0019228 0.42449 1.5795 1.5774 16.0096 144.9816 0.00025815 -85.401 0.34236
1.4464 0.98803 5.5166e-05 3.8182 0.012031 1.9028e-05 0.0011543 0.16957 0.00065861 0.17022 0.15565 0 0.035778 0.0389 0 0.92429 0.26199 0.071407 0.0098939 4.3845 0.061748 7.4455e-05 0.82833 0.0054049 0.0061442 0.0014451 0.98618 0.99121 3.1239e-06 1.2496e-05 0.13295 0.83565 0.85757 0.0014279 0.93041 0.52764 0.0019225 0.42451 1.5806 1.5786 16.0096 144.9816 0.0002577 -85.4028 0.34336
1.4474 0.98803 5.5166e-05 3.8182 0.012031 1.9041e-05 0.0011543 0.16962 0.00065861 0.17028 0.1557 0 0.035775 0.0389 0 0.92438 0.26202 0.071421 0.0098956 4.385 0.061758 7.4469e-05 0.82832 0.0054054 0.0061447 0.0014447 0.98619 0.99121 3.1229e-06 1.2491e-05 0.13295 0.83612 0.85784 0.0014276 0.93083 0.5278 0.0019222 0.42452 1.5818 1.5797 16.0096 144.9816 0.00025726 -85.4047 0.34436
1.4484 0.98803 5.5166e-05 3.8182 0.012031 1.9054e-05 0.0011543 0.16967 0.00065861 0.17033 0.15575 0 0.035772 0.0389 0 0.92446 0.26206 0.071435 0.0098972 4.3854 0.061768 7.4482e-05 0.82831 0.0054059 0.0061452 0.0014442 0.98619 0.99121 3.1219e-06 1.2487e-05 0.13295 0.83658 0.85812 0.0014274 0.93125 0.52796 0.0019219 0.42453 1.583 1.5809 16.0096 144.9817 0.00025682 -85.4065 0.34536
1.4494 0.98803 5.5166e-05 3.8182 0.012031 1.9068e-05 0.0011543 0.16973 0.00065862 0.17038 0.1558 0 0.035769 0.0389 0 0.92455 0.2621 0.071448 0.0098988 4.3859 0.061778 7.4495e-05 0.8283 0.0054064 0.0061456 0.0014438 0.9862 0.99122 3.1209e-06 1.2483e-05 0.13296 0.83703 0.85839 0.0014272 0.93167 0.52813 0.0019216 0.42454 1.5841 1.5821 16.0096 144.9817 0.00025638 -85.4083 0.34636
1.4504 0.98803 5.5166e-05 3.8182 0.012031 1.9081e-05 0.0011543 0.16978 0.00065862 0.17043 0.15585 0 0.035765 0.0389 0 0.92463 0.26214 0.071462 0.0099005 4.3864 0.061789 7.4508e-05 0.82829 0.0054068 0.0061461 0.0014433 0.9862 0.99122 3.1199e-06 1.2479e-05 0.13296 0.83749 0.85867 0.001427 0.93209 0.52829 0.0019213 0.42455 1.5853 1.5832 16.0096 144.9817 0.00025594 -85.4101 0.34736
1.4514 0.98803 5.5166e-05 3.8182 0.012031 1.9094e-05 0.0011543 0.16983 0.00065862 0.17049 0.15589 0 0.035762 0.0389 0 0.92472 0.26217 0.071475 0.0099021 4.3869 0.061799 7.4521e-05 0.82828 0.0054073 0.0061466 0.0014429 0.98621 0.99122 3.1189e-06 1.2476e-05 0.13297 0.83794 0.85894 0.0014267 0.9325 0.52845 0.001921 0.42457 1.5864 1.5844 16.0096 144.9817 0.0002555 -85.4119 0.34836
1.4524 0.98803 5.5166e-05 3.8182 0.012031 1.9107e-05 0.0011543 0.16989 0.00065862 0.17054 0.15594 0 0.035759 0.0389 0 0.9248 0.26221 0.071489 0.0099038 4.3874 0.061809 7.4535e-05 0.82827 0.0054078 0.0061471 0.0014425 0.98621 0.99123 3.1179e-06 1.2472e-05 0.13297 0.8384 0.85921 0.0014265 0.93291 0.52862 0.0019207 0.42458 1.5875 1.5855 16.0096 144.9817 0.00025507 -85.4137 0.34936
1.4534 0.98803 5.5166e-05 3.8182 0.012031 1.912e-05 0.0011543 0.16994 0.00065862 0.17059 0.15599 0 0.035756 0.0389 0 0.92489 0.26225 0.071503 0.0099054 4.3879 0.061819 7.4548e-05 0.82826 0.0054082 0.0061476 0.0014421 0.98622 0.99123 3.1169e-06 1.2468e-05 0.13297 0.83885 0.85948 0.0014263 0.93332 0.52878 0.0019204 0.42459 1.5887 1.5867 16.0096 144.9818 0.00025464 -85.4154 0.35036
1.4544 0.98803 5.5166e-05 3.8182 0.012031 1.9133e-05 0.0011543 0.16999 0.00065862 0.17064 0.15604 0 0.035753 0.0389 0 0.92497 0.26229 0.071516 0.0099071 4.3884 0.061829 7.4561e-05 0.82825 0.0054087 0.006148 0.0014416 0.98622 0.99124 3.116e-06 1.2464e-05 0.13298 0.8393 0.85975 0.0014261 0.93372 0.52894 0.0019201 0.4246 1.5898 1.5878 16.0096 144.9818 0.00025421 -85.4172 0.35136
1.4554 0.98803 5.5165e-05 3.8182 0.012031 1.9146e-05 0.0011543 0.17004 0.00065862 0.1707 0.15609 0 0.035749 0.0389 0 0.92506 0.26233 0.07153 0.0099087 4.3889 0.061839 7.4574e-05 0.82824 0.0054092 0.0061485 0.0014412 0.98623 0.99124 3.115e-06 1.246e-05 0.13298 0.83975 0.86002 0.0014259 0.93413 0.5291 0.0019199 0.42461 1.591 1.5889 16.0096 144.9818 0.00025378 -85.4189 0.35236
1.4564 0.98803 5.5165e-05 3.8182 0.012031 1.9159e-05 0.0011543 0.1701 0.00065862 0.17075 0.15614 0 0.035746 0.0389 0 0.92514 0.26236 0.071544 0.0099103 4.3893 0.06185 7.4587e-05 0.82822 0.0054097 0.006149 0.0014408 0.98624 0.99124 3.1141e-06 1.2456e-05 0.13299 0.8402 0.86029 0.0014256 0.93453 0.52927 0.0019196 0.42462 1.5921 1.5901 16.0096 144.9818 0.00025335 -85.4206 0.35336
1.4574 0.98803 5.5165e-05 3.8182 0.012031 1.9173e-05 0.0011543 0.17015 0.00065862 0.1708 0.15619 0 0.035743 0.0389 0 0.92523 0.2624 0.071557 0.009912 4.3898 0.06186 7.4601e-05 0.82821 0.0054101 0.0061495 0.0014404 0.98624 0.99125 3.1131e-06 1.2452e-05 0.13299 0.84065 0.86055 0.0014254 0.93492 0.52943 0.0019193 0.42464 1.5932 1.5912 16.0096 144.9818 0.00025293 -85.4223 0.35436
1.4584 0.98803 5.5165e-05 3.8182 0.01203 1.9186e-05 0.0011543 0.1702 0.00065862 0.17085 0.15624 0 0.03574 0.0389 0 0.92531 0.26244 0.071571 0.0099136 4.3903 0.06187 7.4614e-05 0.8282 0.0054106 0.00615 0.00144 0.98625 0.99125 3.1122e-06 1.2449e-05 0.13299 0.84109 0.86082 0.0014252 0.93532 0.52959 0.001919 0.42465 1.5943 1.5924 16.0096 144.9819 0.00025251 -85.424 0.35536
1.4594 0.98803 5.5165e-05 3.8182 0.01203 1.9199e-05 0.0011543 0.17025 0.00065862 0.17091 0.15629 0 0.035737 0.0389 0 0.9254 0.26248 0.071585 0.0099153 4.3908 0.06188 7.4627e-05 0.82819 0.0054111 0.0061505 0.0014396 0.98625 0.99125 3.1112e-06 1.2445e-05 0.133 0.84154 0.86108 0.001425 0.93571 0.52976 0.0019187 0.42466 1.5955 1.5935 16.0096 144.9819 0.00025208 -85.4257 0.35636
1.4604 0.98803 5.5165e-05 3.8182 0.01203 1.9212e-05 0.0011543 0.1703 0.00065862 0.17096 0.15634 0 0.035734 0.0389 0 0.92548 0.26251 0.071598 0.0099169 4.3913 0.061891 7.464e-05 0.82818 0.0054116 0.0061509 0.0014392 0.98626 0.99126 3.1103e-06 1.2441e-05 0.133 0.84198 0.86134 0.0014248 0.9361 0.52992 0.0019185 0.42467 1.5966 1.5946 16.0096 144.9819 0.00025166 -85.4274 0.35736
1.4614 0.98803 5.5165e-05 3.8182 0.01203 1.9225e-05 0.0011543 0.17036 0.00065862 0.17101 0.15639 0 0.03573 0.0389 0 0.92557 0.26255 0.071612 0.0099186 4.3918 0.061901 7.4653e-05 0.82817 0.005412 0.0061514 0.0014388 0.98626 0.99126 3.1094e-06 1.2438e-05 0.13301 0.84242 0.8616 0.0014246 0.93649 0.53008 0.0019182 0.42468 1.5977 1.5957 16.0096 144.9819 0.00025125 -85.4291 0.35836
1.4624 0.98803 5.5165e-05 3.8182 0.01203 1.9238e-05 0.0011543 0.17041 0.00065863 0.17106 0.15644 0 0.035727 0.0389 0 0.92565 0.26259 0.071626 0.0099202 4.3923 0.061911 7.4667e-05 0.82816 0.0054125 0.0061519 0.0014384 0.98627 0.99126 3.1085e-06 1.2434e-05 0.13301 0.84286 0.86187 0.0014244 0.93688 0.53024 0.0019179 0.4247 1.5988 1.5969 16.0097 144.9819 0.00025083 -85.4307 0.35936
1.4634 0.98803 5.5165e-05 3.8182 0.01203 1.9251e-05 0.0011543 0.17046 0.00065863 0.17112 0.15649 0 0.035724 0.0389 0 0.92574 0.26263 0.071639 0.0099219 4.3928 0.061921 7.468e-05 0.82815 0.005413 0.0061524 0.001438 0.98627 0.99127 3.1076e-06 1.243e-05 0.13301 0.8433 0.86212 0.0014242 0.93726 0.53041 0.0019177 0.42471 1.5999 1.598 16.0097 144.9819 0.00025042 -85.4324 0.36036
1.4644 0.98803 5.5165e-05 3.8182 0.01203 1.9264e-05 0.0011543 0.17051 0.00065863 0.17117 0.15653 0 0.035721 0.0389 0 0.92582 0.26267 0.071653 0.0099235 4.3933 0.061931 7.4693e-05 0.82814 0.0054135 0.0061529 0.0014376 0.98628 0.99127 3.1067e-06 1.2427e-05 0.13302 0.84373 0.86238 0.001424 0.93764 0.53057 0.0019174 0.42472 1.601 1.5991 16.0097 144.982 0.00025001 -85.434 0.36136
1.4654 0.98803 5.5165e-05 3.8182 0.01203 1.9278e-05 0.0011543 0.17057 0.00065863 0.17122 0.15658 0 0.035718 0.0389 0 0.92591 0.2627 0.071667 0.0099252 4.3938 0.061942 7.4706e-05 0.82813 0.0054139 0.0061534 0.0014372 0.98628 0.99127 3.1058e-06 1.2423e-05 0.13302 0.84417 0.86264 0.0014238 0.93802 0.53073 0.0019171 0.42473 1.6021 1.6002 16.0097 144.982 0.0002496 -85.4356 0.36236
1.4664 0.98803 5.5165e-05 3.8182 0.01203 1.9291e-05 0.0011543 0.17062 0.00065863 0.17127 0.15663 0 0.035715 0.0389 0 0.92599 0.26274 0.07168 0.0099268 4.3942 0.061952 7.472e-05 0.82812 0.0054144 0.0061539 0.0014368 0.98629 0.99128 3.1049e-06 1.242e-05 0.13303 0.8446 0.8629 0.0014236 0.9384 0.53089 0.0019169 0.42474 1.6032 1.6013 16.0097 144.982 0.00024919 -85.4372 0.36336
1.4674 0.98803 5.5165e-05 3.8182 0.01203 1.9304e-05 0.0011543 0.17067 0.00065863 0.17132 0.15668 0 0.035712 0.0389 0 0.92608 0.26278 0.071694 0.0099285 4.3947 0.061962 7.4733e-05 0.82811 0.0054149 0.0061543 0.0014365 0.98629 0.99128 3.104e-06 1.2416e-05 0.13303 0.84504 0.86315 0.0014234 0.93877 0.53105 0.0019166 0.42476 1.6043 1.6024 16.0097 144.982 0.00024878 -85.4388 0.36436
1.4684 0.98803 5.5165e-05 3.8182 0.01203 1.9317e-05 0.0011543 0.17072 0.00065863 0.17138 0.15673 0 0.035708 0.0389 0 0.92616 0.26282 0.071708 0.0099301 4.3952 0.061972 7.4746e-05 0.8281 0.0054154 0.0061548 0.0014361 0.9863 0.99128 3.1032e-06 1.2413e-05 0.13303 0.84547 0.86341 0.0014232 0.93914 0.53122 0.0019164 0.42477 1.6054 1.6035 16.0097 144.982 0.00024837 -85.4404 0.36536
1.4694 0.98803 5.5165e-05 3.8182 0.01203 1.933e-05 0.0011543 0.17077 0.00065863 0.17143 0.15678 0 0.035705 0.0389 0 0.92625 0.26286 0.071721 0.0099317 4.3957 0.061982 7.4759e-05 0.82809 0.0054159 0.0061553 0.0014357 0.9863 0.99129 3.1023e-06 1.2409e-05 0.13304 0.8459 0.86366 0.001423 0.93951 0.53138 0.0019161 0.42478 1.6065 1.6046 16.0097 144.9821 0.00024797 -85.442 0.36636
1.4704 0.98803 5.5165e-05 3.8182 0.01203 1.9343e-05 0.0011543 0.17083 0.00065863 0.17148 0.15683 0 0.035702 0.0389 0 0.92633 0.26289 0.071735 0.0099334 4.3962 0.061993 7.4773e-05 0.82808 0.0054163 0.0061558 0.0014353 0.98631 0.99129 3.1015e-06 1.2406e-05 0.13304 0.84633 0.86391 0.0014228 0.93988 0.53154 0.0019158 0.42479 1.6076 1.6057 16.0097 144.9821 0.00024757 -85.4435 0.36736
1.4714 0.98803 5.5164e-05 3.8182 0.01203 1.9356e-05 0.0011543 0.17088 0.00065863 0.17153 0.15688 0 0.035699 0.0389 0 0.92642 0.26293 0.071749 0.009935 4.3967 0.062003 7.4786e-05 0.82807 0.0054168 0.0061563 0.001435 0.98631 0.99129 3.1006e-06 1.2402e-05 0.13305 0.84676 0.86416 0.0014226 0.94025 0.5317 0.0019156 0.42481 1.6087 1.6068 16.0097 144.9821 0.00024717 -85.4451 0.36836
1.4724 0.98803 5.5164e-05 3.8182 0.01203 1.9369e-05 0.0011543 0.17093 0.00065863 0.17158 0.15693 0 0.035696 0.0389 0 0.9265 0.26297 0.071763 0.0099367 4.3972 0.062013 7.4799e-05 0.82806 0.0054173 0.0061568 0.0014346 0.98632 0.9913 3.0998e-06 1.2399e-05 0.13305 0.84718 0.86441 0.0014224 0.94061 0.53186 0.0019153 0.42482 1.6098 1.6079 16.0097 144.9821 0.00024677 -85.4466 0.36936
1.4734 0.98803 5.5164e-05 3.8182 0.01203 1.9383e-05 0.0011543 0.17098 0.00065863 0.17164 0.15697 0 0.035693 0.0389 0 0.92659 0.26301 0.071776 0.0099383 4.3977 0.062023 7.4812e-05 0.82805 0.0054178 0.0061573 0.0014342 0.98632 0.9913 3.0989e-06 1.2396e-05 0.13305 0.84761 0.86466 0.0014222 0.94097 0.53203 0.0019151 0.42483 1.6109 1.609 16.0097 144.9821 0.00024637 -85.4481 0.37036
1.4744 0.98803 5.5164e-05 3.8182 0.01203 1.9396e-05 0.0011543 0.17103 0.00065863 0.17169 0.15702 0 0.03569 0.0389 0 0.92667 0.26305 0.07179 0.00994 4.3982 0.062034 7.4826e-05 0.82804 0.0054182 0.0061578 0.0014339 0.98633 0.9913 3.0981e-06 1.2392e-05 0.13306 0.84803 0.86491 0.001422 0.94133 0.53219 0.0019148 0.42484 1.6119 1.6101 16.0097 144.9822 0.00024598 -85.4497 0.37136
1.4754 0.98803 5.5164e-05 3.8182 0.01203 1.9409e-05 0.0011543 0.17108 0.00065864 0.17174 0.15707 0 0.035687 0.0389 0 0.92676 0.26308 0.071804 0.0099416 4.3987 0.062044 7.4839e-05 0.82803 0.0054187 0.0061582 0.0014335 0.98633 0.99131 3.0973e-06 1.2389e-05 0.13306 0.84845 0.86515 0.0014218 0.94168 0.53235 0.0019146 0.42485 1.613 1.6111 16.0097 144.9822 0.00024559 -85.4512 0.37236
1.4764 0.98803 5.5164e-05 3.8182 0.01203 1.9422e-05 0.0011543 0.17114 0.00065864 0.17179 0.15712 0 0.035684 0.0389 0 0.92684 0.26312 0.071817 0.0099433 4.3992 0.062054 7.4852e-05 0.82802 0.0054192 0.0061587 0.0014331 0.98634 0.99131 3.0964e-06 1.2386e-05 0.13307 0.84887 0.8654 0.0014217 0.94204 0.53251 0.0019144 0.42487 1.6141 1.6122 16.0097 144.9822 0.0002452 -85.4527 0.37336
1.4774 0.98803 5.5164e-05 3.8182 0.01203 1.9435e-05 0.0011543 0.17119 0.00065864 0.17184 0.15717 0 0.03568 0.0389 0 0.92693 0.26316 0.071831 0.009945 4.3997 0.062064 7.4866e-05 0.82801 0.0054197 0.0061592 0.0014328 0.98634 0.99131 3.0956e-06 1.2383e-05 0.13307 0.84929 0.86564 0.0014215 0.94239 0.53267 0.0019141 0.42488 1.6152 1.6133 16.0097 144.9822 0.00024481 -85.4542 0.37436
1.4784 0.98803 5.5164e-05 3.8182 0.01203 1.9448e-05 0.0011543 0.17124 0.00065864 0.17189 0.15722 0 0.035677 0.0389 0 0.92701 0.2632 0.071845 0.0099466 4.4002 0.062075 7.4879e-05 0.828 0.0054202 0.0061597 0.0014324 0.98635 0.99131 3.0948e-06 1.2379e-05 0.13307 0.84971 0.86589 0.0014213 0.94274 0.53283 0.0019139 0.42489 1.6162 1.6144 16.0097 144.9822 0.00024442 -85.4556 0.37536
1.4794 0.98803 5.5164e-05 3.8182 0.01203 1.9461e-05 0.0011543 0.17129 0.00065864 0.17195 0.15727 0 0.035674 0.0389 0 0.9271 0.26324 0.071859 0.0099483 4.4007 0.062085 7.4892e-05 0.82799 0.0054206 0.0061602 0.0014321 0.98635 0.99132 3.094e-06 1.2376e-05 0.13308 0.85013 0.86613 0.0014211 0.94308 0.533 0.0019136 0.4249 1.6173 1.6154 16.0097 144.9822 0.00024403 -85.4571 0.37636
1.4804 0.98803 5.5164e-05 3.8182 0.01203 1.9474e-05 0.0011543 0.17134 0.00065864 0.172 0.15731 0 0.035671 0.0389 0 0.92718 0.26327 0.071872 0.0099499 4.4012 0.062095 7.4905e-05 0.82798 0.0054211 0.0061607 0.0014317 0.98635 0.99132 3.0932e-06 1.2373e-05 0.13308 0.85055 0.86637 0.0014209 0.94343 0.53316 0.0019134 0.42491 1.6184 1.6165 16.0097 144.9823 0.00024365 -85.4586 0.37736
1.4814 0.98803 5.5164e-05 3.8182 0.01203 1.9488e-05 0.0011543 0.17139 0.00065864 0.17205 0.15736 0 0.035668 0.0389 0 0.92727 0.26331 0.071886 0.0099516 4.4017 0.062105 7.4919e-05 0.82797 0.0054216 0.0061612 0.0014314 0.98636 0.99132 3.0924e-06 1.237e-05 0.13308 0.85096 0.86661 0.0014207 0.94377 0.53332 0.0019132 0.42493 1.6194 1.6176 16.0097 144.9823 0.00024326 -85.46 0.37836
1.4824 0.98803 5.5164e-05 3.8182 0.01203 1.9501e-05 0.0011543 0.17145 0.00065864 0.1721 0.15741 0 0.035665 0.0389 0 0.92735 0.26335 0.0719 0.0099532 4.4022 0.062116 7.4932e-05 0.82796 0.0054221 0.0061617 0.001431 0.98636 0.99133 3.0916e-06 1.2367e-05 0.13309 0.85137 0.86685 0.0014206 0.94411 0.53348 0.0019129 0.42494 1.6205 1.6186 16.0097 144.9823 0.00024288 -85.4614 0.37936
1.4834 0.98803 5.5164e-05 3.8182 0.01203 1.9514e-05 0.0011543 0.1715 0.00065864 0.17215 0.15746 0 0.035662 0.0389 0 0.92744 0.26339 0.071913 0.0099549 4.4027 0.062126 7.4945e-05 0.82795 0.0054226 0.0061622 0.0014307 0.98637 0.99133 3.0909e-06 1.2363e-05 0.13309 0.85179 0.86709 0.0014204 0.94445 0.53364 0.0019127 0.42495 1.6215 1.6197 16.0097 144.9823 0.0002425 -85.4629 0.38036
1.4844 0.98803 5.5164e-05 3.8182 0.01203 1.9527e-05 0.0011543 0.17155 0.00065864 0.1722 0.15751 0 0.035659 0.0389 0 0.92753 0.26343 0.071927 0.0099565 4.4032 0.062136 7.4959e-05 0.82794 0.0054231 0.0061627 0.0014304 0.98637 0.99133 3.0901e-06 1.236e-05 0.1331 0.8522 0.86733 0.0014202 0.94479 0.5338 0.0019125 0.42496 1.6226 1.6207 16.0097 144.9823 0.00024212 -85.4643 0.38136
1.4854 0.98803 5.5164e-05 3.8182 0.01203 1.954e-05 0.0011543 0.1716 0.00065864 0.17225 0.15756 0 0.035656 0.0389 0 0.92761 0.26347 0.071941 0.0099582 4.4037 0.062146 7.4972e-05 0.82793 0.0054235 0.0061632 0.00143 0.98638 0.99134 3.0893e-06 1.2357e-05 0.1331 0.85261 0.86757 0.00142 0.94512 0.53396 0.0019122 0.42498 1.6236 1.6218 16.0097 144.9824 0.00024174 -85.4657 0.38236
1.4864 0.98803 5.5164e-05 3.8182 0.01203 1.9553e-05 0.0011543 0.17165 0.00065864 0.1723 0.1576 0 0.035653 0.0389 0 0.9277 0.2635 0.071955 0.0099598 4.4042 0.062157 7.4985e-05 0.82792 0.005424 0.0061637 0.0014297 0.98638 0.99134 3.0886e-06 1.2354e-05 0.1331 0.85301 0.8678 0.0014199 0.94545 0.53413 0.001912 0.42499 1.6247 1.6228 16.0097 144.9824 0.00024137 -85.4671 0.38336
1.4874 0.98803 5.5163e-05 3.8182 0.01203 1.9566e-05 0.0011543 0.1717 0.00065864 0.17236 0.15765 0 0.03565 0.0389 0 0.92778 0.26354 0.071968 0.0099615 4.4047 0.062167 7.4999e-05 0.82791 0.0054245 0.0061641 0.0014294 0.98639 0.99134 3.0878e-06 1.2351e-05 0.13311 0.85342 0.86804 0.0014197 0.94578 0.53429 0.0019118 0.425 1.6257 1.6239 16.0097 144.9824 0.000241 -85.4685 0.38436
1.4884 0.98803 5.5163e-05 3.8182 0.01203 1.9579e-05 0.0011543 0.17175 0.00065865 0.17241 0.1577 0 0.035646 0.0389 0 0.92787 0.26358 0.071982 0.0099631 4.4052 0.062177 7.5012e-05 0.8279 0.005425 0.0061646 0.001429 0.98639 0.99134 3.087e-06 1.2348e-05 0.13311 0.85383 0.86827 0.0014195 0.94611 0.53445 0.0019116 0.42501 1.6267 1.6249 16.0097 144.9824 0.00024062 -85.4698 0.38536
1.4894 0.98803 5.5163e-05 3.8182 0.01203 1.9593e-05 0.0011543 0.1718 0.00065865 0.17246 0.15775 0 0.035643 0.0389 0 0.92795 0.26362 0.071996 0.0099648 4.4057 0.062187 7.5025e-05 0.82789 0.0054255 0.0061651 0.0014287 0.98639 0.99135 3.0863e-06 1.2345e-05 0.13312 0.85423 0.8685 0.0014193 0.94644 0.53461 0.0019113 0.42503 1.6278 1.626 16.0097 144.9824 0.00024025 -85.4712 0.38636
1.4904 0.98803 5.5163e-05 3.8182 0.01203 1.9606e-05 0.0011543 0.17186 0.00065865 0.17251 0.1578 0 0.03564 0.0389 0 0.92804 0.26366 0.07201 0.0099665 4.4062 0.062198 7.5039e-05 0.82788 0.005426 0.0061656 0.0014284 0.9864 0.99135 3.0856e-06 1.2342e-05 0.13312 0.85463 0.86874 0.0014192 0.94676 0.53477 0.0019111 0.42504 1.6288 1.627 16.0097 144.9825 0.00023988 -85.4726 0.38736
1.4914 0.98803 5.5163e-05 3.8182 0.01203 1.9619e-05 0.0011543 0.17191 0.00065865 0.17256 0.15784 0 0.035637 0.0389 0 0.92812 0.26369 0.072024 0.0099681 4.4067 0.062208 7.5052e-05 0.82787 0.0054264 0.0061661 0.0014281 0.9864 0.99135 3.0848e-06 1.2339e-05 0.13312 0.85504 0.86897 0.001419 0.94708 0.53493 0.0019109 0.42505 1.6298 1.628 16.0097 144.9825 0.00023952 -85.4739 0.38836
1.4924 0.98803 5.5163e-05 3.8182 0.01203 1.9632e-05 0.0011543 0.17196 0.00065865 0.17261 0.15789 0 0.035634 0.0389 0 0.92821 0.26373 0.072037 0.0099698 4.4072 0.062218 7.5065e-05 0.82786 0.0054269 0.0061666 0.0014277 0.98641 0.99135 3.0841e-06 1.2336e-05 0.13313 0.85544 0.8692 0.0014188 0.9474 0.53509 0.0019107 0.42506 1.6309 1.6291 16.0097 144.9825 0.00023915 -85.4753 0.38936
1.4934 0.98803 5.5163e-05 3.8182 0.01203 1.9645e-05 0.0011543 0.17201 0.00065865 0.17266 0.15794 0 0.035631 0.0389 0 0.9283 0.26377 0.072051 0.0099714 4.4077 0.062229 7.5079e-05 0.82785 0.0054274 0.0061671 0.0014274 0.98641 0.99136 3.0834e-06 1.2333e-05 0.13313 0.85584 0.86943 0.0014187 0.94772 0.53525 0.0019105 0.42507 1.6319 1.6301 16.0097 144.9825 0.00023878 -85.4766 0.39036
1.4944 0.98803 5.5163e-05 3.8182 0.01203 1.9658e-05 0.0011543 0.17206 0.00065865 0.17271 0.15799 0 0.035628 0.0389 0 0.92838 0.26381 0.072065 0.0099731 4.4082 0.062239 7.5092e-05 0.82784 0.0054279 0.0061676 0.0014271 0.98641 0.99136 3.0827e-06 1.2331e-05 0.13314 0.85623 0.86965 0.0014185 0.94804 0.53541 0.0019103 0.42509 1.6329 1.6311 16.0097 144.9825 0.00023842 -85.4779 0.39136
1.4954 0.98803 5.5163e-05 3.8182 0.01203 1.9671e-05 0.0011543 0.17211 0.00065865 0.17276 0.15803 0 0.035625 0.0389 0 0.92847 0.26385 0.072079 0.0099747 4.4087 0.062249 7.5105e-05 0.82783 0.0054284 0.0061681 0.0014268 0.98642 0.99136 3.0819e-06 1.2328e-05 0.13314 0.85663 0.86988 0.0014184 0.94835 0.53558 0.00191 0.4251 1.6339 1.6322 16.0097 144.9826 0.00023806 -85.4792 0.39236
1.4964 0.98803 5.5163e-05 3.8182 0.01203 1.9684e-05 0.0011543 0.17216 0.00065865 0.17281 0.15808 0 0.035622 0.0389 0 0.92855 0.26389 0.072092 0.0099764 4.4092 0.062259 7.5119e-05 0.82782 0.0054289 0.0061686 0.0014265 0.98642 0.99137 3.0812e-06 1.2325e-05 0.13315 0.85703 0.87011 0.0014182 0.94867 0.53574 0.0019098 0.42511 1.6349 1.6332 16.0097 144.9826 0.0002377 -85.4805 0.39336
1.4974 0.98803 5.5163e-05 3.8182 0.01203 1.9698e-05 0.0011543 0.17221 0.00065865 0.17287 0.15813 0 0.035619 0.0389 0 0.92864 0.26392 0.072106 0.009978 4.4098 0.06227 7.5132e-05 0.82781 0.0054294 0.0061691 0.0014262 0.98643 0.99137 3.0805e-06 1.2322e-05 0.13315 0.85742 0.87033 0.001418 0.94898 0.5359 0.0019096 0.42512 1.6359 1.6342 16.0097 144.9826 0.00023734 -85.4818 0.39436
1.4984 0.98803 5.5163e-05 3.8182 0.01203 1.9711e-05 0.0011543 0.17226 0.00065865 0.17292 0.15818 0 0.035616 0.0389 0 0.92872 0.26396 0.07212 0.0099797 4.4103 0.06228 7.5145e-05 0.8278 0.0054298 0.0061696 0.0014259 0.98643 0.99137 3.0798e-06 1.2319e-05 0.13315 0.85782 0.87056 0.0014179 0.94928 0.53606 0.0019094 0.42514 1.637 1.6352 16.0097 144.9826 0.00023698 -85.4831 0.39536
1.4994 0.98803 5.5163e-05 3.8182 0.01203 1.9724e-05 0.0011543 0.17231 0.00065865 0.17297 0.15823 0 0.035613 0.0389 0 0.92881 0.264 0.072134 0.0099814 4.4108 0.06229 7.5159e-05 0.82778 0.0054303 0.0061701 0.0014256 0.98643 0.99137 3.0791e-06 1.2316e-05 0.13316 0.85821 0.87078 0.0014177 0.94959 0.53622 0.0019092 0.42515 1.638 1.6362 16.0097 144.9826 0.00023663 -85.4844 0.39636
1.5004 0.98803 5.5163e-05 3.8182 0.01203 1.9737e-05 0.0011543 0.17236 0.00065865 0.17302 0.15827 0 0.03561 0.0389 0 0.92889 0.26404 0.072148 0.009983 4.4113 0.062301 7.5172e-05 0.82777 0.0054308 0.0061706 0.0014253 0.98644 0.99138 3.0784e-06 1.2314e-05 0.13316 0.8586 0.871 0.0014176 0.94989 0.53638 0.001909 0.42516 1.639 1.6372 16.0097 144.9826 0.00023628 -85.4856 0.39736
1.5014 0.98803 5.5163e-05 3.8182 0.01203 1.975e-05 0.0011543 0.17241 0.00065865 0.17307 0.15832 0 0.035607 0.0389 0 0.92898 0.26408 0.072161 0.0099847 4.4118 0.062311 7.5185e-05 0.82776 0.0054313 0.0061711 0.001425 0.98644 0.99138 3.0778e-06 1.2311e-05 0.13317 0.85899 0.87123 0.0014174 0.9502 0.53654 0.0019088 0.42517 1.64 1.6382 16.0096 144.9827 0.00023592 -85.4869 0.39836
1.5024 0.98803 5.5163e-05 3.8182 0.01203 1.9763e-05 0.0011543 0.17246 0.00065866 0.17312 0.15837 0 0.035604 0.0389 0 0.92907 0.26412 0.072175 0.0099863 4.4123 0.062321 7.5199e-05 0.82775 0.0054318 0.0061716 0.0014247 0.98645 0.99138 3.0771e-06 1.2308e-05 0.13317 0.85938 0.87145 0.0014172 0.9505 0.5367 0.0019086 0.42519 1.641 1.6392 16.0096 144.9827 0.00023557 -85.4881 0.39936
1.5034 0.98803 5.5162e-05 3.8182 0.01203 1.9776e-05 0.0011543 0.17252 0.00065866 0.17317 0.15842 0 0.035601 0.0389 0 0.92915 0.26415 0.072189 0.009988 4.4128 0.062332 7.5212e-05 0.82774 0.0054323 0.0061721 0.0014244 0.98645 0.99138 3.0764e-06 1.2306e-05 0.13317 0.85976 0.87167 0.0014171 0.9508 0.53686 0.0019084 0.4252 1.642 1.6402 16.0096 144.9827 0.00023522 -85.4894 0.40036
1.5044 0.98803 5.5162e-05 3.8182 0.01203 1.9789e-05 0.0011543 0.17257 0.00065866 0.17322 0.15846 0 0.035598 0.0389 0 0.92924 0.26419 0.072203 0.0099897 4.4133 0.062342 7.5225e-05 0.82773 0.0054328 0.0061726 0.0014241 0.98645 0.99139 3.0757e-06 1.2303e-05 0.13318 0.86015 0.87189 0.0014169 0.95109 0.53702 0.0019082 0.42521 1.643 1.6412 16.0096 144.9827 0.00023487 -85.4906 0.40136
1.5054 0.98803 5.5162e-05 3.8182 0.01203 1.9802e-05 0.0011543 0.17262 0.00065866 0.17327 0.15851 0 0.035595 0.0389 0 0.92932 0.26423 0.072217 0.0099913 4.4138 0.062352 7.5239e-05 0.82772 0.0054333 0.0061731 0.0014238 0.98646 0.99139 3.0751e-06 1.23e-05 0.13318 0.86053 0.87211 0.0014168 0.95139 0.53718 0.001908 0.42522 1.644 1.6422 16.0096 144.9827 0.00023453 -85.4918 0.40236
1.5064 0.98803 5.5162e-05 3.8182 0.01203 1.9816e-05 0.0011543 0.17267 0.00065866 0.17332 0.15856 0 0.035592 0.0389 0 0.92941 0.26427 0.07223 0.009993 4.4143 0.062362 7.5252e-05 0.82771 0.0054337 0.0061736 0.0014235 0.98646 0.99139 3.0744e-06 1.2298e-05 0.13319 0.86092 0.87232 0.0014166 0.95168 0.53734 0.0019078 0.42524 1.6449 1.6432 16.0096 144.9828 0.00023418 -85.493 0.40336
1.5074 0.98803 5.5162e-05 3.8182 0.01203 1.9829e-05 0.0011543 0.17272 0.00065866 0.17337 0.15861 0 0.035589 0.0389 0 0.9295 0.26431 0.072244 0.0099946 4.4148 0.062373 7.5266e-05 0.8277 0.0054342 0.0061741 0.0014232 0.98647 0.99139 3.0737e-06 1.2295e-05 0.13319 0.8613 0.87254 0.0014165 0.95197 0.5375 0.0019076 0.42525 1.6459 1.6442 16.0096 144.9828 0.00023384 -85.4942 0.40436
1.5084 0.98803 5.5162e-05 3.8182 0.01203 1.9842e-05 0.0011543 0.17277 0.00065866 0.17342 0.15865 0 0.035586 0.0389 0 0.92958 0.26435 0.072258 0.0099963 4.4154 0.062383 7.5279e-05 0.82769 0.0054347 0.0061746 0.0014229 0.98647 0.9914 3.0731e-06 1.2292e-05 0.13319 0.86168 0.87275 0.0014163 0.95226 0.53766 0.0019074 0.42526 1.6469 1.6452 16.0096 144.9828 0.0002335 -85.4954 0.40536
1.5094 0.98803 5.5162e-05 3.8182 0.01203 1.9855e-05 0.0011543 0.17282 0.00065866 0.17347 0.1587 0 0.035583 0.0389 0 0.92967 0.26438 0.072272 0.009998 4.4159 0.062393 7.5292e-05 0.82768 0.0054352 0.0061751 0.0014227 0.98647 0.9914 3.0724e-06 1.229e-05 0.1332 0.86206 0.87297 0.0014162 0.95255 0.53782 0.0019072 0.42527 1.6479 1.6462 16.0096 144.9828 0.00023315 -85.4966 0.40636
1.5104 0.98803 5.5162e-05 3.8182 0.01203 1.9868e-05 0.0011543 0.17287 0.00065866 0.17352 0.15875 0 0.03558 0.0389 0 0.92975 0.26442 0.072286 0.0099996 4.4164 0.062404 7.5306e-05 0.82767 0.0054357 0.0061756 0.0014224 0.98648 0.9914 3.0718e-06 1.2287e-05 0.1332 0.86244 0.87318 0.001416 0.95283 0.53798 0.001907 0.42529 1.6489 1.6472 16.0096 144.9828 0.00023281 -85.4978 0.40736
1.5114 0.98803 5.5162e-05 3.8182 0.01203 1.9881e-05 0.0011543 0.17292 0.00065866 0.17357 0.15879 0 0.035577 0.0389 0 0.92984 0.26446 0.0723 0.010001 4.4169 0.062414 7.5319e-05 0.82766 0.0054362 0.0061761 0.0014221 0.98648 0.9914 3.0712e-06 1.2285e-05 0.13321 0.86282 0.8734 0.0014159 0.95312 0.53814 0.0019068 0.4253 1.6498 1.6482 16.0096 144.9829 0.00023248 -85.499 0.40836
1.5124 0.98803 5.5162e-05 3.8182 0.01203 1.9894e-05 0.0011543 0.17297 0.00065866 0.17362 0.15884 0 0.035574 0.0389 0 0.92993 0.2645 0.072313 0.010003 4.4174 0.062424 7.5333e-05 0.82765 0.0054367 0.0061766 0.0014218 0.98648 0.9914 3.0705e-06 1.2282e-05 0.13321 0.86319 0.87361 0.0014158 0.9534 0.5383 0.0019066 0.42531 1.6508 1.6491 16.0096 144.9829 0.00023214 -85.5001 0.40936
1.5134 0.98803 5.5162e-05 3.8182 0.01203 1.9907e-05 0.0011544 0.17302 0.00065866 0.17367 0.15889 0 0.035571 0.0389 0 0.93001 0.26454 0.072327 0.010005 4.4179 0.062435 7.5346e-05 0.82764 0.0054372 0.0061771 0.0014216 0.98649 0.99141 3.0699e-06 1.228e-05 0.13321 0.86357 0.87382 0.0014156 0.95368 0.53846 0.0019065 0.42532 1.6518 1.6501 16.0096 144.9829 0.0002318 -85.5013 0.41036
1.5144 0.98803 5.5162e-05 3.8182 0.01203 1.9921e-05 0.0011544 0.17307 0.00065866 0.17372 0.15894 0 0.035568 0.0389 0 0.9301 0.26458 0.072341 0.010006 4.4184 0.062445 7.5359e-05 0.82763 0.0054377 0.0061776 0.0014213 0.98649 0.99141 3.0693e-06 1.2277e-05 0.13322 0.86394 0.87403 0.0014155 0.95396 0.53862 0.0019063 0.42534 1.6528 1.6511 16.0096 144.9829 0.00023147 -85.5025 0.41136
1.5154 0.98803 5.5162e-05 3.8182 0.01203 1.9934e-05 0.0011544 0.17312 0.00065867 0.17377 0.15898 0 0.035565 0.0389 0 0.93018 0.26461 0.072355 0.010008 4.419 0.062455 7.5373e-05 0.82762 0.0054382 0.0061781 0.001421 0.98649 0.99141 3.0687e-06 1.2275e-05 0.13322 0.86432 0.87424 0.0014153 0.95424 0.53878 0.0019061 0.42535 1.6537 1.6521 16.0096 144.9829 0.00023114 -85.5036 0.41236
1.5164 0.98803 5.5162e-05 3.8182 0.01203 1.9947e-05 0.0011544 0.17317 0.00065867 0.17382 0.15903 0 0.035562 0.0389 0 0.93027 0.26465 0.072369 0.01001 4.4195 0.062466 7.5386e-05 0.82761 0.0054387 0.0061786 0.0014207 0.9865 0.99141 3.0681e-06 1.2272e-05 0.13323 0.86469 0.87445 0.0014152 0.95451 0.53894 0.0019059 0.42536 1.6547 1.653 16.0096 144.983 0.00023081 -85.5047 0.41336
1.5174 0.98803 5.5162e-05 3.8182 0.01203 1.996e-05 0.0011544 0.17322 0.00065867 0.17387 0.15908 0 0.035559 0.0389 0 0.93036 0.26469 0.072383 0.010011 4.42 0.062476 7.54e-05 0.8276 0.0054391 0.0061791 0.0014205 0.9865 0.99142 3.0674e-06 1.227e-05 0.13323 0.86506 0.87466 0.0014151 0.95479 0.5391 0.0019057 0.42537 1.6556 1.654 16.0096 144.983 0.00023048 -85.5058 0.41436
1.5184 0.98803 5.5161e-05 3.8182 0.01203 1.9973e-05 0.0011544 0.17327 0.00065867 0.17392 0.15912 0 0.035556 0.0389 0 0.93044 0.26473 0.072397 0.010013 4.4205 0.062486 7.5413e-05 0.82759 0.0054396 0.0061796 0.0014202 0.9865 0.99142 3.0668e-06 1.2267e-05 0.13323 0.86543 0.87487 0.0014149 0.95506 0.53926 0.0019055 0.42539 1.6566 1.655 16.0096 144.983 0.00023015 -85.507 0.41536
1.5194 0.98803 5.5161e-05 3.8182 0.01203 1.9986e-05 0.0011544 0.17332 0.00065867 0.17397 0.15917 0 0.035553 0.0389 0 0.93053 0.26477 0.07241 0.010015 4.421 0.062497 7.5426e-05 0.82758 0.0054401 0.0061801 0.00142 0.98651 0.99142 3.0662e-06 1.2265e-05 0.13324 0.8658 0.87507 0.0014148 0.95533 0.53942 0.0019054 0.4254 1.6576 1.6559 16.0096 144.983 0.00022982 -85.5081 0.41636
1.5204 0.98803 5.5161e-05 3.8182 0.01203 1.9999e-05 0.0011544 0.17337 0.00065867 0.17402 0.15922 0 0.03555 0.0389 0 0.93061 0.26481 0.072424 0.010016 4.4215 0.062507 7.544e-05 0.82757 0.0054406 0.0061806 0.0014197 0.98651 0.99142 3.0656e-06 1.2263e-05 0.13324 0.86616 0.87528 0.0014146 0.9556 0.53958 0.0019052 0.42541 1.6585 1.6569 16.0096 144.983 0.00022949 -85.5092 0.41736
1.5214 0.98803 5.5161e-05 3.8182 0.01203 2.0012e-05 0.0011544 0.17342 0.00065867 0.17407 0.15926 0 0.035547 0.0389 0 0.9307 0.26484 0.072438 0.010018 4.4221 0.062517 7.5453e-05 0.82756 0.0054411 0.0061811 0.0014194 0.98651 0.99143 3.065e-06 1.226e-05 0.13325 0.86653 0.87548 0.0014145 0.95586 0.53974 0.001905 0.42542 1.6595 1.6578 16.0096 144.983 0.00022917 -85.5103 0.41836
1.5224 0.98803 5.5161e-05 3.8182 0.01203 2.0026e-05 0.0011544 0.17347 0.00065867 0.17412 0.15931 0 0.035544 0.0389 0 0.93079 0.26488 0.072452 0.01002 4.4226 0.062528 7.5467e-05 0.82755 0.0054416 0.0061816 0.0014192 0.98652 0.99143 3.0645e-06 1.2258e-05 0.13325 0.8669 0.87569 0.0014144 0.95613 0.5399 0.0019048 0.42544 1.6604 1.6588 16.0096 144.9831 0.00022885 -85.5114 0.41936
1.5234 0.98803 5.5161e-05 3.8182 0.01203 2.0039e-05 0.0011544 0.17352 0.00065867 0.17417 0.15936 0 0.035541 0.0389 0 0.93087 0.26492 0.072466 0.010021 4.4231 0.062538 7.548e-05 0.82754 0.0054421 0.0061821 0.0014189 0.98652 0.99143 3.0639e-06 1.2255e-05 0.13325 0.86726 0.87589 0.0014142 0.95639 0.54006 0.0019047 0.42545 1.6614 1.6597 16.0096 144.9831 0.00022852 -85.5124 0.42036
1.5244 0.98803 5.5161e-05 3.8182 0.01203 2.0052e-05 0.0011544 0.17357 0.00065867 0.17422 0.15941 0 0.035538 0.0389 0 0.93096 0.26496 0.07248 0.010023 4.4236 0.062548 7.5493e-05 0.82753 0.0054426 0.0061826 0.0014187 0.98652 0.99143 3.0633e-06 1.2253e-05 0.13326 0.86762 0.87609 0.0014141 0.95665 0.54022 0.0019045 0.42546 1.6623 1.6607 16.0096 144.9831 0.0002282 -85.5135 0.42136
1.5254 0.98803 5.5161e-05 3.8182 0.01203 2.0065e-05 0.0011544 0.17362 0.00065867 0.17427 0.15945 0 0.035535 0.0389 0 0.93104 0.265 0.072494 0.010025 4.4241 0.062559 7.5507e-05 0.82752 0.0054431 0.0061831 0.0014184 0.98653 0.99143 3.0627e-06 1.2251e-05 0.13326 0.86798 0.87629 0.001414 0.95691 0.54038 0.0019043 0.42547 1.6632 1.6616 16.0095 144.9831 0.00022788 -85.5146 0.42236
1.5264 0.98803 5.5161e-05 3.8182 0.01203 2.0078e-05 0.0011544 0.17367 0.00065867 0.17432 0.1595 0 0.035532 0.0389 0 0.93113 0.26504 0.072508 0.010026 4.4247 0.062569 7.552e-05 0.82751 0.0054436 0.0061836 0.0014182 0.98653 0.99144 3.0621e-06 1.2249e-05 0.13327 0.86834 0.87649 0.0014138 0.95717 0.54054 0.0019041 0.42549 1.6642 1.6626 16.0095 144.9831 0.00022756 -85.5156 0.42336
1.5274 0.98803 5.5161e-05 3.8182 0.01203 2.0091e-05 0.0011544 0.17372 0.00065867 0.17437 0.15955 0 0.035529 0.0389 0 0.93122 0.26508 0.072521 0.010028 4.4252 0.062579 7.5534e-05 0.8275 0.0054441 0.0061842 0.0014179 0.98653 0.99144 3.0616e-06 1.2246e-05 0.13327 0.8687 0.87669 0.0014137 0.95743 0.5407 0.001904 0.4255 1.6651 1.6635 16.0095 144.9832 0.00022725 -85.5167 0.42436
1.5284 0.98803 5.5161e-05 3.8182 0.01203 2.0104e-05 0.0011544 0.17377 0.00065867 0.17442 0.15959 0 0.035526 0.0389 0 0.9313 0.26511 0.072535 0.01003 4.4257 0.06259 7.5547e-05 0.82749 0.0054446 0.0061847 0.0014177 0.98654 0.99144 3.061e-06 1.2244e-05 0.13328 0.86906 0.87689 0.0014136 0.95768 0.54085 0.0019038 0.42551 1.666 1.6644 16.0095 144.9832 0.00022693 -85.5177 0.42536
1.5294 0.98803 5.5161e-05 3.8182 0.01203 2.0117e-05 0.0011544 0.17382 0.00065868 0.17447 0.15964 0 0.035523 0.0389 0 0.93139 0.26515 0.072549 0.010031 4.4262 0.0626 7.5561e-05 0.82748 0.0054451 0.0061852 0.0014174 0.98654 0.99144 3.0604e-06 1.2242e-05 0.13328 0.86942 0.87709 0.0014135 0.95794 0.54101 0.0019036 0.42553 1.667 1.6654 16.0095 144.9832 0.00022662 -85.5188 0.42636
1.5304 0.98803 5.5161e-05 3.8182 0.01203 2.0131e-05 0.0011544 0.17386 0.00065868 0.17452 0.15968 0 0.03552 0.0389 0 0.93148 0.26519 0.072563 0.010033 4.4267 0.062611 7.5574e-05 0.82747 0.0054456 0.0061857 0.0014172 0.98654 0.99144 3.0599e-06 1.224e-05 0.13328 0.86977 0.87729 0.0014133 0.95819 0.54117 0.0019035 0.42554 1.6679 1.6663 16.0095 144.9832 0.00022631 -85.5198 0.42736
1.5314 0.98803 5.5161e-05 3.8182 0.012029 2.0144e-05 0.0011544 0.17391 0.00065868 0.17457 0.15973 0 0.035517 0.0389 0 0.93156 0.26523 0.072577 0.010035 4.4273 0.062621 7.5588e-05 0.82745 0.0054461 0.0061862 0.0014169 0.98655 0.99145 3.0593e-06 1.2237e-05 0.13329 0.87013 0.87749 0.0014132 0.95844 0.54133 0.0019033 0.42555 1.6688 1.6672 16.0095 144.9832 0.00022599 -85.5208 0.42836
1.5324 0.98803 5.5161e-05 3.8182 0.012029 2.0157e-05 0.0011544 0.17396 0.00065868 0.17462 0.15978 0 0.035514 0.0389 0 0.93165 0.26527 0.072591 0.010036 4.4278 0.062631 7.5601e-05 0.82744 0.0054466 0.0061867 0.0014167 0.98655 0.99145 3.0588e-06 1.2235e-05 0.13329 0.87048 0.87768 0.0014131 0.95869 0.54149 0.0019031 0.42556 1.6697 1.6682 16.0095 144.9833 0.00022568 -85.5218 0.42936
1.5334 0.98803 5.5161e-05 3.8182 0.012029 2.017e-05 0.0011544 0.17401 0.00065868 0.17467 0.15982 0 0.035511 0.0389 0 0.93173 0.26531 0.072605 0.010038 4.4283 0.062642 7.5614e-05 0.82743 0.0054471 0.0061872 0.0014165 0.98655 0.99145 3.0582e-06 1.2233e-05 0.1333 0.87084 0.87788 0.001413 0.95893 0.54165 0.001903 0.42558 1.6707 1.6691 16.0095 144.9833 0.00022537 -85.5228 0.43036
1.5344 0.98803 5.516e-05 3.8182 0.012029 2.0183e-05 0.0011544 0.17406 0.00065868 0.17472 0.15987 0 0.035508 0.0389 0 0.93182 0.26535 0.072619 0.01004 4.4288 0.062652 7.5628e-05 0.82742 0.0054476 0.0061877 0.0014162 0.98656 0.99145 3.0577e-06 1.2231e-05 0.1333 0.87119 0.87807 0.0014128 0.95918 0.54181 0.0019028 0.42559 1.6716 1.67 16.0095 144.9833 0.00022507 -85.5238 0.43136
1.5354 0.98803 5.516e-05 3.8182 0.012029 2.0196e-05 0.0011544 0.17411 0.00065868 0.17477 0.15992 0 0.035505 0.0389 0 0.93191 0.26538 0.072633 0.010041 4.4294 0.062662 7.5641e-05 0.82741 0.0054481 0.0061882 0.001416 0.98656 0.99145 3.0572e-06 1.2229e-05 0.1333 0.87154 0.87826 0.0014127 0.95942 0.54197 0.0019027 0.4256 1.6725 1.6709 16.0095 144.9833 0.00022476 -85.5248 0.43236
1.5364 0.98803 5.516e-05 3.8182 0.012029 2.0209e-05 0.0011544 0.17416 0.00065868 0.17481 0.15996 0 0.035502 0.0389 0 0.93199 0.26542 0.072647 0.010043 4.4299 0.062673 7.5655e-05 0.8274 0.0054486 0.0061887 0.0014158 0.98656 0.99146 3.0566e-06 1.2226e-05 0.13331 0.87189 0.87846 0.0014126 0.95967 0.54213 0.0019025 0.42561 1.6734 1.6719 16.0095 144.9833 0.00022445 -85.5258 0.43336
1.5374 0.98803 5.516e-05 3.8182 0.012029 2.0222e-05 0.0011544 0.17421 0.00065868 0.17486 0.16001 0 0.035499 0.0389 0 0.93208 0.26546 0.07266 0.010045 4.4304 0.062683 7.5668e-05 0.82739 0.0054491 0.0061892 0.0014155 0.98657 0.99146 3.0561e-06 1.2224e-05 0.13331 0.87224 0.87865 0.0014125 0.95991 0.54229 0.0019023 0.42563 1.6743 1.6728 16.0095 144.9834 0.00022415 -85.5268 0.43436
1.5384 0.98803 5.516e-05 3.8182 0.012029 2.0235e-05 0.0011544 0.17426 0.00065868 0.17491 0.16006 0 0.035496 0.0389 0 0.93217 0.2655 0.072674 0.010046 4.4309 0.062693 7.5682e-05 0.82738 0.0054496 0.0061897 0.0014153 0.98657 0.99146 3.0556e-06 1.2222e-05 0.13332 0.87258 0.87884 0.0014123 0.96015 0.54244 0.0019022 0.42564 1.6752 1.6737 16.0095 144.9834 0.00022385 -85.5277 0.43536
1.5394 0.98803 5.516e-05 3.8182 0.012029 2.0249e-05 0.0011544 0.17431 0.00065868 0.17496 0.1601 0 0.035494 0.0389 0 0.93225 0.26554 0.072688 0.010048 4.4315 0.062704 7.5695e-05 0.82737 0.0054501 0.0061903 0.0014151 0.98657 0.99146 3.0551e-06 1.222e-05 0.13332 0.87293 0.87903 0.0014122 0.96038 0.5426 0.001902 0.42565 1.6761 1.6746 16.0095 144.9834 0.00022354 -85.5287 0.43636
1.5404 0.98803 5.516e-05 3.8182 0.012029 2.0262e-05 0.0011544 0.17436 0.00065868 0.17501 0.16015 0 0.035491 0.0389 0 0.93234 0.26558 0.072702 0.01005 4.432 0.062714 7.5709e-05 0.82736 0.0054506 0.0061908 0.0014148 0.98657 0.99146 3.0545e-06 1.2218e-05 0.13332 0.87327 0.87922 0.0014121 0.96062 0.54276 0.0019019 0.42566 1.677 1.6755 16.0094 144.9834 0.00022324 -85.5297 0.43736
1.5414 0.98803 5.516e-05 3.8182 0.012029 2.0275e-05 0.0011544 0.17441 0.00065868 0.17506 0.16019 0 0.035488 0.0389 0 0.93243 0.26562 0.072716 0.010051 4.4325 0.062725 7.5722e-05 0.82735 0.0054511 0.0061913 0.0014146 0.98658 0.99147 3.054e-06 1.2216e-05 0.13333 0.87362 0.87941 0.001412 0.96086 0.54292 0.0019017 0.42568 1.6779 1.6764 16.0094 144.9834 0.00022294 -85.5306 0.43836
1.5424 0.98803 5.516e-05 3.8182 0.012029 2.0288e-05 0.0011544 0.17446 0.00065868 0.17511 0.16024 0 0.035485 0.0389 0 0.93251 0.26566 0.07273 0.010053 4.433 0.062735 7.5736e-05 0.82734 0.0054516 0.0061918 0.0014144 0.98658 0.99147 3.0535e-06 1.2214e-05 0.13333 0.87396 0.8796 0.0014119 0.96109 0.54308 0.0019016 0.42569 1.6788 1.6773 16.0094 144.9835 0.00022265 -85.5316 0.43936
1.5434 0.98803 5.516e-05 3.8182 0.012029 2.0301e-05 0.0011544 0.1745 0.00065868 0.17516 0.16029 0 0.035482 0.0389 0 0.9326 0.26569 0.072744 0.010055 4.4336 0.062745 7.5749e-05 0.82733 0.0054521 0.0061923 0.0014142 0.98658 0.99147 3.053e-06 1.2212e-05 0.13334 0.8743 0.87979 0.0014118 0.96132 0.54324 0.0019014 0.4257 1.6797 1.6782 16.0094 144.9835 0.00022235 -85.5325 0.44036
1.5444 0.98803 5.516e-05 3.8182 0.012029 2.0314e-05 0.0011544 0.17455 0.00065869 0.17521 0.16033 0 0.035479 0.0389 0 0.93269 0.26573 0.072758 0.010056 4.4341 0.062756 7.5763e-05 0.82732 0.0054526 0.0061928 0.001414 0.98659 0.99147 3.0525e-06 1.221e-05 0.13334 0.87464 0.87997 0.0014116 0.96155 0.5434 0.0019013 0.42572 1.6806 1.6791 16.0094 144.9835 0.00022205 -85.5334 0.44136
1.5454 0.98803 5.516e-05 3.8182 0.012029 2.0327e-05 0.0011544 0.1746 0.00065869 0.17526 0.16038 0 0.035476 0.0389 0 0.93277 0.26577 0.072772 0.010058 4.4346 0.062766 7.5776e-05 0.82731 0.0054531 0.0061933 0.0014137 0.98659 0.99147 3.052e-06 1.2208e-05 0.13335 0.87498 0.88016 0.0014115 0.96178 0.54355 0.0019011 0.42573 1.6815 1.68 16.0094 144.9835 0.00022176 -85.5344 0.44236
1.5464 0.98803 5.516e-05 3.8182 0.012029 2.034e-05 0.0011544 0.17465 0.00065869 0.1753 0.16042 0 0.035473 0.0389 0 0.93286 0.26581 0.072786 0.01006 4.4352 0.062777 7.579e-05 0.8273 0.0054536 0.0061938 0.0014135 0.98659 0.99148 3.0515e-06 1.2206e-05 0.13335 0.87532 0.88035 0.0014114 0.96201 0.54371 0.001901 0.42574 1.6824 1.6809 16.0094 144.9835 0.00022147 -85.5353 0.44336
1.5474 0.98803 5.516e-05 3.8182 0.012029 2.0354e-05 0.0011544 0.1747 0.00065869 0.17535 0.16047 0 0.03547 0.0389 0 0.93295 0.26585 0.0728 0.010061 4.4357 0.062787 7.5803e-05 0.82729 0.0054541 0.0061944 0.0014133 0.98659 0.99148 3.051e-06 1.2204e-05 0.13335 0.87566 0.88053 0.0014113 0.96223 0.54387 0.0019008 0.42575 1.6833 1.6818 16.0094 144.9836 0.00022117 -85.5362 0.44436
1.5484 0.98803 5.516e-05 3.8182 0.012029 2.0367e-05 0.0011544 0.17475 0.00065869 0.1754 0.16052 0 0.035467 0.0389 0 0.93303 0.26589 0.072814 0.010063 4.4362 0.062797 7.5817e-05 0.82728 0.0054546 0.0061949 0.0014131 0.9866 0.99148 3.0505e-06 1.2202e-05 0.13336 0.876 0.88071 0.0014112 0.96246 0.54403 0.0019007 0.42577 1.6842 1.6827 16.0094 144.9836 0.00022088 -85.5371 0.44536
1.5494 0.98803 5.5159e-05 3.8182 0.012029 2.038e-05 0.0011544 0.1748 0.00065869 0.17545 0.16056 0 0.035464 0.0389 0 0.93312 0.26593 0.072828 0.010065 4.4367 0.062808 7.583e-05 0.82727 0.0054551 0.0061954 0.0014129 0.9866 0.99148 3.05e-06 1.22e-05 0.13336 0.87633 0.8809 0.0014111 0.96268 0.54419 0.0019005 0.42578 1.6851 1.6836 16.0094 144.9836 0.00022059 -85.538 0.44636
1.5504 0.98803 5.5159e-05 3.8182 0.012029 2.0393e-05 0.0011544 0.17485 0.00065869 0.1755 0.16061 0 0.035462 0.0389 0 0.93321 0.26596 0.072842 0.010066 4.4373 0.062818 7.5844e-05 0.82726 0.0054556 0.0061959 0.0014127 0.9866 0.99148 3.0495e-06 1.2198e-05 0.13337 0.87667 0.88108 0.001411 0.9629 0.54434 0.0019004 0.42579 1.6859 1.6844 16.0094 144.9836 0.0002203 -85.5389 0.44736
1.5514 0.98803 5.5159e-05 3.8182 0.012029 2.0406e-05 0.0011544 0.17489 0.00065869 0.17555 0.16065 0 0.035459 0.0389 0 0.93329 0.266 0.072856 0.010068 4.4378 0.062829 7.5857e-05 0.82725 0.0054561 0.0061964 0.0014125 0.98661 0.99148 3.0491e-06 1.2196e-05 0.13337 0.877 0.88126 0.0014109 0.96313 0.5445 0.0019002 0.4258 1.6868 1.6853 16.0094 144.9836 0.00022002 -85.5398 0.44836
1.5524 0.98803 5.5159e-05 3.8182 0.012029 2.0419e-05 0.0011544 0.17494 0.00065869 0.1756 0.1607 0 0.035456 0.0389 0 0.93338 0.26604 0.07287 0.01007 4.4383 0.062839 7.5871e-05 0.82724 0.0054566 0.0061969 0.0014122 0.98661 0.99149 3.0486e-06 1.2194e-05 0.13337 0.87733 0.88144 0.0014107 0.96334 0.54466 0.0019001 0.42582 1.6877 1.6862 16.0094 144.9837 0.00021973 -85.5407 0.44936
1.5534 0.98803 5.5159e-05 3.8182 0.012029 2.0432e-05 0.0011544 0.17499 0.00065869 0.17565 0.16074 0 0.035453 0.0389 0 0.93347 0.26608 0.072884 0.010071 4.4389 0.062849 7.5884e-05 0.82723 0.0054571 0.0061974 0.001412 0.98661 0.99149 3.0481e-06 1.2192e-05 0.13338 0.87766 0.88162 0.0014106 0.96356 0.54482 0.0018999 0.42583 1.6886 1.6871 16.0093 144.9837 0.00021944 -85.5416 0.45036
1.5544 0.98803 5.5159e-05 3.8182 0.012029 2.0445e-05 0.0011544 0.17504 0.00065869 0.17569 0.16079 0 0.03545 0.0389 0 0.93355 0.26612 0.072898 0.010073 4.4394 0.06286 7.5898e-05 0.82722 0.0054576 0.006198 0.0014118 0.98661 0.99149 3.0476e-06 1.2191e-05 0.13338 0.87799 0.8818 0.0014105 0.96378 0.54498 0.0018998 0.42584 1.6894 1.688 16.0093 144.9837 0.00021916 -85.5424 0.45136
1.5554 0.98803 5.5159e-05 3.8182 0.012029 2.0459e-05 0.0011544 0.17509 0.00065869 0.17574 0.16084 0 0.035447 0.0389 0 0.93364 0.26616 0.072912 0.010075 4.4399 0.06287 7.5911e-05 0.82721 0.0054581 0.0061985 0.0014116 0.98662 0.99149 3.0472e-06 1.2189e-05 0.13339 0.87832 0.88198 0.0014104 0.96399 0.54513 0.0018997 0.42586 1.6903 1.6888 16.0093 144.9837 0.00021888 -85.5433 0.45236
1.5564 0.98803 5.5159e-05 3.8182 0.012029 2.0472e-05 0.0011544 0.17514 0.00065869 0.17579 0.16088 0 0.035444 0.0389 0 0.93373 0.2662 0.072926 0.010076 4.4405 0.062881 7.5925e-05 0.8272 0.0054586 0.006199 0.0014114 0.98662 0.99149 3.0467e-06 1.2187e-05 0.13339 0.87865 0.88216 0.0014103 0.96421 0.54529 0.0018995 0.42587 1.6912 1.6897 16.0093 144.9837 0.0002186 -85.5442 0.45336
1.5574 0.98803 5.5159e-05 3.8182 0.012029 2.0485e-05 0.0011544 0.17519 0.00065869 0.17584 0.16093 0 0.035441 0.0389 0 0.93381 0.26624 0.07294 0.010078 4.441 0.062891 7.5938e-05 0.82718 0.0054591 0.0061995 0.0014112 0.98662 0.99149 3.0463e-06 1.2185e-05 0.1334 0.87898 0.88234 0.0014102 0.96442 0.54545 0.0018994 0.42588 1.692 1.6906 16.0093 144.9838 0.00021831 -85.545 0.45436
1.5584 0.98803 5.5159e-05 3.8182 0.012029 2.0498e-05 0.0011544 0.17523 0.0006587 0.17589 0.16097 0 0.035438 0.0389 0 0.9339 0.26628 0.072954 0.01008 4.4415 0.062901 7.5952e-05 0.82717 0.0054596 0.0062 0.001411 0.98662 0.9915 3.0458e-06 1.2183e-05 0.1334 0.8793 0.88252 0.0014101 0.96463 0.54561 0.0018993 0.42589 1.6929 1.6914 16.0093 144.9838 0.00021803 -85.5459 0.45536
1.5594 0.98803 5.5159e-05 3.8182 0.012029 2.0511e-05 0.0011544 0.17528 0.0006587 0.17594 0.16102 0 0.035436 0.0389 0 0.93399 0.26631 0.072968 0.010081 4.4421 0.062912 7.5965e-05 0.82716 0.0054601 0.0062005 0.0014108 0.98663 0.9915 3.0453e-06 1.2181e-05 0.1334 0.87963 0.88269 0.00141 0.96484 0.54577 0.0018991 0.42591 1.6937 1.6923 16.0093 144.9838 0.00021776 -85.5467 0.45636
1.5604 0.98803 5.5159e-05 3.8182 0.012029 2.0524e-05 0.0011544 0.17533 0.0006587 0.17598 0.16106 0 0.035433 0.0389 0 0.93407 0.26635 0.072982 0.010083 4.4426 0.062922 7.5979e-05 0.82715 0.0054606 0.006201 0.0014106 0.98663 0.9915 3.0449e-06 1.218e-05 0.13341 0.87995 0.88287 0.0014099 0.96505 0.54592 0.001899 0.42592 1.6946 1.6932 16.0093 144.9838 0.00021748 -85.5475 0.45736
1.5614 0.98803 5.5159e-05 3.8182 0.012029 2.0537e-05 0.0011544 0.17538 0.0006587 0.17603 0.16111 0 0.03543 0.0389 0 0.93416 0.26639 0.072996 0.010085 4.4432 0.062933 7.5993e-05 0.82714 0.0054611 0.0062016 0.0014104 0.98663 0.9915 3.0444e-06 1.2178e-05 0.13341 0.88028 0.88304 0.0014098 0.96525 0.54608 0.0018989 0.42593 1.6955 1.694 16.0093 144.9838 0.0002172 -85.5484 0.45836
1.5624 0.98803 5.5159e-05 3.8182 0.012029 2.055e-05 0.0011544 0.17543 0.0006587 0.17608 0.16115 0 0.035427 0.0389 0 0.93425 0.26643 0.07301 0.010086 4.4437 0.062943 7.6006e-05 0.82713 0.0054616 0.0062021 0.0014102 0.98663 0.9915 3.044e-06 1.2176e-05 0.13342 0.8806 0.88322 0.0014097 0.96546 0.54624 0.0018987 0.42594 1.6963 1.6949 16.0093 144.9838 0.00021693 -85.5492 0.45936
1.5634 0.98803 5.5159e-05 3.8182 0.012029 2.0563e-05 0.0011544 0.17547 0.0006587 0.17613 0.1612 0 0.035424 0.0389 0 0.93433 0.26647 0.073024 0.010088 4.4442 0.062954 7.602e-05 0.82712 0.0054621 0.0062026 0.0014101 0.98664 0.9915 3.0436e-06 1.2174e-05 0.13342 0.88092 0.88339 0.0014096 0.96566 0.5464 0.0018986 0.42596 1.6972 1.6957 16.0092 144.9839 0.00021665 -85.55 0.46036
1.5644 0.98803 5.5159e-05 3.8182 0.012029 2.0577e-05 0.0011544 0.17552 0.0006587 0.17618 0.16124 0 0.035421 0.0389 0 0.93442 0.26651 0.073038 0.01009 4.4448 0.062964 7.6033e-05 0.82711 0.0054626 0.0062031 0.0014099 0.98664 0.99151 3.0431e-06 1.2172e-05 0.13342 0.88124 0.88356 0.0014095 0.96587 0.54655 0.0018985 0.42597 1.698 1.6966 16.0092 144.9839 0.00021638 -85.5508 0.46136
1.5654 0.98803 5.5158e-05 3.8182 0.012029 2.059e-05 0.0011544 0.17557 0.0006587 0.17623 0.16129 0 0.035418 0.0389 0 0.93451 0.26655 0.073052 0.010092 4.4453 0.062974 7.6047e-05 0.8271 0.0054631 0.0062036 0.0014097 0.98664 0.99151 3.0427e-06 1.2171e-05 0.13343 0.88156 0.88374 0.0014094 0.96607 0.54671 0.0018983 0.42598 1.6988 1.6974 16.0092 144.9839 0.00021611 -85.5516 0.46236
1.5664 0.98803 5.5158e-05 3.8182 0.012029 2.0603e-05 0.0011544 0.17562 0.0006587 0.17627 0.16133 0 0.035416 0.0389 0 0.9346 0.26659 0.073066 0.010093 4.4458 0.062985 7.606e-05 0.82709 0.0054637 0.0062042 0.0014095 0.98664 0.99151 3.0423e-06 1.2169e-05 0.13343 0.88188 0.88391 0.0014093 0.96627 0.54687 0.0018982 0.426 1.6997 1.6983 16.0092 144.9839 0.00021584 -85.5524 0.46336
1.5674 0.98803 5.5158e-05 3.8182 0.012029 2.0616e-05 0.0011544 0.17567 0.0006587 0.17632 0.16138 0 0.035413 0.0389 0 0.93468 0.26662 0.07308 0.010095 4.4464 0.062995 7.6074e-05 0.82708 0.0054642 0.0062047 0.0014093 0.98665 0.99151 3.0418e-06 1.2167e-05 0.13344 0.8822 0.88408 0.0014092 0.96647 0.54702 0.0018981 0.42601 1.7005 1.6991 16.0092 144.9839 0.00021557 -85.5532 0.46436
1.5684 0.98803 5.5158e-05 3.8182 0.012029 2.0629e-05 0.0011544 0.17572 0.0006587 0.17637 0.16142 0 0.03541 0.0389 0 0.93477 0.26666 0.073094 0.010097 4.4469 0.063006 7.6087e-05 0.82707 0.0054647 0.0062052 0.0014091 0.98665 0.99151 3.0414e-06 1.2166e-05 0.13344 0.88251 0.88425 0.0014091 0.96667 0.54718 0.0018979 0.42602 1.7014 1.7 16.0092 144.984 0.0002153 -85.554 0.46536
1.5694 0.98803 5.5158e-05 3.8182 0.012029 2.0642e-05 0.0011544 0.17576 0.0006587 0.17642 0.16147 0 0.035407 0.0389 0 0.93486 0.2667 0.073108 0.010098 4.4475 0.063016 7.6101e-05 0.82706 0.0054652 0.0062057 0.0014089 0.98665 0.99151 3.041e-06 1.2164e-05 0.13345 0.88283 0.88442 0.001409 0.96686 0.54734 0.0018978 0.42603 1.7022 1.7008 16.0092 144.984 0.00021503 -85.5548 0.46636
1.5704 0.98803 5.5158e-05 3.8182 0.012029 2.0655e-05 0.0011544 0.17581 0.0006587 0.17646 0.16152 0 0.035404 0.0389 0 0.93494 0.26674 0.073122 0.0101 4.448 0.063027 7.6115e-05 0.82705 0.0054657 0.0062062 0.0014087 0.98665 0.99152 3.0406e-06 1.2162e-05 0.13345 0.88314 0.88459 0.0014089 0.96706 0.5475 0.0018977 0.42605 1.703 1.7017 16.0092 144.984 0.00021476 -85.5556 0.46736
1.5714 0.98803 5.5158e-05 3.8182 0.012029 2.0668e-05 0.0011544 0.17586 0.0006587 0.17651 0.16156 0 0.035401 0.0389 0 0.93503 0.26678 0.073136 0.010102 4.4485 0.063037 7.6128e-05 0.82704 0.0054662 0.0062068 0.0014086 0.98666 0.99152 3.0401e-06 1.2161e-05 0.13345 0.88345 0.88475 0.0014088 0.96725 0.54765 0.0018976 0.42606 1.7039 1.7025 16.0092 144.984 0.0002145 -85.5564 0.46836
1.5724 0.98803 5.5158e-05 3.8182 0.012029 2.0682e-05 0.0011544 0.17591 0.0006587 0.17656 0.16161 0 0.035399 0.0389 0 0.93512 0.26682 0.07315 0.010103 4.4491 0.063047 7.6142e-05 0.82703 0.0054667 0.0062073 0.0014084 0.98666 0.99152 3.0397e-06 1.2159e-05 0.13346 0.88377 0.88492 0.0014087 0.96744 0.54781 0.0018974 0.42607 1.7047 1.7033 16.0092 144.984 0.00021423 -85.5571 0.46936
1.5734 0.98803 5.5158e-05 3.8182 0.012029 2.0695e-05 0.0011544 0.17595 0.00065871 0.17661 0.16165 0 0.035396 0.0389 0 0.9352 0.26686 0.073164 0.010105 4.4496 0.063058 7.6155e-05 0.82702 0.0054672 0.0062078 0.0014082 0.98666 0.99152 3.0393e-06 1.2157e-05 0.13346 0.88408 0.88509 0.0014086 0.96764 0.54797 0.0018973 0.42609 1.7055 1.7042 16.0091 144.9841 0.00021397 -85.5579 0.47036
1.5744 0.98803 5.5158e-05 3.8182 0.012029 2.0708e-05 0.0011544 0.176 0.00065871 0.17666 0.16169 0 0.035393 0.0389 0 0.93529 0.2669 0.073178 0.010107 4.4502 0.063068 7.6169e-05 0.82701 0.0054677 0.0062083 0.001408 0.98666 0.99152 3.0389e-06 1.2156e-05 0.13347 0.88439 0.88526 0.0014085 0.96783 0.54812 0.0018972 0.4261 1.7064 1.705 16.0091 144.9841 0.00021371 -85.5587 0.47136
1.5754 0.98803 5.5158e-05 3.8182 0.012029 2.0721e-05 0.0011544 0.17605 0.00065871 0.1767 0.16174 0 0.03539 0.0389 0 0.93538 0.26694 0.073192 0.010108 4.4507 0.063079 7.6182e-05 0.827 0.0054682 0.0062088 0.0014078 0.98667 0.99152 3.0385e-06 1.2154e-05 0.13347 0.8847 0.88542 0.0014084 0.96802 0.54828 0.0018971 0.42611 1.7072 1.7058 16.0091 144.9841 0.00021345 -85.5594 0.47236
1.5764 0.98803 5.5158e-05 3.8182 0.012029 2.0734e-05 0.0011544 0.1761 0.00065871 0.17675 0.16178 0 0.035387 0.0389 0 0.93547 0.26698 0.073206 0.01011 4.4513 0.063089 7.6196e-05 0.82699 0.0054687 0.0062094 0.0014077 0.98667 0.99152 3.0381e-06 1.2152e-05 0.13348 0.88501 0.88559 0.0014083 0.9682 0.54844 0.0018969 0.42612 1.708 1.7066 16.0091 144.9841 0.00021319 -85.5602 0.47336
1.5774 0.98803 5.5158e-05 3.8182 0.012029 2.0747e-05 0.0011544 0.17615 0.00065871 0.1768 0.16183 0 0.035384 0.0389 0 0.93555 0.26701 0.07322 0.010112 4.4518 0.0631 7.621e-05 0.82698 0.0054692 0.0062099 0.0014075 0.98667 0.99153 3.0377e-06 1.2151e-05 0.13348 0.88531 0.88575 0.0014083 0.96839 0.54859 0.0018968 0.42614 1.7088 1.7075 16.0091 144.9841 0.00021293 -85.5609 0.47436
1.5784 0.98803 5.5158e-05 3.8182 0.012029 2.076e-05 0.0011544 0.17619 0.00065871 0.17685 0.16187 0 0.035382 0.0389 0 0.93564 0.26705 0.073234 0.010113 4.4523 0.06311 7.6223e-05 0.82697 0.0054698 0.0062104 0.0014073 0.98667 0.99153 3.0373e-06 1.2149e-05 0.13348 0.88562 0.88591 0.0014082 0.96858 0.54875 0.0018967 0.42615 1.7096 1.7083 16.0091 144.9842 0.00021267 -85.5616 0.47536
1.5794 0.98803 5.5158e-05 3.8182 0.012029 2.0773e-05 0.0011544 0.17624 0.00065871 0.17689 0.16192 0 0.035379 0.0389 0 0.93573 0.26709 0.073248 0.010115 4.4529 0.063121 7.6237e-05 0.82696 0.0054703 0.0062109 0.0014071 0.98667 0.99153 3.0369e-06 1.2148e-05 0.13349 0.88593 0.88608 0.0014081 0.96876 0.54891 0.0018966 0.42616 1.7105 1.7091 16.0091 144.9842 0.00021241 -85.5624 0.47636
1.5804 0.98803 5.5158e-05 3.8182 0.012029 2.0786e-05 0.0011544 0.17629 0.00065871 0.17694 0.16196 0 0.035376 0.0389 0 0.93582 0.26713 0.073262 0.010117 4.4534 0.063131 7.625e-05 0.82695 0.0054708 0.0062115 0.001407 0.98668 0.99153 3.0365e-06 1.2146e-05 0.13349 0.88623 0.88624 0.001408 0.96894 0.54906 0.0018965 0.42618 1.7113 1.7099 16.0091 144.9842 0.00021215 -85.5631 0.47736
1.5814 0.98803 5.5157e-05 3.8182 0.012029 2.08e-05 0.0011544 0.17634 0.00065871 0.17699 0.16201 0 0.035373 0.0389 0 0.9359 0.26717 0.073276 0.010118 4.454 0.063142 7.6264e-05 0.82693 0.0054713 0.006212 0.0014068 0.98668 0.99153 3.0361e-06 1.2144e-05 0.1335 0.88653 0.8864 0.0014079 0.96913 0.54922 0.0018964 0.42619 1.7121 1.7107 16.0091 144.9842 0.0002119 -85.5638 0.47836
1.5824 0.98803 5.5157e-05 3.8182 0.012029 2.0813e-05 0.0011544 0.17638 0.00065871 0.17704 0.16205 0 0.03537 0.0389 0 0.93599 0.26721 0.07329 0.01012 4.4545 0.063152 7.6278e-05 0.82692 0.0054718 0.0062125 0.0014066 0.98668 0.99153 3.0357e-06 1.2143e-05 0.1335 0.88684 0.88656 0.0014078 0.96931 0.54938 0.0018962 0.4262 1.7129 1.7115 16.009 144.9842 0.00021164 -85.5646 0.47936
1.5834 0.98803 5.5157e-05 3.8182 0.012029 2.0826e-05 0.0011544 0.17643 0.00065871 0.17708 0.1621 0 0.035368 0.0389 0 0.93608 0.26725 0.073304 0.010122 4.4551 0.063162 7.6291e-05 0.82691 0.0054723 0.006213 0.0014065 0.98668 0.99153 3.0354e-06 1.2141e-05 0.1335 0.88714 0.88672 0.0014077 0.96949 0.54953 0.0018961 0.42621 1.7137 1.7124 16.009 144.9843 0.00021139 -85.5653 0.48036
1.5844 0.98803 5.5157e-05 3.8182 0.012029 2.0839e-05 0.0011544 0.17648 0.00065871 0.17713 0.16214 0 0.035365 0.0389 0 0.93616 0.26729 0.073318 0.010123 4.4556 0.063173 7.6305e-05 0.8269 0.0054728 0.0062136 0.0014063 0.98669 0.99154 3.035e-06 1.214e-05 0.13351 0.88744 0.88688 0.0014076 0.96967 0.54969 0.001896 0.42623 1.7145 1.7132 16.009 144.9843 0.00021114 -85.566 0.48136
1.5854 0.98803 5.5157e-05 3.8182 0.012029 2.0852e-05 0.0011544 0.17652 0.00065871 0.17718 0.16219 0 0.035362 0.0389 0 0.93625 0.26733 0.073332 0.010125 4.4562 0.063183 7.6318e-05 0.82689 0.0054733 0.0062141 0.0014061 0.98669 0.99154 3.0346e-06 1.2138e-05 0.13351 0.88774 0.88704 0.0014075 0.96984 0.54985 0.0018959 0.42624 1.7153 1.714 16.009 144.9843 0.00021089 -85.5667 0.48236
1.5864 0.98803 5.5157e-05 3.8182 0.012029 2.0865e-05 0.0011544 0.17657 0.00065871 0.17723 0.16223 0 0.035359 0.0389 0 0.93634 0.26737 0.073346 0.010127 4.4567 0.063194 7.6332e-05 0.82688 0.0054739 0.0062146 0.001406 0.98669 0.99154 3.0342e-06 1.2137e-05 0.13352 0.88804 0.8872 0.0014075 0.97002 0.55 0.0018958 0.42625 1.7161 1.7148 16.009 144.9843 0.00021064 -85.5674 0.48336
1.5874 0.98803 5.5157e-05 3.8182 0.012029 2.0878e-05 0.0011544 0.17662 0.00065871 0.17727 0.16228 0 0.035356 0.0389 0 0.93643 0.2674 0.073361 0.010129 4.4573 0.063204 7.6346e-05 0.82687 0.0054744 0.0062151 0.0014058 0.98669 0.99154 3.0338e-06 1.2135e-05 0.13352 0.88834 0.88736 0.0014074 0.97019 0.55016 0.0018957 0.42627 1.7169 1.7156 16.009 144.9843 0.00021039 -85.5681 0.48436
1.5884 0.98803 5.5157e-05 3.8182 0.012029 2.0891e-05 0.0011544 0.17667 0.00065872 0.17732 0.16232 0 0.035354 0.0389 0 0.93651 0.26744 0.073375 0.01013 4.4578 0.063215 7.6359e-05 0.82686 0.0054749 0.0062157 0.0014056 0.98669 0.99154 3.0335e-06 1.2134e-05 0.13353 0.88863 0.88752 0.0014073 0.97037 0.55031 0.0018956 0.42628 1.7177 1.7164 16.009 144.9844 0.00021014 -85.5688 0.48536
1.5894 0.98803 5.5157e-05 3.8182 0.012029 2.0905e-05 0.0011544 0.17671 0.00065872 0.17737 0.16236 0 0.035351 0.0389 0 0.9366 0.26748 0.073389 0.010132 4.4584 0.063225 7.6373e-05 0.82685 0.0054754 0.0062162 0.0014055 0.9867 0.99154 3.0331e-06 1.2132e-05 0.13353 0.88893 0.88768 0.0014072 0.97054 0.55047 0.0018955 0.42629 1.7185 1.7172 16.009 144.9844 0.00020989 -85.5695 0.48636
1.5904 0.98803 5.5157e-05 3.8182 0.012029 2.0918e-05 0.0011544 0.17676 0.00065872 0.17741 0.16241 0 0.035348 0.0389 0 0.93669 0.26752 0.073403 0.010134 4.4589 0.063236 7.6386e-05 0.82684 0.0054759 0.0062167 0.0014053 0.9867 0.99154 3.0327e-06 1.2131e-05 0.13353 0.88922 0.88783 0.0014071 0.97071 0.55063 0.0018953 0.4263 1.7193 1.718 16.0089 144.9844 0.00020964 -85.5701 0.48736
1.5914 0.98803 5.5157e-05 3.8182 0.012029 2.0931e-05 0.0011544 0.17681 0.00065872 0.17746 0.16245 0 0.035345 0.0389 0 0.93678 0.26756 0.073417 0.010135 4.4595 0.063246 7.64e-05 0.82683 0.0054764 0.0062172 0.0014052 0.9867 0.99155 3.0324e-06 1.2129e-05 0.13354 0.88952 0.88799 0.001407 0.97088 0.55078 0.0018952 0.42632 1.7201 1.7188 16.0089 144.9844 0.0002094 -85.5708 0.48836
1.5924 0.98803 5.5157e-05 3.8182 0.012029 2.0944e-05 0.0011544 0.17685 0.00065872 0.17751 0.1625 0 0.035342 0.0389 0 0.93686 0.2676 0.073431 0.010137 4.46 0.063257 7.6414e-05 0.82682 0.0054769 0.0062178 0.001405 0.9867 0.99155 3.032e-06 1.2128e-05 0.13354 0.88981 0.88814 0.0014069 0.97105 0.55094 0.0018951 0.42633 1.7209 1.7196 16.0089 144.9844 0.00020915 -85.5715 0.48936
1.5934 0.98803 5.5157e-05 3.8182 0.012029 2.0957e-05 0.0011544 0.1769 0.00065872 0.17756 0.16254 0 0.03534 0.0389 0 0.93695 0.26764 0.073445 0.010139 4.4606 0.063267 7.6427e-05 0.82681 0.0054775 0.0062183 0.0014049 0.9867 0.99155 3.0317e-06 1.2127e-05 0.13355 0.8901 0.8883 0.0014069 0.97122 0.55109 0.001895 0.42634 1.7217 1.7204 16.0089 144.9845 0.00020891 -85.5722 0.49036
1.5944 0.98803 5.5157e-05 3.8182 0.012029 2.097e-05 0.0011544 0.17695 0.00065872 0.1776 0.16259 0 0.035337 0.0389 0 0.93704 0.26768 0.073459 0.01014 4.4611 0.063278 7.6441e-05 0.8268 0.005478 0.0062188 0.0014047 0.98671 0.99155 3.0313e-06 1.2125e-05 0.13355 0.8904 0.88845 0.0014068 0.97139 0.55125 0.0018949 0.42636 1.7224 1.7211 16.0089 144.9845 0.00020867 -85.5728 0.49136
1.5954 0.98803 5.5157e-05 3.8182 0.012029 2.0983e-05 0.0011544 0.177 0.00065872 0.17765 0.16263 0 0.035334 0.0389 0 0.93713 0.26772 0.073473 0.010142 4.4617 0.063288 7.6455e-05 0.82679 0.0054785 0.0062194 0.0014045 0.98671 0.99155 3.031e-06 1.2124e-05 0.13356 0.89069 0.8886 0.0014067 0.97156 0.55141 0.0018948 0.42637 1.7232 1.7219 16.0089 144.9845 0.00020843 -85.5735 0.49236
1.5964 0.98803 5.5156e-05 3.8182 0.012029 2.0996e-05 0.0011544 0.17704 0.00065872 0.1777 0.16267 0 0.035331 0.0389 0 0.93721 0.26776 0.073487 0.010144 4.4622 0.063299 7.6468e-05 0.82678 0.005479 0.0062199 0.0014044 0.98671 0.99155 3.0306e-06 1.2122e-05 0.13356 0.89098 0.88876 0.0014066 0.97172 0.55156 0.0018947 0.42638 1.724 1.7227 16.0089 144.9845 0.00020818 -85.5741 0.49336
1.5974 0.98803 5.5156e-05 3.8182 0.012029 2.1009e-05 0.0011544 0.17709 0.00065872 0.17774 0.16272 0 0.035329 0.0389 0 0.9373 0.2678 0.073501 0.010145 4.4628 0.063309 7.6482e-05 0.82677 0.0054795 0.0062204 0.0014042 0.98671 0.99155 3.0303e-06 1.2121e-05 0.13356 0.89127 0.88891 0.0014065 0.97189 0.55172 0.0018946 0.42639 1.7248 1.7235 16.0089 144.9845 0.00020794 -85.5748 0.49436
1.5984 0.98803 5.5156e-05 3.8182 0.012029 2.1023e-05 0.0011544 0.17714 0.00065872 0.17779 0.16276 0 0.035326 0.0389 0 0.93739 0.26783 0.073516 0.010147 4.4633 0.06332 7.6496e-05 0.82676 0.00548 0.0062209 0.0014041 0.98671 0.99155 3.0299e-06 1.212e-05 0.13357 0.89155 0.88906 0.0014065 0.97205 0.55187 0.0018945 0.42641 1.7256 1.7243 16.0088 144.9846 0.00020771 -85.5754 0.49536
1.5994 0.98803 5.5156e-05 3.8182 0.012029 2.1036e-05 0.0011544 0.17718 0.00065872 0.17784 0.16281 0 0.035323 0.0389 0 0.93748 0.26787 0.07353 0.010149 4.4639 0.06333 7.6509e-05 0.82675 0.0054806 0.0062215 0.0014039 0.98672 0.99156 3.0296e-06 1.2118e-05 0.13357 0.89184 0.88921 0.0014064 0.97221 0.55203 0.0018944 0.42642 1.7263 1.7251 16.0088 144.9846 0.00020747 -85.5761 0.49636
1.6004 0.98803 5.5156e-05 3.8182 0.012029 2.1049e-05 0.0011544 0.17723 0.00065872 0.17788 0.16285 0 0.03532 0.0389 0 0.93756 0.26791 0.073544 0.01015 4.4644 0.063341 7.6523e-05 0.82674 0.0054811 0.006222 0.0014038 0.98672 0.99156 3.0292e-06 1.2117e-05 0.13358 0.89213 0.88936 0.0014063 0.97237 0.55218 0.0018943 0.42643 1.7271 1.7258 16.0088 144.9846 0.00020723 -85.5767 0.49736
1.6014 0.98803 5.5156e-05 3.8182 0.012029 2.1062e-05 0.0011544 0.17728 0.00065872 0.17793 0.16289 0 0.035317 0.0389 0 0.93765 0.26795 0.073558 0.010152 4.465 0.063351 7.6536e-05 0.82673 0.0054816 0.0062225 0.0014036 0.98672 0.99156 3.0289e-06 1.2115e-05 0.13358 0.89241 0.88951 0.0014062 0.97253 0.55234 0.0018942 0.42645 1.7279 1.7266 16.0088 144.9846 0.00020699 -85.5773 0.49836
1.6024 0.98803 5.5156e-05 3.8182 0.012029 2.1075e-05 0.0011544 0.17732 0.00065872 0.17798 0.16294 0 0.035315 0.0389 0 0.93774 0.26799 0.073572 0.010154 4.4655 0.063362 7.655e-05 0.82671 0.0054821 0.0062231 0.0014035 0.98672 0.99156 3.0285e-06 1.2114e-05 0.13359 0.8927 0.88966 0.0014062 0.97269 0.5525 0.0018941 0.42646 1.7286 1.7274 16.0088 144.9846 0.00020676 -85.578 0.49936
1.6034 0.98803 5.5156e-05 3.8182 0.012029 2.1088e-05 0.0011544 0.17737 0.00065872 0.17802 0.16298 0 0.035312 0.0389 0 0.93783 0.26803 0.073586 0.010155 4.4661 0.063372 7.6564e-05 0.8267 0.0054826 0.0062236 0.0014033 0.98672 0.99156 3.0282e-06 1.2113e-05 0.13359 0.89298 0.88981 0.0014061 0.97285 0.55265 0.001894 0.42647 1.7294 1.7282 16.0088 144.9847 0.00020652 -85.5786 0.50036
1.6044 0.98803 5.5156e-05 3.8182 0.012028 2.1101e-05 0.0011544 0.17742 0.00065873 0.17807 0.16303 0 0.035309 0.0389 0 0.93791 0.26807 0.0736 0.010157 4.4666 0.063383 7.6577e-05 0.82669 0.0054831 0.0062241 0.0014032 0.98673 0.99156 3.0279e-06 1.2111e-05 0.13359 0.89326 0.88996 0.001406 0.97301 0.55281 0.0018939 0.42648 1.7302 1.7289 16.0088 144.9847 0.00020629 -85.5792 0.50136
1.6054 0.98803 5.5156e-05 3.8182 0.012028 2.1114e-05 0.0011544 0.17746 0.00065873 0.17812 0.16307 0 0.035306 0.0389 0 0.938 0.26811 0.073614 0.010159 4.4672 0.063393 7.6591e-05 0.82668 0.0054837 0.0062247 0.0014031 0.98673 0.99156 3.0276e-06 1.211e-05 0.1336 0.89354 0.89011 0.0014059 0.97316 0.55296 0.0018938 0.4265 1.7309 1.7297 16.0087 144.9847 0.00020606 -85.5798 0.50236
1.6064 0.98803 5.5156e-05 3.8182 0.012028 2.1128e-05 0.0011544 0.17751 0.00065873 0.17816 0.16311 0 0.035304 0.0389 0 0.93809 0.26815 0.073629 0.010161 4.4678 0.063404 7.6605e-05 0.82667 0.0054842 0.0062252 0.0014029 0.98673 0.99156 3.0272e-06 1.2109e-05 0.1336 0.89383 0.89025 0.0014058 0.97332 0.55312 0.0018937 0.42651 1.7317 1.7305 16.0087 144.9847 0.00020583 -85.5804 0.50336
1.6074 0.98803 5.5156e-05 3.8182 0.012028 2.1141e-05 0.0011544 0.17756 0.00065873 0.17821 0.16316 0 0.035301 0.0389 0 0.93818 0.26819 0.073643 0.010162 4.4683 0.063414 7.6618e-05 0.82666 0.0054847 0.0062257 0.0014028 0.98673 0.99157 3.0269e-06 1.2108e-05 0.13361 0.89411 0.8904 0.0014058 0.97347 0.55327 0.0018936 0.42652 1.7325 1.7312 16.0087 144.9847 0.0002056 -85.581 0.50436
1.6084 0.98803 5.5156e-05 3.8182 0.012028 2.1154e-05 0.0011544 0.1776 0.00065873 0.17826 0.1632 0 0.035298 0.0389 0 0.93827 0.26823 0.073657 0.010164 4.4689 0.063425 7.6632e-05 0.82665 0.0054852 0.0062262 0.0014026 0.98673 0.99157 3.0266e-06 1.2106e-05 0.13361 0.89438 0.89055 0.0014057 0.97363 0.55343 0.0018935 0.42654 1.7332 1.732 16.0087 144.9848 0.00020537 -85.5816 0.50536
1.6094 0.98803 5.5156e-05 3.8182 0.012028 2.1167e-05 0.0011544 0.17765 0.00065873 0.1783 0.16324 0 0.035296 0.0389 0 0.93835 0.26827 0.073671 0.010166 4.4694 0.063435 7.6646e-05 0.82664 0.0054857 0.0062268 0.0014025 0.98673 0.99157 3.0263e-06 1.2105e-05 0.13362 0.89466 0.89069 0.0014056 0.97378 0.55358 0.0018934 0.42655 1.734 1.7327 16.0087 144.9848 0.00020514 -85.5822 0.50636
1.6104 0.98803 5.5156e-05 3.8182 0.012028 2.118e-05 0.0011544 0.1777 0.00065873 0.17835 0.16329 0 0.035293 0.0389 0 0.93844 0.26831 0.073685 0.010167 4.47 0.063446 7.6659e-05 0.82663 0.0054863 0.0062273 0.0014024 0.98674 0.99157 3.0259e-06 1.2104e-05 0.13362 0.89494 0.89084 0.0014056 0.97393 0.55374 0.0018933 0.42656 1.7347 1.7335 16.0087 144.9848 0.00020491 -85.5828 0.50736
1.6114 0.98803 5.5156e-05 3.8182 0.012028 2.1193e-05 0.0011544 0.17774 0.00065873 0.1784 0.16333 0 0.03529 0.0389 0 0.93853 0.26834 0.073699 0.010169 4.4705 0.063456 7.6673e-05 0.82662 0.0054868 0.0062278 0.0014022 0.98674 0.99157 3.0256e-06 1.2102e-05 0.13362 0.89522 0.89098 0.0014055 0.97408 0.55389 0.0018932 0.42657 1.7355 1.7342 16.0087 144.9848 0.00020468 -85.5834 0.50836
1.6124 0.98803 5.5155e-05 3.8182 0.012028 2.1206e-05 0.0011544 0.17779 0.00065873 0.17844 0.16338 0 0.035287 0.0389 0 0.93862 0.26838 0.073713 0.010171 4.4711 0.063467 7.6687e-05 0.82661 0.0054873 0.0062284 0.0014021 0.98674 0.99157 3.0253e-06 1.2101e-05 0.13363 0.89549 0.89113 0.0014054 0.97423 0.55405 0.0018931 0.42659 1.7362 1.735 16.0086 144.9848 0.00020445 -85.584 0.50936
1.6134 0.98803 5.5155e-05 3.8182 0.012028 2.1219e-05 0.0011544 0.17783 0.00065873 0.17849 0.16342 0 0.035285 0.0389 0 0.9387 0.26842 0.073728 0.010172 4.4717 0.063477 7.6701e-05 0.8266 0.0054878 0.0062289 0.0014019 0.98674 0.99157 3.025e-06 1.21e-05 0.13363 0.89577 0.89127 0.0014053 0.97438 0.5542 0.001893 0.4266 1.737 1.7357 16.0086 144.9849 0.00020423 -85.5846 0.51036
1.6144 0.98803 5.5155e-05 3.8182 0.012028 2.1232e-05 0.0011544 0.17788 0.00065873 0.17853 0.16346 0 0.035282 0.0389 0 0.93879 0.26846 0.073742 0.010174 4.4722 0.063488 7.6714e-05 0.82659 0.0054883 0.0062294 0.0014018 0.98674 0.99157 3.0247e-06 1.2099e-05 0.13364 0.89604 0.89141 0.0014053 0.97453 0.55436 0.0018929 0.42661 1.7377 1.7365 16.0086 144.9849 0.000204 -85.5852 0.51136
1.6154 0.98803 5.5155e-05 3.8182 0.012028 2.1246e-05 0.0011544 0.17793 0.00065873 0.17858 0.16351 0 0.035279 0.0389 0 0.93888 0.2685 0.073756 0.010176 4.4728 0.063498 7.6728e-05 0.82658 0.0054889 0.00623 0.0014017 0.98674 0.99158 3.0244e-06 1.2097e-05 0.13364 0.89631 0.89155 0.0014052 0.97467 0.55451 0.0018928 0.42663 1.7385 1.7372 16.0086 144.9849 0.00020378 -85.5857 0.51236
1.6164 0.98803 5.5155e-05 3.8182 0.012028 2.1259e-05 0.0011544 0.17797 0.00065873 0.17863 0.16355 0 0.035276 0.0389 0 0.93897 0.26854 0.07377 0.010177 4.4733 0.063509 7.6741e-05 0.82657 0.0054894 0.0062305 0.0014015 0.98675 0.99158 3.0241e-06 1.2096e-05 0.13365 0.89659 0.8917 0.0014051 0.97482 0.55467 0.0018927 0.42664 1.7392 1.738 16.0086 144.9849 0.00020356 -85.5863 0.51336
1.6174 0.98803 5.5155e-05 3.8182 0.012028 2.1272e-05 0.0011544 0.17802 0.00065873 0.17867 0.16359 0 0.035274 0.0389 0 0.93906 0.26858 0.073784 0.010179 4.4739 0.063519 7.6756e-05 0.82656 0.0054899 0.0062311 0.0014014 0.98675 0.99158 3.0238e-06 1.2095e-05 0.13365 0.89686 0.89184 0.0014051 0.97496 0.55482 0.0018926 0.42665 1.7399 1.7387 16.0086 144.9849 0.00020333 -85.5869 0.51436
1.6184 0.98803 5.5155e-05 3.8182 0.012028 2.1285e-05 0.0011544 0.17806 0.00065873 0.17872 0.16364 0 0.035271 0.0389 0 0.93914 0.26862 0.073798 0.010181 4.4745 0.06353 7.6769e-05 0.82655 0.0054904 0.0062316 0.0014013 0.98675 0.99158 3.0235e-06 1.2094e-05 0.13365 0.89713 0.89198 0.001405 0.97511 0.55498 0.0018926 0.42666 1.7407 1.7395 16.0086 144.985 0.00020311 -85.5874 0.51536
1.6194 0.98803 5.5155e-05 3.8182 0.012028 2.1298e-05 0.0011544 0.17811 0.00065873 0.17877 0.16368 0 0.035268 0.0389 0 0.93923 0.26866 0.073813 0.010183 4.475 0.06354 7.6782e-05 0.82654 0.005491 0.0062321 0.0014011 0.98675 0.99158 3.0232e-06 1.2093e-05 0.13366 0.8974 0.89212 0.0014049 0.97525 0.55513 0.0018925 0.42668 1.7414 1.7402 16.0085 144.985 0.00020289 -85.588 0.51636
1.6204 0.98803 5.5155e-05 3.8182 0.012028 2.1311e-05 0.0011544 0.17816 0.00065874 0.17881 0.16372 0 0.035266 0.0389 0 0.93932 0.2687 0.073827 0.010184 4.4756 0.063551 7.6796e-05 0.82653 0.0054915 0.0062327 0.001401 0.98675 0.99158 3.0229e-06 1.2091e-05 0.13366 0.89767 0.89226 0.0014048 0.97539 0.55529 0.0018924 0.42669 1.7422 1.741 16.0085 144.985 0.00020267 -85.5886 0.51736
1.6214 0.98803 5.5155e-05 3.8182 0.012028 2.1324e-05 0.0011544 0.1782 0.00065874 0.17886 0.16377 0 0.035263 0.0389 0 0.93941 0.26874 0.073841 0.010186 4.4762 0.063562 7.681e-05 0.82652 0.005492 0.0062332 0.0014009 0.98676 0.99158 3.0226e-06 1.209e-05 0.13367 0.89794 0.8924 0.0014048 0.97553 0.55544 0.0018923 0.4267 1.7429 1.7417 16.0085 144.985 0.00020245 -85.5891 0.51836
1.6224 0.98803 5.5155e-05 3.8182 0.012028 2.1337e-05 0.0011544 0.17825 0.00065874 0.1789 0.16381 0 0.03526 0.0389 0 0.9395 0.26878 0.073855 0.010188 4.4767 0.063572 7.6824e-05 0.8265 0.0054925 0.0062337 0.0014008 0.98676 0.99158 3.0223e-06 1.2089e-05 0.13367 0.8982 0.89253 0.0014047 0.97567 0.55559 0.0018922 0.42672 1.7436 1.7424 16.0085 144.985 0.00020224 -85.5897 0.51936
1.6234 0.98803 5.5155e-05 3.8182 0.012028 2.1351e-05 0.0011544 0.17829 0.00065874 0.17895 0.16385 0 0.035257 0.0389 0 0.93958 0.26882 0.073869 0.010189 4.4773 0.063583 7.6837e-05 0.82649 0.005493 0.0062343 0.0014006 0.98676 0.99158 3.022e-06 1.2088e-05 0.13368 0.89847 0.89267 0.0014046 0.97581 0.55575 0.0018921 0.42673 1.7443 1.7432 16.0085 144.9851 0.00020202 -85.5902 0.52036
1.6244 0.98803 5.5155e-05 3.8182 0.012028 2.1364e-05 0.0011544 0.17834 0.00065874 0.17899 0.1639 0 0.035255 0.0389 0 0.93967 0.26886 0.073884 0.010191 4.4779 0.063593 7.6852e-05 0.82648 0.0054936 0.0062348 0.0014005 0.98676 0.99158 3.0217e-06 1.2087e-05 0.13368 0.89873 0.89281 0.0014046 0.97595 0.5559 0.001892 0.42674 1.7451 1.7439 16.0085 144.9851 0.0002018 -85.5908 0.52136
1.6254 0.98803 5.5155e-05 3.8182 0.012028 2.1377e-05 0.0011544 0.17839 0.00065874 0.17904 0.16394 0 0.035252 0.0389 0 0.93976 0.2689 0.073898 0.010193 4.4784 0.063604 7.6865e-05 0.82647 0.0054941 0.0062353 0.0014004 0.98676 0.99159 3.0214e-06 1.2086e-05 0.13368 0.899 0.89295 0.0014045 0.97609 0.55606 0.0018919 0.42675 1.7458 1.7446 16.0085 144.9851 0.00020159 -85.5913 0.52236
1.6264 0.98803 5.5155e-05 3.8182 0.012028 2.139e-05 0.0011544 0.17843 0.00065874 0.17909 0.16398 0 0.035249 0.0389 0 0.93985 0.26894 0.073912 0.010194 4.479 0.063614 7.6878e-05 0.82646 0.0054946 0.0062359 0.0014002 0.98676 0.99159 3.0211e-06 1.2084e-05 0.13369 0.89926 0.89308 0.0014044 0.97622 0.55621 0.0018919 0.42677 1.7465 1.7453 16.0084 144.9851 0.00020137 -85.5918 0.52336
1.6274 0.98803 5.5155e-05 3.8182 0.012028 2.1403e-05 0.0011544 0.17848 0.00065874 0.17913 0.16402 0 0.035247 0.0389 0 0.93994 0.26897 0.073926 0.010196 4.4796 0.063625 7.6892e-05 0.82645 0.0054951 0.0062364 0.0014001 0.98676 0.99159 3.0208e-06 1.2083e-05 0.13369 0.89953 0.89322 0.0014044 0.97636 0.55637 0.0018918 0.42678 1.7472 1.7461 16.0084 144.9851 0.00020116 -85.5924 0.52436
1.6284 0.98803 5.5154e-05 3.8182 0.012028 2.1416e-05 0.0011544 0.17852 0.00065874 0.17918 0.16407 0 0.035244 0.0389 0 0.94002 0.26901 0.07394 0.010198 4.4801 0.063635 7.6906e-05 0.82644 0.0054957 0.006237 0.0014 0.98677 0.99159 3.0206e-06 1.2082e-05 0.1337 0.89979 0.89335 0.0014043 0.97649 0.55652 0.0018917 0.42679 1.748 1.7468 16.0084 144.9852 0.00020095 -85.5929 0.52536
1.6294 0.98803 5.5154e-05 3.8182 0.012028 2.1429e-05 0.0011544 0.17857 0.00065874 0.17922 0.16411 0 0.035241 0.0389 0 0.94011 0.26905 0.073955 0.010199 4.4807 0.063646 7.692e-05 0.82643 0.0054962 0.0062375 0.0013999 0.98677 0.99159 3.0203e-06 1.2081e-05 0.1337 0.90005 0.89349 0.0014043 0.97663 0.55667 0.0018916 0.42681 1.7487 1.7475 16.0084 144.9852 0.00020073 -85.5934 0.52636
1.6304 0.98803 5.5154e-05 3.8182 0.012028 2.1442e-05 0.0011544 0.17862 0.00065874 0.17927 0.16415 0 0.035239 0.0389 0 0.9402 0.26909 0.073969 0.010201 4.4813 0.063656 7.6934e-05 0.82642 0.0054967 0.006238 0.0013998 0.98677 0.99159 3.02e-06 1.208e-05 0.13371 0.90031 0.89362 0.0014042 0.97676 0.55683 0.0018915 0.42682 1.7494 1.7482 16.0084 144.9852 0.00020052 -85.5939 0.52736
1.6314 0.98803 5.5154e-05 3.8182 0.012028 2.1455e-05 0.0011544 0.17866 0.00065874 0.17931 0.1642 0 0.035236 0.0389 0 0.94029 0.26913 0.073983 0.010203 4.4818 0.063667 7.6947e-05 0.82641 0.0054972 0.0062386 0.0013996 0.98677 0.99159 3.0197e-06 1.2079e-05 0.13371 0.90057 0.89376 0.0014041 0.97689 0.55698 0.0018914 0.42683 1.7501 1.7489 16.0084 144.9852 0.00020031 -85.5944 0.52836
1.6324 0.98803 5.5154e-05 3.8182 0.012028 2.1469e-05 0.0011544 0.17871 0.00065874 0.17936 0.16424 0 0.035233 0.0389 0 0.94038 0.26917 0.073997 0.010205 4.4824 0.063678 7.6961e-05 0.8264 0.0054978 0.0062391 0.0013995 0.98677 0.99159 3.0195e-06 1.2078e-05 0.13372 0.90083 0.89389 0.0014041 0.97702 0.55714 0.0018914 0.42684 1.7508 1.7497 16.0083 144.9852 0.0002001 -85.595 0.52936
1.6334 0.98803 5.5154e-05 3.8182 0.012028 2.1482e-05 0.0011544 0.17875 0.00065874 0.17941 0.16428 0 0.035231 0.0389 0 0.94046 0.26921 0.074011 0.010206 4.483 0.063688 7.6975e-05 0.82639 0.0054983 0.0062397 0.0013994 0.98677 0.99159 3.0192e-06 1.2077e-05 0.13372 0.90109 0.89402 0.001404 0.97715 0.55729 0.0018913 0.42686 1.7515 1.7504 16.0083 144.9853 0.00019989 -85.5955 0.53036
1.6344 0.98803 5.5154e-05 3.8182 0.012028 2.1495e-05 0.0011544 0.1788 0.00065874 0.17945 0.16433 0 0.035228 0.0389 0 0.94055 0.26925 0.074026 0.010208 4.4835 0.063699 7.6989e-05 0.82638 0.0054988 0.0062402 0.0013993 0.98678 0.9916 3.0189e-06 1.2076e-05 0.13372 0.90135 0.89416 0.0014039 0.97728 0.55744 0.0018912 0.42687 1.7522 1.7511 16.0083 144.9853 0.00019968 -85.596 0.53136
1.6354 0.98803 5.5154e-05 3.8182 0.012028 2.1508e-05 0.0011544 0.17884 0.00065874 0.1795 0.16437 0 0.035225 0.0389 0 0.94064 0.26929 0.07404 0.01021 4.4841 0.063709 7.7002e-05 0.82637 0.0054993 0.0062407 0.0013992 0.98678 0.9916 3.0186e-06 1.2074e-05 0.13373 0.9016 0.89429 0.0014039 0.97741 0.5576 0.0018911 0.42688 1.753 1.7518 16.0083 144.9853 0.00019948 -85.5965 0.53236
1.6364 0.98803 5.5154e-05 3.8182 0.012028 2.1521e-05 0.0011544 0.17889 0.00065875 0.17954 0.16441 0 0.035223 0.0389 0 0.94073 0.26933 0.074054 0.010211 4.4847 0.06372 7.7016e-05 0.82636 0.0054999 0.0062413 0.001399 0.98678 0.9916 3.0184e-06 1.2073e-05 0.13373 0.90186 0.89442 0.0014038 0.97754 0.55775 0.001891 0.4269 1.7537 1.7525 16.0083 144.9853 0.00019927 -85.597 0.53336
1.6374 0.98803 5.5154e-05 3.8182 0.012028 2.1534e-05 0.0011544 0.17893 0.00065875 0.17959 0.16445 0 0.03522 0.0389 0 0.94082 0.26937 0.074068 0.010213 4.4852 0.06373 7.703e-05 0.82635 0.0055004 0.0062418 0.0013989 0.98678 0.9916 3.0181e-06 1.2072e-05 0.13374 0.90211 0.89455 0.0014038 0.97767 0.5579 0.0018909 0.42691 1.7544 1.7532 16.0083 144.9853 0.00019906 -85.5975 0.53436
1.6384 0.98803 5.5154e-05 3.8182 0.012028 2.1547e-05 0.0011544 0.17898 0.00065875 0.17963 0.1645 0 0.035217 0.0389 0 0.94091 0.26941 0.074082 0.010215 4.4858 0.063741 7.7044e-05 0.82634 0.0055009 0.0062424 0.0013988 0.98678 0.9916 3.0178e-06 1.2071e-05 0.13374 0.90237 0.89468 0.0014037 0.97779 0.55806 0.0018909 0.42692 1.7551 1.7539 16.0082 144.9854 0.00019886 -85.598 0.53536
1.6394 0.98803 5.5154e-05 3.8182 0.012028 2.156e-05 0.0011544 0.17902 0.00065875 0.17968 0.16454 0 0.035215 0.0389 0 0.94099 0.26945 0.074097 0.010216 4.4864 0.063751 7.7057e-05 0.82633 0.0055015 0.0062429 0.0013987 0.98678 0.9916 3.0176e-06 1.207e-05 0.13375 0.90262 0.89481 0.0014036 0.97792 0.55821 0.0018908 0.42693 1.7558 1.7546 16.0082 144.9854 0.00019865 -85.5984 0.53636
1.6404 0.98803 5.5154e-05 3.8182 0.012028 2.1574e-05 0.0011544 0.17907 0.00065875 0.17972 0.16458 0 0.035212 0.0389 0 0.94108 0.26949 0.074111 0.010218 4.487 0.063762 7.7071e-05 0.82632 0.005502 0.0062434 0.0013986 0.98678 0.9916 3.0173e-06 1.2069e-05 0.13375 0.90287 0.89494 0.0014036 0.97804 0.55837 0.0018907 0.42695 1.7565 1.7553 16.0082 144.9854 0.00019845 -85.5989 0.53736
1.6414 0.98803 5.5154e-05 3.8182 0.012028 2.1587e-05 0.0011544 0.17911 0.00065875 0.17977 0.16462 0 0.035209 0.0389 0 0.94117 0.26953 0.074125 0.01022 4.4875 0.063773 7.7085e-05 0.8263 0.0055025 0.006244 0.0013985 0.98679 0.9916 3.0171e-06 1.2068e-05 0.13375 0.90312 0.89507 0.0014035 0.97817 0.55852 0.0018906 0.42696 1.7572 1.756 16.0082 144.9854 0.00019825 -85.5994 0.53836
1.6424 0.98803 5.5154e-05 3.8182 0.012028 2.16e-05 0.0011544 0.17916 0.00065875 0.17981 0.16467 0 0.035207 0.0389 0 0.94126 0.26957 0.074139 0.010222 4.4881 0.063783 7.7099e-05 0.82629 0.005503 0.0062445 0.0013984 0.98679 0.9916 3.0168e-06 1.2067e-05 0.13376 0.90338 0.8952 0.0014035 0.97829 0.55867 0.0018906 0.42697 1.7579 1.7567 16.0082 144.9854 0.00019804 -85.5999 0.53936
1.6434 0.98803 5.5153e-05 3.8182 0.012028 2.1613e-05 0.0011544 0.1792 0.00065875 0.17986 0.16471 0 0.035204 0.0389 0 0.94135 0.26961 0.074154 0.010223 4.4887 0.063794 7.7112e-05 0.82628 0.0055036 0.0062451 0.0013983 0.98679 0.9916 3.0166e-06 1.2066e-05 0.13376 0.90363 0.89533 0.0014034 0.97841 0.55883 0.0018905 0.42699 1.7586 1.7574 16.0082 144.9855 0.00019784 -85.6004 0.54036
1.6444 0.98803 5.5153e-05 3.8182 0.012028 2.1626e-05 0.0011544 0.17925 0.00065875 0.1799 0.16475 0 0.035201 0.0389 0 0.94144 0.26965 0.074168 0.010225 4.4892 0.063804 7.7126e-05 0.82627 0.0055041 0.0062456 0.0013981 0.98679 0.9916 3.0163e-06 1.2065e-05 0.13377 0.90388 0.89545 0.0014033 0.97853 0.55898 0.0018904 0.427 1.7592 1.7581 16.0081 144.9855 0.00019764 -85.6008 0.54136
1.6454 0.98803 5.5153e-05 3.8182 0.012028 2.1639e-05 0.0011544 0.1793 0.00065875 0.17995 0.16479 0 0.035199 0.0389 0 0.94152 0.26969 0.074182 0.010227 4.4898 0.063815 7.714e-05 0.82626 0.0055046 0.0062462 0.001398 0.98679 0.99161 3.0161e-06 1.2064e-05 0.13377 0.90412 0.89558 0.0014033 0.97865 0.55913 0.0018903 0.42701 1.7599 1.7588 16.0081 144.9855 0.00019744 -85.6013 0.54236
1.6464 0.98803 5.5153e-05 3.8182 0.012028 2.1652e-05 0.0011544 0.17934 0.00065875 0.17999 0.16484 0 0.035196 0.0389 0 0.94161 0.26972 0.074196 0.010228 4.4904 0.063825 7.7154e-05 0.82625 0.0055052 0.0062467 0.0013979 0.98679 0.99161 3.0158e-06 1.2063e-05 0.13378 0.90437 0.89571 0.0014032 0.97877 0.55929 0.0018903 0.42702 1.7606 1.7595 16.0081 144.9855 0.00019724 -85.6018 0.54336
1.6474 0.98803 5.5153e-05 3.8182 0.012028 2.1665e-05 0.0011544 0.17939 0.00065875 0.18004 0.16488 0 0.035193 0.0389 0 0.9417 0.26976 0.074211 0.01023 4.491 0.063836 7.7167e-05 0.82624 0.0055057 0.0062472 0.0013978 0.98679 0.99161 3.0156e-06 1.2062e-05 0.13378 0.90462 0.89583 0.0014032 0.97889 0.55944 0.0018902 0.42704 1.7613 1.7602 16.0081 144.9855 0.00019705 -85.6022 0.54436
1.6484 0.98803 5.5153e-05 3.8182 0.012028 2.1678e-05 0.0011544 0.17943 0.00065875 0.18008 0.16492 0 0.035191 0.0389 0 0.94179 0.2698 0.074225 0.010232 4.4915 0.063847 7.7181e-05 0.82623 0.0055062 0.0062478 0.0013977 0.9868 0.99161 3.0153e-06 1.2061e-05 0.13379 0.90487 0.89596 0.0014031 0.97901 0.55959 0.0018901 0.42705 1.762 1.7609 16.0081 144.9856 0.00019685 -85.6027 0.54536
1.6494 0.98803 5.5153e-05 3.8182 0.012028 2.1692e-05 0.0011544 0.17948 0.00065875 0.18013 0.16496 0 0.035188 0.0389 0 0.94188 0.26984 0.074239 0.010233 4.4921 0.063857 7.7195e-05 0.82622 0.0055068 0.0062483 0.0013976 0.9868 0.99161 3.0151e-06 1.206e-05 0.13379 0.90511 0.89609 0.0014031 0.97913 0.55975 0.00189 0.42706 1.7627 1.7616 16.0081 144.9856 0.00019665 -85.6032 0.54636
1.6504 0.98803 5.5153e-05 3.8182 0.012028 2.1705e-05 0.0011544 0.17952 0.00065875 0.18017 0.16501 0 0.035185 0.0389 0 0.94197 0.26988 0.074253 0.010235 4.4927 0.063868 7.7209e-05 0.82621 0.0055073 0.0062489 0.0013975 0.9868 0.99161 3.0148e-06 1.2059e-05 0.13379 0.90536 0.89621 0.001403 0.97925 0.5599 0.00189 0.42708 1.7634 1.7623 16.008 144.9856 0.00019646 -85.6036 0.54736
1.6514 0.98803 5.5153e-05 3.8182 0.012028 2.1718e-05 0.0011544 0.17956 0.00065875 0.18022 0.16505 0 0.035183 0.0389 0 0.94205 0.26992 0.074268 0.010237 4.4933 0.063878 7.7223e-05 0.8262 0.0055078 0.0062494 0.0013974 0.9868 0.99161 3.0146e-06 1.2058e-05 0.1338 0.9056 0.89633 0.0014029 0.97936 0.56005 0.0018899 0.42709 1.764 1.7629 16.008 144.9856 0.00019626 -85.6041 0.54836
1.6524 0.98803 5.5153e-05 3.8182 0.012028 2.1731e-05 0.0011544 0.17961 0.00065876 0.18026 0.16509 0 0.03518 0.0389 0 0.94214 0.26996 0.074282 0.010239 4.4939 0.063889 7.7236e-05 0.82619 0.0055084 0.00625 0.0013973 0.9868 0.99161 3.0144e-06 1.2057e-05 0.1338 0.90584 0.89646 0.0014029 0.97948 0.5602 0.0018898 0.4271 1.7647 1.7636 16.008 144.9856 0.00019606 -85.6045 0.54936
1.6534 0.98803 5.5153e-05 3.8182 0.012028 2.1744e-05 0.0011544 0.17965 0.00065876 0.18031 0.16513 0 0.035178 0.0389 0 0.94223 0.27 0.074296 0.01024 4.4944 0.0639 7.725e-05 0.82618 0.0055089 0.0062505 0.0013972 0.9868 0.99161 3.0141e-06 1.2056e-05 0.13381 0.90609 0.89658 0.0014028 0.97959 0.56036 0.0018897 0.42711 1.7654 1.7643 16.008 144.9857 0.00019587 -85.605 0.55036
1.6544 0.98803 5.5153e-05 3.8182 0.012028 2.1757e-05 0.0011544 0.1797 0.00065876 0.18035 0.16517 0 0.035175 0.0389 0 0.94232 0.27004 0.07431 0.010242 4.495 0.06391 7.7264e-05 0.82617 0.0055094 0.0062511 0.0013971 0.9868 0.99161 3.0139e-06 1.2055e-05 0.13381 0.90633 0.8967 0.0014028 0.97971 0.56051 0.0018897 0.42713 1.7661 1.765 16.008 144.9857 0.00019568 -85.6054 0.55136
1.6554 0.98803 5.5153e-05 3.8182 0.012028 2.177e-05 0.0011544 0.17974 0.00065876 0.1804 0.16522 0 0.035172 0.0389 0 0.94241 0.27008 0.074325 0.010244 4.4956 0.063921 7.7278e-05 0.82616 0.0055099 0.0062516 0.001397 0.98681 0.99161 3.0136e-06 1.2054e-05 0.13382 0.90657 0.89683 0.0014027 0.97982 0.56066 0.0018896 0.42714 1.7667 1.7657 16.008 144.9857 0.00019549 -85.6058 0.55236
1.6564 0.98803 5.5153e-05 3.8182 0.012028 2.1783e-05 0.0011544 0.17979 0.00065876 0.18044 0.16526 0 0.03517 0.0389 0 0.9425 0.27012 0.074339 0.010245 4.4962 0.063931 7.7292e-05 0.82615 0.0055105 0.0062522 0.0013969 0.98681 0.99162 3.0134e-06 1.2054e-05 0.13382 0.90681 0.89695 0.0014027 0.97993 0.56082 0.0018895 0.42715 1.7674 1.7663 16.0079 144.9857 0.00019529 -85.6063 0.55336
1.6574 0.98803 5.5153e-05 3.8182 0.012028 2.1796e-05 0.0011544 0.17983 0.00065876 0.18049 0.1653 0 0.035167 0.0389 0 0.94259 0.27016 0.074353 0.010247 4.4968 0.063942 7.7305e-05 0.82614 0.005511 0.0062527 0.0013968 0.98681 0.99162 3.0132e-06 1.2053e-05 0.13382 0.90705 0.89707 0.0014026 0.98004 0.56097 0.0018895 0.42717 1.7681 1.767 16.0079 144.9857 0.0001951 -85.6067 0.55436
1.6584 0.98803 5.5153e-05 3.8182 0.012028 2.181e-05 0.0011544 0.17988 0.00065876 0.18053 0.16534 0 0.035165 0.0389 0 0.94267 0.2702 0.074368 0.010249 4.4973 0.063953 7.7319e-05 0.82612 0.0055115 0.0062533 0.0013967 0.98681 0.99162 3.013e-06 1.2052e-05 0.13383 0.90729 0.89719 0.0014026 0.98015 0.56112 0.0018894 0.42718 1.7688 1.7677 16.0079 144.9858 0.00019491 -85.6071 0.55536
1.6594 0.98803 5.5152e-05 3.8182 0.012028 2.1823e-05 0.0011544 0.17992 0.00065876 0.18058 0.16538 0 0.035162 0.0389 0 0.94276 0.27024 0.074382 0.01025 4.4979 0.063963 7.7333e-05 0.82611 0.0055121 0.0062538 0.0013966 0.98681 0.99162 3.0127e-06 1.2051e-05 0.13383 0.90753 0.89731 0.0014025 0.98026 0.56127 0.0018893 0.42719 1.7694 1.7683 16.0079 144.9858 0.00019472 -85.6076 0.55636
1.6604 0.98803 5.5152e-05 3.8182 0.012028 2.1836e-05 0.0011544 0.17997 0.00065876 0.18062 0.16543 0 0.035159 0.0389 0 0.94285 0.27028 0.074396 0.010252 4.4985 0.063974 7.7347e-05 0.8261 0.0055126 0.0062543 0.0013965 0.98681 0.99162 3.0125e-06 1.205e-05 0.13384 0.90776 0.89743 0.0014025 0.98037 0.56143 0.0018893 0.4272 1.7701 1.769 16.0079 144.9858 0.00019453 -85.608 0.55736
1.6614 0.98803 5.5152e-05 3.8182 0.012028 2.1849e-05 0.0011544 0.18001 0.00065876 0.18067 0.16547 0 0.035157 0.0389 0 0.94294 0.27032 0.07441 0.010254 4.4991 0.063984 7.736e-05 0.82609 0.0055131 0.0062549 0.0013964 0.98681 0.99162 3.0123e-06 1.2049e-05 0.13384 0.908 0.89755 0.0014024 0.98048 0.56158 0.0018892 0.42722 1.7708 1.7697 16.0078 144.9858 0.00019435 -85.6084 0.55836
1.6624 0.98803 5.5152e-05 3.8182 0.012028 2.1862e-05 0.0011544 0.18006 0.00065876 0.18071 0.16551 0 0.035154 0.0389 0 0.94303 0.27036 0.074425 0.010256 4.4997 0.063995 7.7374e-05 0.82608 0.0055137 0.0062554 0.0013963 0.98681 0.99162 3.012e-06 1.2048e-05 0.13385 0.90824 0.89767 0.0014024 0.98059 0.56173 0.0018891 0.42723 1.7714 1.7703 16.0078 144.9858 0.00019416 -85.6088 0.55936
1.6634 0.98803 5.5152e-05 3.8182 0.012028 2.1875e-05 0.0011544 0.1801 0.00065876 0.18075 0.16555 0 0.035151 0.0389 0 0.94312 0.2704 0.074439 0.010257 4.5002 0.064006 7.7388e-05 0.82607 0.0055142 0.006256 0.0013962 0.98682 0.99162 3.0118e-06 1.2047e-05 0.13385 0.90847 0.89779 0.0014023 0.9807 0.56188 0.0018891 0.42724 1.7721 1.771 16.0078 144.9859 0.00019397 -85.6092 0.56036
1.6644 0.98803 5.5152e-05 3.8182 0.012028 2.1888e-05 0.0011544 0.18014 0.00065876 0.1808 0.16559 0 0.035149 0.0389 0 0.94321 0.27044 0.074453 0.010259 4.5008 0.064016 7.7402e-05 0.82606 0.0055148 0.0062565 0.0013961 0.98682 0.99162 3.0116e-06 1.2046e-05 0.13386 0.90871 0.89791 0.0014023 0.98081 0.56203 0.001889 0.42726 1.7727 1.7717 16.0078 144.9859 0.00019378 -85.6097 0.56136
1.6654 0.98803 5.5152e-05 3.8182 0.012028 2.1901e-05 0.0011544 0.18019 0.00065876 0.18084 0.16564 0 0.035146 0.0389 0 0.94329 0.27048 0.074468 0.010261 4.5014 0.064027 7.7415e-05 0.82605 0.0055153 0.0062571 0.001396 0.98682 0.99162 3.0114e-06 1.2045e-05 0.13386 0.90894 0.89803 0.0014022 0.98091 0.56219 0.0018889 0.42727 1.7734 1.7723 16.0078 144.9859 0.0001936 -85.6101 0.56236
1.6664 0.98803 5.5152e-05 3.8182 0.012028 2.1914e-05 0.0011544 0.18023 0.00065876 0.18089 0.16568 0 0.035144 0.0389 0 0.94338 0.27052 0.074482 0.010262 4.502 0.064037 7.743e-05 0.82604 0.0055158 0.0062576 0.0013959 0.98682 0.99162 3.0112e-06 1.2045e-05 0.13386 0.90917 0.89814 0.0014022 0.98102 0.56234 0.0018889 0.42728 1.774 1.773 16.0078 144.9859 0.00019341 -85.6105 0.56336
1.6674 0.98803 5.5152e-05 3.8182 0.012028 2.1928e-05 0.0011544 0.18028 0.00065876 0.18093 0.16572 0 0.035141 0.0389 0 0.94347 0.27056 0.074496 0.010264 4.5026 0.064048 7.7444e-05 0.82603 0.0055164 0.0062582 0.0013958 0.98682 0.99162 3.011e-06 1.2044e-05 0.13387 0.9094 0.89826 0.0014021 0.98112 0.56249 0.0018888 0.42729 1.7747 1.7736 16.0077 144.9859 0.00019323 -85.6109 0.56436
1.6684 0.98803 5.5152e-05 3.8182 0.012028 2.1941e-05 0.0011544 0.18032 0.00065876 0.18098 0.16576 0 0.035139 0.0389 0 0.94356 0.2706 0.074511 0.010266 4.5032 0.064059 7.7457e-05 0.82602 0.0055169 0.0062587 0.0013957 0.98682 0.99162 3.0107e-06 1.2043e-05 0.13387 0.90964 0.89838 0.0014021 0.98123 0.56264 0.0018887 0.42731 1.7754 1.7743 16.0077 144.986 0.00019305 -85.6113 0.56536
1.6694 0.98803 5.5152e-05 3.8182 0.012028 2.1954e-05 0.0011544 0.18037 0.00065877 0.18102 0.1658 0 0.035136 0.0389 0 0.94365 0.27064 0.074525 0.010268 4.5037 0.064069 7.7471e-05 0.82601 0.0055174 0.0062593 0.0013956 0.98682 0.99163 3.0105e-06 1.2042e-05 0.13388 0.90987 0.89849 0.001402 0.98133 0.5628 0.0018887 0.42732 1.776 1.775 16.0077 144.986 0.00019286 -85.6117 0.56636
1.6704 0.98803 5.5152e-05 3.8182 0.012028 2.1967e-05 0.0011545 0.18041 0.00065877 0.18106 0.16584 0 0.035133 0.0389 0 0.94374 0.27068 0.074539 0.010269 4.5043 0.06408 7.7485e-05 0.826 0.005518 0.0062598 0.0013955 0.98682 0.99163 3.0103e-06 1.2041e-05 0.13388 0.9101 0.89861 0.001402 0.98143 0.56295 0.0018886 0.42733 1.7767 1.7756 16.0077 144.986 0.00019268 -85.6121 0.56736
1.6714 0.98803 5.5152e-05 3.8182 0.012028 2.198e-05 0.0011545 0.18045 0.00065877 0.18111 0.16589 0 0.035131 0.0389 0 0.94383 0.27072 0.074554 0.010271 4.5049 0.06409 7.7499e-05 0.82599 0.0055185 0.0062604 0.0013954 0.98683 0.99163 3.0101e-06 1.204e-05 0.13389 0.91033 0.89873 0.0014019 0.98153 0.5631 0.0018885 0.42735 1.7773 1.7763 16.0077 144.986 0.0001925 -85.6125 0.56836
1.6724 0.98803 5.5152e-05 3.8182 0.012028 2.1993e-05 0.0011545 0.1805 0.00065877 0.18115 0.16593 0 0.035128 0.0389 0 0.94392 0.27076 0.074568 0.010273 4.5055 0.064101 7.7513e-05 0.82598 0.005519 0.0062609 0.0013953 0.98683 0.99163 3.0099e-06 1.204e-05 0.13389 0.91055 0.89884 0.0014019 0.98163 0.56325 0.0018885 0.42736 1.7779 1.7769 16.0076 144.986 0.00019232 -85.6129 0.56936
1.6734 0.98803 5.5152e-05 3.8182 0.012028 2.2006e-05 0.0011545 0.18054 0.00065877 0.1812 0.16597 0 0.035126 0.0389 0 0.944 0.2708 0.074582 0.010274 4.5061 0.064112 7.7526e-05 0.82597 0.0055196 0.0062615 0.0013953 0.98683 0.99163 3.0097e-06 1.2039e-05 0.1339 0.91078 0.89896 0.0014018 0.98174 0.5634 0.0018884 0.42737 1.7786 1.7776 16.0076 144.9861 0.00019214 -85.6133 0.57036
1.6744 0.98803 5.5151e-05 3.8182 0.012028 2.2019e-05 0.0011545 0.18059 0.00065877 0.18124 0.16601 0 0.035123 0.0389 0 0.94409 0.27084 0.074597 0.010276 4.5067 0.064122 7.754e-05 0.82596 0.0055201 0.0062621 0.0013952 0.98683 0.99163 3.0095e-06 1.2038e-05 0.1339 0.91101 0.89907 0.0014018 0.98184 0.56356 0.0018884 0.42738 1.7792 1.7782 16.0076 144.9861 0.00019196 -85.6136 0.57136
1.6754 0.98803 5.5151e-05 3.8182 0.012028 2.2033e-05 0.0011545 0.18063 0.00065877 0.18129 0.16605 0 0.03512 0.0389 0 0.94418 0.27088 0.074611 0.010278 4.5073 0.064133 7.7554e-05 0.82594 0.0055207 0.0062626 0.0013951 0.98683 0.99163 3.0093e-06 1.2037e-05 0.1339 0.91124 0.89918 0.0014017 0.98194 0.56371 0.0018883 0.4274 1.7799 1.7788 16.0076 144.9861 0.00019178 -85.614 0.57236
1.6764 0.98803 5.5151e-05 3.8182 0.012027 2.2046e-05 0.0011545 0.18068 0.00065877 0.18133 0.16609 0 0.035118 0.0389 0 0.94427 0.27092 0.074625 0.010279 4.5079 0.064144 7.7568e-05 0.82593 0.0055212 0.0062632 0.001395 0.98683 0.99163 3.0091e-06 1.2036e-05 0.13391 0.91146 0.8993 0.0014017 0.98203 0.56386 0.0018882 0.42741 1.7805 1.7795 16.0076 144.9861 0.0001916 -85.6144 0.57336
1.6774 0.98803 5.5151e-05 3.8182 0.012027 2.2059e-05 0.0011545 0.18072 0.00065877 0.18137 0.16613 0 0.035115 0.0389 0 0.94436 0.27096 0.07464 0.010281 4.5084 0.064154 7.7582e-05 0.82592 0.0055217 0.0062637 0.0013949 0.98683 0.99163 3.0089e-06 1.2035e-05 0.13391 0.91169 0.89941 0.0014016 0.98213 0.56401 0.0018882 0.42742 1.7812 1.7801 16.0075 144.9861 0.00019143 -85.6148 0.57436
1.6784 0.98803 5.5151e-05 3.8182 0.012027 2.2072e-05 0.0011545 0.18076 0.00065877 0.18142 0.16618 0 0.035113 0.0389 0 0.94445 0.271 0.074654 0.010283 4.509 0.064165 7.7596e-05 0.82591 0.0055223 0.0062643 0.0013948 0.98683 0.99163 3.0087e-06 1.2035e-05 0.13392 0.91191 0.89952 0.0014016 0.98223 0.56416 0.0018881 0.42744 1.7818 1.7808 16.0075 144.9862 0.00019125 -85.6152 0.57536
1.6794 0.98803 5.5151e-05 3.8182 0.012027 2.2085e-05 0.0011545 0.18081 0.00065877 0.18146 0.16622 0 0.03511 0.0389 0 0.94454 0.27104 0.074668 0.010285 4.5096 0.064175 7.761e-05 0.8259 0.0055228 0.0062648 0.0013947 0.98683 0.99163 3.0085e-06 1.2034e-05 0.13392 0.91214 0.89963 0.0014015 0.98233 0.56431 0.001888 0.42745 1.7824 1.7814 16.0075 144.9862 0.00019107 -85.6155 0.57636
1.6804 0.98803 5.5151e-05 3.8182 0.012027 2.2098e-05 0.0011545 0.18085 0.00065877 0.1815 0.16626 0 0.035108 0.0389 0 0.94463 0.27108 0.074683 0.010286 4.5102 0.064186 7.7623e-05 0.82589 0.0055234 0.0062654 0.0013946 0.98684 0.99163 3.0083e-06 1.2033e-05 0.13393 0.91236 0.89975 0.0014015 0.98242 0.56446 0.001888 0.42746 1.7831 1.782 16.0075 144.9862 0.0001909 -85.6159 0.57736
1.6814 0.98803 5.5151e-05 3.8182 0.012027 2.2111e-05 0.0011545 0.18089 0.00065877 0.18155 0.1663 0 0.035105 0.0389 0 0.94472 0.27111 0.074697 0.010288 4.5108 0.064197 7.7637e-05 0.82588 0.0055239 0.0062659 0.0013945 0.98684 0.99163 3.0081e-06 1.2032e-05 0.13393 0.91258 0.89986 0.0014014 0.98252 0.56462 0.0018879 0.42747 1.7837 1.7827 16.0075 144.9862 0.00019072 -85.6163 0.57836
1.6824 0.98803 5.5151e-05 3.8182 0.012027 2.2124e-05 0.0011545 0.18094 0.00065877 0.18159 0.16634 0 0.035103 0.0389 0 0.9448 0.27115 0.074711 0.01029 4.5114 0.064207 7.7651e-05 0.82587 0.0055244 0.0062665 0.0013945 0.98684 0.99164 3.0079e-06 1.2031e-05 0.13394 0.9128 0.89997 0.0014014 0.98261 0.56477 0.0018879 0.42749 1.7843 1.7833 16.0074 144.9862 0.00019055 -85.6166 0.57936
1.6834 0.98803 5.5151e-05 3.8182 0.012027 2.2137e-05 0.0011545 0.18098 0.00065877 0.18164 0.16638 0 0.0351 0.0389 0 0.94489 0.27119 0.074726 0.010291 4.512 0.064218 7.7665e-05 0.82586 0.005525 0.006267 0.0013944 0.98684 0.99164 3.0077e-06 1.2031e-05 0.13394 0.91302 0.90008 0.0014014 0.98271 0.56492 0.0018878 0.4275 1.785 1.7839 16.0074 144.9863 0.00019038 -85.617 0.58036
1.6844 0.98803 5.5151e-05 3.8182 0.012027 2.2151e-05 0.0011545 0.18103 0.00065877 0.18168 0.16642 0 0.035097 0.0389 0 0.94498 0.27123 0.07474 0.010293 4.5126 0.064229 7.7679e-05 0.82585 0.0055255 0.0062676 0.0013943 0.98684 0.99164 3.0075e-06 1.203e-05 0.13394 0.91324 0.90019 0.0014013 0.9828 0.56507 0.0018878 0.42751 1.7856 1.7846 16.0074 144.9863 0.0001902 -85.6174 0.58136
1.6854 0.98803 5.5151e-05 3.8182 0.012027 2.2164e-05 0.0011545 0.18107 0.00065877 0.18172 0.16646 0 0.035095 0.0389 0 0.94507 0.27127 0.074754 0.010295 4.5132 0.064239 7.7693e-05 0.82584 0.0055261 0.0062681 0.0013942 0.98684 0.99164 3.0073e-06 1.2029e-05 0.13395 0.91346 0.9003 0.0014013 0.9829 0.56522 0.0018877 0.42753 1.7862 1.7852 16.0074 144.9863 0.00019003 -85.6177 0.58236
1.6864 0.98803 5.5151e-05 3.8182 0.012027 2.2177e-05 0.0011545 0.18111 0.00065877 0.18177 0.16651 0 0.035092 0.0389 0 0.94516 0.27131 0.074769 0.010297 4.5138 0.06425 7.7707e-05 0.82583 0.0055266 0.0062687 0.0013941 0.98684 0.99164 3.0071e-06 1.2028e-05 0.13395 0.91368 0.90041 0.0014012 0.98299 0.56537 0.0018876 0.42754 1.7868 1.7858 16.0074 144.9863 0.00018986 -85.6181 0.58336
1.6874 0.98803 5.5151e-05 3.8182 0.012027 2.219e-05 0.0011545 0.18116 0.00065878 0.18181 0.16655 0 0.03509 0.0389 0 0.94525 0.27135 0.074783 0.010298 4.5144 0.064261 7.772e-05 0.82582 0.0055271 0.0062693 0.001394 0.98684 0.99164 3.0069e-06 1.2028e-05 0.13396 0.9139 0.90052 0.0014012 0.98308 0.56552 0.0018876 0.42755 1.7875 1.7865 16.0074 144.9863 0.00018969 -85.6184 0.58436
1.6884 0.98803 5.5151e-05 3.8182 0.012027 2.2203e-05 0.0011545 0.1812 0.00065878 0.18185 0.16659 0 0.035087 0.0389 0 0.94534 0.27139 0.074797 0.0103 4.515 0.064271 7.7734e-05 0.82581 0.0055277 0.0062698 0.001394 0.98684 0.99164 3.0067e-06 1.2027e-05 0.13396 0.91412 0.90063 0.0014011 0.98317 0.56567 0.0018875 0.42756 1.7881 1.7871 16.0073 144.9864 0.00018952 -85.6188 0.58536
1.6894 0.98803 5.5151e-05 3.8182 0.012027 2.2216e-05 0.0011545 0.18124 0.00065878 0.1819 0.16663 0 0.035085 0.0389 0 0.94543 0.27143 0.074812 0.010302 4.5156 0.064282 7.7748e-05 0.8258 0.0055282 0.0062704 0.0013939 0.98685 0.99164 3.0066e-06 1.2026e-05 0.13397 0.91433 0.90073 0.0014011 0.98326 0.56583 0.0018875 0.42758 1.7887 1.7877 16.0073 144.9864 0.00018935 -85.6191 0.58636
1.6904 0.98803 5.515e-05 3.8182 0.012027 2.2229e-05 0.0011545 0.18129 0.00065878 0.18194 0.16667 0 0.035082 0.0389 0 0.94552 0.27147 0.074826 0.010303 4.5161 0.064293 7.7762e-05 0.82579 0.0055288 0.0062709 0.0013938 0.98685 0.99164 3.0064e-06 1.2025e-05 0.13397 0.91455 0.90084 0.0014011 0.98335 0.56598 0.0018874 0.42759 1.7893 1.7883 16.0073 144.9864 0.00018918 -85.6195 0.58736
1.6914 0.98803 5.515e-05 3.8182 0.012027 2.2242e-05 0.0011545 0.18133 0.00065878 0.18198 0.16671 0 0.03508 0.0389 0 0.94561 0.27151 0.074841 0.010305 4.5167 0.064303 7.7776e-05 0.82577 0.0055293 0.0062715 0.0013937 0.98685 0.99164 3.0062e-06 1.2025e-05 0.13398 0.91477 0.90095 0.001401 0.98344 0.56613 0.0018874 0.4276 1.7899 1.789 16.0073 144.9864 0.00018901 -85.6198 0.58836
1.6924 0.98803 5.515e-05 3.8182 0.012027 2.2255e-05 0.0011545 0.18137 0.00065878 0.18203 0.16675 0 0.035077 0.0389 0 0.9457 0.27155 0.074855 0.010307 4.5173 0.064314 7.779e-05 0.82576 0.0055298 0.006272 0.0013936 0.98685 0.99164 3.006e-06 1.2024e-05 0.13398 0.91498 0.90106 0.001401 0.98353 0.56628 0.0018873 0.42762 1.7906 1.7896 16.0072 144.9864 0.00018884 -85.6202 0.58936
1.6934 0.98803 5.515e-05 3.8182 0.012027 2.2269e-05 0.0011545 0.18142 0.00065878 0.18207 0.16679 0 0.035075 0.0389 0 0.94578 0.27159 0.074869 0.010309 4.5179 0.064324 7.7804e-05 0.82575 0.0055304 0.0062726 0.0013936 0.98685 0.99164 3.0058e-06 1.2023e-05 0.13399 0.91519 0.90116 0.0014009 0.98362 0.56643 0.0018872 0.42763 1.7912 1.7902 16.0072 144.9865 0.00018867 -85.6205 0.59036
1.6944 0.98803 5.515e-05 3.8182 0.012027 2.2282e-05 0.0011545 0.18146 0.00065878 0.18211 0.16683 0 0.035072 0.0389 0 0.94587 0.27163 0.074884 0.01031 4.5185 0.064335 7.7818e-05 0.82574 0.0055309 0.0062732 0.0013935 0.98685 0.99164 3.0056e-06 1.2022e-05 0.13399 0.91541 0.90127 0.0014009 0.98371 0.56658 0.0018872 0.42764 1.7918 1.7908 16.0072 144.9865 0.00018851 -85.6209 0.59136
1.6954 0.98803 5.515e-05 3.8182 0.012027 2.2295e-05 0.0011545 0.1815 0.00065878 0.18216 0.16687 0 0.03507 0.0389 0 0.94596 0.27167 0.074898 0.010312 4.5191 0.064346 7.7832e-05 0.82573 0.0055315 0.0062737 0.0013934 0.98685 0.99164 3.0055e-06 1.2022e-05 0.13399 0.91562 0.90137 0.0014008 0.98379 0.56673 0.0018871 0.42765 1.7924 1.7914 16.0072 144.9865 0.00018834 -85.6212 0.59236
1.6964 0.98803 5.515e-05 3.8182 0.012027 2.2308e-05 0.0011545 0.18155 0.00065878 0.1822 0.16691 0 0.035067 0.0389 0 0.94605 0.27171 0.074912 0.010314 4.5197 0.064356 7.7845e-05 0.82572 0.005532 0.0062743 0.0013933 0.98685 0.99164 3.0053e-06 1.2021e-05 0.134 0.91583 0.90148 0.0014008 0.98388 0.56688 0.0018871 0.42767 1.793 1.792 16.0072 144.9865 0.00018818 -85.6215 0.59336
1.6974 0.98803 5.515e-05 3.8182 0.012027 2.2321e-05 0.0011545 0.18159 0.00065878 0.18224 0.16695 0 0.035065 0.0389 0 0.94614 0.27175 0.074927 0.010315 4.5203 0.064367 7.7859e-05 0.82571 0.0055326 0.0062748 0.0013933 0.98685 0.99165 3.0051e-06 1.202e-05 0.134 0.91604 0.90158 0.0014008 0.98397 0.56703 0.001887 0.42768 1.7936 1.7926 16.0071 144.9865 0.00018801 -85.6219 0.59436
1.6984 0.98803 5.515e-05 3.8182 0.012027 2.2334e-05 0.0011545 0.18163 0.00065878 0.18229 0.167 0 0.035062 0.0389 0 0.94623 0.27179 0.074941 0.010317 4.5209 0.064378 7.7873e-05 0.8257 0.0055331 0.0062754 0.0013932 0.98685 0.99165 3.0049e-06 1.202e-05 0.13401 0.91625 0.90169 0.0014007 0.98405 0.56718 0.001887 0.42769 1.7942 1.7933 16.0071 144.9866 0.00018785 -85.6222 0.59536
1.6994 0.98803 5.515e-05 3.8182 0.012027 2.2347e-05 0.0011545 0.18168 0.00065878 0.18233 0.16704 0 0.035059 0.0389 0 0.94632 0.27183 0.074956 0.010319 4.5215 0.064388 7.7887e-05 0.82569 0.0055337 0.006276 0.0013931 0.98686 0.99165 3.0048e-06 1.2019e-05 0.13401 0.91646 0.90179 0.0014007 0.98414 0.56733 0.0018869 0.42771 1.7948 1.7939 16.0071 144.9866 0.00018768 -85.6225 0.59636
1.7004 0.98803 5.515e-05 3.8182 0.012027 2.236e-05 0.0011545 0.18172 0.00065878 0.18237 0.16708 0 0.035057 0.0389 0 0.94641 0.27187 0.07497 0.01032 4.5221 0.064399 7.7901e-05 0.82568 0.0055342 0.0062765 0.001393 0.98686 0.99165 3.0046e-06 1.2018e-05 0.13402 0.91667 0.9019 0.0014006 0.98422 0.56748 0.0018869 0.42772 1.7954 1.7945 16.0071 144.9866 0.00018752 -85.6228 0.59736
1.7014 0.98803 5.515e-05 3.8182 0.012027 2.2373e-05 0.0011545 0.18176 0.00065878 0.18242 0.16712 0 0.035054 0.0389 0 0.9465 0.27191 0.074984 0.010322 4.5227 0.06441 7.7915e-05 0.82567 0.0055347 0.0062771 0.0013929 0.98686 0.99165 3.0044e-06 1.2018e-05 0.13402 0.91688 0.902 0.0014006 0.98431 0.56763 0.0018868 0.42773 1.796 1.7951 16.0071 144.9866 0.00018736 -85.6232 0.59836
1.7024 0.98803 5.515e-05 3.8182 0.012027 2.2387e-05 0.0011545 0.18181 0.00065878 0.18246 0.16716 0 0.035052 0.0389 0 0.94659 0.27195 0.074999 0.010324 4.5233 0.06442 7.7929e-05 0.82566 0.0055353 0.0062776 0.0013929 0.98686 0.99165 3.0043e-06 1.2017e-05 0.13403 0.91709 0.9021 0.0014006 0.98439 0.56778 0.0018868 0.42774 1.7966 1.7957 16.007 144.9866 0.0001872 -85.6235 0.59936
1.7034 0.98803 5.515e-05 3.8182 0.012027 2.24e-05 0.0011545 0.18185 0.00065878 0.1825 0.1672 0 0.035049 0.0389 0 0.94668 0.27199 0.075013 0.010326 4.5239 0.064431 7.7943e-05 0.82565 0.0055358 0.0062782 0.0013928 0.98686 0.99165 3.0041e-06 1.2016e-05 0.13403 0.9173 0.90221 0.0014005 0.98447 0.56793 0.0018867 0.42776 1.7972 1.7963 16.007 144.9867 0.00018703 -85.6238 0.60036
1.7044 0.98803 5.515e-05 3.8182 0.012027 2.2413e-05 0.0011545 0.18189 0.00065879 0.18255 0.16724 0 0.035047 0.0389 0 0.94677 0.27203 0.075028 0.010327 4.5245 0.064442 7.7957e-05 0.82564 0.0055364 0.0062788 0.0013927 0.98686 0.99165 3.0039e-06 1.2016e-05 0.13403 0.91751 0.90231 0.0014005 0.98456 0.56809 0.0018867 0.42777 1.7978 1.7969 16.007 144.9867 0.00018687 -85.6241 0.60136
1.7054 0.98803 5.5149e-05 3.8182 0.012027 2.2426e-05 0.0011545 0.18194 0.00065879 0.18259 0.16728 0 0.035044 0.0389 0 0.94686 0.27207 0.075042 0.010329 4.5251 0.064452 7.797e-05 0.82563 0.0055369 0.0062793 0.0013927 0.98686 0.99165 3.0037e-06 1.2015e-05 0.13404 0.91771 0.90241 0.0014004 0.98464 0.56824 0.0018866 0.42778 1.7984 1.7975 16.007 144.9867 0.00018671 -85.6244 0.60236
1.7064 0.98803 5.5149e-05 3.8182 0.012027 2.2439e-05 0.0011545 0.18198 0.00065879 0.18263 0.16732 0 0.035042 0.0389 0 0.94694 0.27211 0.075056 0.010331 4.5257 0.064463 7.7984e-05 0.82561 0.0055375 0.0062799 0.0013926 0.98686 0.99165 3.0036e-06 1.2014e-05 0.13404 0.91792 0.90251 0.0014004 0.98472 0.56839 0.0018866 0.42779 1.799 1.7981 16.007 144.9867 0.00018655 -85.6247 0.60336
1.7074 0.98803 5.5149e-05 3.8182 0.012027 2.2452e-05 0.0011545 0.18202 0.00065879 0.18268 0.16736 0 0.035039 0.0389 0 0.94703 0.27215 0.075071 0.010332 4.5263 0.064474 7.7998e-05 0.8256 0.005538 0.0062804 0.0013925 0.98686 0.99165 3.0034e-06 1.2014e-05 0.13405 0.91812 0.90261 0.0014004 0.9848 0.56854 0.0018865 0.42781 1.7996 1.7987 16.0069 144.9867 0.00018639 -85.625 0.60436
1.7084 0.98803 5.5149e-05 3.8182 0.012027 2.2465e-05 0.0011545 0.18206 0.00065879 0.18272 0.1674 0 0.035037 0.0389 0 0.94712 0.27219 0.075085 0.010334 4.5269 0.064484 7.8012e-05 0.82559 0.0055386 0.006281 0.0013924 0.98686 0.99165 3.0033e-06 1.2013e-05 0.13405 0.91833 0.90271 0.0014003 0.98488 0.56869 0.0018865 0.42782 1.8002 1.7993 16.0069 144.9868 0.00018624 -85.6254 0.60536
1.7094 0.98803 5.5149e-05 3.8182 0.012027 2.2478e-05 0.0011545 0.18211 0.00065879 0.18276 0.16744 0 0.035034 0.0389 0 0.94721 0.27223 0.0751 0.010336 4.5275 0.064495 7.8026e-05 0.82558 0.0055391 0.0062816 0.0013924 0.98687 0.99165 3.0031e-06 1.2012e-05 0.13406 0.91853 0.90281 0.0014003 0.98496 0.56884 0.0018864 0.42783 1.8008 1.7999 16.0069 144.9868 0.00018608 -85.6257 0.60636
1.7104 0.98803 5.5149e-05 3.8182 0.012027 2.2491e-05 0.0011545 0.18215 0.00065879 0.1828 0.16748 0 0.035032 0.0389 0 0.9473 0.27227 0.075114 0.010338 4.5281 0.064506 7.804e-05 0.82557 0.0055397 0.0062821 0.0013923 0.98687 0.99165 3.0029e-06 1.2012e-05 0.13406 0.91873 0.90291 0.0014003 0.98504 0.56899 0.0018864 0.42785 1.8014 1.8005 16.0069 144.9868 0.00018592 -85.626 0.60736
1.7114 0.98803 5.5149e-05 3.8182 0.012027 2.2505e-05 0.0011545 0.18219 0.00065879 0.18285 0.16752 0 0.03503 0.0389 0 0.94739 0.27231 0.075129 0.010339 4.5287 0.064517 7.8054e-05 0.82556 0.0055402 0.0062827 0.0013922 0.98687 0.99165 3.0028e-06 1.2011e-05 0.13407 0.91894 0.90301 0.0014002 0.98512 0.56914 0.0018863 0.42786 1.802 1.8011 16.0069 144.9868 0.00018576 -85.6263 0.60836
1.7124 0.98803 5.5149e-05 3.8182 0.012027 2.2518e-05 0.0011545 0.18223 0.00065879 0.18289 0.16756 0 0.035027 0.0389 0 0.94748 0.27235 0.075143 0.010341 4.5294 0.064527 7.8068e-05 0.82555 0.0055408 0.0062833 0.0013922 0.98687 0.99165 3.0026e-06 1.201e-05 0.13407 0.91914 0.90311 0.0014002 0.9852 0.56929 0.0018863 0.42787 1.8026 1.8017 16.0068 144.9868 0.00018561 -85.6266 0.60936
1.7134 0.98803 5.5149e-05 3.8182 0.012027 2.2531e-05 0.0011545 0.18228 0.00065879 0.18293 0.1676 0 0.035025 0.0389 0 0.94757 0.27239 0.075157 0.010343 4.53 0.064538 7.8082e-05 0.82554 0.0055413 0.0062838 0.0013921 0.98687 0.99166 3.0025e-06 1.201e-05 0.13408 0.91934 0.90321 0.0014001 0.98527 0.56944 0.0018862 0.42788 1.8032 1.8022 16.0068 144.9869 0.00018545 -85.6269 0.61036
1.7144 0.98803 5.5149e-05 3.8182 0.012027 2.2544e-05 0.0011545 0.18232 0.00065879 0.18297 0.16764 0 0.035022 0.0389 0 0.94766 0.27243 0.075172 0.010344 4.5306 0.064549 7.8096e-05 0.82553 0.0055419 0.0062844 0.001392 0.98687 0.99166 3.0023e-06 1.2009e-05 0.13408 0.91954 0.90331 0.0014001 0.98535 0.56958 0.0018862 0.4279 1.8038 1.8028 16.0068 144.9869 0.0001853 -85.6272 0.61136
1.7154 0.98803 5.5149e-05 3.8182 0.012027 2.2557e-05 0.0011545 0.18236 0.00065879 0.18302 0.16768 0 0.03502 0.0389 0 0.94775 0.27247 0.075186 0.010346 4.5312 0.064559 7.811e-05 0.82552 0.0055424 0.0062849 0.0013919 0.98687 0.99166 3.0021e-06 1.2008e-05 0.13408 0.91974 0.90341 0.0014001 0.98543 0.56973 0.0018861 0.42791 1.8043 1.8034 16.0068 144.9869 0.00018514 -85.6275 0.61236
1.7164 0.98803 5.5149e-05 3.8182 0.012027 2.257e-05 0.0011545 0.18241 0.00065879 0.18306 0.16772 0 0.035017 0.0389 0 0.94784 0.27251 0.075201 0.010348 4.5318 0.06457 7.8124e-05 0.82551 0.0055429 0.0062855 0.0013919 0.98687 0.99166 3.002e-06 1.2008e-05 0.13409 0.91994 0.90351 0.0014 0.98551 0.56988 0.0018861 0.42792 1.8049 1.804 16.0067 144.9869 0.00018499 -85.6277 0.61336
1.7174 0.98803 5.5149e-05 3.8182 0.012027 2.2583e-05 0.0011545 0.18245 0.00065879 0.1831 0.16776 0 0.035015 0.0389 0 0.94793 0.27255 0.075215 0.01035 4.5324 0.064581 7.8138e-05 0.8255 0.0055435 0.0062861 0.0013918 0.98687 0.99166 3.0018e-06 1.2007e-05 0.13409 0.92014 0.90361 0.0014 0.98558 0.57003 0.001886 0.42793 1.8055 1.8046 16.0067 144.9869 0.00018484 -85.628 0.61436
1.7184 0.98803 5.5149e-05 3.8182 0.012027 2.2596e-05 0.0011545 0.18249 0.00065879 0.18314 0.1678 0 0.035012 0.0389 0 0.94802 0.27259 0.07523 0.010351 4.533 0.064591 7.8152e-05 0.82549 0.005544 0.0062866 0.0013917 0.98687 0.99166 3.0017e-06 1.2007e-05 0.1341 0.92034 0.9037 0.0014 0.98566 0.57018 0.001886 0.42795 1.8061 1.8052 16.0067 144.987 0.00018468 -85.6283 0.61536
1.7194 0.98803 5.5149e-05 3.8182 0.012027 2.261e-05 0.0011545 0.18253 0.00065879 0.18319 0.16784 0 0.03501 0.0389 0 0.94811 0.27264 0.075244 0.010353 4.5336 0.064602 7.8166e-05 0.82548 0.0055446 0.0062872 0.0013917 0.98687 0.99166 3.0015e-06 1.2006e-05 0.1341 0.92053 0.9038 0.0013999 0.98573 0.57033 0.001886 0.42796 1.8067 1.8057 16.0067 144.987 0.00018453 -85.6286 0.61636
1.7204 0.98803 5.5149e-05 3.8182 0.012027 2.2623e-05 0.0011545 0.18258 0.00065879 0.18323 0.16788 0 0.035007 0.0389 0 0.9482 0.27268 0.075259 0.010355 4.5342 0.064613 7.818e-05 0.82547 0.0055451 0.0062878 0.0013916 0.98687 0.99166 3.0014e-06 1.2005e-05 0.13411 0.92073 0.9039 0.0013999 0.98581 0.57048 0.0018859 0.42797 1.8072 1.8063 16.0067 144.987 0.00018438 -85.6289 0.61736
1.7214 0.98803 5.5148e-05 3.8182 0.012027 2.2636e-05 0.0011545 0.18262 0.00065879 0.18327 0.16792 0 0.035005 0.0389 0 0.94829 0.27272 0.075273 0.010357 4.5348 0.064623 7.8194e-05 0.82545 0.0055457 0.0062883 0.0013915 0.98688 0.99166 3.0012e-06 1.2005e-05 0.13411 0.92093 0.90399 0.0013999 0.98588 0.57063 0.0018859 0.42799 1.8078 1.8069 16.0066 144.987 0.00018423 -85.6292 0.61836
1.7224 0.98803 5.5148e-05 3.8182 0.012027 2.2649e-05 0.0011545 0.18266 0.0006588 0.18331 0.16796 0 0.035002 0.0389 0 0.94838 0.27276 0.075288 0.010358 4.5354 0.064634 7.8207e-05 0.82544 0.0055462 0.0062889 0.0013915 0.98688 0.99166 3.0011e-06 1.2004e-05 0.13412 0.92112 0.90409 0.0013998 0.98595 0.57078 0.0018858 0.428 1.8084 1.8075 16.0066 144.987 0.00018408 -85.6295 0.61936
1.7234 0.98803 5.5148e-05 3.8182 0.012027 2.2662e-05 0.0011545 0.1827 0.0006588 0.18336 0.168 0 0.035 0.0389 0 0.94847 0.2728 0.075302 0.01036 4.536 0.064645 7.8221e-05 0.82543 0.0055468 0.0062895 0.0013914 0.98688 0.99166 3.0009e-06 1.2004e-05 0.13412 0.92132 0.90418 0.0013998 0.98603 0.57093 0.0018858 0.42801 1.809 1.8081 16.0066 144.9871 0.00018393 -85.6297 0.62036
1.7244 0.98803 5.5148e-05 3.8182 0.012027 2.2675e-05 0.0011545 0.18274 0.0006588 0.1834 0.16804 0 0.034997 0.0389 0 0.94856 0.27284 0.075316 0.010362 4.5366 0.064656 7.8235e-05 0.82542 0.0055474 0.00629 0.0013914 0.98688 0.99166 3.0008e-06 1.2003e-05 0.13413 0.92151 0.90428 0.0013998 0.9861 0.57108 0.0018857 0.42802 1.8095 1.8086 16.0066 144.9871 0.00018378 -85.63 0.62136
1.7254 0.98803 5.5148e-05 3.8182 0.012027 2.2688e-05 0.0011545 0.18279 0.0006588 0.18344 0.16808 0 0.034995 0.0389 0 0.94865 0.27288 0.075331 0.010363 4.5373 0.064666 7.8249e-05 0.82541 0.0055479 0.0062906 0.0013913 0.98688 0.99166 3.0006e-06 1.2002e-05 0.13413 0.9217 0.90437 0.0013997 0.98617 0.57123 0.0018857 0.42804 1.8101 1.8092 16.0065 144.9871 0.00018363 -85.6303 0.62236
1.7264 0.98803 5.5148e-05 3.8182 0.012027 2.2701e-05 0.0011545 0.18283 0.0006588 0.18348 0.16812 0 0.034992 0.0389 0 0.94873 0.27292 0.075345 0.010365 4.5379 0.064677 7.8263e-05 0.8254 0.0055485 0.0062912 0.0013912 0.98688 0.99166 3.0005e-06 1.2002e-05 0.13413 0.9219 0.90447 0.0013997 0.98624 0.57138 0.0018856 0.42805 1.8107 1.8098 16.0065 144.9871 0.00018348 -85.6306 0.62336
1.7274 0.98803 5.5148e-05 3.8182 0.012027 2.2714e-05 0.0011545 0.18287 0.0006588 0.18353 0.16816 0 0.03499 0.0389 0 0.94882 0.27296 0.07536 0.010367 4.5385 0.064688 7.8277e-05 0.82539 0.005549 0.0062917 0.0013912 0.98688 0.99166 3.0003e-06 1.2001e-05 0.13414 0.92209 0.90456 0.0013997 0.98631 0.57153 0.0018856 0.42806 1.8112 1.8103 16.0065 144.9872 0.00018333 -85.6308 0.62436
1.7284 0.98803 5.5148e-05 3.8182 0.012027 2.2728e-05 0.0011545 0.18291 0.0006588 0.18357 0.1682 0 0.034988 0.0389 0 0.94891 0.273 0.075374 0.010369 4.5391 0.064698 7.8291e-05 0.82538 0.0055496 0.0062923 0.0013911 0.98688 0.99166 3.0002e-06 1.2001e-05 0.13414 0.92228 0.90466 0.0013996 0.98638 0.57168 0.0018856 0.42807 1.8118 1.8109 16.0065 144.9872 0.00018318 -85.6311 0.62536
1.7294 0.98803 5.5148e-05 3.8182 0.012027 2.2741e-05 0.0011545 0.18296 0.0006588 0.18361 0.16824 0 0.034985 0.0389 0 0.949 0.27304 0.075389 0.01037 4.5397 0.064709 7.8305e-05 0.82537 0.0055501 0.0062929 0.001391 0.98688 0.99166 3.0001e-06 1.2e-05 0.13415 0.92247 0.90475 0.0013996 0.98645 0.57182 0.0018855 0.42809 1.8124 1.8115 16.0065 144.9872 0.00018304 -85.6314 0.62636
1.7304 0.98803 5.5148e-05 3.8182 0.012027 2.2754e-05 0.0011545 0.183 0.0006588 0.18365 0.16828 0 0.034983 0.0389 0 0.94909 0.27308 0.075403 0.010372 4.5403 0.06472 7.8319e-05 0.82536 0.0055507 0.0062934 0.001391 0.98688 0.99166 2.9999e-06 1.2e-05 0.13415 0.92266 0.90484 0.0013996 0.98652 0.57197 0.0018855 0.4281 1.8129 1.8121 16.0064 144.9872 0.00018289 -85.6316 0.62736
1.7314 0.98803 5.5148e-05 3.8182 0.012027 2.2767e-05 0.0011545 0.18304 0.0006588 0.18369 0.16832 0 0.03498 0.0389 0 0.94918 0.27312 0.075418 0.010374 4.5409 0.06473 7.8333e-05 0.82535 0.0055512 0.006294 0.0013909 0.98688 0.99166 2.9998e-06 1.1999e-05 0.13416 0.92285 0.90494 0.0013995 0.98659 0.57212 0.0018854 0.42811 1.8135 1.8126 16.0064 144.9872 0.00018275 -85.6319 0.62836
1.7324 0.98803 5.5148e-05 3.8182 0.012027 2.278e-05 0.0011545 0.18308 0.0006588 0.18374 0.16836 0 0.034978 0.0389 0 0.94927 0.27316 0.075432 0.010375 4.5415 0.064741 7.8347e-05 0.82534 0.0055518 0.0062946 0.0013909 0.98688 0.99167 2.9996e-06 1.1998e-05 0.13416 0.92304 0.90503 0.0013995 0.98666 0.57227 0.0018854 0.42813 1.8141 1.8132 16.0064 144.9873 0.0001826 -85.6322 0.62936
1.7334 0.98803 5.5148e-05 3.8182 0.012027 2.2793e-05 0.0011545 0.18312 0.0006588 0.18378 0.1684 0 0.034975 0.0389 0 0.94936 0.2732 0.075447 0.010377 4.5422 0.064752 7.8361e-05 0.82533 0.0055523 0.0062952 0.0013908 0.98689 0.99167 2.9995e-06 1.1998e-05 0.13417 0.92323 0.90512 0.0013995 0.98673 0.57242 0.0018853 0.42814 1.8146 1.8137 16.0064 144.9873 0.00018246 -85.6324 0.63036
1.7344 0.98803 5.5148e-05 3.8182 0.012027 2.2806e-05 0.0011545 0.18317 0.0006588 0.18382 0.16844 0 0.034973 0.0389 0 0.94945 0.27324 0.075461 0.010379 4.5428 0.064763 7.8375e-05 0.82532 0.0055529 0.0062957 0.0013907 0.98689 0.99167 2.9994e-06 1.1997e-05 0.13417 0.92342 0.90521 0.0013994 0.9868 0.57257 0.0018853 0.42815 1.8152 1.8143 16.0063 144.9873 0.00018231 -85.6327 0.63136
1.7354 0.98803 5.5148e-05 3.8182 0.012027 2.2819e-05 0.0011545 0.18321 0.0006588 0.18386 0.16848 0 0.034971 0.0389 0 0.94954 0.27328 0.075476 0.010381 4.5434 0.064773 7.8389e-05 0.82531 0.0055534 0.0062963 0.0013907 0.98689 0.99167 2.9992e-06 1.1997e-05 0.13418 0.92361 0.90531 0.0013994 0.98686 0.57272 0.0018853 0.42816 1.8157 1.8149 16.0063 144.9873 0.00018217 -85.6329 0.63236
1.7364 0.98803 5.5147e-05 3.8182 0.012027 2.2832e-05 0.0011545 0.18325 0.0006588 0.1839 0.16852 0 0.034968 0.0389 0 0.94963 0.27332 0.07549 0.010382 4.544 0.064784 7.8403e-05 0.82529 0.005554 0.0062969 0.0013906 0.98689 0.99167 2.9991e-06 1.1996e-05 0.13418 0.9238 0.9054 0.0013994 0.98693 0.57287 0.0018852 0.42818 1.8163 1.8154 16.0063 144.9873 0.00018202 -85.6332 0.63336
1.7374 0.98803 5.5147e-05 3.8182 0.012027 2.2846e-05 0.0011545 0.18329 0.0006588 0.18395 0.16856 0 0.034966 0.0389 0 0.94972 0.27336 0.075505 0.010384 4.5446 0.064795 7.8417e-05 0.82528 0.0055545 0.0062974 0.0013906 0.98689 0.99167 2.999e-06 1.1996e-05 0.13418 0.92398 0.90549 0.0013993 0.987 0.57301 0.0018852 0.42819 1.8169 1.816 16.0063 144.9874 0.00018188 -85.6334 0.63436
1.7384 0.98803 5.5147e-05 3.8182 0.012027 2.2859e-05 0.0011545 0.18333 0.0006588 0.18399 0.1686 0 0.034963 0.0389 0 0.94981 0.2734 0.075519 0.010386 4.5452 0.064805 7.8431e-05 0.82527 0.0055551 0.006298 0.0013905 0.98689 0.99167 2.9988e-06 1.1995e-05 0.13419 0.92417 0.90558 0.0013993 0.98706 0.57316 0.0018851 0.4282 1.8174 1.8165 16.0063 144.9874 0.00018174 -85.6337 0.63536
1.7394 0.98803 5.5147e-05 3.8182 0.012027 2.2872e-05 0.0011545 0.18338 0.0006588 0.18403 0.16864 0 0.034961 0.0389 0 0.9499 0.27344 0.075534 0.010387 4.5459 0.064816 7.8445e-05 0.82526 0.0055556 0.0062986 0.0013904 0.98689 0.99167 2.9987e-06 1.1995e-05 0.13419 0.92435 0.90567 0.0013993 0.98713 0.57331 0.0018851 0.42821 1.818 1.8171 16.0062 144.9874 0.0001816 -85.6339 0.63636
1.7404 0.98803 5.5147e-05 3.8182 0.012027 2.2885e-05 0.0011545 0.18342 0.0006588 0.18407 0.16868 0 0.034958 0.0389 0 0.94999 0.27348 0.075548 0.010389 4.5465 0.064827 7.8459e-05 0.82525 0.0055562 0.0062991 0.0013904 0.98689 0.99167 2.9986e-06 1.1994e-05 0.1342 0.92454 0.90576 0.0013993 0.98719 0.57346 0.0018851 0.42823 1.8185 1.8176 16.0062 144.9874 0.00018146 -85.6342 0.63736
1.7414 0.98803 5.5147e-05 3.8182 0.012027 2.2898e-05 0.0011545 0.18346 0.00065881 0.18411 0.16871 0 0.034956 0.0389 0 0.95008 0.27352 0.075563 0.010391 4.5471 0.064838 7.8473e-05 0.82524 0.0055568 0.0062997 0.0013903 0.98689 0.99167 2.9984e-06 1.1994e-05 0.1342 0.92472 0.90585 0.0013992 0.98726 0.57361 0.001885 0.42824 1.8191 1.8182 16.0062 144.9874 0.00018132 -85.6344 0.63836
1.7424 0.98803 5.5147e-05 3.8182 0.012027 2.2911e-05 0.0011545 0.1835 0.00065881 0.18415 0.16875 0 0.034954 0.0389 0 0.95017 0.27356 0.075577 0.010393 4.5477 0.064848 7.8487e-05 0.82523 0.0055573 0.0063003 0.0013903 0.98689 0.99167 2.9983e-06 1.1993e-05 0.13421 0.92491 0.90594 0.0013992 0.98732 0.57376 0.001885 0.42825 1.8196 1.8188 16.0062 144.9875 0.00018117 -85.6347 0.63936
1.7434 0.98803 5.5147e-05 3.8182 0.012027 2.2924e-05 0.0011545 0.18354 0.00065881 0.1842 0.16879 0 0.034951 0.0389 0 0.95026 0.2736 0.075592 0.010394 4.5483 0.064859 7.8501e-05 0.82522 0.0055579 0.0063009 0.0013902 0.98689 0.99167 2.9982e-06 1.1993e-05 0.13421 0.92509 0.90603 0.0013992 0.98739 0.57391 0.0018849 0.42827 1.8202 1.8193 16.0061 144.9875 0.00018104 -85.6349 0.64036
1.7444 0.98803 5.5147e-05 3.8182 0.012027 2.2937e-05 0.0011545 0.18358 0.00065881 0.18424 0.16883 0 0.034949 0.0389 0 0.95035 0.27364 0.075606 0.010396 4.549 0.06487 7.8515e-05 0.82521 0.0055584 0.0063014 0.0013902 0.98689 0.99167 2.998e-06 1.1992e-05 0.13422 0.92527 0.90612 0.0013991 0.98745 0.57405 0.0018849 0.42828 1.8207 1.8199 16.0061 144.9875 0.0001809 -85.6352 0.64136
1.7454 0.98803 5.5147e-05 3.8182 0.012027 2.295e-05 0.0011545 0.18363 0.00065881 0.18428 0.16887 0 0.034946 0.0389 0 0.95044 0.27368 0.075621 0.010398 4.5496 0.064881 7.8529e-05 0.8252 0.005559 0.006302 0.0013901 0.98689 0.99167 2.9979e-06 1.1992e-05 0.13422 0.92545 0.9062 0.0013991 0.98751 0.5742 0.0018849 0.42829 1.8213 1.8204 16.0061 144.9875 0.00018076 -85.6354 0.64236
1.7464 0.98803 5.5147e-05 3.8182 0.012027 2.2964e-05 0.0011545 0.18367 0.00065881 0.18432 0.16891 0 0.034944 0.0389 0 0.95053 0.27372 0.075635 0.010399 4.5502 0.064891 7.8543e-05 0.82519 0.0055595 0.0063026 0.00139 0.98689 0.99167 2.9978e-06 1.1991e-05 0.13423 0.92564 0.90629 0.0013991 0.98758 0.57435 0.0018848 0.4283 1.8218 1.8209 16.0061 144.9875 0.00018062 -85.6356 0.64336
1.7474 0.98804 5.5147e-05 3.8182 0.012027 2.2977e-05 0.0011545 0.18371 0.00065881 0.18436 0.16895 0 0.034942 0.0389 0 0.95062 0.27376 0.07565 0.010401 4.5508 0.064902 7.8557e-05 0.82518 0.0055601 0.0063031 0.00139 0.9869 0.99167 2.9977e-06 1.1991e-05 0.13423 0.92582 0.90638 0.001399 0.98764 0.5745 0.0018848 0.42832 1.8223 1.8215 16.006 144.9876 0.00018048 -85.6359 0.64436
1.7484 0.98804 5.5147e-05 3.8182 0.012027 2.299e-05 0.0011545 0.18375 0.00065881 0.1844 0.16899 0 0.034939 0.0389 0 0.95071 0.2738 0.075664 0.010403 4.5514 0.064913 7.8571e-05 0.82517 0.0055607 0.0063037 0.0013899 0.9869 0.99167 2.9975e-06 1.199e-05 0.13424 0.926 0.90647 0.001399 0.9877 0.57465 0.0018847 0.42833 1.8229 1.822 16.006 144.9876 0.00018034 -85.6361 0.64536
1.7494 0.98804 5.5147e-05 3.8182 0.012026 2.3003e-05 0.0011545 0.18379 0.00065881 0.18445 0.16903 0 0.034937 0.0389 0 0.9508 0.27384 0.075679 0.010405 4.5521 0.064924 7.8585e-05 0.82516 0.0055612 0.0063043 0.0013899 0.9869 0.99167 2.9974e-06 1.199e-05 0.13424 0.92618 0.90655 0.001399 0.98776 0.57479 0.0018847 0.42834 1.8234 1.8226 16.006 144.9876 0.00018021 -85.6363 0.64636
1.7504 0.98804 5.5147e-05 3.8182 0.012026 2.3016e-05 0.0011545 0.18383 0.00065881 0.18449 0.16907 0 0.034934 0.0389 0 0.95089 0.27388 0.075693 0.010406 4.5527 0.064934 7.8599e-05 0.82514 0.0055618 0.0063049 0.0013898 0.9869 0.99167 2.9973e-06 1.1989e-05 0.13424 0.92636 0.90664 0.001399 0.98782 0.57494 0.0018847 0.42835 1.824 1.8231 16.006 144.9876 0.00018007 -85.6366 0.64736
1.7514 0.98804 5.5147e-05 3.8182 0.012026 2.3029e-05 0.0011545 0.18387 0.00065881 0.18453 0.16911 0 0.034932 0.0389 0 0.95098 0.27392 0.075708 0.010408 4.5533 0.064945 7.8613e-05 0.82513 0.0055623 0.0063054 0.0013898 0.9869 0.99167 2.9972e-06 1.1989e-05 0.13425 0.92653 0.90673 0.0013989 0.98789 0.57509 0.0018846 0.42837 1.8245 1.8237 16.006 144.9876 0.00017994 -85.6368 0.64836
1.7524 0.98804 5.5146e-05 3.8182 0.012026 2.3042e-05 0.0011545 0.18392 0.00065881 0.18457 0.16915 0 0.03493 0.0389 0 0.95107 0.27396 0.075722 0.01041 4.5539 0.064956 7.8627e-05 0.82512 0.0055629 0.006306 0.0013897 0.9869 0.99167 2.997e-06 1.1988e-05 0.13425 0.92671 0.90681 0.0013989 0.98795 0.57524 0.0018846 0.42838 1.825 1.8242 16.0059 144.9877 0.0001798 -85.637 0.64936
1.7534 0.98804 5.5146e-05 3.8182 0.012026 2.3055e-05 0.0011545 0.18396 0.00065881 0.18461 0.16918 0 0.034927 0.0389 0 0.95116 0.274 0.075737 0.010412 4.5545 0.064966 7.8641e-05 0.82511 0.0055634 0.0063066 0.0013897 0.9869 0.99168 2.9969e-06 1.1988e-05 0.13426 0.92689 0.9069 0.0013989 0.98801 0.57539 0.0018846 0.42839 1.8256 1.8247 16.0059 144.9877 0.00017966 -85.6373 0.65036
1.7544 0.98804 5.5146e-05 3.8182 0.012026 2.3068e-05 0.0011545 0.184 0.00065881 0.18465 0.16922 0 0.034925 0.0389 0 0.95125 0.27404 0.075751 0.010413 4.5552 0.064977 7.8655e-05 0.8251 0.005564 0.0063072 0.0013896 0.9869 0.99168 2.9968e-06 1.1987e-05 0.13426 0.92707 0.90698 0.0013988 0.98806 0.57553 0.0018845 0.4284 1.8261 1.8253 16.0059 144.9877 0.00017953 -85.6375 0.65136
1.7554 0.98804 5.5146e-05 3.8182 0.012026 2.3082e-05 0.0011545 0.18404 0.00065881 0.18469 0.16926 0 0.034922 0.0389 0 0.95134 0.27409 0.075766 0.010415 4.5558 0.064988 7.8669e-05 0.82509 0.0055646 0.0063077 0.0013896 0.9869 0.99168 2.9967e-06 1.1987e-05 0.13427 0.92724 0.90707 0.0013988 0.98812 0.57568 0.0018845 0.42842 1.8266 1.8258 16.0059 144.9877 0.0001794 -85.6377 0.65236
1.7564 0.98804 5.5146e-05 3.8182 0.012026 2.3095e-05 0.0011545 0.18408 0.00065881 0.18474 0.1693 0 0.03492 0.0389 0 0.95143 0.27413 0.075781 0.010417 4.5564 0.064999 7.8683e-05 0.82508 0.0055651 0.0063083 0.0013895 0.9869 0.99168 2.9966e-06 1.1986e-05 0.13427 0.92742 0.90715 0.0013988 0.98818 0.57583 0.0018845 0.42843 1.8272 1.8263 16.0058 144.9877 0.00017926 -85.6379 0.65336
1.7574 0.98804 5.5146e-05 3.8182 0.012026 2.3108e-05 0.0011545 0.18412 0.00065881 0.18478 0.16934 0 0.034918 0.0389 0 0.95152 0.27417 0.075795 0.010418 4.557 0.065009 7.8697e-05 0.82507 0.0055657 0.0063089 0.0013895 0.9869 0.99168 2.9965e-06 1.1986e-05 0.13428 0.9276 0.90724 0.0013988 0.98824 0.57598 0.0018844 0.42844 1.8277 1.8269 16.0058 144.9878 0.00017913 -85.6382 0.65436
1.7584 0.98804 5.5146e-05 3.8182 0.012026 2.3121e-05 0.0011545 0.18416 0.00065881 0.18482 0.16938 0 0.034915 0.0389 0 0.95161 0.27421 0.07581 0.01042 4.5577 0.06502 7.8711e-05 0.82506 0.0055662 0.0063095 0.0013894 0.9869 0.99168 2.9963e-06 1.1985e-05 0.13428 0.92777 0.90732 0.0013987 0.9883 0.57612 0.0018844 0.42845 1.8282 1.8274 16.0058 144.9878 0.000179 -85.6384 0.65536
1.7594 0.98804 5.5146e-05 3.8182 0.012026 2.3134e-05 0.0011545 0.1842 0.00065881 0.18486 0.16942 0 0.034913 0.0389 0 0.9517 0.27425 0.075824 0.010422 4.5583 0.065031 7.8726e-05 0.82505 0.0055668 0.0063101 0.0013894 0.9869 0.99168 2.9962e-06 1.1985e-05 0.13429 0.92794 0.90741 0.0013987 0.98836 0.57627 0.0018844 0.42847 1.8288 1.8279 16.0058 144.9878 0.00017887 -85.6386 0.65636
1.7604 0.98804 5.5146e-05 3.8182 0.012026 2.3147e-05 0.0011545 0.18425 0.00065882 0.1849 0.16946 0 0.034911 0.0389 0 0.95179 0.27429 0.075839 0.010424 4.5589 0.065042 7.8739e-05 0.82504 0.0055674 0.0063106 0.0013893 0.9869 0.99168 2.9961e-06 1.1984e-05 0.13429 0.92812 0.90749 0.0013987 0.98841 0.57642 0.0018843 0.42848 1.8293 1.8285 16.0057 144.9878 0.00017873 -85.6388 0.65736
1.7614 0.98804 5.5146e-05 3.8182 0.012026 2.316e-05 0.0011545 0.18429 0.00065882 0.18494 0.16949 0 0.034908 0.0389 0 0.95188 0.27433 0.075853 0.010425 4.5596 0.065052 7.8753e-05 0.82503 0.0055679 0.0063112 0.0013893 0.98691 0.99168 2.996e-06 1.1984e-05 0.1343 0.92829 0.90758 0.0013987 0.98847 0.57657 0.0018843 0.42849 1.8298 1.829 16.0057 144.9878 0.0001786 -85.639 0.65836
1.7624 0.98804 5.5146e-05 3.8182 0.012026 2.3173e-05 0.0011545 0.18433 0.00065882 0.18498 0.16953 0 0.034906 0.0389 0 0.95197 0.27437 0.075868 0.010427 4.5602 0.065063 7.8768e-05 0.82502 0.0055685 0.0063118 0.0013892 0.98691 0.99168 2.9959e-06 1.1983e-05 0.1343 0.92846 0.90766 0.0013986 0.98853 0.57671 0.0018842 0.42851 1.8303 1.8295 16.0057 144.9879 0.00017847 -85.6392 0.65936
1.7634 0.98804 5.5146e-05 3.8182 0.012026 2.3186e-05 0.0011545 0.18437 0.00065882 0.18502 0.16957 0 0.034903 0.0389 0 0.95206 0.27441 0.075882 0.010429 4.5608 0.065074 7.8782e-05 0.825 0.005569 0.0063124 0.0013892 0.98691 0.99168 2.9958e-06 1.1983e-05 0.1343 0.92864 0.90774 0.0013986 0.98858 0.57686 0.0018842 0.42852 1.8309 1.8301 16.0057 144.9879 0.00017834 -85.6395 0.66036
1.7644 0.98804 5.5146e-05 3.8182 0.012026 2.32e-05 0.0011545 0.18441 0.00065882 0.18506 0.16961 0 0.034901 0.0389 0 0.95215 0.27445 0.075897 0.010431 4.5614 0.065085 7.8796e-05 0.82499 0.0055696 0.0063129 0.0013891 0.98691 0.99168 2.9957e-06 1.1983e-05 0.13431 0.92881 0.90782 0.0013986 0.98864 0.57701 0.0018842 0.42853 1.8314 1.8306 16.0056 144.9879 0.00017821 -85.6397 0.66136
1.7654 0.98804 5.5146e-05 3.8182 0.012026 2.3213e-05 0.0011545 0.18445 0.00065882 0.1851 0.16965 0 0.034899 0.0389 0 0.95224 0.27449 0.075912 0.010432 4.5621 0.065095 7.881e-05 0.82498 0.0055702 0.0063135 0.0013891 0.98691 0.99168 2.9955e-06 1.1982e-05 0.13431 0.92898 0.90791 0.0013986 0.9887 0.57715 0.0018841 0.42854 1.8319 1.8311 16.0056 144.9879 0.00017808 -85.6399 0.66236
1.7664 0.98804 5.5146e-05 3.8182 0.012026 2.3226e-05 0.0011545 0.18449 0.00065882 0.18515 0.16969 0 0.034896 0.0389 0 0.95233 0.27453 0.075926 0.010434 4.5627 0.065106 7.8824e-05 0.82497 0.0055707 0.0063141 0.001389 0.98691 0.99168 2.9954e-06 1.1982e-05 0.13432 0.92915 0.90799 0.0013985 0.98875 0.5773 0.0018841 0.42856 1.8324 1.8316 16.0056 144.9879 0.00017795 -85.6401 0.66336
1.7674 0.98804 5.5146e-05 3.8182 0.012026 2.3239e-05 0.0011545 0.18453 0.00065882 0.18519 0.16973 0 0.034894 0.0389 0 0.95242 0.27457 0.075941 0.010436 4.5633 0.065117 7.8838e-05 0.82496 0.0055713 0.0063147 0.001389 0.98691 0.99168 2.9953e-06 1.1981e-05 0.13432 0.92932 0.90807 0.0013985 0.98881 0.57745 0.0018841 0.42857 1.833 1.8321 16.0056 144.988 0.00017783 -85.6403 0.66436
1.7684 0.98804 5.5145e-05 3.8182 0.012026 2.3252e-05 0.0011545 0.18457 0.00065882 0.18523 0.16976 0 0.034892 0.0389 0 0.95251 0.27461 0.075955 0.010437 4.564 0.065128 7.8852e-05 0.82495 0.0055719 0.0063153 0.0013889 0.98691 0.99168 2.9952e-06 1.1981e-05 0.13433 0.92949 0.90815 0.0013985 0.98886 0.5776 0.001884 0.42858 1.8335 1.8327 16.0055 144.988 0.0001777 -85.6405 0.66536
1.7694 0.98804 5.5145e-05 3.8182 0.012026 2.3265e-05 0.0011545 0.18461 0.00065882 0.18527 0.1698 0 0.034889 0.0389 0 0.9526 0.27465 0.07597 0.010439 4.5646 0.065139 7.8866e-05 0.82494 0.0055724 0.0063158 0.0013889 0.98691 0.99168 2.9951e-06 1.198e-05 0.13433 0.92966 0.90823 0.0013985 0.98891 0.57774 0.001884 0.42859 1.834 1.8332 16.0055 144.988 0.00017757 -85.6407 0.66636
1.7704 0.98804 5.5145e-05 3.8182 0.012026 2.3278e-05 0.0011545 0.18465 0.00065882 0.18531 0.16984 0 0.034887 0.0389 0 0.95269 0.27469 0.075984 0.010441 4.5652 0.065149 7.888e-05 0.82493 0.005573 0.0063164 0.0013888 0.98691 0.99168 2.995e-06 1.198e-05 0.13434 0.92982 0.90831 0.0013984 0.98897 0.57789 0.001884 0.42861 1.8345 1.8337 16.0055 144.988 0.00017744 -85.6409 0.66736
1.7714 0.98804 5.5145e-05 3.8182 0.012026 2.3291e-05 0.0011545 0.1847 0.00065882 0.18535 0.16988 0 0.034885 0.0389 0 0.95278 0.27473 0.075999 0.010443 4.5658 0.06516 7.8894e-05 0.82492 0.0055735 0.006317 0.0013888 0.98691 0.99168 2.9949e-06 1.1979e-05 0.13434 0.92999 0.90839 0.0013984 0.98902 0.57804 0.0018839 0.42862 1.835 1.8342 16.0055 144.988 0.00017732 -85.6411 0.66836
1.7724 0.98804 5.5145e-05 3.8182 0.012026 2.3304e-05 0.0011545 0.18474 0.00065882 0.18539 0.16992 0 0.034882 0.0389 0 0.95288 0.27477 0.076014 0.010444 4.5665 0.065171 7.8908e-05 0.82491 0.0055741 0.0063176 0.0013887 0.98691 0.99168 2.9948e-06 1.1979e-05 0.13435 0.93016 0.90847 0.0013984 0.98907 0.57818 0.0018839 0.42863 1.8355 1.8347 16.0054 144.9881 0.00017719 -85.6413 0.66936
1.7734 0.98804 5.5145e-05 3.8182 0.012026 2.3317e-05 0.0011545 0.18478 0.00065882 0.18543 0.16996 0 0.03488 0.0389 0 0.95297 0.27481 0.076028 0.010446 4.5671 0.065182 7.8922e-05 0.8249 0.0055747 0.0063182 0.0013887 0.98691 0.99168 2.9947e-06 1.1979e-05 0.13435 0.93033 0.90855 0.0013984 0.98913 0.57833 0.0018839 0.42864 1.8361 1.8353 16.0054 144.9881 0.00017707 -85.6415 0.67036
1.7744 0.98804 5.5145e-05 3.8182 0.012026 2.3331e-05 0.0011545 0.18482 0.00065882 0.18547 0.16999 0 0.034878 0.0389 0 0.95306 0.27485 0.076043 0.010448 4.5677 0.065192 7.8936e-05 0.82489 0.0055752 0.0063187 0.0013886 0.98691 0.99168 2.9946e-06 1.1978e-05 0.13436 0.93049 0.90863 0.0013983 0.98918 0.57848 0.0018839 0.42866 1.8366 1.8358 16.0054 144.9881 0.00017694 -85.6417 0.67136
1.7754 0.98804 5.5145e-05 3.8182 0.012026 2.3344e-05 0.0011545 0.18486 0.00065882 0.18551 0.17003 0 0.034875 0.0389 0 0.95315 0.27489 0.076057 0.01045 4.5684 0.065203 7.895e-05 0.82488 0.0055758 0.0063193 0.0013886 0.98691 0.99168 2.9945e-06 1.1978e-05 0.13436 0.93066 0.90871 0.0013983 0.98923 0.57862 0.0018838 0.42867 1.8371 1.8363 16.0054 144.9881 0.00017682 -85.6419 0.67236
1.7764 0.98804 5.5145e-05 3.8182 0.012026 2.3357e-05 0.0011545 0.1849 0.00065882 0.18555 0.17007 0 0.034873 0.0389 0 0.95324 0.27494 0.076072 0.010451 4.569 0.065214 7.8964e-05 0.82487 0.0055764 0.0063199 0.0013885 0.98691 0.99168 2.9944e-06 1.1977e-05 0.13436 0.93082 0.90879 0.0013983 0.98928 0.57877 0.0018838 0.42868 1.8376 1.8368 16.0053 144.9881 0.00017669 -85.6421 0.67336
1.7774 0.98804 5.5145e-05 3.8182 0.012026 2.337e-05 0.0011545 0.18494 0.00065882 0.18559 0.17011 0 0.03487 0.0389 0 0.95333 0.27498 0.076087 0.010453 4.5697 0.065225 7.8978e-05 0.82485 0.0055769 0.0063205 0.0013885 0.98691 0.99169 2.9943e-06 1.1977e-05 0.13437 0.93099 0.90887 0.0013983 0.98933 0.57892 0.0018838 0.42869 1.8381 1.8373 16.0053 144.9882 0.00017657 -85.6423 0.67436
1.7784 0.98804 5.5145e-05 3.8182 0.012026 2.3383e-05 0.0011545 0.18498 0.00065882 0.18563 0.17015 0 0.034868 0.0389 0 0.95342 0.27502 0.076101 0.010455 4.5703 0.065235 7.8993e-05 0.82484 0.0055775 0.0063211 0.0013885 0.98692 0.99169 2.9942e-06 1.1977e-05 0.13437 0.93115 0.90895 0.0013982 0.98938 0.57906 0.0018837 0.42871 1.8386 1.8378 16.0053 144.9882 0.00017644 -85.6425 0.67536
1.7794 0.98804 5.5145e-05 3.8182 0.012026 2.3396e-05 0.0011545 0.18502 0.00065883 0.18567 0.17019 0 0.034866 0.0389 0 0.95351 0.27506 0.076116 0.010456 4.5709 0.065246 7.9007e-05 0.82483 0.0055781 0.0063216 0.0013884 0.98692 0.99169 2.9941e-06 1.1976e-05 0.13438 0.93132 0.90903 0.0013982 0.98944 0.57921 0.0018837 0.42872 1.8391 1.8383 16.0053 144.9882 0.00017632 -85.6427 0.67636
1.7804 0.98804 5.5145e-05 3.8182 0.012026 2.3409e-05 0.0011545 0.18506 0.00065883 0.18571 0.17022 0 0.034863 0.0389 0 0.9536 0.2751 0.07613 0.010458 4.5716 0.065257 7.9021e-05 0.82482 0.0055786 0.0063222 0.0013884 0.98692 0.99169 2.994e-06 1.1976e-05 0.13438 0.93148 0.90911 0.0013982 0.98949 0.57936 0.0018837 0.42873 1.8396 1.8388 16.0052 144.9882 0.0001762 -85.6429 0.67736
1.7814 0.98804 5.5145e-05 3.8182 0.012026 2.3422e-05 0.0011545 0.1851 0.00065883 0.18576 0.17026 0 0.034861 0.0389 0 0.95369 0.27514 0.076145 0.01046 4.5722 0.065268 7.9035e-05 0.82481 0.0055792 0.0063228 0.0013883 0.98692 0.99169 2.9939e-06 1.1975e-05 0.13439 0.93164 0.90918 0.0013982 0.98954 0.5795 0.0018836 0.42874 1.8401 1.8393 16.0052 144.9882 0.00017608 -85.6431 0.67836
1.7824 0.98804 5.5145e-05 3.8182 0.012026 2.3435e-05 0.0011545 0.18514 0.00065883 0.1858 0.1703 0 0.034859 0.0389 0 0.95378 0.27518 0.07616 0.010462 4.5728 0.065279 7.9049e-05 0.8248 0.0055797 0.0063234 0.0013883 0.98692 0.99169 2.9938e-06 1.1975e-05 0.13439 0.9318 0.90926 0.0013981 0.98959 0.57965 0.0018836 0.42876 1.8406 1.8398 16.0052 144.9883 0.00017595 -85.6432 0.67936
1.7834 0.98804 5.5144e-05 3.8182 0.012026 2.3449e-05 0.0011545 0.18518 0.00065883 0.18584 0.17034 0 0.034857 0.0389 0 0.95387 0.27522 0.076174 0.010463 4.5735 0.065289 7.9063e-05 0.82479 0.0055803 0.006324 0.0013882 0.98692 0.99169 2.9937e-06 1.1975e-05 0.1344 0.93197 0.90934 0.0013981 0.98963 0.57979 0.0018836 0.42877 1.8411 1.8403 16.0052 144.9883 0.00017583 -85.6434 0.68036
1.7844 0.98804 5.5144e-05 3.8182 0.012026 2.3462e-05 0.0011545 0.18522 0.00065883 0.18588 0.17038 0 0.034854 0.0389 0 0.95396 0.27526 0.076189 0.010465 4.5741 0.0653 7.9077e-05 0.82478 0.0055809 0.0063246 0.0013882 0.98692 0.99169 2.9936e-06 1.1974e-05 0.1344 0.93213 0.90942 0.0013981 0.98968 0.57994 0.0018835 0.42878 1.8416 1.8408 16.0051 144.9883 0.00017571 -85.6436 0.68136
1.7854 0.98804 5.5144e-05 3.8182 0.012026 2.3475e-05 0.0011545 0.18526 0.00065883 0.18592 0.17041 0 0.034852 0.0389 0 0.95405 0.2753 0.076203 0.010467 4.5747 0.065311 7.9091e-05 0.82477 0.0055814 0.0063251 0.0013882 0.98692 0.99169 2.9935e-06 1.1974e-05 0.13441 0.93229 0.90949 0.0013981 0.98973 0.58009 0.0018835 0.42879 1.8421 1.8413 16.0051 144.9883 0.00017559 -85.6438 0.68236
1.7864 0.98804 5.5144e-05 3.8182 0.012026 2.3488e-05 0.0011545 0.1853 0.00065883 0.18596 0.17045 0 0.03485 0.0389 0 0.95414 0.27534 0.076218 0.010469 4.5754 0.065322 7.9105e-05 0.82476 0.005582 0.0063257 0.0013881 0.98692 0.99169 2.9934e-06 1.1973e-05 0.13441 0.93245 0.90957 0.0013981 0.98978 0.58023 0.0018835 0.42881 1.8426 1.8418 16.0051 144.9884 0.00017547 -85.644 0.68336
1.7874 0.98804 5.5144e-05 3.8182 0.012026 2.3501e-05 0.0011545 0.18534 0.00065883 0.186 0.17049 0 0.034847 0.0389 0 0.95423 0.27538 0.076233 0.01047 4.576 0.065333 7.9119e-05 0.82475 0.0055826 0.0063263 0.0013881 0.98692 0.99169 2.9933e-06 1.1973e-05 0.13442 0.93261 0.90965 0.001398 0.98983 0.58038 0.0018835 0.42882 1.8431 1.8423 16.0051 144.9884 0.00017535 -85.6442 0.68436
1.7884 0.98804 5.5144e-05 3.8182 0.012026 2.3514e-05 0.0011545 0.18538 0.00065883 0.18604 0.17053 0 0.034845 0.0389 0 0.95432 0.27542 0.076247 0.010472 4.5767 0.065343 7.9133e-05 0.82474 0.0055831 0.0063269 0.001388 0.98692 0.99169 2.9932e-06 1.1973e-05 0.13442 0.93277 0.90972 0.001398 0.98988 0.58053 0.0018834 0.42883 1.8436 1.8428 16.005 144.9884 0.00017523 -85.6443 0.68536
1.7894 0.98804 5.5144e-05 3.8182 0.012026 2.3527e-05 0.0011545 0.18542 0.00065883 0.18608 0.17057 0 0.034843 0.0389 0 0.95441 0.27546 0.076262 0.010474 4.5773 0.065354 7.9147e-05 0.82473 0.0055837 0.0063275 0.001388 0.98692 0.99169 2.9931e-06 1.1972e-05 0.13443 0.93293 0.9098 0.001398 0.98992 0.58067 0.0018834 0.42884 1.8441 1.8433 16.005 144.9884 0.00017511 -85.6445 0.68636
1.7904 0.98804 5.5144e-05 3.8182 0.012026 2.354e-05 0.0011545 0.18546 0.00065883 0.18612 0.1706 0 0.03484 0.0389 0 0.9545 0.2755 0.076277 0.010475 4.5779 0.065365 7.9162e-05 0.82471 0.0055843 0.0063281 0.0013879 0.98692 0.99169 2.993e-06 1.1972e-05 0.13443 0.93308 0.90987 0.001398 0.98997 0.58082 0.0018834 0.42886 1.8446 1.8438 16.005 144.9884 0.00017499 -85.6447 0.68736
1.7914 0.98804 5.5144e-05 3.8182 0.012026 2.3553e-05 0.0011545 0.1855 0.00065883 0.18616 0.17064 0 0.034838 0.0389 0 0.95459 0.27554 0.076291 0.010477 4.5786 0.065376 7.9176e-05 0.8247 0.0055849 0.0063286 0.0013879 0.98692 0.99169 2.9929e-06 1.1971e-05 0.13444 0.93324 0.90995 0.0013979 0.99002 0.58096 0.0018833 0.42887 1.8451 1.8443 16.005 144.9885 0.00017488 -85.6449 0.68836
1.7924 0.98804 5.5144e-05 3.8182 0.012026 2.3567e-05 0.0011545 0.18554 0.00065883 0.1862 0.17068 0 0.034836 0.0389 0 0.95468 0.27559 0.076306 0.010479 4.5792 0.065386 7.919e-05 0.82469 0.0055854 0.0063292 0.0013879 0.98692 0.99169 2.9928e-06 1.1971e-05 0.13444 0.9334 0.91002 0.0013979 0.99006 0.58111 0.0018833 0.42888 1.8456 1.8448 16.0049 144.9885 0.00017476 -85.6451 0.68936
1.7934 0.98804 5.5144e-05 3.8182 0.012026 2.358e-05 0.0011545 0.18558 0.00065883 0.18624 0.17072 0 0.034833 0.0389 0 0.95478 0.27563 0.07632 0.010481 4.5799 0.065397 7.9204e-05 0.82468 0.005586 0.0063298 0.0013878 0.98692 0.99169 2.9927e-06 1.1971e-05 0.13444 0.93355 0.9101 0.0013979 0.99011 0.58125 0.0018833 0.42889 1.8461 1.8453 16.0049 144.9885 0.00017464 -85.6452 0.69036
1.7944 0.98804 5.5144e-05 3.8182 0.012026 2.3593e-05 0.0011545 0.18562 0.00065883 0.18628 0.17075 0 0.034831 0.0389 0 0.95487 0.27567 0.076335 0.010482 4.5805 0.065408 7.9218e-05 0.82467 0.0055866 0.0063304 0.0013878 0.98692 0.99169 2.9926e-06 1.197e-05 0.13445 0.93371 0.91017 0.0013979 0.99016 0.5814 0.0018833 0.42891 1.8466 1.8458 16.0049 144.9885 0.00017453 -85.6454 0.69136
1.7954 0.98804 5.5144e-05 3.8182 0.012026 2.3606e-05 0.0011545 0.18566 0.00065883 0.18632 0.17079 0 0.034829 0.0389 0 0.95496 0.27571 0.07635 0.010484 4.5811 0.065419 7.9232e-05 0.82466 0.0055871 0.006331 0.0013877 0.98692 0.99169 2.9925e-06 1.197e-05 0.13445 0.93387 0.91025 0.0013979 0.9902 0.58155 0.0018832 0.42892 1.8471 1.8463 16.0049 144.9885 0.00017441 -85.6456 0.69236
1.7964 0.98804 5.5144e-05 3.8182 0.012026 2.3619e-05 0.0011545 0.1857 0.00065883 0.18636 0.17083 0 0.034826 0.0389 0 0.95505 0.27575 0.076364 0.010486 4.5818 0.06543 7.9246e-05 0.82465 0.0055877 0.0063316 0.0013877 0.98693 0.99169 2.9924e-06 1.197e-05 0.13446 0.93402 0.91032 0.0013978 0.99025 0.58169 0.0018832 0.42893 1.8475 1.8468 16.0048 144.9886 0.00017429 -85.6457 0.69336
1.7974 0.98804 5.5144e-05 3.8182 0.012026 2.3632e-05 0.0011545 0.18574 0.00065883 0.1864 0.17087 0 0.034824 0.0389 0 0.95514 0.27579 0.076379 0.010488 4.5824 0.06544 7.9261e-05 0.82464 0.0055883 0.0063322 0.0013877 0.98693 0.99169 2.9923e-06 1.1969e-05 0.13446 0.93418 0.91039 0.0013978 0.99029 0.58184 0.0018832 0.42894 1.848 1.8473 16.0048 144.9886 0.00017418 -85.6459 0.69436
1.7984 0.98804 5.5144e-05 3.8182 0.012026 2.3645e-05 0.0011545 0.18578 0.00065883 0.18644 0.1709 0 0.034822 0.0389 0 0.95523 0.27583 0.076394 0.010489 4.5831 0.065451 7.9275e-05 0.82463 0.0055888 0.0063328 0.0013876 0.98693 0.99169 2.9923e-06 1.1969e-05 0.13447 0.93433 0.91047 0.0013978 0.99034 0.58198 0.0018832 0.42896 1.8485 1.8478 16.0048 144.9886 0.00017406 -85.6461 0.69536
1.7994 0.98804 5.5143e-05 3.8182 0.012026 2.3658e-05 0.0011545 0.18582 0.00065884 0.18648 0.17094 0 0.03482 0.0389 0 0.95532 0.27587 0.076408 0.010491 4.5837 0.065462 7.9289e-05 0.82462 0.0055894 0.0063333 0.0013876 0.98693 0.99169 2.9922e-06 1.1969e-05 0.13447 0.93448 0.91054 0.0013978 0.99038 0.58213 0.0018831 0.42897 1.849 1.8483 16.0048 144.9886 0.00017395 -85.6462 0.69636
1.8004 0.98804 5.5143e-05 3.8182 0.012026 2.3671e-05 0.0011545 0.18586 0.00065884 0.18652 0.17098 0 0.034817 0.0389 0 0.95541 0.27591 0.076423 0.010493 4.5844 0.065473 7.9303e-05 0.82461 0.00559 0.0063339 0.0013876 0.98693 0.99169 2.9921e-06 1.1968e-05 0.13448 0.93464 0.91061 0.0013978 0.99043 0.58227 0.0018831 0.42898 1.8495 1.8487 16.0047 144.9886 0.00017383 -85.6464 0.69736
1.8014 0.98804 5.5143e-05 3.8182 0.012026 2.3685e-05 0.0011545 0.1859 0.00065884 0.18656 0.17102 0 0.034815 0.0389 0 0.9555 0.27595 0.076438 0.010495 4.585 0.065484 7.9317e-05 0.8246 0.0055905 0.0063345 0.0013875 0.98693 0.99169 2.992e-06 1.1968e-05 0.13448 0.93479 0.91069 0.0013977 0.99047 0.58242 0.0018831 0.42899 1.85 1.8492 16.0047 144.9887 0.00017372 -85.6466 0.69836
1.8024 0.98804 5.5143e-05 3.8182 0.012026 2.3698e-05 0.0011545 0.18594 0.00065884 0.1866 0.17105 0 0.034813 0.0389 0 0.95559 0.27599 0.076452 0.010496 4.5857 0.065494 7.9331e-05 0.82458 0.0055911 0.0063351 0.0013875 0.98693 0.99169 2.9919e-06 1.1968e-05 0.13449 0.93494 0.91076 0.0013977 0.99051 0.58256 0.001883 0.42901 1.8505 1.8497 16.0047 144.9887 0.00017361 -85.6467 0.69936
1.8034 0.98804 5.5143e-05 3.8182 0.012026 2.3711e-05 0.0011545 0.18598 0.00065884 0.18664 0.17109 0 0.03481 0.0389 0 0.95568 0.27603 0.076467 0.010498 4.5863 0.065505 7.9345e-05 0.82457 0.0055917 0.0063357 0.0013874 0.98693 0.99169 2.9918e-06 1.1967e-05 0.13449 0.93509 0.91083 0.0013977 0.99056 0.58271 0.001883 0.42902 1.8509 1.8502 16.0047 144.9887 0.00017349 -85.6469 0.70036
1.8044 0.98804 5.5143e-05 3.8182 0.012026 2.3724e-05 0.0011545 0.18602 0.00065884 0.18668 0.17113 0 0.034808 0.0389 0 0.95577 0.27607 0.076482 0.0105 4.587 0.065516 7.9359e-05 0.82456 0.0055923 0.0063363 0.0013874 0.98693 0.99169 2.9917e-06 1.1967e-05 0.1345 0.93525 0.9109 0.0013977 0.9906 0.58285 0.001883 0.42903 1.8514 1.8507 16.0046 144.9887 0.00017338 -85.6471 0.70136
1.8054 0.98804 5.5143e-05 3.8182 0.012026 2.3737e-05 0.0011545 0.18606 0.00065884 0.18672 0.17117 0 0.034806 0.0389 0 0.95586 0.27611 0.076496 0.010501 4.5876 0.065527 7.9373e-05 0.82455 0.0055928 0.0063369 0.0013874 0.98693 0.99169 2.9917e-06 1.1967e-05 0.1345 0.9354 0.91097 0.0013977 0.99064 0.583 0.001883 0.42904 1.8519 1.8512 16.0046 144.9887 0.00017327 -85.6472 0.70236
1.8064 0.98804 5.5143e-05 3.8182 0.012026 2.375e-05 0.0011545 0.1861 0.00065884 0.18675 0.1712 0 0.034804 0.0389 0 0.95595 0.27616 0.076511 0.010503 4.5882 0.065538 7.9388e-05 0.82454 0.0055934 0.0063375 0.0013873 0.98693 0.99169 2.9916e-06 1.1966e-05 0.13451 0.93555 0.91104 0.0013976 0.99069 0.58315 0.0018829 0.42906 1.8524 1.8516 16.0046 144.9888 0.00017315 -85.6474 0.70336
1.8074 0.98804 5.5143e-05 3.8182 0.012026 2.3763e-05 0.0011546 0.18614 0.00065884 0.18679 0.17124 0 0.034801 0.0389 0 0.95605 0.2762 0.076526 0.010505 4.5889 0.065549 7.9402e-05 0.82453 0.005594 0.006338 0.0013873 0.98693 0.9917 2.9915e-06 1.1966e-05 0.13451 0.9357 0.91112 0.0013976 0.99073 0.58329 0.0018829 0.42907 1.8529 1.8521 16.0046 144.9888 0.00017304 -85.6475 0.70436
1.8084 0.98804 5.5143e-05 3.8182 0.012026 2.3776e-05 0.0011546 0.18618 0.00065884 0.18683 0.17128 0 0.034799 0.0389 0 0.95614 0.27624 0.07654 0.010507 4.5895 0.065559 7.9416e-05 0.82452 0.0055945 0.0063386 0.0013873 0.98693 0.9917 2.9914e-06 1.1966e-05 0.13452 0.93585 0.91119 0.0013976 0.99077 0.58344 0.0018829 0.42908 1.8533 1.8526 16.0045 144.9888 0.00017293 -85.6477 0.70536
1.8094 0.98804 5.5143e-05 3.8182 0.012026 2.3789e-05 0.0011546 0.18622 0.00065884 0.18687 0.17132 0 0.034797 0.0389 0 0.95623 0.27628 0.076555 0.010508 4.5902 0.06557 7.943e-05 0.82451 0.0055951 0.0063392 0.0013872 0.98693 0.9917 2.9913e-06 1.1965e-05 0.13452 0.936 0.91126 0.0013976 0.99081 0.58358 0.0018829 0.42909 1.8538 1.8531 16.0045 144.9888 0.00017282 -85.6479 0.70636
1.8104 0.98804 5.5143e-05 3.8182 0.012026 2.3803e-05 0.0011546 0.18626 0.00065884 0.18691 0.17135 0 0.034795 0.0389 0 0.95632 0.27632 0.07657 0.01051 4.5908 0.065581 7.9444e-05 0.8245 0.0055957 0.0063398 0.0013872 0.98693 0.9917 2.9912e-06 1.1965e-05 0.13452 0.93614 0.91133 0.0013976 0.99085 0.58372 0.0018828 0.42911 1.8543 1.8535 16.0045 144.9888 0.00017271 -85.648 0.70736
1.8114 0.98804 5.5143e-05 3.8182 0.012026 2.3816e-05 0.0011546 0.1863 0.00065884 0.18695 0.17139 0 0.034792 0.0389 0 0.95641 0.27636 0.076584 0.010512 4.5915 0.065592 7.9458e-05 0.82449 0.0055963 0.0063404 0.0013871 0.98693 0.9917 2.9912e-06 1.1965e-05 0.13453 0.93629 0.9114 0.0013975 0.99089 0.58387 0.0018828 0.42912 1.8547 1.854 16.0044 144.9889 0.0001726 -85.6482 0.70836
1.8124 0.98804 5.5143e-05 3.8182 0.012026 2.3829e-05 0.0011546 0.18634 0.00065884 0.18699 0.17143 0 0.03479 0.0389 0 0.9565 0.2764 0.076599 0.010514 4.5921 0.065603 7.9472e-05 0.82448 0.0055968 0.006341 0.0013871 0.98693 0.9917 2.9911e-06 1.1964e-05 0.13453 0.93644 0.91147 0.0013975 0.99093 0.58401 0.0018828 0.42913 1.8552 1.8545 16.0044 144.9889 0.00017249 -85.6483 0.70936
1.8134 0.98804 5.5143e-05 3.8182 0.012026 2.3842e-05 0.0011546 0.18638 0.00065884 0.18703 0.17146 0 0.034788 0.0389 0 0.95659 0.27644 0.076614 0.010515 4.5928 0.065613 7.9487e-05 0.82447 0.0055974 0.0063416 0.0013871 0.98693 0.9917 2.991e-06 1.1964e-05 0.13454 0.93659 0.91154 0.0013975 0.99098 0.58416 0.0018828 0.42914 1.8557 1.855 16.0044 144.9889 0.00017238 -85.6485 0.71036
1.8144 0.98804 5.5142e-05 3.8182 0.012026 2.3855e-05 0.0011546 0.18642 0.00065884 0.18707 0.1715 0 0.034786 0.0389 0 0.95668 0.27648 0.076628 0.010517 4.5934 0.065624 7.9501e-05 0.82446 0.005598 0.0063422 0.001387 0.98693 0.9917 2.9909e-06 1.1964e-05 0.13454 0.93673 0.91161 0.0013975 0.99102 0.5843 0.0018827 0.42916 1.8562 1.8554 16.0044 144.9889 0.00017227 -85.6486 0.71136
1.8154 0.98804 5.5142e-05 3.8182 0.012026 2.3868e-05 0.0011546 0.18646 0.00065884 0.18711 0.17154 0 0.034783 0.0389 0 0.95677 0.27652 0.076643 0.010519 4.5941 0.065635 7.9515e-05 0.82444 0.0055986 0.0063428 0.001387 0.98693 0.9917 2.9908e-06 1.1963e-05 0.13455 0.93688 0.91168 0.0013975 0.99106 0.58445 0.0018827 0.42917 1.8566 1.8559 16.0043 144.9889 0.00017216 -85.6488 0.71236
1.8164 0.98804 5.5142e-05 3.8182 0.012026 2.3881e-05 0.0011546 0.1865 0.00065884 0.18715 0.17158 0 0.034781 0.0389 0 0.95686 0.27656 0.076658 0.010521 4.5947 0.065646 7.9529e-05 0.82443 0.0055991 0.0063434 0.001387 0.98693 0.9917 2.9908e-06 1.1963e-05 0.13455 0.93703 0.91174 0.0013974 0.9911 0.58459 0.0018827 0.42918 1.8571 1.8564 16.0043 144.989 0.00017206 -85.6489 0.71336
1.8174 0.98804 5.5142e-05 3.8182 0.012026 2.3894e-05 0.0011546 0.18653 0.00065884 0.18719 0.17161 0 0.034779 0.0389 0 0.95695 0.2766 0.076672 0.010522 4.5954 0.065657 7.9543e-05 0.82442 0.0055997 0.006344 0.0013869 0.98693 0.9917 2.9907e-06 1.1963e-05 0.13456 0.93717 0.91181 0.0013974 0.99113 0.58474 0.0018827 0.42919 1.8576 1.8568 16.0043 144.989 0.00017195 -85.6491 0.71436
1.8184 0.98804 5.5142e-05 3.8182 0.012026 2.3907e-05 0.0011546 0.18657 0.00065884 0.18723 0.17165 0 0.034777 0.0389 0 0.95705 0.27665 0.076687 0.010524 4.5961 0.065668 7.9557e-05 0.82441 0.0056003 0.0063446 0.0013869 0.98694 0.9917 2.9906e-06 1.1962e-05 0.13456 0.93732 0.91188 0.0013974 0.99117 0.58488 0.0018827 0.4292 1.858 1.8573 16.0043 144.989 0.00017184 -85.6492 0.71536
1.8194 0.98804 5.5142e-05 3.8182 0.012026 2.392e-05 0.0011546 0.18661 0.00065885 0.18727 0.17169 0 0.034774 0.0389 0 0.95714 0.27669 0.076702 0.010526 4.5967 0.065678 7.9571e-05 0.8244 0.0056009 0.0063451 0.0013869 0.98694 0.9917 2.9905e-06 1.1962e-05 0.13457 0.93746 0.91195 0.0013974 0.99121 0.58503 0.0018826 0.42922 1.8585 1.8578 16.0042 144.989 0.00017173 -85.6494 0.71636
1.8204 0.98804 5.5142e-05 3.8182 0.012026 2.3934e-05 0.0011546 0.18665 0.00065885 0.18731 0.17172 0 0.034772 0.0389 0 0.95723 0.27673 0.076716 0.010527 4.5974 0.065689 7.9586e-05 0.82439 0.0056014 0.0063457 0.0013868 0.98694 0.9917 2.9904e-06 1.1962e-05 0.13457 0.9376 0.91202 0.0013974 0.99125 0.58517 0.0018826 0.42923 1.859 1.8582 16.0042 144.989 0.00017163 -85.6495 0.71736
1.8214 0.98804 5.5142e-05 3.8182 0.012025 2.3947e-05 0.0011546 0.18669 0.00065885 0.18735 0.17176 0 0.03477 0.0389 0 0.95732 0.27677 0.076731 0.010529 4.598 0.0657 7.96e-05 0.82438 0.005602 0.0063463 0.0013868 0.98694 0.9917 2.9904e-06 1.1961e-05 0.13458 0.93775 0.91208 0.0013974 0.99129 0.58532 0.0018826 0.42924 1.8594 1.8587 16.0042 144.9891 0.00017152 -85.6496 0.71836
1.8224 0.98804 5.5142e-05 3.8182 0.012025 2.396e-05 0.0011546 0.18673 0.00065885 0.18738 0.1718 0 0.034768 0.0389 0 0.95741 0.27681 0.076746 0.010531 4.5987 0.065711 7.9614e-05 0.82437 0.0056026 0.0063469 0.0013868 0.98694 0.9917 2.9903e-06 1.1961e-05 0.13458 0.93789 0.91215 0.0013973 0.99133 0.58546 0.0018826 0.42925 1.8599 1.8592 16.0042 144.9891 0.00017141 -85.6498 0.71936
1.8234 0.98804 5.5142e-05 3.8182 0.012025 2.3973e-05 0.0011546 0.18677 0.00065885 0.18742 0.17183 0 0.034765 0.0389 0 0.9575 0.27685 0.076761 0.010533 4.5993 0.065722 7.9628e-05 0.82436 0.0056032 0.0063475 0.0013867 0.98694 0.9917 2.9902e-06 1.1961e-05 0.13459 0.93803 0.91222 0.0013973 0.99137 0.5856 0.0018825 0.42927 1.8603 1.8596 16.0041 144.9891 0.00017131 -85.6499 0.72036
1.8244 0.98804 5.5142e-05 3.8182 0.012025 2.3986e-05 0.0011546 0.18681 0.00065885 0.18746 0.17187 0 0.034763 0.0389 0 0.95759 0.27689 0.076775 0.010534 4.6 0.065733 7.9642e-05 0.82435 0.0056037 0.0063481 0.0013867 0.98694 0.9917 2.9901e-06 1.196e-05 0.13459 0.93818 0.91229 0.0013973 0.9914 0.58575 0.0018825 0.42928 1.8608 1.8601 16.0041 144.9891 0.0001712 -85.6501 0.72136
1.8254 0.98804 5.5142e-05 3.8182 0.012025 2.3999e-05 0.0011546 0.18685 0.00065885 0.1875 0.17191 0 0.034761 0.0389 0 0.95768 0.27693 0.07679 0.010536 4.6006 0.065743 7.9656e-05 0.82434 0.0056043 0.0063487 0.0013867 0.98694 0.9917 2.9901e-06 1.196e-05 0.1346 0.93832 0.91235 0.0013973 0.99144 0.58589 0.0018825 0.42929 1.8613 1.8606 16.0041 144.9891 0.0001711 -85.6502 0.72236
1.8264 0.98804 5.5142e-05 3.8182 0.012025 2.4012e-05 0.0011546 0.18689 0.00065885 0.18754 0.17194 0 0.034759 0.0389 0 0.95777 0.27697 0.076805 0.010538 4.6013 0.065754 7.9671e-05 0.82433 0.0056049 0.0063493 0.0013866 0.98694 0.9917 2.99e-06 1.196e-05 0.1346 0.93846 0.91242 0.0013973 0.99148 0.58604 0.0018825 0.4293 1.8617 1.861 16.004 144.9892 0.00017099 -85.6504 0.72336
1.8274 0.98804 5.5142e-05 3.8182 0.012025 2.4025e-05 0.0011546 0.18693 0.00065885 0.18758 0.17198 0 0.034756 0.0389 0 0.95786 0.27701 0.076819 0.01054 4.602 0.065765 7.9685e-05 0.82431 0.0056055 0.0063499 0.0013866 0.98694 0.9917 2.9899e-06 1.196e-05 0.13461 0.9386 0.91249 0.0013973 0.99152 0.58618 0.0018824 0.42932 1.8622 1.8615 16.004 144.9892 0.00017089 -85.6505 0.72436
1.8284 0.98804 5.5142e-05 3.8182 0.012025 2.4038e-05 0.0011546 0.18696 0.00065885 0.18762 0.17202 0 0.034754 0.0389 0 0.95796 0.27705 0.076834 0.010541 4.6026 0.065776 7.9699e-05 0.8243 0.005606 0.0063505 0.0013866 0.98694 0.9917 2.9899e-06 1.1959e-05 0.13461 0.93874 0.91255 0.0013972 0.99155 0.58632 0.0018824 0.42933 1.8626 1.8619 16.004 144.9892 0.00017079 -85.6506 0.72536
1.8294 0.98804 5.5141e-05 3.8182 0.012025 2.4052e-05 0.0011546 0.187 0.00065885 0.18766 0.17205 0 0.034752 0.0389 0 0.95805 0.2771 0.076849 0.010543 4.6033 0.065787 7.9713e-05 0.82429 0.0056066 0.0063511 0.0013865 0.98694 0.9917 2.9898e-06 1.1959e-05 0.13461 0.93888 0.91262 0.0013972 0.99159 0.58647 0.0018824 0.42934 1.8631 1.8624 16.004 144.9892 0.00017068 -85.6508 0.72636
1.8304 0.98804 5.5141e-05 3.8182 0.012025 2.4065e-05 0.0011546 0.18704 0.00065885 0.1877 0.17209 0 0.03475 0.0389 0 0.95814 0.27714 0.076864 0.010545 4.6039 0.065798 7.9727e-05 0.82428 0.0056072 0.0063517 0.0013865 0.98694 0.9917 2.9897e-06 1.1959e-05 0.13462 0.93902 0.91268 0.0013972 0.99163 0.58661 0.0018824 0.42935 1.8636 1.8629 16.0039 144.9892 0.00017058 -85.6509 0.72736
1.8314 0.98804 5.5141e-05 3.8182 0.012025 2.4078e-05 0.0011546 0.18708 0.00065885 0.18773 0.17213 0 0.034747 0.0389 0 0.95823 0.27718 0.076878 0.010547 4.6046 0.065808 7.9742e-05 0.82427 0.0056078 0.0063523 0.0013865 0.98694 0.9917 2.9896e-06 1.1958e-05 0.13462 0.93916 0.91275 0.0013972 0.99166 0.58676 0.0018824 0.42937 1.864 1.8633 16.0039 144.9893 0.00017048 -85.651 0.72836
1.8324 0.98804 5.5141e-05 3.8182 0.012025 2.4091e-05 0.0011546 0.18712 0.00065885 0.18777 0.17216 0 0.034745 0.0389 0 0.95832 0.27722 0.076893 0.010548 4.6052 0.065819 7.9756e-05 0.82426 0.0056083 0.0063529 0.0013865 0.98694 0.9917 2.9896e-06 1.1958e-05 0.13463 0.9393 0.91281 0.0013972 0.9917 0.5869 0.0018823 0.42938 1.8645 1.8638 16.0039 144.9893 0.00017037 -85.6512 0.72936
1.8334 0.98804 5.5141e-05 3.8182 0.012025 2.4104e-05 0.0011546 0.18716 0.00065885 0.18781 0.1722 0 0.034743 0.0389 0 0.95841 0.27726 0.076908 0.01055 4.6059 0.06583 7.977e-05 0.82425 0.0056089 0.0063535 0.0013864 0.98694 0.9917 2.9895e-06 1.1958e-05 0.13463 0.93944 0.91288 0.0013972 0.99173 0.58704 0.0018823 0.42939 1.8649 1.8642 16.0039 144.9893 0.00017027 -85.6513 0.73036
1.8344 0.98804 5.5141e-05 3.8182 0.012025 2.4117e-05 0.0011546 0.1872 0.00065885 0.18785 0.17224 0 0.034741 0.0389 0 0.9585 0.2773 0.076922 0.010552 4.6066 0.065841 7.9784e-05 0.82424 0.0056095 0.0063541 0.0013864 0.98694 0.9917 2.9894e-06 1.1958e-05 0.13464 0.93957 0.91294 0.0013971 0.99177 0.58719 0.0018823 0.4294 1.8654 1.8647 16.0038 144.9893 0.00017017 -85.6514 0.73136
1.8354 0.98804 5.5141e-05 3.8182 0.012025 2.413e-05 0.0011546 0.18724 0.00065885 0.18789 0.17227 0 0.034739 0.0389 0 0.95859 0.27734 0.076937 0.010554 4.6072 0.065852 7.9798e-05 0.82423 0.0056101 0.0063547 0.0013864 0.98694 0.9917 2.9894e-06 1.1957e-05 0.13464 0.93971 0.91301 0.0013971 0.9918 0.58733 0.0018823 0.42941 1.8658 1.8651 16.0038 144.9894 0.00017007 -85.6516 0.73236
1.8364 0.98804 5.5141e-05 3.8182 0.012025 2.4143e-05 0.0011546 0.18727 0.00065885 0.18793 0.17231 0 0.034736 0.0389 0 0.95868 0.27738 0.076952 0.010555 4.6079 0.065863 7.9812e-05 0.82422 0.0056107 0.0063553 0.0013863 0.98694 0.9917 2.9893e-06 1.1957e-05 0.13465 0.93985 0.91307 0.0013971 0.99184 0.58747 0.0018823 0.42943 1.8663 1.8656 16.0038 144.9894 0.00016997 -85.6517 0.73336
1.8374 0.98804 5.5141e-05 3.8182 0.012025 2.4156e-05 0.0011546 0.18731 0.00065885 0.18797 0.17235 0 0.034734 0.0389 0 0.95878 0.27742 0.076967 0.010557 4.6085 0.065873 7.9827e-05 0.82421 0.0056112 0.0063559 0.0013863 0.98694 0.9917 2.9892e-06 1.1957e-05 0.13465 0.93998 0.91314 0.0013971 0.99187 0.58762 0.0018822 0.42944 1.8667 1.866 16.0037 144.9894 0.00016987 -85.6518 0.73436
1.8384 0.98804 5.5141e-05 3.8182 0.012025 2.417e-05 0.0011546 0.18735 0.00065885 0.18801 0.17238 0 0.034732 0.0389 0 0.95887 0.27746 0.076981 0.010559 4.6092 0.065884 7.9841e-05 0.8242 0.0056118 0.0063565 0.0013863 0.98694 0.9917 2.9892e-06 1.1957e-05 0.13466 0.94012 0.9132 0.0013971 0.99191 0.58776 0.0018822 0.42945 1.8672 1.8665 16.0037 144.9894 0.00016977 -85.6519 0.73536
1.8394 0.98804 5.5141e-05 3.8182 0.012025 2.4183e-05 0.0011546 0.18739 0.00065885 0.18804 0.17242 0 0.03473 0.0389 0 0.95896 0.2775 0.076996 0.010561 4.6099 0.065895 7.9855e-05 0.82418 0.0056124 0.0063571 0.0013862 0.98694 0.9917 2.9891e-06 1.1956e-05 0.13466 0.94026 0.91326 0.0013971 0.99194 0.58791 0.0018822 0.42946 1.8676 1.8669 16.0037 144.9894 0.00016967 -85.6521 0.73636
1.8404 0.98804 5.5141e-05 3.8182 0.012025 2.4196e-05 0.0011546 0.18743 0.00065886 0.18808 0.17246 0 0.034728 0.0389 0 0.95905 0.27755 0.077011 0.010562 4.6105 0.065906 7.9869e-05 0.82417 0.005613 0.0063577 0.0013862 0.98694 0.9917 2.989e-06 1.1956e-05 0.13467 0.94039 0.91333 0.001397 0.99198 0.58805 0.0018822 0.42948 1.8681 1.8674 16.0037 144.9895 0.00016957 -85.6522 0.73736
1.8414 0.98804 5.5141e-05 3.8182 0.012025 2.4209e-05 0.0011546 0.18747 0.00065886 0.18812 0.17249 0 0.034725 0.0389 0 0.95914 0.27759 0.077026 0.010564 4.6112 0.065917 7.9883e-05 0.82416 0.0056136 0.0063583 0.0013862 0.98694 0.9917 2.989e-06 1.1956e-05 0.13467 0.94053 0.91339 0.001397 0.99201 0.58819 0.0018822 0.42949 1.8685 1.8678 16.0036 144.9895 0.00016947 -85.6523 0.73836
1.8424 0.98804 5.5141e-05 3.8182 0.012025 2.4222e-05 0.0011546 0.18751 0.00065886 0.18816 0.17253 0 0.034723 0.0389 0 0.95923 0.27763 0.07704 0.010566 4.6119 0.065928 7.9898e-05 0.82415 0.0056141 0.0063589 0.0013862 0.98695 0.9917 2.9889e-06 1.1955e-05 0.13468 0.94066 0.91345 0.001397 0.99204 0.58834 0.0018821 0.4295 1.8689 1.8683 16.0036 144.9895 0.00016937 -85.6525 0.73936
1.8434 0.98804 5.5141e-05 3.8182 0.012025 2.4235e-05 0.0011546 0.18754 0.00065886 0.1882 0.17256 0 0.034721 0.0389 0 0.95932 0.27767 0.077055 0.010567 4.6125 0.065939 7.9912e-05 0.82414 0.0056147 0.0063595 0.0013861 0.98695 0.9917 2.9888e-06 1.1955e-05 0.13468 0.94079 0.91352 0.001397 0.99208 0.58848 0.0018821 0.42951 1.8694 1.8687 16.0036 144.9895 0.00016927 -85.6526 0.74036
1.8444 0.98804 5.5141e-05 3.8182 0.012025 2.4248e-05 0.0011546 0.18758 0.00065886 0.18824 0.1726 0 0.034719 0.0389 0 0.95941 0.27771 0.07707 0.010569 4.6132 0.065949 7.9926e-05 0.82413 0.0056153 0.0063601 0.0013861 0.98695 0.99171 2.9888e-06 1.1955e-05 0.13469 0.94093 0.91358 0.001397 0.99211 0.58862 0.0018821 0.42952 1.8698 1.8691 16.0036 144.9895 0.00016917 -85.6527 0.74136
1.8454 0.98804 5.514e-05 3.8182 0.012025 2.4261e-05 0.0011546 0.18762 0.00065886 0.18827 0.17264 0 0.034717 0.0389 0 0.95951 0.27775 0.077085 0.010571 4.6139 0.06596 7.994e-05 0.82412 0.0056159 0.0063607 0.0013861 0.98695 0.99171 2.9887e-06 1.1955e-05 0.13469 0.94106 0.91364 0.001397 0.99214 0.58877 0.0018821 0.42954 1.8703 1.8696 16.0035 144.9896 0.00016907 -85.6528 0.74236
1.8464 0.98804 5.514e-05 3.8182 0.012025 2.4274e-05 0.0011546 0.18766 0.00065886 0.18831 0.17267 0 0.034714 0.0389 0 0.9596 0.27779 0.077099 0.010573 4.6145 0.065971 7.9954e-05 0.82411 0.0056165 0.0063613 0.001386 0.98695 0.99171 2.9886e-06 1.1954e-05 0.1347 0.94119 0.9137 0.001397 0.99218 0.58891 0.0018821 0.42955 1.8707 1.87 16.0035 144.9896 0.00016898 -85.6529 0.74336
1.8474 0.98804 5.514e-05 3.8182 0.012025 2.4287e-05 0.0011546 0.1877 0.00065886 0.18835 0.17271 0 0.034712 0.0389 0 0.95969 0.27783 0.077114 0.010574 4.6152 0.065982 7.9969e-05 0.8241 0.005617 0.0063619 0.001386 0.98695 0.99171 2.9886e-06 1.1954e-05 0.1347 0.94133 0.91377 0.0013969 0.99221 0.58905 0.001882 0.42956 1.8711 1.8705 16.0035 144.9896 0.00016888 -85.6531 0.74436
1.8484 0.98804 5.514e-05 3.8182 0.012025 2.4301e-05 0.0011546 0.18774 0.00065886 0.18839 0.17275 0 0.03471 0.0389 0 0.95978 0.27787 0.077129 0.010576 4.6159 0.065993 7.9983e-05 0.82409 0.0056176 0.0063625 0.001386 0.98695 0.99171 2.9885e-06 1.1954e-05 0.13471 0.94146 0.91383 0.0013969 0.99224 0.58919 0.001882 0.42957 1.8716 1.8709 16.0034 144.9896 0.00016878 -85.6532 0.74536
1.8494 0.98804 5.514e-05 3.8182 0.012025 2.4314e-05 0.0011546 0.18777 0.00065886 0.18843 0.17278 0 0.034708 0.0389 0 0.95987 0.27792 0.077144 0.010578 4.6165 0.066004 7.9997e-05 0.82408 0.0056182 0.0063631 0.001386 0.98695 0.99171 2.9884e-06 1.1954e-05 0.13471 0.94159 0.91389 0.0013969 0.99227 0.58934 0.001882 0.42959 1.872 1.8714 16.0034 144.9896 0.00016868 -85.6533 0.74636
1.8504 0.98804 5.514e-05 3.8182 0.012025 2.4327e-05 0.0011546 0.18781 0.00065886 0.18847 0.17282 0 0.034706 0.0389 0 0.95996 0.27796 0.077158 0.01058 4.6172 0.066015 8.0011e-05 0.82407 0.0056188 0.0063637 0.0013859 0.98695 0.99171 2.9884e-06 1.1953e-05 0.13472 0.94172 0.91395 0.0013969 0.99231 0.58948 0.001882 0.4296 1.8725 1.8718 16.0034 144.9897 0.00016859 -85.6534 0.74736
1.8514 0.98804 5.514e-05 3.8182 0.012025 2.434e-05 0.0011546 0.18785 0.00065886 0.1885 0.17285 0 0.034703 0.0389 0 0.96005 0.278 0.077173 0.010581 4.6179 0.066025 8.0026e-05 0.82405 0.0056194 0.0063643 0.0013859 0.98695 0.99171 2.9883e-06 1.1953e-05 0.13472 0.94185 0.91401 0.0013969 0.99234 0.58962 0.001882 0.42961 1.8729 1.8722 16.0034 144.9897 0.00016849 -85.6535 0.74836
1.8524 0.98804 5.514e-05 3.8182 0.012025 2.4353e-05 0.0011546 0.18789 0.00065886 0.18854 0.17289 0 0.034701 0.0389 0 0.96015 0.27804 0.077188 0.010583 4.6185 0.066036 8.004e-05 0.82404 0.00562 0.0063649 0.0013859 0.98695 0.99171 2.9883e-06 1.1953e-05 0.13472 0.94198 0.91407 0.0013969 0.99237 0.58977 0.0018819 0.42962 1.8733 1.8727 16.0033 144.9897 0.0001684 -85.6537 0.74936
1.8534 0.98804 5.514e-05 3.8182 0.012025 2.4366e-05 0.0011546 0.18793 0.00065886 0.18858 0.17293 0 0.034699 0.0389 0 0.96024 0.27808 0.077203 0.010585 4.6192 0.066047 8.0054e-05 0.82403 0.0056205 0.0063655 0.0013858 0.98695 0.99171 2.9882e-06 1.1953e-05 0.13473 0.94211 0.91413 0.0013969 0.9924 0.58991 0.0018819 0.42964 1.8738 1.8731 16.0033 144.9897 0.0001683 -85.6538 0.75036
1.8544 0.98804 5.514e-05 3.8182 0.012025 2.4379e-05 0.0011546 0.18796 0.00065886 0.18862 0.17296 0 0.034697 0.0389 0 0.96033 0.27812 0.077218 0.010587 4.6199 0.066058 8.0068e-05 0.82402 0.0056211 0.0063661 0.0013858 0.98695 0.99171 2.9881e-06 1.1952e-05 0.13473 0.94224 0.91419 0.0013968 0.99243 0.59005 0.0018819 0.42965 1.8742 1.8735 16.0033 144.9897 0.00016821 -85.6539 0.75136
1.8554 0.98804 5.514e-05 3.8182 0.012025 2.4392e-05 0.0011546 0.188 0.00065886 0.18866 0.173 0 0.034695 0.0389 0 0.96042 0.27816 0.077232 0.010588 4.6205 0.066069 8.0083e-05 0.82401 0.0056217 0.0063667 0.0013858 0.98695 0.99171 2.9881e-06 1.1952e-05 0.13474 0.94237 0.91425 0.0013968 0.99246 0.59019 0.0018819 0.42966 1.8746 1.874 16.0032 144.9898 0.00016811 -85.654 0.75236
1.8564 0.98804 5.514e-05 3.8182 0.012025 2.4405e-05 0.0011546 0.18804 0.00065886 0.1887 0.17303 0 0.034693 0.0389 0 0.96051 0.2782 0.077247 0.01059 4.6212 0.06608 8.0097e-05 0.824 0.0056223 0.0063673 0.0013858 0.98695 0.99171 2.988e-06 1.1952e-05 0.13474 0.9425 0.91431 0.0013968 0.99249 0.59034 0.0018819 0.42967 1.8751 1.8744 16.0032 144.9898 0.00016802 -85.6541 0.75336
1.8574 0.98804 5.514e-05 3.8182 0.012025 2.4419e-05 0.0011546 0.18808 0.00065886 0.18873 0.17307 0 0.03469 0.0389 0 0.9606 0.27824 0.077262 0.010592 4.6219 0.066091 8.0111e-05 0.82399 0.0056229 0.0063679 0.0013857 0.98695 0.99171 2.9879e-06 1.1952e-05 0.13475 0.94263 0.91437 0.0013968 0.99252 0.59048 0.0018819 0.42968 1.8755 1.8748 16.0032 144.9898 0.00016792 -85.6542 0.75436
1.8584 0.98804 5.514e-05 3.8182 0.012025 2.4432e-05 0.0011546 0.18812 0.00065886 0.18877 0.17311 0 0.034688 0.0389 0 0.96069 0.27828 0.077277 0.010594 4.6225 0.066102 8.0125e-05 0.82398 0.0056235 0.0063685 0.0013857 0.98695 0.99171 2.9879e-06 1.1951e-05 0.13475 0.94275 0.91443 0.0013968 0.99255 0.59062 0.0018818 0.4297 1.8759 1.8753 16.0032 144.9898 0.00016783 -85.6543 0.75536
1.8594 0.98804 5.514e-05 3.8182 0.012025 2.4445e-05 0.0011546 0.18815 0.00065886 0.18881 0.17314 0 0.034686 0.0389 0 0.96079 0.27833 0.077291 0.010595 4.6232 0.066112 8.0139e-05 0.82397 0.005624 0.0063691 0.0013857 0.98695 0.99171 2.9878e-06 1.1951e-05 0.13476 0.94288 0.91449 0.0013968 0.99258 0.59076 0.0018818 0.42971 1.8764 1.8757 16.0031 144.9898 0.00016774 -85.6544 0.75636
1.8604 0.98804 5.5139e-05 3.8182 0.012025 2.4458e-05 0.0011546 0.18819 0.00065886 0.18885 0.17318 0 0.034684 0.0389 0 0.96088 0.27837 0.077306 0.010597 4.6239 0.066123 8.0154e-05 0.82396 0.0056246 0.0063697 0.0013857 0.98695 0.99171 2.9878e-06 1.1951e-05 0.13476 0.94301 0.91455 0.0013968 0.99261 0.59091 0.0018818 0.42972 1.8768 1.8761 16.0031 144.9899 0.00016764 -85.6546 0.75736
1.8614 0.98804 5.5139e-05 3.8182 0.012025 2.4471e-05 0.0011546 0.18823 0.00065886 0.18888 0.17321 0 0.034682 0.0389 0 0.96097 0.27841 0.077321 0.010599 4.6246 0.066134 8.0168e-05 0.82395 0.0056252 0.0063703 0.0013856 0.98695 0.99171 2.9877e-06 1.1951e-05 0.13477 0.94314 0.91461 0.0013967 0.99264 0.59105 0.0018818 0.42973 1.8772 1.8766 16.0031 144.9899 0.00016755 -85.6547 0.75836
1.8624 0.98804 5.5139e-05 3.8182 0.012025 2.4484e-05 0.0011546 0.18827 0.00065887 0.18892 0.17325 0 0.03468 0.0389 0 0.96106 0.27845 0.077336 0.010601 4.6252 0.066145 8.0182e-05 0.82394 0.0056258 0.0063709 0.0013856 0.98695 0.99171 2.9877e-06 1.1951e-05 0.13477 0.94326 0.91467 0.0013967 0.99267 0.59119 0.0018818 0.42975 1.8776 1.877 16.0031 144.9899 0.00016746 -85.6548 0.75936
1.8634 0.98804 5.5139e-05 3.8182 0.012025 2.4497e-05 0.0011546 0.18831 0.00065887 0.18896 0.17328 0 0.034677 0.0389 0 0.96115 0.27849 0.077351 0.010602 4.6259 0.066156 8.0196e-05 0.82392 0.0056264 0.0063715 0.0013856 0.98695 0.99171 2.9876e-06 1.195e-05 0.13478 0.94339 0.91473 0.0013967 0.9927 0.59133 0.0018817 0.42976 1.8781 1.8774 16.003 144.9899 0.00016737 -85.6549 0.76036
1.8644 0.98804 5.5139e-05 3.8182 0.012025 2.451e-05 0.0011546 0.18834 0.00065887 0.189 0.17332 0 0.034675 0.0389 0 0.96124 0.27853 0.077365 0.010604 4.6266 0.066167 8.0211e-05 0.82391 0.005627 0.0063721 0.0013856 0.98695 0.99171 2.9875e-06 1.195e-05 0.13478 0.94351 0.91479 0.0013967 0.99273 0.59148 0.0018817 0.42977 1.8785 1.8778 16.003 144.9899 0.00016727 -85.655 0.76136
1.8654 0.98804 5.5139e-05 3.8182 0.012025 2.4523e-05 0.0011546 0.18838 0.00065887 0.18904 0.17335 0 0.034673 0.0389 0 0.96134 0.27857 0.07738 0.010606 4.6273 0.066178 8.0225e-05 0.8239 0.0056275 0.0063727 0.0013855 0.98695 0.99171 2.9875e-06 1.195e-05 0.13479 0.94364 0.91484 0.0013967 0.99276 0.59162 0.0018817 0.42978 1.8789 1.8783 16.003 144.99 0.00016718 -85.6551 0.76236
1.8664 0.98804 5.5139e-05 3.8182 0.012025 2.4537e-05 0.0011546 0.18842 0.00065887 0.18907 0.17339 0 0.034671 0.0389 0 0.96143 0.27861 0.077395 0.010608 4.6279 0.066189 8.0239e-05 0.82389 0.0056281 0.0063733 0.0013855 0.98695 0.99171 2.9874e-06 1.195e-05 0.13479 0.94376 0.9149 0.0013967 0.99279 0.59176 0.0018817 0.42979 1.8793 1.8787 16.0029 144.99 0.00016709 -85.6552 0.76336
1.8674 0.98804 5.5139e-05 3.8182 0.012025 2.455e-05 0.0011546 0.18846 0.00065887 0.18911 0.17343 0 0.034669 0.0389 0 0.96152 0.27866 0.07741 0.010609 4.6286 0.066199 8.0253e-05 0.82388 0.0056287 0.0063739 0.0013855 0.98695 0.99171 2.9874e-06 1.1949e-05 0.1348 0.94389 0.91496 0.0013967 0.99282 0.5919 0.0018817 0.42981 1.8798 1.8791 16.0029 144.99 0.000167 -85.6553 0.76436
1.8684 0.98804 5.5139e-05 3.8182 0.012025 2.4563e-05 0.0011546 0.18849 0.00065887 0.18915 0.17346 0 0.034667 0.0389 0 0.96161 0.2787 0.077425 0.010611 4.6293 0.06621 8.0268e-05 0.82387 0.0056293 0.0063745 0.0013855 0.98695 0.99171 2.9873e-06 1.1949e-05 0.1348 0.94401 0.91502 0.0013967 0.99285 0.59204 0.0018817 0.42982 1.8802 1.8795 16.0029 144.99 0.00016691 -85.6554 0.76536
1.8694 0.98804 5.5139e-05 3.8182 0.012025 2.4576e-05 0.0011546 0.18853 0.00065887 0.18919 0.1735 0 0.034665 0.0389 0 0.9617 0.27874 0.077439 0.010613 4.63 0.066221 8.0282e-05 0.82386 0.0056299 0.0063751 0.0013854 0.98695 0.99171 2.9873e-06 1.1949e-05 0.13481 0.94414 0.91508 0.0013966 0.99287 0.59219 0.0018816 0.42983 1.8806 1.88 16.0029 144.99 0.00016682 -85.6555 0.76636
1.8704 0.98804 5.5139e-05 3.8182 0.012025 2.4589e-05 0.0011546 0.18857 0.00065887 0.18922 0.17353 0 0.034662 0.0389 0 0.96179 0.27878 0.077454 0.010615 4.6306 0.066232 8.0296e-05 0.82385 0.0056305 0.0063757 0.0013854 0.98695 0.99171 2.9872e-06 1.1949e-05 0.13481 0.94426 0.91513 0.0013966 0.9929 0.59233 0.0018816 0.42984 1.881 1.8804 16.0028 144.9901 0.00016673 -85.6556 0.76736
1.8714 0.98804 5.5139e-05 3.8182 0.012025 2.4602e-05 0.0011546 0.18861 0.00065887 0.18926 0.17357 0 0.03466 0.0389 0 0.96189 0.27882 0.077469 0.010616 4.6313 0.066243 8.031e-05 0.82384 0.0056311 0.0063763 0.0013854 0.98695 0.99171 2.9872e-06 1.1949e-05 0.13482 0.94438 0.91519 0.0013966 0.99293 0.59247 0.0018816 0.42985 1.8814 1.8808 16.0028 144.9901 0.00016664 -85.6557 0.76836
1.8724 0.98804 5.5139e-05 3.8182 0.012025 2.4615e-05 0.0011546 0.18865 0.00065887 0.1893 0.1736 0 0.034658 0.0389 0 0.96198 0.27886 0.077484 0.010618 4.632 0.066254 8.0325e-05 0.82383 0.0056317 0.0063769 0.0013854 0.98696 0.99171 2.9871e-06 1.1948e-05 0.13482 0.9445 0.91525 0.0013966 0.99296 0.59261 0.0018816 0.42987 1.8819 1.8812 16.0028 144.9901 0.00016655 -85.6558 0.76936
1.8734 0.98804 5.5139e-05 3.8182 0.012025 2.4628e-05 0.0011546 0.18868 0.00065887 0.18934 0.17364 0 0.034656 0.0389 0 0.96207 0.2789 0.077499 0.01062 4.6327 0.066265 8.0339e-05 0.82382 0.0056322 0.0063775 0.0013854 0.98696 0.99171 2.9871e-06 1.1948e-05 0.13483 0.94463 0.9153 0.0013966 0.99298 0.59275 0.0018816 0.42988 1.8823 1.8816 16.0027 144.9901 0.00016646 -85.6559 0.77036
1.8744 0.98804 5.5139e-05 3.8182 0.012025 2.4641e-05 0.0011546 0.18872 0.00065887 0.18937 0.17367 0 0.034654 0.0389 0 0.96216 0.27894 0.077514 0.010621 4.6333 0.066276 8.0353e-05 0.8238 0.0056328 0.0063782 0.0013853 0.98696 0.99171 2.987e-06 1.1948e-05 0.13483 0.94475 0.91536 0.0013966 0.99301 0.5929 0.0018816 0.42989 1.8827 1.8821 16.0027 144.9901 0.00016637 -85.656 0.77136
1.8754 0.98804 5.5139e-05 3.8182 0.012025 2.4654e-05 0.0011546 0.18876 0.00065887 0.18941 0.17371 0 0.034652 0.0389 0 0.96225 0.27898 0.077528 0.010623 4.634 0.066287 8.0367e-05 0.82379 0.0056334 0.0063788 0.0013853 0.98696 0.99171 2.9869e-06 1.1948e-05 0.13484 0.94487 0.91542 0.0013966 0.99304 0.59304 0.0018815 0.4299 1.8831 1.8825 16.0027 144.9902 0.00016628 -85.6561 0.77236
1.8764 0.98804 5.5138e-05 3.8182 0.012025 2.4668e-05 0.0011546 0.1888 0.00065887 0.18945 0.17374 0 0.03465 0.0389 0 0.96234 0.27903 0.077543 0.010625 4.6347 0.066297 8.0382e-05 0.82378 0.005634 0.0063794 0.0013853 0.98696 0.99171 2.9869e-06 1.1947e-05 0.13484 0.94499 0.91547 0.0013966 0.99307 0.59318 0.0018815 0.42992 1.8835 1.8829 16.0027 144.9902 0.0001662 -85.6562 0.77336
1.8774 0.98804 5.5138e-05 3.8182 0.012025 2.4681e-05 0.0011546 0.18883 0.00065887 0.18949 0.17378 0 0.034647 0.0389 0 0.96244 0.27907 0.077558 0.010627 4.6354 0.066308 8.0396e-05 0.82377 0.0056346 0.00638 0.0013853 0.98696 0.99171 2.9868e-06 1.1947e-05 0.13485 0.94511 0.91553 0.0013965 0.99309 0.59332 0.0018815 0.42993 1.8839 1.8833 16.0026 144.9902 0.00016611 -85.6563 0.77436
1.8784 0.98804 5.5138e-05 3.8182 0.012025 2.4694e-05 0.0011546 0.18887 0.00065887 0.18952 0.17382 0 0.034645 0.0389 0 0.96253 0.27911 0.077573 0.010628 4.6361 0.066319 8.041e-05 0.82376 0.0056352 0.0063806 0.0013852 0.98696 0.99171 2.9868e-06 1.1947e-05 0.13485 0.94523 0.91558 0.0013965 0.99312 0.59346 0.0018815 0.42994 1.8844 1.8837 16.0026 144.9902 0.00016602 -85.6564 0.77536
1.8794 0.98804 5.5138e-05 3.8182 0.012025 2.4707e-05 0.0011546 0.18891 0.00065887 0.18956 0.17385 0 0.034643 0.0389 0 0.96262 0.27915 0.077588 0.01063 4.6367 0.06633 8.0425e-05 0.82375 0.0056358 0.0063812 0.0013852 0.98696 0.99171 2.9867e-06 1.1947e-05 0.13486 0.94535 0.91564 0.0013965 0.99315 0.5936 0.0018815 0.42995 1.8848 1.8841 16.0026 144.9903 0.00016593 -85.6565 0.77636
1.8804 0.98804 5.5138e-05 3.8182 0.012025 2.472e-05 0.0011546 0.18894 0.00065887 0.1896 0.17389 0 0.034641 0.0389 0 0.96271 0.27919 0.077603 0.010632 4.6374 0.066341 8.044e-05 0.82374 0.0056364 0.0063818 0.0013852 0.98696 0.99171 2.9867e-06 1.1947e-05 0.13486 0.94547 0.91569 0.0013965 0.99317 0.59374 0.0018815 0.42996 1.8852 1.8846 16.0025 144.9903 0.00016585 -85.6566 0.77736
1.8814 0.98804 5.5138e-05 3.8182 0.012025 2.4733e-05 0.0011546 0.18898 0.00065887 0.18964 0.17392 0 0.034639 0.0389 0 0.9628 0.27923 0.077617 0.010634 4.6381 0.066352 8.0452e-05 0.82373 0.0056369 0.0063824 0.0013852 0.98696 0.99171 2.9866e-06 1.1946e-05 0.13486 0.94559 0.91575 0.0013965 0.9932 0.59389 0.0018815 0.42998 1.8856 1.885 16.0025 144.9903 0.00016576 -85.6567 0.77836
1.8824 0.98804 5.5138e-05 3.8182 0.012025 2.4746e-05 0.0011546 0.18902 0.00065887 0.18967 0.17396 0 0.034637 0.0389 0 0.96289 0.27927 0.077632 0.010635 4.6388 0.066363 8.0466e-05 0.82372 0.0056375 0.006383 0.0013851 0.98696 0.99171 2.9866e-06 1.1946e-05 0.13487 0.94571 0.9158 0.0013965 0.99322 0.59403 0.0018814 0.42999 1.886 1.8854 16.0025 144.9903 0.00016567 -85.6568 0.77936
1.8834 0.98804 5.5138e-05 3.8182 0.012025 2.4759e-05 0.0011546 0.18906 0.00065887 0.18971 0.17399 0 0.034635 0.0389 0 0.96299 0.27932 0.077647 0.010637 4.6395 0.066374 8.0484e-05 0.82371 0.0056381 0.0063836 0.0013851 0.98696 0.99171 2.9865e-06 1.1946e-05 0.13487 0.94582 0.91586 0.0013965 0.99325 0.59417 0.0018814 0.43 1.8864 1.8858 16.0024 144.9903 0.00016559 -85.6569 0.78036
1.8844 0.98804 5.5138e-05 3.8182 0.012025 2.4772e-05 0.0011546 0.18909 0.00065888 0.18975 0.17403 0 0.034633 0.0389 0 0.96308 0.27936 0.077662 0.010639 4.6401 0.066385 8.0496e-05 0.8237 0.0056387 0.0063842 0.0013851 0.98696 0.99171 2.9865e-06 1.1946e-05 0.13488 0.94594 0.91591 0.0013965 0.99327 0.59431 0.0018814 0.43001 1.8868 1.8862 16.0024 144.9904 0.0001655 -85.657 0.78136
1.8854 0.98804 5.5138e-05 3.8182 0.012025 2.4786e-05 0.0011546 0.18913 0.00065888 0.18979 0.17406 0 0.03463 0.0389 0 0.96317 0.2794 0.077677 0.010641 4.6408 0.066396 8.0508e-05 0.82368 0.0056393 0.0063848 0.0013851 0.98696 0.99171 2.9864e-06 1.1946e-05 0.13488 0.94606 0.91597 0.0013965 0.9933 0.59445 0.0018814 0.43002 1.8872 1.8866 16.0024 144.9904 0.00016542 -85.6571 0.78236
1.8864 0.98804 5.5138e-05 3.8182 0.012025 2.4799e-05 0.0011546 0.18917 0.00065888 0.18982 0.1741 0 0.034628 0.0389 0 0.96326 0.27944 0.077692 0.010642 4.6415 0.066406 8.0526e-05 0.82367 0.0056399 0.0063855 0.0013851 0.98696 0.99171 2.9864e-06 1.1945e-05 0.13489 0.94618 0.91602 0.0013964 0.99333 0.59459 0.0018814 0.43004 1.8876 1.887 16.0024 144.9904 0.00016533 -85.6572 0.78336
1.8874 0.98804 5.5138e-05 3.8182 0.012025 2.4812e-05 0.0011546 0.18921 0.00065888 0.18986 0.17413 0 0.034626 0.0389 0 0.96335 0.27948 0.077706 0.010644 4.6422 0.066417 8.054e-05 0.82366 0.0056405 0.0063861 0.001385 0.98696 0.99171 2.9863e-06 1.1945e-05 0.13489 0.94629 0.91608 0.0013964 0.99335 0.59473 0.0018814 0.43005 1.888 1.8874 16.0023 144.9904 0.00016524 -85.6573 0.78436
1.8884 0.98804 5.5138e-05 3.8182 0.012025 2.4825e-05 0.0011546 0.18924 0.00065888 0.1899 0.17417 0 0.034624 0.0389 0 0.96345 0.27952 0.077721 0.010646 4.6429 0.066428 8.0551e-05 0.82365 0.0056411 0.0063867 0.001385 0.98696 0.99171 2.9863e-06 1.1945e-05 0.1349 0.94641 0.91613 0.0013964 0.99338 0.59487 0.0018814 0.43006 1.8884 1.8878 16.0023 144.9904 0.00016516 -85.6574 0.78536
1.8894 0.98804 5.5138e-05 3.8182 0.012025 2.4838e-05 0.0011546 0.18928 0.00065888 0.18993 0.1742 0 0.034622 0.0389 0 0.96354 0.27956 0.077736 0.010648 4.6436 0.066439 8.0568e-05 0.82364 0.0056417 0.0063873 0.001385 0.98696 0.99171 2.9862e-06 1.1945e-05 0.1349 0.94653 0.91618 0.0013964 0.9934 0.59502 0.0018813 0.43007 1.8889 1.8882 16.0023 144.9905 0.00016508 -85.6574 0.78636
1.8904 0.98804 5.5138e-05 3.8182 0.012025 2.4851e-05 0.0011546 0.18932 0.00065888 0.18997 0.17424 0 0.03462 0.0389 0 0.96363 0.2796 0.077751 0.010649 4.6443 0.06645 8.0582e-05 0.82363 0.0056423 0.0063879 0.001385 0.98696 0.99171 2.9862e-06 1.1945e-05 0.13491 0.94664 0.91624 0.0013964 0.99342 0.59516 0.0018813 0.43008 1.8893 1.8886 16.0022 144.9905 0.00016499 -85.6575 0.78736
1.8914 0.98804 5.5137e-05 3.8182 0.012025 2.4864e-05 0.0011546 0.18935 0.00065888 0.19001 0.17427 0 0.034618 0.0389 0 0.96372 0.27965 0.077766 0.010651 4.6449 0.066461 8.0596e-05 0.82362 0.0056429 0.0063885 0.001385 0.98696 0.99171 2.9862e-06 1.1945e-05 0.13491 0.94676 0.91629 0.0013964 0.99345 0.5953 0.0018813 0.4301 1.8897 1.889 16.0022 144.9905 0.00016491 -85.6576 0.78836
1.8924 0.98804 5.5137e-05 3.8182 0.012025 2.4877e-05 0.0011546 0.18939 0.00065888 0.19004 0.17431 0 0.034616 0.0389 0 0.96381 0.27969 0.077781 0.010653 4.6456 0.066472 8.061e-05 0.82361 0.0056434 0.0063891 0.0013849 0.98696 0.99171 2.9861e-06 1.1944e-05 0.13492 0.94687 0.91634 0.0013964 0.99347 0.59544 0.0018813 0.43011 1.8901 1.8895 16.0022 144.9905 0.00016482 -85.6577 0.78936
1.8934 0.98804 5.5137e-05 3.8182 0.012024 2.489e-05 0.0011546 0.18943 0.00065888 0.19008 0.17434 0 0.034614 0.0389 0 0.9639 0.27973 0.077796 0.010655 4.6463 0.066483 8.0625e-05 0.8236 0.005644 0.0063897 0.0013849 0.98696 0.99171 2.9861e-06 1.1944e-05 0.13492 0.94699 0.9164 0.0013964 0.9935 0.59558 0.0018813 0.43012 1.8905 1.8899 16.0022 144.9905 0.00016474 -85.6578 0.79036
1.8944 0.98804 5.5137e-05 3.8182 0.012024 2.4903e-05 0.0011546 0.18946 0.00065888 0.19012 0.17438 0 0.034612 0.0389 0 0.964 0.27977 0.07781 0.010656 4.647 0.066494 8.0639e-05 0.82359 0.0056446 0.0063903 0.0013849 0.98696 0.99172 2.986e-06 1.1944e-05 0.13493 0.9471 0.91645 0.0013964 0.99352 0.59572 0.0018813 0.43013 1.8909 1.8903 16.0021 144.9906 0.00016466 -85.6579 0.79136
1.8954 0.98804 5.5137e-05 3.8182 0.012024 2.4917e-05 0.0011546 0.1895 0.00065888 0.19016 0.17441 0 0.034609 0.0389 0 0.96409 0.27981 0.077825 0.010658 4.6477 0.066505 8.0653e-05 0.82358 0.0056452 0.006391 0.0013849 0.98696 0.99172 2.986e-06 1.1944e-05 0.13493 0.94721 0.9165 0.0013963 0.99354 0.59586 0.0018813 0.43014 1.8913 1.8907 16.0021 144.9906 0.00016458 -85.658 0.79236
1.8964 0.98804 5.5137e-05 3.8182 0.012024 2.493e-05 0.0011546 0.18954 0.00065888 0.19019 0.17444 0 0.034607 0.0389 0 0.96418 0.27985 0.07784 0.01066 4.6484 0.066516 8.0667e-05 0.82357 0.0056458 0.0063916 0.0013849 0.98696 0.99172 2.9859e-06 1.1944e-05 0.13494 0.94733 0.91655 0.0013963 0.99357 0.596 0.0018812 0.43016 1.8917 1.8911 16.0021 144.9906 0.00016449 -85.6581 0.79336
1.8974 0.98804 5.5137e-05 3.8182 0.012024 2.4943e-05 0.0011546 0.18957 0.00065888 0.19023 0.17448 0 0.034605 0.0389 0 0.96427 0.27989 0.077855 0.010662 4.6491 0.066526 8.0682e-05 0.82355 0.0056464 0.0063922 0.0013848 0.98696 0.99172 2.9859e-06 1.1943e-05 0.13494 0.94744 0.91661 0.0013963 0.99359 0.59614 0.0018812 0.43017 1.8921 1.8915 16.002 144.9906 0.00016441 -85.6581 0.79436
1.8984 0.98804 5.5137e-05 3.8182 0.012024 2.4956e-05 0.0011546 0.18961 0.00065888 0.19027 0.17451 0 0.034603 0.0389 0 0.96436 0.27994 0.07787 0.010663 4.6498 0.066537 8.0696e-05 0.82354 0.005647 0.0063928 0.0013848 0.98696 0.99172 2.9858e-06 1.1943e-05 0.13495 0.94755 0.91666 0.0013963 0.99362 0.59628 0.0018812 0.43018 1.8925 1.8919 16.002 144.9906 0.00016433 -85.6582 0.79536
1.8994 0.98804 5.5137e-05 3.8182 0.012024 2.4969e-05 0.0011546 0.18965 0.00065888 0.1903 0.17455 0 0.034601 0.0389 0 0.96446 0.27998 0.077885 0.010665 4.6504 0.066548 8.071e-05 0.82353 0.0056476 0.0063934 0.0013848 0.98696 0.99172 2.9858e-06 1.1943e-05 0.13495 0.94767 0.91671 0.0013963 0.99364 0.59642 0.0018812 0.43019 1.8929 1.8923 16.002 144.9907 0.00016425 -85.6583 0.79636
1.9004 0.98804 5.5137e-05 3.8182 0.012024 2.4982e-05 0.0011546 0.18968 0.00065888 0.19034 0.17458 0 0.034599 0.0389 0 0.96455 0.28002 0.0779 0.010667 4.6511 0.066559 8.0725e-05 0.82352 0.0056482 0.006394 0.0013848 0.98696 0.99172 2.9857e-06 1.1943e-05 0.13496 0.94778 0.91676 0.0013963 0.99366 0.59656 0.0018812 0.4302 1.8933 1.8927 16.0019 144.9907 0.00016417 -85.6584 0.79736
1.9014 0.98804 5.5137e-05 3.8182 0.012024 2.4995e-05 0.0011546 0.18972 0.00065888 0.19038 0.17462 0 0.034597 0.0389 0 0.96464 0.28006 0.077914 0.010669 4.6518 0.06657 8.0739e-05 0.82351 0.0056488 0.0063946 0.0013848 0.98696 0.99172 2.9857e-06 1.1943e-05 0.13496 0.94789 0.91681 0.0013963 0.99368 0.5967 0.0018812 0.43022 1.8937 1.8931 16.0019 144.9907 0.00016408 -85.6585 0.79836
1.9024 0.98804 5.5137e-05 3.8182 0.012024 2.5008e-05 0.0011546 0.18976 0.00065888 0.19041 0.17465 0 0.034595 0.0389 0 0.96473 0.2801 0.077929 0.01067 4.6525 0.066581 8.0753e-05 0.8235 0.0056494 0.0063952 0.0013847 0.98696 0.99172 2.9857e-06 1.1943e-05 0.13497 0.948 0.91687 0.0013963 0.99371 0.59684 0.0018812 0.43023 1.894 1.8934 16.0019 144.9907 0.000164 -85.6586 0.79936
1.9034 0.98804 5.5137e-05 3.8182 0.012024 2.5021e-05 0.0011546 0.18979 0.00065888 0.19045 0.17469 0 0.034593 0.0389 0 0.96482 0.28014 0.077944 0.010672 4.6532 0.066592 8.0768e-05 0.82349 0.00565 0.0063959 0.0013847 0.98696 0.99172 2.9856e-06 1.1942e-05 0.13497 0.94811 0.91692 0.0013963 0.99373 0.59698 0.0018811 0.43024 1.8944 1.8938 16.0019 144.9907 0.00016392 -85.6586 0.80036
1.9044 0.98804 5.5137e-05 3.8182 0.012024 2.5034e-05 0.0011546 0.18983 0.00065888 0.19049 0.17472 0 0.034591 0.0389 0 0.96492 0.28018 0.077959 0.010674 4.6539 0.066603 8.0782e-05 0.82348 0.0056506 0.0063965 0.0013847 0.98696 0.99172 2.9856e-06 1.1942e-05 0.13498 0.94822 0.91697 0.0013963 0.99375 0.59712 0.0018811 0.43025 1.8948 1.8942 16.0018 144.9908 0.00016384 -85.6587 0.80136
1.9054 0.98804 5.5137e-05 3.8182 0.012024 2.5048e-05 0.0011546 0.18987 0.00065888 0.19052 0.17476 0 0.034589 0.0389 0 0.96501 0.28022 0.077974 0.010676 4.6546 0.066614 8.0796e-05 0.82347 0.0056512 0.0063971 0.0013847 0.98696 0.99172 2.9855e-06 1.1942e-05 0.13498 0.94833 0.91702 0.0013962 0.99377 0.59726 0.0018811 0.43026 1.8952 1.8946 16.0018 144.9908 0.00016376 -85.6588 0.80236
1.9064 0.98804 5.5137e-05 3.8182 0.012024 2.5061e-05 0.0011546 0.1899 0.00065889 0.19056 0.17479 0 0.034586 0.0389 0 0.9651 0.28027 0.077989 0.010677 4.6553 0.066625 8.0811e-05 0.82346 0.0056518 0.0063977 0.0013847 0.98696 0.99172 2.9855e-06 1.1942e-05 0.13499 0.94844 0.91707 0.0013962 0.9938 0.5974 0.0018811 0.43028 1.8956 1.895 16.0018 144.9908 0.00016368 -85.6589 0.80336
1.9074 0.98804 5.5136e-05 3.8182 0.012024 2.5074e-05 0.0011546 0.18994 0.00065889 0.1906 0.17483 0 0.034584 0.0389 0 0.96519 0.28031 0.078004 0.010679 4.656 0.066636 8.0825e-05 0.82345 0.0056523 0.0063983 0.0013846 0.98696 0.99172 2.9854e-06 1.1942e-05 0.13499 0.94855 0.91712 0.0013962 0.99382 0.59754 0.0018811 0.43029 1.896 1.8954 16.0017 144.9908 0.0001636 -85.659 0.80436
1.9084 0.98804 5.5136e-05 3.8182 0.012024 2.5087e-05 0.0011546 0.18998 0.00065889 0.19063 0.17486 0 0.034582 0.0389 0 0.96529 0.28035 0.078019 0.010681 4.6567 0.066647 8.0839e-05 0.82343 0.0056529 0.0063989 0.0013846 0.98696 0.99172 2.9854e-06 1.1942e-05 0.135 0.94866 0.91717 0.0013962 0.99384 0.59768 0.0018811 0.4303 1.8964 1.8958 16.0017 144.9908 0.00016352 -85.659 0.80536
1.9094 0.98804 5.5136e-05 3.8182 0.012024 2.51e-05 0.0011546 0.19001 0.00065889 0.19067 0.17489 0 0.03458 0.0389 0 0.96538 0.28039 0.078034 0.010683 4.6574 0.066658 8.0854e-05 0.82342 0.0056535 0.0063996 0.0013846 0.98696 0.99172 2.9854e-06 1.1941e-05 0.135 0.94877 0.91722 0.0013962 0.99386 0.59782 0.0018811 0.43031 1.8968 1.8962 16.0017 144.9909 0.00016345 -85.6591 0.80636
1.9104 0.98804 5.5136e-05 3.8182 0.012024 2.5113e-05 0.0011546 0.19005 0.00065889 0.1907 0.17493 0 0.034578 0.0389 0 0.96547 0.28043 0.078048 0.010684 4.6581 0.066668 8.0868e-05 0.82341 0.0056541 0.0064002 0.0013846 0.98697 0.99172 2.9853e-06 1.1941e-05 0.13501 0.94888 0.91727 0.0013962 0.99388 0.59796 0.0018811 0.43032 1.8972 1.8966 16.0017 144.9909 0.00016337 -85.6592 0.80736
1.9114 0.98804 5.5136e-05 3.8182 0.012024 2.5126e-05 0.0011546 0.19009 0.00065889 0.19074 0.17496 0 0.034576 0.0389 0 0.96556 0.28047 0.078063 0.010686 4.6588 0.066679 8.0882e-05 0.8234 0.0056547 0.0064008 0.0013846 0.98697 0.99172 2.9853e-06 1.1941e-05 0.13501 0.94899 0.91732 0.0013962 0.9939 0.5981 0.001881 0.43034 1.8976 1.897 16.0016 144.9909 0.00016329 -85.6593 0.80836
1.9124 0.98804 5.5136e-05 3.8182 0.012024 2.5139e-05 0.0011546 0.19012 0.00065889 0.19078 0.175 0 0.034574 0.0389 0 0.96565 0.28051 0.078078 0.010688 4.6594 0.06669 8.0897e-05 0.82339 0.0056553 0.0064014 0.0013846 0.98697 0.99172 2.9852e-06 1.1941e-05 0.13502 0.9491 0.91737 0.0013962 0.99393 0.59824 0.001881 0.43035 1.898 1.8974 16.0016 144.9909 0.00016321 -85.6593 0.80936
1.9134 0.98804 5.5136e-05 3.8182 0.012024 2.5152e-05 0.0011546 0.19016 0.00065889 0.19081 0.17503 0 0.034572 0.0389 0 0.96575 0.28056 0.078093 0.01069 4.6601 0.066701 8.091e-05 0.82338 0.0056559 0.006402 0.0013845 0.98697 0.99172 2.9852e-06 1.1941e-05 0.13502 0.9492 0.91742 0.0013962 0.99395 0.59838 0.001881 0.43036 1.8983 1.8978 16.0016 144.9909 0.00016313 -85.6594 0.81036
1.9144 0.98804 5.5136e-05 3.8182 0.012024 2.5166e-05 0.0011546 0.1902 0.00065889 0.19085 0.17507 0 0.03457 0.0389 0 0.96584 0.2806 0.078108 0.010691 4.6608 0.066712 8.0925e-05 0.82337 0.0056565 0.0064026 0.0013845 0.98697 0.99172 2.9852e-06 1.1941e-05 0.13503 0.94931 0.91747 0.0013962 0.99397 0.59852 0.001881 0.43037 1.8987 1.8982 16.0015 144.991 0.00016306 -85.6595 0.81136
1.9154 0.98804 5.5136e-05 3.8182 0.012024 2.5179e-05 0.0011546 0.19023 0.00065889 0.19089 0.1751 0 0.034568 0.0389 0 0.96593 0.28064 0.078123 0.010693 4.6615 0.066723 8.094e-05 0.82336 0.0056571 0.0064033 0.0013845 0.98697 0.99172 2.9851e-06 1.194e-05 0.13503 0.94942 0.91752 0.0013961 0.99399 0.59866 0.001881 0.43038 1.8991 1.8985 16.0015 144.991 0.00016298 -85.6596 0.81236
1.9164 0.98804 5.5136e-05 3.8182 0.012024 2.5192e-05 0.0011546 0.19027 0.00065889 0.19092 0.17513 0 0.034566 0.0389 0 0.96602 0.28068 0.078138 0.010695 4.6622 0.066734 8.0954e-05 0.82335 0.0056577 0.0064039 0.0013845 0.98697 0.99172 2.9851e-06 1.194e-05 0.13504 0.94953 0.91757 0.0013961 0.99401 0.5988 0.001881 0.4304 1.8995 1.8989 16.0015 144.991 0.0001629 -85.6596 0.81336
1.9174 0.98804 5.5136e-05 3.8182 0.012024 2.5205e-05 0.0011546 0.1903 0.00065889 0.19096 0.17517 0 0.034564 0.0389 0 0.96611 0.28072 0.078153 0.010697 4.6629 0.066745 8.0967e-05 0.82334 0.0056583 0.0064045 0.0013845 0.98697 0.99172 2.985e-06 1.194e-05 0.13504 0.94963 0.91762 0.0013961 0.99403 0.59894 0.001881 0.43041 1.8999 1.8993 16.0014 144.991 0.00016282 -85.6597 0.81436
1.9184 0.98804 5.5136e-05 3.8182 0.012024 2.5218e-05 0.0011546 0.19034 0.00065889 0.19099 0.1752 0 0.034562 0.0389 0 0.96621 0.28076 0.078168 0.010698 4.6636 0.066756 8.0984e-05 0.82333 0.0056589 0.0064051 0.0013845 0.98697 0.99172 2.985e-06 1.194e-05 0.13505 0.94974 0.91766 0.0013961 0.99405 0.59908 0.001881 0.43042 1.9003 1.8997 16.0014 144.9911 0.00016275 -85.6598 0.81536
1.9194 0.98804 5.5136e-05 3.8182 0.012024 2.5231e-05 0.0011546 0.19038 0.00065889 0.19103 0.17524 0 0.03456 0.0389 0 0.9663 0.28081 0.078183 0.0107 4.6643 0.066767 8.0998e-05 0.82331 0.0056595 0.0064057 0.0013844 0.98697 0.99172 2.985e-06 1.194e-05 0.13505 0.94984 0.91771 0.0013961 0.99407 0.59922 0.001881 0.43043 1.9007 1.9001 16.0014 144.9911 0.00016267 -85.6599 0.81636
1.9204 0.98804 5.5136e-05 3.8182 0.012024 2.5244e-05 0.0011546 0.19041 0.00065889 0.19107 0.17527 0 0.034558 0.0389 0 0.96639 0.28085 0.078198 0.010702 4.665 0.066778 8.1011e-05 0.8233 0.0056601 0.0064063 0.0013844 0.98697 0.99172 2.9849e-06 1.194e-05 0.13506 0.94995 0.91776 0.0013961 0.99409 0.59936 0.0018809 0.43044 1.901 1.9005 16.0014 144.9911 0.00016259 -85.6599 0.81736
1.9214 0.98804 5.5136e-05 3.8182 0.012024 2.5257e-05 0.0011546 0.19045 0.00065889 0.1911 0.1753 0 0.034556 0.0389 0 0.96648 0.28089 0.078212 0.010704 4.6657 0.066789 8.1029e-05 0.82329 0.0056607 0.006407 0.0013844 0.98697 0.99172 2.9849e-06 1.1939e-05 0.13506 0.95005 0.91781 0.0013961 0.99411 0.5995 0.0018809 0.43046 1.9014 1.9008 16.0013 144.9911 0.00016252 -85.66 0.81836
1.9224 0.98804 5.5135e-05 3.8182 0.012024 2.527e-05 0.0011546 0.19049 0.00065889 0.19114 0.17534 0 0.034554 0.0389 0 0.96658 0.28093 0.078227 0.010705 4.6664 0.0668 8.1042e-05 0.82328 0.0056613 0.0064076 0.0013844 0.98697 0.99172 2.9849e-06 1.1939e-05 0.13507 0.95016 0.91786 0.0013961 0.99413 0.59964 0.0018809 0.43047 1.9018 1.9012 16.0013 144.9911 0.00016244 -85.6601 0.81936
1.9234 0.98804 5.5135e-05 3.8182 0.012024 2.5283e-05 0.0011546 0.19052 0.00065889 0.19118 0.17537 0 0.034552 0.0389 0 0.96667 0.28097 0.078242 0.010707 4.6671 0.066811 8.1048e-05 0.82327 0.0056619 0.0064082 0.0013844 0.98697 0.99172 2.9848e-06 1.1939e-05 0.13507 0.95026 0.91791 0.0013961 0.99415 0.59978 0.0018809 0.43048 1.9022 1.9016 16.0013 144.9912 0.00016237 -85.6602 0.82036
1.9244 0.98804 5.5135e-05 3.8182 0.012024 2.5297e-05 0.0011546 0.19056 0.00065889 0.19121 0.17541 0 0.034549 0.0389 0 0.96676 0.28101 0.078257 0.010709 4.6678 0.066822 8.1069e-05 0.82326 0.0056625 0.0064088 0.0013844 0.98697 0.99172 2.9848e-06 1.1939e-05 0.13508 0.95037 0.91795 0.0013961 0.99417 0.59992 0.0018809 0.43049 1.9026 1.902 16.0012 144.9912 0.00016229 -85.6602 0.82136
1.9254 0.98804 5.5135e-05 3.8182 0.012024 2.531e-05 0.0011546 0.19059 0.00065889 0.19125 0.17544 0 0.034547 0.0389 0 0.96685 0.28105 0.078272 0.010711 4.6685 0.066832 8.1093e-05 0.82325 0.0056631 0.0064094 0.0013843 0.98697 0.99172 2.9847e-06 1.1939e-05 0.13508 0.95047 0.918 0.0013961 0.99419 0.60006 0.0018809 0.4305 1.9029 1.9024 16.0012 144.9912 0.00016222 -85.6603 0.82236
1.9264 0.98804 5.5135e-05 3.8182 0.012024 2.5323e-05 0.0011546 0.19063 0.00065889 0.19128 0.17547 0 0.034545 0.0389 0 0.96695 0.2811 0.078287 0.010712 4.6692 0.066843 8.1097e-05 0.82324 0.0056637 0.0064101 0.0013843 0.98697 0.99172 2.9847e-06 1.1939e-05 0.13509 0.95057 0.91805 0.0013961 0.99421 0.6002 0.0018809 0.43052 1.9033 1.9027 16.0012 144.9912 0.00016214 -85.6604 0.82336
1.9274 0.98804 5.5135e-05 3.8182 0.012024 2.5336e-05 0.0011546 0.19066 0.00065889 0.19132 0.17551 0 0.034543 0.0389 0 0.96704 0.28114 0.078302 0.010714 4.6699 0.066854 8.1107e-05 0.82323 0.0056643 0.0064107 0.0013843 0.98697 0.99172 2.9847e-06 1.1939e-05 0.13509 0.95068 0.91809 0.001396 0.99423 0.60034 0.0018809 0.43053 1.9037 1.9031 16.0011 144.9912 0.00016207 -85.6604 0.82436
1.9284 0.98804 5.5135e-05 3.8182 0.012024 2.5349e-05 0.0011546 0.1907 0.00065889 0.19136 0.17554 0 0.034541 0.0389 0 0.96713 0.28118 0.078317 0.010716 4.6706 0.066865 8.1131e-05 0.82322 0.0056649 0.0064113 0.0013843 0.98697 0.99172 2.9846e-06 1.1938e-05 0.1351 0.95078 0.91814 0.001396 0.99425 0.60048 0.0018808 0.43054 1.9041 1.9035 16.0011 144.9913 0.000162 -85.6605 0.82536
1.9294 0.98804 5.5135e-05 3.8182 0.012024 2.5362e-05 0.0011546 0.19074 0.00065889 0.19139 0.17558 0 0.034539 0.0389 0 0.96722 0.28122 0.078332 0.010718 4.6713 0.066876 8.1142e-05 0.8232 0.0056655 0.0064119 0.0013843 0.98697 0.99172 2.9846e-06 1.1938e-05 0.1351 0.95088 0.91819 0.001396 0.99427 0.60062 0.0018808 0.43055 1.9045 1.9039 16.0011 144.9913 0.00016192 -85.6606 0.82636
1.9304 0.98804 5.5135e-05 3.8182 0.012024 2.5375e-05 0.0011547 0.19077 0.0006589 0.19143 0.17561 0 0.034537 0.0389 0 0.96731 0.28126 0.078347 0.010719 4.672 0.066887 8.1149e-05 0.82319 0.0056661 0.0064125 0.0013843 0.98697 0.99172 2.9846e-06 1.1938e-05 0.13511 0.95098 0.91824 0.001396 0.99429 0.60075 0.0018808 0.43056 1.9048 1.9043 16.001 144.9913 0.00016185 -85.6606 0.82736
1.9314 0.98804 5.5135e-05 3.8182 0.012024 2.5388e-05 0.0011547 0.19081 0.0006589 0.19146 0.17564 0 0.034535 0.0389 0 0.96741 0.2813 0.078362 0.010721 4.6727 0.066898 8.1171e-05 0.82318 0.0056667 0.0064132 0.0013842 0.98697 0.99172 2.9845e-06 1.1938e-05 0.13511 0.95109 0.91828 0.001396 0.99431 0.60089 0.0018808 0.43057 1.9052 1.9046 16.001 144.9913 0.00016177 -85.6607 0.82836
1.9324 0.98804 5.5135e-05 3.8182 0.012024 2.5401e-05 0.0011547 0.19084 0.0006589 0.1915 0.17568 0 0.034533 0.0389 0 0.9675 0.28135 0.078377 0.010723 4.6735 0.066909 8.1187e-05 0.82317 0.0056673 0.0064138 0.0013842 0.98697 0.99172 2.9845e-06 1.1938e-05 0.13512 0.95119 0.91833 0.001396 0.99432 0.60103 0.0018808 0.43059 1.9056 1.905 16.001 144.9913 0.0001617 -85.6608 0.82936
1.9334 0.98804 5.5135e-05 3.8182 0.012024 2.5414e-05 0.0011547 0.19088 0.0006589 0.19153 0.17571 0 0.034531 0.0389 0 0.96759 0.28139 0.078392 0.010725 4.6742 0.06692 8.1193e-05 0.82316 0.0056679 0.0064144 0.0013842 0.98697 0.99172 2.9845e-06 1.1938e-05 0.13512 0.95129 0.91837 0.001396 0.99434 0.60117 0.0018808 0.4306 1.9059 1.9054 16.001 144.9914 0.00016163 -85.6608 0.83036
1.9344 0.98804 5.5135e-05 3.8182 0.012024 2.5428e-05 0.0011547 0.19092 0.0006589 0.19157 0.17574 0 0.034529 0.0389 0 0.96768 0.28143 0.078407 0.010726 4.6749 0.066931 8.1212e-05 0.82315 0.0056685 0.006415 0.0013842 0.98697 0.99172 2.9844e-06 1.1938e-05 0.13513 0.95139 0.91842 0.001396 0.99436 0.60131 0.0018808 0.43061 1.9063 1.9058 16.0009 144.9914 0.00016156 -85.6609 0.83136
1.9354 0.98804 5.5135e-05 3.8182 0.012024 2.5441e-05 0.0011547 0.19095 0.0006589 0.19161 0.17578 0 0.034527 0.0389 0 0.96778 0.28147 0.078422 0.010728 4.6756 0.066942 8.1231e-05 0.82314 0.0056691 0.0064156 0.0013842 0.98697 0.99172 2.9844e-06 1.1937e-05 0.13513 0.95149 0.91847 0.001396 0.99438 0.60145 0.0018808 0.43062 1.9067 1.9061 16.0009 144.9914 0.00016148 -85.661 0.83236
1.9364 0.98804 5.5135e-05 3.8182 0.012024 2.5454e-05 0.0011547 0.19099 0.0006589 0.19164 0.17581 0 0.034525 0.0389 0 0.96787 0.28151 0.078436 0.01073 4.6763 0.066953 8.1238e-05 0.82313 0.0056697 0.0064163 0.0013842 0.98697 0.99172 2.9844e-06 1.1937e-05 0.13514 0.95159 0.91851 0.001396 0.9944 0.60159 0.0018808 0.43063 1.9071 1.9065 16.0009 144.9914 0.00016141 -85.661 0.83336
1.9374 0.98804 5.5134e-05 3.8182 0.012024 2.5467e-05 0.0011547 0.19102 0.0006589 0.19168 0.17585 0 0.034523 0.0389 0 0.96796 0.28155 0.078451 0.010732 4.677 0.066964 8.1253e-05 0.82312 0.0056703 0.0064169 0.0013842 0.98697 0.99172 2.9843e-06 1.1937e-05 0.13514 0.95169 0.91856 0.001396 0.99442 0.60173 0.0018808 0.43065 1.9074 1.9069 16.0008 144.9914 0.00016134 -85.6611 0.83436
1.9384 0.98804 5.5134e-05 3.8182 0.012024 2.548e-05 0.0011547 0.19106 0.0006589 0.19171 0.17588 0 0.034521 0.0389 0 0.96805 0.2816 0.078466 0.010733 4.6777 0.066975 8.1273e-05 0.82311 0.0056709 0.0064175 0.0013841 0.98697 0.99172 2.9843e-06 1.1937e-05 0.13514 0.95179 0.9186 0.001396 0.99443 0.60186 0.0018807 0.43066 1.9078 1.9072 16.0008 144.9915 0.00016127 -85.6612 0.83536
1.9394 0.98804 5.5134e-05 3.8182 0.012024 2.5493e-05 0.0011547 0.19109 0.0006589 0.19175 0.17591 0 0.034519 0.0389 0 0.96815 0.28164 0.078481 0.010735 4.6784 0.066986 8.1284e-05 0.8231 0.0056715 0.0064181 0.0013841 0.98697 0.99172 2.9843e-06 1.1937e-05 0.13515 0.95189 0.91865 0.0013959 0.99445 0.602 0.0018807 0.43067 1.9082 1.9076 16.0008 144.9915 0.0001612 -85.6612 0.83636
1.9404 0.98804 5.5134e-05 3.8182 0.012024 2.5506e-05 0.0011547 0.19113 0.0006589 0.19178 0.17595 0 0.034517 0.0389 0 0.96824 0.28168 0.078496 0.010737 4.6791 0.066997 8.1295e-05 0.82308 0.0056721 0.0064188 0.0013841 0.98697 0.99172 2.9842e-06 1.1937e-05 0.13515 0.95199 0.91869 0.0013959 0.99447 0.60214 0.0018807 0.43068 1.9085 1.908 16.0007 144.9915 0.00016113 -85.6613 0.83736
1.9414 0.98804 5.5134e-05 3.8182 0.012024 2.5519e-05 0.0011547 0.19116 0.0006589 0.19182 0.17598 0 0.034515 0.0389 0 0.96833 0.28172 0.078511 0.010739 4.6798 0.067008 8.1315e-05 0.82307 0.0056727 0.0064194 0.0013841 0.98697 0.99172 2.9842e-06 1.1937e-05 0.13516 0.95209 0.91874 0.0013959 0.99449 0.60228 0.0018807 0.43069 1.9089 1.9084 16.0007 144.9915 0.00016105 -85.6613 0.83836
1.9424 0.98804 5.5134e-05 3.8182 0.012024 2.5532e-05 0.0011547 0.1912 0.0006589 0.19185 0.17601 0 0.034513 0.0389 0 0.96842 0.28176 0.078526 0.010741 4.6805 0.067019 8.1328e-05 0.82306 0.0056733 0.00642 0.0013841 0.98697 0.99172 2.9842e-06 1.1937e-05 0.13516 0.95218 0.91878 0.0013959 0.9945 0.60242 0.0018807 0.4307 1.9093 1.9087 16.0007 144.9915 0.00016098 -85.6614 0.83936
1.9434 0.98804 5.5134e-05 3.8182 0.012024 2.5546e-05 0.0011547 0.19124 0.0006589 0.19189 0.17605 0 0.034511 0.0389 0 0.96852 0.2818 0.078541 0.010742 4.6812 0.06703 8.1338e-05 0.82305 0.0056739 0.0064206 0.0013841 0.98697 0.99172 2.9841e-06 1.1936e-05 0.13517 0.95228 0.91883 0.0013959 0.99452 0.60256 0.0018807 0.43072 1.9096 1.9091 16.0007 144.9916 0.00016091 -85.6615 0.84036
1.9444 0.98804 5.5134e-05 3.8182 0.012024 2.5559e-05 0.0011547 0.19127 0.0006589 0.19193 0.17608 0 0.034509 0.0389 0 0.96861 0.28185 0.078556 0.010744 4.6819 0.067041 8.1357e-05 0.82304 0.0056745 0.0064213 0.0013841 0.98697 0.99172 2.9841e-06 1.1936e-05 0.13517 0.95238 0.91887 0.0013959 0.99454 0.60269 0.0018807 0.43073 1.91 1.9095 16.0006 144.9916 0.00016084 -85.6615 0.84136
1.9454 0.98804 5.5134e-05 3.8182 0.012024 2.5572e-05 0.0011547 0.19131 0.0006589 0.19196 0.17611 0 0.034507 0.0389 0 0.9687 0.28189 0.078571 0.010746 4.6826 0.067052 8.1373e-05 0.82303 0.0056751 0.0064219 0.001384 0.98697 0.99172 2.9841e-06 1.1936e-05 0.13518 0.95248 0.91892 0.0013959 0.99456 0.60283 0.0018807 0.43074 1.9104 1.9098 16.0006 144.9916 0.00016077 -85.6616 0.84236
1.9464 0.98804 5.5134e-05 3.8182 0.012024 2.5585e-05 0.0011547 0.19134 0.0006589 0.192 0.17615 0 0.034505 0.0389 0 0.96879 0.28193 0.078586 0.010748 4.6834 0.067062 8.1382e-05 0.82302 0.0056757 0.0064225 0.001384 0.98697 0.99172 2.984e-06 1.1936e-05 0.13518 0.95257 0.91896 0.0013959 0.99457 0.60297 0.0018807 0.43075 1.9107 1.9102 16.0006 144.9916 0.0001607 -85.6616 0.84336
1.9474 0.98804 5.5134e-05 3.8182 0.012024 2.5598e-05 0.0011547 0.19138 0.0006589 0.19203 0.17618 0 0.034503 0.0389 0 0.96889 0.28197 0.078601 0.010749 4.6841 0.067073 8.1398e-05 0.82301 0.0056763 0.0064231 0.001384 0.98697 0.99172 2.984e-06 1.1936e-05 0.13519 0.95267 0.91901 0.0013959 0.99459 0.60311 0.0018807 0.43076 1.9111 1.9106 16.0005 144.9916 0.00016063 -85.6617 0.84436
1.9484 0.98804 5.5134e-05 3.8182 0.012024 2.5611e-05 0.0011547 0.19141 0.0006589 0.19207 0.17621 0 0.034501 0.0389 0 0.96898 0.28201 0.078616 0.010751 4.6848 0.067084 8.1416e-05 0.823 0.0056769 0.0064238 0.001384 0.98697 0.99172 2.984e-06 1.1936e-05 0.13519 0.95277 0.91905 0.0013959 0.99461 0.60325 0.0018806 0.43078 1.9115 1.9109 16.0005 144.9917 0.00016056 -85.6618 0.84536
1.9494 0.98804 5.5134e-05 3.8182 0.012024 2.5624e-05 0.0011547 0.19145 0.0006589 0.1921 0.17625 0 0.034499 0.0389 0 0.96907 0.28205 0.078631 0.010753 4.6855 0.067095 8.1427e-05 0.82299 0.0056775 0.0064244 0.001384 0.98697 0.99172 2.9839e-06 1.1936e-05 0.1352 0.95286 0.91909 0.0013959 0.99462 0.60339 0.0018806 0.43079 1.9118 1.9113 16.0005 144.9917 0.00016049 -85.6618 0.84636
1.9504 0.98804 5.5134e-05 3.8182 0.012024 2.5637e-05 0.0011547 0.19148 0.0006589 0.19214 0.17628 0 0.034497 0.0389 0 0.96916 0.2821 0.078646 0.010755 4.6862 0.067106 8.1441e-05 0.82298 0.0056781 0.006425 0.001384 0.98697 0.99172 2.9839e-06 1.1936e-05 0.1352 0.95296 0.91914 0.0013959 0.99464 0.60352 0.0018806 0.4308 1.9122 1.9117 16.0004 144.9917 0.00016043 -85.6619 0.84736
1.9514 0.98804 5.5134e-05 3.8182 0.012024 2.565e-05 0.0011547 0.19152 0.0006589 0.19217 0.17631 0 0.034495 0.0389 0 0.96926 0.28214 0.078661 0.010756 4.6869 0.067117 8.1458e-05 0.82296 0.0056787 0.0064256 0.001384 0.98697 0.99172 2.9839e-06 1.1935e-05 0.13521 0.95305 0.91918 0.0013959 0.99466 0.60366 0.0018806 0.43081 1.9126 1.912 16.0004 144.9917 0.00016036 -85.6619 0.84836
1.9524 0.98804 5.5134e-05 3.8182 0.012024 2.5663e-05 0.0011547 0.19155 0.0006589 0.19221 0.17635 0 0.034493 0.0389 0 0.96935 0.28218 0.078676 0.010758 4.6876 0.067128 8.1471e-05 0.82295 0.0056793 0.0064263 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13521 0.95315 0.91923 0.0013959 0.99467 0.6038 0.0018806 0.43082 1.9129 1.9124 16.0004 144.9917 0.00016029 -85.662 0.84936
1.9534 0.98804 5.5133e-05 3.8182 0.012024 2.5677e-05 0.0011547 0.19159 0.0006589 0.19224 0.17638 0 0.034491 0.0389 0 0.96944 0.28222 0.078691 0.01076 4.6883 0.067139 8.1484e-05 0.82294 0.0056799 0.0064269 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13522 0.95325 0.91927 0.0013958 0.99469 0.60394 0.0018806 0.43083 1.9133 1.9127 16.0003 144.9918 0.00016022 -85.6621 0.85036
1.9544 0.98804 5.5133e-05 3.8182 0.012024 2.569e-05 0.0011547 0.19162 0.00065891 0.19228 0.17641 0 0.034489 0.0389 0 0.96953 0.28226 0.078706 0.010762 4.6891 0.06715 8.1501e-05 0.82293 0.0056806 0.0064275 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13522 0.95334 0.91931 0.0013958 0.99471 0.60408 0.0018806 0.43085 1.9136 1.9131 16.0003 144.9918 0.00016015 -85.6621 0.85136
1.9554 0.98804 5.5133e-05 3.8182 0.012024 2.5703e-05 0.0011547 0.19166 0.00065891 0.19231 0.17645 0 0.034487 0.0389 0 0.96963 0.2823 0.078721 0.010763 4.6898 0.067161 8.1515e-05 0.82292 0.0056812 0.0064281 0.0013839 0.98697 0.99172 2.9838e-06 1.1935e-05 0.13523 0.95343 0.91936 0.0013958 0.99472 0.60421 0.0018806 0.43086 1.914 1.9135 16.0003 144.9918 0.00016009 -85.6622 0.85236
1.9564 0.98804 5.5133e-05 3.8182 0.012024 2.5716e-05 0.0011547 0.19169 0.00065891 0.19235 0.17648 0 0.034485 0.0389 0 0.96972 0.28235 0.078736 0.010765 4.6905 0.067172 8.1527e-05 0.82291 0.0056818 0.0064288 0.0013839 0.98697 0.99172 2.9837e-06 1.1935e-05 0.13523 0.95353 0.9194 0.0013958 0.99474 0.60435 0.0018806 0.43087 1.9144 1.9138 16.0002 144.9918 0.00016002 -85.6622 0.85336
1.9574 0.98804 5.5133e-05 3.8182 0.012024 2.5729e-05 0.0011547 0.19173 0.00065891 0.19238 0.17651 0 0.034483 0.0389 0 0.96981 0.28239 0.078751 0.010767 4.6912 0.067183 8.1543e-05 0.8229 0.0056824 0.0064294 0.0013839 0.98697 0.99172 2.9837e-06 1.1935e-05 0.13524 0.95362 0.91944 0.0013958 0.99475 0.60449 0.0018806 0.43088 1.9147 1.9142 16.0002 144.9919 0.00015995 -85.6623 0.85436
1.9584 0.98804 5.5133e-05 3.8182 0.012024 2.5742e-05 0.0011547 0.19176 0.00065891 0.19242 0.17655 0 0.034481 0.0389 0 0.96991 0.28243 0.078766 0.010769 4.6919 0.067194 8.1559e-05 0.82289 0.005683 0.00643 0.0013839 0.98697 0.99172 2.9837e-06 1.1935e-05 0.13524 0.95372 0.91948 0.0013958 0.99477 0.60463 0.0018806 0.43089 1.9151 1.9145 16.0002 144.9919 0.00015988 -85.6623 0.85536
1.9594 0.98804 5.5133e-05 3.8182 0.012024 2.5755e-05 0.0011547 0.1918 0.00065891 0.19245 0.17658 0 0.034479 0.0389 0 0.97 0.28247 0.078781 0.01077 4.6926 0.067205 8.1571e-05 0.82288 0.0056836 0.0064306 0.0013839 0.98697 0.99172 2.9836e-06 1.1934e-05 0.13525 0.95381 0.91953 0.0013958 0.99478 0.60476 0.0018805 0.4309 1.9154 1.9149 16.0002 144.9919 0.00015982 -85.6624 0.85636
1.9604 0.98804 5.5133e-05 3.8182 0.012024 2.5768e-05 0.0011547 0.19183 0.00065891 0.19249 0.17661 0 0.034477 0.0389 0 0.97009 0.28251 0.078796 0.010772 4.6934 0.067216 8.1586e-05 0.82287 0.0056842 0.0064313 0.0013838 0.98697 0.99172 2.9836e-06 1.1934e-05 0.13525 0.9539 0.91957 0.0013958 0.9948 0.6049 0.0018805 0.43092 1.9158 1.9153 16.0001 144.9919 0.00015975 -85.6624 0.85736
1.9614 0.98804 5.5133e-05 3.8182 0.012024 2.5781e-05 0.0011547 0.19187 0.00065891 0.19252 0.17664 0 0.034475 0.0389 0 0.97018 0.28255 0.078811 0.010774 4.6941 0.067227 8.1602e-05 0.82285 0.0056848 0.0064319 0.0013838 0.98697 0.99172 2.9836e-06 1.1934e-05 0.13526 0.95399 0.91961 0.0013958 0.99482 0.60504 0.0018805 0.43093 1.9161 1.9156 16.0001 144.9919 0.00015968 -85.6625 0.85836
1.9624 0.98804 5.5133e-05 3.8182 0.012024 2.5794e-05 0.0011547 0.1919 0.00065891 0.19256 0.17668 0 0.034473 0.0389 0 0.97028 0.2826 0.078826 0.010776 4.6948 0.067238 8.1615e-05 0.82284 0.0056854 0.0064325 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13526 0.95409 0.91965 0.0013958 0.99483 0.60518 0.0018805 0.43094 1.9165 1.916 16.0001 144.992 0.00015962 -85.6625 0.85936
1.9634 0.98804 5.5133e-05 3.8182 0.012024 2.5808e-05 0.0011547 0.19194 0.00065891 0.19259 0.17671 0 0.034471 0.0389 0 0.97037 0.28264 0.078841 0.010777 4.6955 0.067249 8.1628e-05 0.82283 0.005686 0.0064332 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13527 0.95418 0.91969 0.0013958 0.99485 0.60531 0.0018805 0.43095 1.9169 1.9163 16 144.992 0.00015955 -85.6626 0.86036
1.9644 0.98804 5.5133e-05 3.8182 0.012023 2.5821e-05 0.0011547 0.19197 0.00065891 0.19263 0.17674 0 0.034469 0.0389 0 0.97046 0.28268 0.078856 0.010779 4.6962 0.06726 8.1645e-05 0.82282 0.0056866 0.0064338 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13527 0.95427 0.91974 0.0013958 0.99486 0.60545 0.0018805 0.43096 1.9172 1.9167 16 144.992 0.00015949 -85.6627 0.86136
1.9654 0.98804 5.5133e-05 3.8182 0.012023 2.5834e-05 0.0011547 0.19201 0.00065891 0.19266 0.17678 0 0.034467 0.0389 0 0.97055 0.28272 0.078871 0.010781 4.6969 0.067271 8.1659e-05 0.82281 0.0056872 0.0064344 0.0013838 0.98698 0.99172 2.9835e-06 1.1934e-05 0.13528 0.95436 0.91978 0.0013958 0.99488 0.60559 0.0018805 0.43097 1.9176 1.917 16 144.992 0.00015942 -85.6627 0.86236
1.9664 0.98804 5.5133e-05 3.8182 0.012023 2.5847e-05 0.0011547 0.19204 0.00065891 0.1927 0.17681 0 0.034465 0.0389 0 0.97065 0.28276 0.078886 0.010783 4.6977 0.067282 8.1672e-05 0.8228 0.0056878 0.006435 0.0013838 0.98698 0.99172 2.9834e-06 1.1934e-05 0.13528 0.95445 0.91982 0.0013958 0.99489 0.60573 0.0018805 0.43099 1.9179 1.9174 15.9999 144.992 0.00015935 -85.6628 0.86336
1.9674 0.98804 5.5133e-05 3.8182 0.012023 2.586e-05 0.0011547 0.19208 0.00065891 0.19273 0.17684 0 0.034464 0.0389 0 0.97074 0.2828 0.078901 0.010784 4.6984 0.067293 8.1687e-05 0.82279 0.0056884 0.0064357 0.0013838 0.98698 0.99172 2.9834e-06 1.1934e-05 0.13529 0.95454 0.91986 0.0013958 0.99491 0.60586 0.0018805 0.431 1.9183 1.9177 15.9999 144.9921 0.00015929 -85.6628 0.86436
1.9684 0.98804 5.5132e-05 3.8182 0.012023 2.5873e-05 0.0011547 0.19211 0.00065891 0.19277 0.17687 0 0.034462 0.0389 0 0.97083 0.28285 0.078916 0.010786 4.6991 0.067304 8.1702e-05 0.82278 0.005689 0.0064363 0.0013837 0.98698 0.99172 2.9834e-06 1.1933e-05 0.13529 0.95463 0.9199 0.0013957 0.99492 0.606 0.0018805 0.43101 1.9186 1.9181 15.9999 144.9921 0.00015922 -85.6629 0.86536
1.9694 0.98804 5.5132e-05 3.8182 0.012023 2.5886e-05 0.0011547 0.19215 0.00065891 0.1928 0.17691 0 0.03446 0.0389 0 0.97093 0.28289 0.078931 0.010788 4.6998 0.067315 8.1715e-05 0.82277 0.0056897 0.0064369 0.0013837 0.98698 0.99172 2.9834e-06 1.1933e-05 0.1353 0.95473 0.91994 0.0013957 0.99494 0.60614 0.0018805 0.43102 1.919 1.9184 15.9998 144.9921 0.00015916 -85.6629 0.86636
1.9704 0.98804 5.5132e-05 3.8182 0.012023 2.5899e-05 0.0011547 0.19218 0.00065891 0.19284 0.17694 0 0.034458 0.0389 0 0.97102 0.28293 0.078946 0.01079 4.7005 0.067326 8.173e-05 0.82276 0.0056903 0.0064376 0.0013837 0.98698 0.99172 2.9833e-06 1.1933e-05 0.1353 0.95482 0.91998 0.0013957 0.99495 0.60627 0.0018805 0.43103 1.9193 1.9188 15.9998 144.9921 0.0001591 -85.663 0.86736
1.9714 0.98804 5.5132e-05 3.8182 0.012023 2.5912e-05 0.0011547 0.19222 0.00065891 0.19287 0.17697 0 0.034456 0.0389 0 0.97111 0.28297 0.078961 0.010791 4.7013 0.067337 8.1746e-05 0.82274 0.0056909 0.0064382 0.0013837 0.98698 0.99172 2.9833e-06 1.1933e-05 0.13531 0.9549 0.92002 0.0013957 0.99496 0.60641 0.0018804 0.43104 1.9197 1.9191 15.9998 144.9921 0.00015903 -85.663 0.86836
1.9724 0.98804 5.5132e-05 3.8182 0.012023 2.5925e-05 0.0011547 0.19225 0.00065891 0.19291 0.17701 0 0.034454 0.0389 0 0.9712 0.28301 0.078976 0.010793 4.702 0.067348 8.1759e-05 0.82273 0.0056915 0.0064388 0.0013837 0.98698 0.99173 2.9833e-06 1.1933e-05 0.13531 0.95499 0.92007 0.0013957 0.99498 0.60655 0.0018804 0.43106 1.92 1.9195 15.9997 144.9922 0.00015897 -85.6631 0.86936
1.9734 0.98804 5.5132e-05 3.8182 0.012023 2.5939e-05 0.0011547 0.19229 0.00065891 0.19294 0.17704 0 0.034452 0.0389 0 0.9713 0.28306 0.078991 0.010795 4.7027 0.067359 8.1773e-05 0.82272 0.0056921 0.0064395 0.0013837 0.98698 0.99173 2.9833e-06 1.1933e-05 0.13532 0.95508 0.92011 0.0013957 0.99499 0.60669 0.0018804 0.43107 1.9204 1.9198 15.9997 144.9922 0.0001589 -85.6631 0.87036
1.9744 0.98804 5.5132e-05 3.8182 0.012023 2.5952e-05 0.0011547 0.19232 0.00065891 0.19298 0.17707 0 0.03445 0.0389 0 0.97139 0.2831 0.079006 0.010797 4.7034 0.06737 8.1789e-05 0.82271 0.0056927 0.0064401 0.0013837 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13532 0.95517 0.92015 0.0013957 0.99501 0.60682 0.0018804 0.43108 1.9207 1.9202 15.9997 144.9922 0.00015884 -85.6632 0.87136
1.9754 0.98804 5.5132e-05 3.8182 0.012023 2.5965e-05 0.0011547 0.19236 0.00065891 0.19301 0.1771 0 0.034448 0.0389 0 0.97148 0.28314 0.079021 0.010798 4.7042 0.067381 8.1802e-05 0.8227 0.0056933 0.0064407 0.0013837 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13533 0.95526 0.92019 0.0013957 0.99502 0.60696 0.0018804 0.43109 1.9211 1.9205 15.9997 144.9922 0.00015878 -85.6632 0.87236
1.9764 0.98804 5.5132e-05 3.8182 0.012023 2.5978e-05 0.0011547 0.19239 0.00065891 0.19304 0.17714 0 0.034446 0.0389 0 0.97158 0.28318 0.079036 0.0108 4.7049 0.067392 8.1816e-05 0.82269 0.0056939 0.0064414 0.0013837 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13533 0.95535 0.92023 0.0013957 0.99504 0.6071 0.0018804 0.4311 1.9214 1.9209 15.9996 144.9922 0.00015871 -85.6633 0.87336
1.9774 0.98804 5.5132e-05 3.8182 0.012023 2.5991e-05 0.0011547 0.19242 0.00065891 0.19308 0.17717 0 0.034444 0.0389 0 0.97167 0.28322 0.079051 0.010802 4.7056 0.067403 8.1832e-05 0.82268 0.0056945 0.006442 0.0013836 0.98698 0.99173 2.9832e-06 1.1933e-05 0.13534 0.95544 0.92027 0.0013957 0.99505 0.60723 0.0018804 0.43111 1.9218 1.9212 15.9996 144.9923 0.00015865 -85.6633 0.87436
1.9784 0.98804 5.5132e-05 3.8182 0.012023 2.6004e-05 0.0011547 0.19246 0.00065892 0.19311 0.1772 0 0.034442 0.0389 0 0.97176 0.28326 0.079066 0.010804 4.7063 0.067414 8.1846e-05 0.82267 0.0056951 0.0064426 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.13534 0.95553 0.92031 0.0013957 0.99506 0.60737 0.0018804 0.43113 1.9221 1.9216 15.9996 144.9923 0.00015859 -85.6633 0.87536
1.9794 0.98804 5.5132e-05 3.8182 0.012023 2.6017e-05 0.0011547 0.19249 0.00065892 0.19315 0.17723 0 0.03444 0.0389 0 0.97185 0.28331 0.079081 0.010806 4.7071 0.067425 8.186e-05 0.82266 0.0056957 0.0064433 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.13535 0.95561 0.92035 0.0013957 0.99508 0.60751 0.0018804 0.43114 1.9224 1.9219 15.9995 144.9923 0.00015853 -85.6634 0.87636
1.9804 0.98804 5.5132e-05 3.8182 0.012023 2.603e-05 0.0011547 0.19253 0.00065892 0.19318 0.17727 0 0.034438 0.0389 0 0.97195 0.28335 0.079096 0.010807 4.7078 0.067436 8.1875e-05 0.82265 0.0056964 0.0064439 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.13535 0.9557 0.92039 0.0013957 0.99509 0.60764 0.0018804 0.43115 1.9228 1.9223 15.9995 144.9923 0.00015846 -85.6634 0.87736
1.9814 0.98804 5.5132e-05 3.8182 0.012023 2.6043e-05 0.0011547 0.19256 0.00065892 0.19322 0.1773 0 0.034436 0.0389 0 0.97204 0.28339 0.079111 0.010809 4.7085 0.067447 8.189e-05 0.82264 0.005697 0.0064445 0.0013836 0.98698 0.99173 2.9831e-06 1.1932e-05 0.13536 0.95579 0.92043 0.0013957 0.9951 0.60778 0.0018804 0.43116 1.9231 1.9226 15.9995 144.9923 0.0001584 -85.6635 0.87836
1.9824 0.98804 5.5132e-05 3.8182 0.012023 2.6056e-05 0.0011547 0.1926 0.00065892 0.19325 0.17733 0 0.034434 0.0389 0 0.97213 0.28343 0.079126 0.010811 4.7092 0.067458 8.1903e-05 0.82262 0.0056976 0.0064451 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13536 0.95587 0.92046 0.0013957 0.99512 0.60792 0.0018804 0.43117 1.9235 1.923 15.9994 144.9924 0.00015834 -85.6635 0.87936
1.9834 0.98804 5.5132e-05 3.8182 0.012023 2.607e-05 0.0011547 0.19263 0.00065892 0.19329 0.17736 0 0.034432 0.0389 0 0.97223 0.28347 0.079141 0.010813 4.71 0.067469 8.1918e-05 0.82261 0.0056982 0.0064458 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13537 0.95596 0.9205 0.0013957 0.99513 0.60805 0.0018804 0.43118 1.9238 1.9233 15.9994 144.9924 0.00015828 -85.6636 0.88036
1.9844 0.98804 5.5131e-05 3.8182 0.012023 2.6083e-05 0.0011547 0.19267 0.00065892 0.19332 0.1774 0 0.03443 0.0389 0 0.97232 0.28352 0.079156 0.010814 4.7107 0.06748 8.1933e-05 0.8226 0.0056988 0.0064464 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13537 0.95605 0.92054 0.0013957 0.99514 0.60819 0.0018804 0.4312 1.9242 1.9236 15.9994 144.9924 0.00015822 -85.6636 0.88136
1.9854 0.98804 5.5131e-05 3.8182 0.012023 2.6096e-05 0.0011547 0.1927 0.00065892 0.19335 0.17743 0 0.034429 0.0389 0 0.97241 0.28356 0.079171 0.010816 4.7114 0.067491 8.1947e-05 0.82259 0.0056994 0.006447 0.0013836 0.98698 0.99173 2.983e-06 1.1932e-05 0.13538 0.95613 0.92058 0.0013956 0.99516 0.60832 0.0018803 0.43121 1.9245 1.924 15.9993 144.9924 0.00015815 -85.6637 0.88236
1.9864 0.98804 5.5131e-05 3.8182 0.012023 2.6109e-05 0.0011547 0.19273 0.00065892 0.19339 0.17746 0 0.034427 0.0389 0 0.97251 0.2836 0.079186 0.010818 4.7121 0.067502 8.1961e-05 0.82258 0.0057 0.0064477 0.0013836 0.98698 0.99173 2.9829e-06 1.1932e-05 0.13539 0.95622 0.92062 0.0013956 0.99517 0.60846 0.0018803 0.43122 1.9248 1.9243 15.9993 144.9924 0.00015809 -85.6637 0.88336
1.9874 0.98804 5.5131e-05 3.8182 0.012023 2.6122e-05 0.0011547 0.19277 0.00065892 0.19342 0.17749 0 0.034425 0.0389 0 0.9726 0.28364 0.079202 0.01082 4.7129 0.067513 8.1976e-05 0.82257 0.0057006 0.0064483 0.0013835 0.98698 0.99173 2.9829e-06 1.1932e-05 0.13539 0.9563 0.92066 0.0013956 0.99518 0.6086 0.0018803 0.43123 1.9252 1.9247 15.9993 144.9925 0.00015803 -85.6638 0.88436
1.9884 0.98804 5.5131e-05 3.8182 0.012023 2.6135e-05 0.0011547 0.1928 0.00065892 0.19346 0.17753 0 0.034423 0.0389 0 0.97269 0.28368 0.079217 0.010821 4.7136 0.067524 8.199e-05 0.82256 0.0057013 0.006449 0.0013835 0.98698 0.99173 2.9829e-06 1.1931e-05 0.1354 0.95639 0.9207 0.0013956 0.9952 0.60873 0.0018803 0.43124 1.9255 1.925 15.9992 144.9925 0.00015797 -85.6638 0.88536
1.9894 0.98804 5.5131e-05 3.8182 0.012023 2.6148e-05 0.0011547 0.19284 0.00065892 0.19349 0.17756 0 0.034421 0.0389 0 0.97278 0.28373 0.079232 0.010823 4.7143 0.067535 8.2004e-05 0.82255 0.0057019 0.0064496 0.0013835 0.98698 0.99173 2.9829e-06 1.1931e-05 0.1354 0.95647 0.92074 0.0013956 0.99521 0.60887 0.0018803 0.43125 1.9259 1.9254 15.9992 144.9925 0.00015791 -85.6638 0.88636
1.9904 0.98804 5.5131e-05 3.8182 0.012023 2.6161e-05 0.0011547 0.19287 0.00065892 0.19353 0.17759 0 0.034419 0.0389 0 0.97288 0.28377 0.079247 0.010825 4.7151 0.067546 8.2019e-05 0.82254 0.0057025 0.0064502 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13541 0.95656 0.92077 0.0013956 0.99522 0.60901 0.0018803 0.43127 1.9262 1.9257 15.9992 144.9925 0.00015785 -85.6639 0.88736
1.9914 0.98804 5.5131e-05 3.8182 0.012023 2.6174e-05 0.0011547 0.19291 0.00065892 0.19356 0.17762 0 0.034417 0.0389 0 0.97297 0.28381 0.079262 0.010827 4.7158 0.067557 8.2034e-05 0.82253 0.0057031 0.0064509 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13541 0.95664 0.92081 0.0013956 0.99523 0.60914 0.0018803 0.43128 1.9265 1.926 15.9991 144.9925 0.00015779 -85.6639 0.88836
1.9924 0.98804 5.5131e-05 3.8182 0.012023 2.6187e-05 0.0011547 0.19294 0.00065892 0.19359 0.17765 0 0.034415 0.0389 0 0.97306 0.28385 0.079277 0.010828 4.7165 0.067568 8.2048e-05 0.82251 0.0057037 0.0064515 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13542 0.95673 0.92085 0.0013956 0.99525 0.60928 0.0018803 0.43129 1.9269 1.9264 15.9991 144.9926 0.00015773 -85.664 0.88936
1.9934 0.98804 5.5131e-05 3.8182 0.012023 2.6201e-05 0.0011547 0.19297 0.00065892 0.19363 0.17769 0 0.034413 0.0389 0 0.97316 0.28389 0.079292 0.01083 4.7173 0.067579 8.2062e-05 0.8225 0.0057043 0.0064521 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13542 0.95681 0.92089 0.0013956 0.99526 0.60941 0.0018803 0.4313 1.9272 1.9267 15.9991 144.9926 0.00015767 -85.664 0.89036
1.9944 0.98804 5.5131e-05 3.8182 0.012023 2.6214e-05 0.0011547 0.19301 0.00065892 0.19366 0.17772 0 0.034411 0.0389 0 0.97325 0.28394 0.079307 0.010832 4.718 0.06759 8.2077e-05 0.82249 0.0057049 0.0064528 0.0013835 0.98698 0.99173 2.9828e-06 1.1931e-05 0.13543 0.95689 0.92093 0.0013956 0.99527 0.60955 0.0018803 0.43131 1.9275 1.927 15.999 144.9926 0.00015761 -85.6641 0.89136
1.9954 0.98804 5.5131e-05 3.8182 0.012023 2.6227e-05 0.0011547 0.19304 0.00065892 0.1937 0.17775 0 0.034409 0.0389 0 0.97334 0.28398 0.079322 0.010834 4.7187 0.067601 8.2091e-05 0.82248 0.0057055 0.0064534 0.0013835 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13543 0.95698 0.92096 0.0013956 0.99528 0.60969 0.0018803 0.43132 1.9279 1.9274 15.999 144.9926 0.00015755 -85.6641 0.89236
1.9964 0.98804 5.5131e-05 3.8182 0.012023 2.624e-05 0.0011547 0.19308 0.00065892 0.19373 0.17778 0 0.034407 0.0389 0 0.97344 0.28402 0.079337 0.010835 4.7195 0.067612 8.2106e-05 0.82247 0.0057062 0.006454 0.0013835 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13544 0.95706 0.921 0.0013956 0.9953 0.60982 0.0018803 0.43133 1.9282 1.9277 15.999 144.9927 0.00015749 -85.6641 0.89336
1.9974 0.98804 5.5131e-05 3.8182 0.012023 2.6253e-05 0.0011547 0.19311 0.00065892 0.19376 0.17781 0 0.034405 0.0389 0 0.97353 0.28406 0.079352 0.010837 4.7202 0.067623 8.2121e-05 0.82246 0.0057068 0.0064547 0.0013834 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13544 0.95714 0.92104 0.0013956 0.99531 0.60996 0.0018803 0.43135 1.9286 1.9281 15.999 144.9927 0.00015743 -85.6642 0.89436
1.9984 0.98804 5.5131e-05 3.8182 0.012023 2.6266e-05 0.0011547 0.19314 0.00065892 0.1938 0.17785 0 0.034404 0.0389 0 0.97362 0.2841 0.079367 0.010839 4.7209 0.067634 8.2135e-05 0.82245 0.0057074 0.0064553 0.0013834 0.98698 0.99173 2.9827e-06 1.1931e-05 0.13545 0.95723 0.92108 0.0013956 0.99532 0.61009 0.0018803 0.43136 1.9289 1.9284 15.9989 144.9927 0.00015737 -85.6642 0.89536
1.9994 0.98804 5.513e-05 3.8182 0.012023 2.6279e-05 0.0011547 0.19318 0.00065892 0.19383 0.17788 0 0.034402 0.0389 0 0.97372 0.28415 0.079382 0.010841 4.7217 0.067645 8.2149e-05 0.82244 0.005708 0.0064559 0.0013834 0.98698 0.99173 2.9826e-06 1.193e-05 0.13545 0.95731 0.92111 0.0013956 0.99533 0.61023 0.0018802 0.43137 1.9292 1.9287 15.9989 144.9927 0.00015732 -85.6643 0.89636
2.0004 0.98804 5.513e-05 3.8182 0.012023 2.6292e-05 0.0011547 0.19321 0.00065892 0.19387 0.17791 0 0.0344 0.0389 0 0.97381 0.28419 0.079397 0.010843 4.7224 0.067656 8.2164e-05 0.82243 0.0057086 0.0064566 0.0013834 0.98698 0.99173 2.9826e-06 1.193e-05 0.13546 0.95739 0.92115 0.0013956 0.99535 0.61036 0.0018802 0.43138 1.9296 1.9291 15.9989 144.9927 0.00015726 -85.6643 0.89736
