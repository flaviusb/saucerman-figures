0 0.98801 5.5258e-005 3.8182 0.01205 0 0.001154 0.02505 0.0006446 0.02569 0.022413 0 0.047063 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0014 0.99 0.99 0 0 0.13 0.96 0.92 0.0014 1 0.613 0.198 0.43 1.92 1.92 16 145 0.000158 -85.66 0.9
0.001 0.98801 5.5256e-005 3.8182 0.01205 1.3187e-008 0.001154 0.025219 0.0006446 0.025859 0.022565 0 0.047046 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013826 0.98919 0.99011 2.9805e-006 1.1922e-005 0.13039 0.96007 0.92005 0.0013952 0.99998 0.61313 0.063153 0.43001 1.9204 1.9201 16 145 0.00015794 -85.6679 0.901
0.002 0.98801 5.5256e-005 3.8182 0.01205 2.6374e-008 0.001154 0.025387 0.00064461 0.026027 0.022717 0 0.047029 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013821 0.98859 0.99022 2.9797e-006 1.1919e-005 0.13043 0.96015 0.92009 0.0013949 0.99996 0.61327 0.021013 0.43002 1.9208 1.9203 15.9999 145 0.00015788 -85.6699 0.902
0.003 0.98801 5.5256e-005 3.8182 0.01205 3.9561e-008 0.001154 0.025556 0.00064462 0.026196 0.022868 0 0.047012 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013821 0.98816 0.99032 2.9796e-006 1.1918e-005 0.13044 0.96022 0.92014 0.0013949 0.99994 0.6134 0.0078539 0.43004 1.9211 1.9206 15.9999 145.0001 0.00015782 -85.67 0.903
0.004 0.98801 5.5256e-005 3.8182 0.01205 5.2748e-008 0.001154 0.025724 0.00064464 0.026364 0.02302 0 0.046995 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013822 0.98785 0.99041 2.9798e-006 1.1919e-005 0.13044 0.96029 0.92018 0.0013949 0.99993 0.61354 0.0037452 0.43005 1.9214 1.921 15.9999 145.0001 0.00015776 -85.6697 0.904
0.005 0.98801 5.5256e-005 3.8182 0.01205 6.5935e-008 0.001154 0.025892 0.00064465 0.026532 0.023171 0 0.046979 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013823 0.98762 0.9905 2.98e-006 1.192e-005 0.13044 0.96037 0.92023 0.001395 0.99991 0.61367 0.0024624 0.43006 1.9218 1.9213 15.9998 145.0001 0.0001577 -85.6693 0.905
0.006 0.98801 5.5256e-005 3.8182 0.01205 7.9122e-008 0.001154 0.02606 0.00064467 0.026701 0.023322 0 0.046962 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013824 0.98745 0.99058 2.9802e-006 1.1921e-005 0.13044 0.96044 0.92027 0.001395 0.99989 0.61381 0.0020617 0.43007 1.9221 1.9216 15.9998 145.0001 0.00015764 -85.6689 0.906
0.007 0.98801 5.5256e-005 3.8182 0.01205 9.2309e-008 0.001154 0.026228 0.00064469 0.026868 0.023473 0 0.046945 0.0389 0 0.8453 0.22699 0.05879 0.0083354 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013824 0.98733 0.99066 2.9804e-006 1.1921e-005 0.13044 0.96051 0.92032 0.0013951 0.99987 0.61394 0.0019367 0.43009 1.9224 1.9219 15.9998 145.0001 0.00015759 -85.6685 0.907
0.008 0.98801 5.5256e-005 3.8182 0.01205 1.055e-007 0.001154 0.026396 0.00064472 0.027036 0.023625 0 0.046928 0.0389 0 0.8453 0.22699 0.05879 0.0083355 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013825 0.98724 0.99073 2.9806e-006 1.1922e-005 0.13044 0.96058 0.92036 0.0013951 0.99986 0.61408 0.0018975 0.4301 1.9228 1.9223 15.9997 145.0002 0.00015753 -85.6682 0.908
0.009 0.98801 5.5256e-005 3.8182 0.01205 1.1868e-007 0.001154 0.026564 0.00064474 0.027204 0.023775 0 0.046912 0.0389 0 0.84531 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013826 0.98717 0.99079 2.9807e-006 1.1923e-005 0.13044 0.96065 0.9204 0.0013951 0.99984 0.61421 0.0018854 0.43011 1.9231 1.9226 15.9997 145.0002 0.00015747 -85.6679 0.909
0.01 0.98801 5.5255e-005 3.8182 0.01205 1.3187e-007 0.001154 0.026731 0.00064477 0.027372 0.023926 0 0.046895 0.0389 0 0.84531 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013826 0.98712 0.99086 2.9808e-006 1.1923e-005 0.13044 0.96073 0.92045 0.0013952 0.99982 0.61434 0.0018815 0.43012 1.9234 1.9229 15.9997 145.0002 0.00015741 -85.6677 0.91
0.011 0.98801 5.5255e-005 3.8182 0.01205 1.4506e-007 0.001154 0.026899 0.00064481 0.027539 0.024077 0 0.046878 0.0389 0 0.84531 0.227 0.058791 0.0083355 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013827 0.98709 0.99091 2.981e-006 1.1924e-005 0.13044 0.9608 0.92049 0.0013952 0.9998 0.61448 0.0018803 0.43013 1.9238 1.9233 15.9996 145.0002 0.00015735 -85.6675 0.911
0.012 0.98801 5.5255e-005 3.8182 0.01205 1.5824e-007 0.001154 0.027066 0.00064484 0.027706 0.024228 0 0.046862 0.0389 0 0.84531 0.227 0.058791 0.0083356 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013827 0.98706 0.99097 2.981e-006 1.1924e-005 0.13044 0.96087 0.92054 0.0013952 0.99979 0.61461 0.0018799 0.43015 1.9241 1.9236 15.9996 145.0002 0.0001573 -85.6673 0.912
0.013 0.98801 5.5255e-005 3.8182 0.01205 1.7143e-007 0.001154 0.027233 0.00064488 0.027873 0.024378 0 0.046845 0.0389 0 0.84531 0.227 0.058792 0.0083356 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013828 0.98704 0.99102 2.9811e-006 1.1924e-005 0.13044 0.96094 0.92058 0.0013952 0.99977 0.61475 0.0018798 0.43016 1.9244 1.9239 15.9996 145.0003 0.00015724 -85.6671 0.913
0.014 0.98801 5.5255e-005 3.8182 0.01205 1.8462e-007 0.001154 0.0274 0.00064491 0.02804 0.024529 0 0.046828 0.0389 0 0.84531 0.227 0.058792 0.0083356 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013828 0.98703 0.99106 2.9812e-006 1.1925e-005 0.13044 0.96101 0.92062 0.0013952 0.99975 0.61488 0.0018798 0.43017 1.9247 1.9243 15.9996 145.0003 0.00015718 -85.667 0.914
0.015 0.98801 5.5255e-005 3.8182 0.01205 1.978e-007 0.001154 0.027567 0.00064495 0.028207 0.024679 0 0.046812 0.0389 0 0.84531 0.227 0.058792 0.0083357 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013828 0.98702 0.99111 2.9812e-006 1.1925e-005 0.13044 0.96108 0.92067 0.0013953 0.99973 0.61502 0.0018798 0.43018 1.9251 1.9246 15.9995 145.0003 0.00015712 -85.6669 0.915
0.016 0.98801 5.5255e-005 3.8182 0.01205 2.1099e-007 0.001154 0.027734 0.00064499 0.028374 0.024829 0 0.046795 0.0389 0 0.84532 0.227 0.058792 0.0083357 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013828 0.98701 0.99115 2.9813e-006 1.1925e-005 0.13044 0.96115 0.92071 0.0013953 0.99972 0.61515 0.0018798 0.43019 1.9254 1.9249 15.9995 145.0003 0.00015707 -85.6668 0.916
0.017 0.98801 5.5255e-005 3.8182 0.01205 2.2418e-007 0.001154 0.0279 0.00064504 0.028541 0.024979 0 0.046779 0.0389 0 0.84532 0.227 0.058793 0.0083358 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.987 0.99119 2.9813e-006 1.1925e-005 0.13044 0.96122 0.92075 0.0013953 0.9997 0.61528 0.0018798 0.43021 1.9257 1.9252 15.9995 145.0003 0.00015701 -85.6667 0.917
0.018 0.98801 5.5255e-005 3.8182 0.01205 2.3736e-007 0.001154 0.028067 0.00064508 0.028707 0.025129 0 0.046762 0.0389 0 0.84532 0.227 0.058793 0.0083358 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.987 0.99122 2.9814e-006 1.1925e-005 0.13044 0.96129 0.92079 0.0013953 0.99968 0.61542 0.0018799 0.43022 1.9261 1.9256 15.9994 145.0004 0.00015695 -85.6667 0.918
0.019 0.98801 5.5255e-005 3.8182 0.01205 2.5055e-007 0.001154 0.028233 0.00064513 0.028874 0.025279 0 0.046746 0.0389 0 0.84532 0.227 0.058794 0.0083358 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.987 0.99126 2.9814e-006 1.1925e-005 0.13044 0.96136 0.92084 0.0013953 0.99967 0.61555 0.0018799 0.43023 1.9264 1.9259 15.9994 145.0004 0.0001569 -85.6666 0.919
0.02 0.98801 5.5255e-005 3.8182 0.01205 2.6374e-007 0.001154 0.028399 0.00064518 0.02904 0.025429 0 0.046729 0.0389 0 0.84533 0.227 0.058794 0.0083359 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99129 2.9814e-006 1.1926e-005 0.13044 0.96143 0.92088 0.0013953 0.99965 0.61568 0.0018799 0.43024 1.9267 1.9262 15.9994 145.0004 0.00015684 -85.6666 0.92
0.021 0.98801 5.5255e-005 3.8182 0.01205 2.7692e-007 0.001154 0.028565 0.00064523 0.029206 0.025578 0 0.046713 0.0389 0 0.84533 0.22701 0.058794 0.0083359 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99132 2.9814e-006 1.1926e-005 0.13044 0.9615 0.92092 0.0013953 0.99964 0.61582 0.0018799 0.43026 1.927 1.9265 15.9993 145.0004 0.00015679 -85.6666 0.921
0.022 0.98801 5.5255e-005 3.8182 0.01205 2.9011e-007 0.001154 0.028731 0.00064528 0.029372 0.025728 0 0.046697 0.0389 0 0.84533 0.22701 0.058795 0.008336 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99134 2.9814e-006 1.1926e-005 0.13044 0.96157 0.92096 0.0013953 0.99962 0.61595 0.0018799 0.43027 1.9274 1.9269 15.9993 145.0005 0.00015673 -85.6666 0.922
0.023 0.98801 5.5255e-005 3.8182 0.01205 3.0329e-007 0.001154 0.028897 0.00064533 0.029538 0.025877 0 0.04668 0.0389 0 0.84533 0.22701 0.058795 0.0083361 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99137 2.9814e-006 1.1926e-005 0.13044 0.96164 0.921 0.0013953 0.9996 0.61609 0.0018799 0.43028 1.9277 1.9272 15.9993 145.0005 0.00015668 -85.6665 0.923
0.024 0.98801 5.5255e-005 3.8182 0.01205 3.1648e-007 0.001154 0.029063 0.00064539 0.029704 0.026027 0 0.046664 0.0389 0 0.84534 0.22701 0.058796 0.0083361 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99139 2.9814e-006 1.1926e-005 0.13044 0.9617 0.92104 0.0013953 0.99959 0.61622 0.0018799 0.43029 1.928 1.9275 15.9992 145.0005 0.00015662 -85.6665 0.924
0.025 0.98801 5.5255e-005 3.8182 0.01205 3.2967e-007 0.001154 0.029228 0.00064544 0.029869 0.026176 0 0.046647 0.0389 0 0.84534 0.22701 0.058796 0.0083362 4.105 0.0526 6.2734e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99142 2.9814e-006 1.1926e-005 0.13044 0.96177 0.92109 0.0013953 0.99957 0.61635 0.0018799 0.4303 1.9283 1.9278 15.9992 145.0005 0.00015656 -85.6665 0.925
0.026 0.98801 5.5254e-005 3.8182 0.01205 3.4285e-007 0.001154 0.029394 0.0006455 0.030035 0.026325 0 0.046631 0.0389 0 0.84534 0.22701 0.058797 0.0083363 4.105 0.052601 6.2735e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99144 2.9814e-006 1.1926e-005 0.13044 0.96184 0.92113 0.0013953 0.99956 0.61649 0.0018799 0.43032 1.9286 1.9282 15.9992 145.0005 0.00015651 -85.6665 0.926
0.027 0.98801 5.5254e-005 3.8182 0.01205 3.5604e-007 0.001154 0.029559 0.00064555 0.0302 0.026474 0 0.046615 0.0389 0 0.84535 0.22701 0.058797 0.0083363 4.105 0.052601 6.2735e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99146 2.9814e-006 1.1926e-005 0.13044 0.96191 0.92117 0.0013953 0.99954 0.61662 0.0018799 0.43033 1.929 1.9285 15.9991 145.0006 0.00015646 -85.6665 0.927
0.028 0.98801 5.5254e-005 3.8182 0.01205 3.6922e-007 0.001154 0.029724 0.00064561 0.030365 0.026623 0 0.046599 0.0389 0 0.84535 0.22702 0.058798 0.0083364 4.105 0.052601 6.2735e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99147 2.9814e-006 1.1926e-005 0.13044 0.96198 0.92121 0.0013953 0.99953 0.61675 0.0018799 0.43034 1.9293 1.9288 15.9991 145.0006 0.0001564 -85.6665 0.928
0.029 0.98801 5.5254e-005 3.8182 0.01205 3.8241e-007 0.001154 0.029889 0.00064567 0.03053 0.026771 0 0.046582 0.0389 0 0.84535 0.22702 0.058798 0.0083365 4.105 0.052601 6.2735e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99149 2.9814e-006 1.1926e-005 0.13044 0.96204 0.92125 0.0013953 0.99951 0.61689 0.0018799 0.43035 1.9296 1.9291 15.9991 145.0006 0.00015635 -85.6666 0.929
0.03 0.98801 5.5254e-005 3.8182 0.01205 3.956e-007 0.001154 0.030054 0.00064573 0.030695 0.02692 0 0.046566 0.0389 0 0.84536 0.22702 0.058799 0.0083365 4.105 0.052601 6.2735e-005 0.83746 0.005103 0.005841 0.0013829 0.98699 0.99151 2.9814e-006 1.1926e-005 0.13044 0.96211 0.92129 0.0013953 0.99949 0.61702 0.0018799 0.43036 1.9299 1.9295 15.999 145.0006 0.00015629 -85.6666 0.93
0.031 0.98801 5.5254e-005 3.8182 0.01205 4.0878e-007 0.001154 0.030219 0.00064579 0.03086 0.027069 0 0.04655 0.0389 0 0.84536 0.22702 0.0588 0.0083366 4.105 0.052601 6.2735e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99152 2.9814e-006 1.1926e-005 0.13044 0.96218 0.92133 0.0013953 0.99948 0.61715 0.0018799 0.43038 1.9303 1.9298 15.999 145.0006 0.00015624 -85.6666 0.931
0.032 0.98801 5.5254e-005 3.8182 0.01205 4.2197e-007 0.001154 0.030383 0.00064585 0.031025 0.027217 0 0.046534 0.0389 0 0.84537 0.22702 0.0588 0.0083367 4.105 0.052601 6.2735e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99154 2.9814e-006 1.1926e-005 0.13044 0.96224 0.92137 0.0013953 0.99946 0.61729 0.0018799 0.43039 1.9306 1.9301 15.999 145.0007 0.00015618 -85.6666 0.932
0.033 0.98801 5.5254e-005 3.8182 0.01205 4.3515e-007 0.001154 0.030548 0.00064591 0.031189 0.027365 0 0.046518 0.0389 0 0.84537 0.22702 0.058801 0.0083368 4.105 0.052601 6.2735e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99155 2.9814e-006 1.1925e-005 0.13044 0.96231 0.92141 0.0013953 0.99945 0.61742 0.0018799 0.4304 1.9309 1.9304 15.9989 145.0007 0.00015613 -85.6666 0.933
0.034 0.98801 5.5254e-005 3.8182 0.01205 4.4834e-007 0.001154 0.030712 0.00064598 0.031353 0.027514 0 0.046501 0.0389 0 0.84537 0.22703 0.058802 0.0083369 4.105 0.052601 6.2735e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99156 2.9814e-006 1.1925e-005 0.13044 0.96238 0.92145 0.0013953 0.99943 0.61755 0.0018799 0.43041 1.9312 1.9307 15.9989 145.0007 0.00015608 -85.6666 0.934
0.035 0.98801 5.5254e-005 3.8182 0.01205 4.6152e-007 0.001154 0.030876 0.00064604 0.031518 0.027662 0 0.046485 0.0389 0 0.84538 0.22703 0.058802 0.008337 4.105 0.052601 6.2736e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99157 2.9814e-006 1.1925e-005 0.13044 0.96244 0.92149 0.0013953 0.99942 0.61769 0.0018799 0.43042 1.9315 1.9311 15.9989 145.0007 0.00015602 -85.6667 0.935
0.036 0.98801 5.5254e-005 3.8182 0.01205 4.7471e-007 0.001154 0.03104 0.0006461 0.031682 0.02781 0 0.046469 0.0389 0 0.84538 0.22703 0.058803 0.0083371 4.105 0.052602 6.2736e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99158 2.9814e-006 1.1925e-005 0.13044 0.96251 0.92153 0.0013953 0.9994 0.61782 0.0018799 0.43044 1.9318 1.9314 15.9988 145.0007 0.00015597 -85.6667 0.936
0.037 0.98801 5.5254e-005 3.8182 0.01205 4.879e-007 0.001154 0.031204 0.00064617 0.031846 0.027958 0 0.046453 0.0389 0 0.84539 0.22703 0.058804 0.0083371 4.105 0.052602 6.2736e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.99159 2.9813e-006 1.1925e-005 0.13044 0.96257 0.92156 0.0013953 0.99939 0.61795 0.0018799 0.43045 1.9322 1.9317 15.9988 145.0008 0.00015592 -85.6667 0.937
0.038 0.98801 5.5254e-005 3.8182 0.012049 5.0108e-007 0.001154 0.031368 0.00064623 0.03201 0.028105 0 0.046437 0.0389 0 0.84539 0.22703 0.058805 0.0083372 4.105 0.052602 6.2736e-005 0.83746 0.0051031 0.0058411 0.0013829 0.98699 0.9916 2.9813e-006 1.1925e-005 0.13044 0.96264 0.9216 0.0013953 0.99938 0.61809 0.0018799 0.43046 1.9325 1.932 15.9988 145.0008 0.00015586 -85.6667 0.938
0.039 0.98801 5.5254e-005 3.8182 0.012049 5.1427e-007 0.001154 0.031532 0.0006463 0.032174 0.028253 0 0.046421 0.0389 0 0.8454 0.22704 0.058805 0.0083373 4.105 0.052602 6.2736e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99161 2.9813e-006 1.1925e-005 0.13044 0.96271 0.92164 0.0013953 0.99936 0.61822 0.0018798 0.43047 1.9328 1.9323 15.9987 145.0008 0.00015581 -85.6668 0.939
0.04 0.98801 5.5254e-005 3.8182 0.012049 5.2745e-007 0.001154 0.031695 0.00064636 0.032337 0.028401 0 0.046405 0.0389 0 0.8454 0.22704 0.058806 0.0083374 4.105 0.052602 6.2737e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99162 2.9813e-006 1.1925e-005 0.13044 0.96277 0.92168 0.0013953 0.99935 0.61835 0.0018798 0.43048 1.9331 1.9326 15.9987 145.0008 0.00015576 -85.6668 0.94
0.041 0.98801 5.5254e-005 3.8182 0.012049 5.4064e-007 0.001154 0.031859 0.00064643 0.032501 0.028548 0 0.046389 0.0389 0 0.84541 0.22704 0.058807 0.0083375 4.105 0.052602 6.2737e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99163 2.9813e-006 1.1925e-005 0.13044 0.96284 0.92172 0.0013953 0.99933 0.61848 0.0018798 0.4305 1.9334 1.933 15.9987 145.0008 0.00015571 -85.6668 0.941
0.042 0.98801 5.5254e-005 3.8182 0.012049 5.5382e-007 0.001154 0.032022 0.00064649 0.032664 0.028695 0 0.046373 0.0389 0 0.84541 0.22704 0.058808 0.0083377 4.105 0.052602 6.2737e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99163 2.9813e-006 1.1925e-005 0.13044 0.9629 0.92176 0.0013953 0.99932 0.61862 0.0018798 0.43051 1.9337 1.9333 15.9986 145.0009 0.00015565 -85.6668 0.942
0.043 0.98801 5.5253e-005 3.8182 0.012049 5.6701e-007 0.001154 0.032185 0.00064656 0.032827 0.028843 0 0.046357 0.0389 0 0.84542 0.22705 0.058809 0.0083378 4.105 0.052603 6.2737e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99164 2.9813e-006 1.1925e-005 0.13044 0.96296 0.9218 0.0013953 0.9993 0.61875 0.0018798 0.43052 1.934 1.9336 15.9986 145.0009 0.0001556 -85.6669 0.943
0.044 0.98801 5.5253e-005 3.8182 0.012049 5.8019e-007 0.001154 0.032348 0.00064663 0.03299 0.02899 0 0.046341 0.0389 0 0.84542 0.22705 0.05881 0.0083379 4.105 0.052603 6.2737e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99165 2.9813e-006 1.1925e-005 0.13044 0.96303 0.92183 0.0013953 0.99929 0.61888 0.0018798 0.43053 1.9344 1.9339 15.9986 145.0009 0.00015555 -85.6669 0.944
0.045 0.98801 5.5253e-005 3.8182 0.012049 5.9338e-007 0.001154 0.032511 0.00064669 0.033153 0.029137 0 0.046326 0.0389 0 0.84543 0.22705 0.05881 0.008338 4.1051 0.052603 6.2738e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99165 2.9812e-006 1.1925e-005 0.13044 0.96309 0.92187 0.0013952 0.99928 0.61901 0.0018798 0.43054 1.9347 1.9342 15.9985 145.0009 0.0001555 -85.6669 0.945
0.046 0.98801 5.5253e-005 3.8182 0.012049 6.0656e-007 0.001154 0.032674 0.00064676 0.033316 0.029284 0 0.04631 0.0389 0 0.84544 0.22705 0.058811 0.0083381 4.1051 0.052603 6.2738e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99166 2.9812e-006 1.1925e-005 0.13044 0.96316 0.92191 0.0013952 0.99926 0.61915 0.0018798 0.43056 1.935 1.9345 15.9985 145.0009 0.00015545 -85.667 0.946
0.047 0.98801 5.5253e-005 3.8182 0.012049 6.1975e-007 0.001154 0.032837 0.00064683 0.033479 0.02943 0 0.046294 0.0389 0 0.84544 0.22706 0.058812 0.0083382 4.1051 0.052603 6.2738e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99166 2.9812e-006 1.1925e-005 0.13044 0.96322 0.92195 0.0013952 0.99925 0.61928 0.0018798 0.43057 1.9353 1.9348 15.9985 145.001 0.0001554 -85.667 0.947
0.048 0.98801 5.5253e-005 3.8182 0.012049 6.3293e-007 0.001154 0.032999 0.00064689 0.033641 0.029577 0 0.046278 0.0389 0 0.84545 0.22706 0.058813 0.0083383 4.1051 0.052604 6.2738e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99167 2.9812e-006 1.1925e-005 0.13044 0.96328 0.92198 0.0013952 0.99924 0.61941 0.0018798 0.43058 1.9356 1.9351 15.9984 145.001 0.00015535 -85.667 0.948
0.049 0.98801 5.5253e-005 3.8182 0.012049 6.4612e-007 0.001154 0.033161 0.00064696 0.033804 0.029724 0 0.046262 0.0389 0 0.84545 0.22706 0.058814 0.0083385 4.1051 0.052604 6.2739e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99167 2.9812e-006 1.1925e-005 0.13044 0.96335 0.92202 0.0013952 0.99922 0.61954 0.0018798 0.43059 1.9359 1.9355 15.9984 145.001 0.00015529 -85.667 0.949
0.05 0.98801 5.5253e-005 3.8182 0.012049 6.593e-007 0.001154 0.033324 0.00064703 0.033966 0.02987 0 0.046247 0.0389 0 0.84546 0.22706 0.058815 0.0083386 4.1051 0.052604 6.2739e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99167 2.9812e-006 1.1925e-005 0.13044 0.96341 0.92206 0.0013952 0.99921 0.61968 0.0018798 0.4306 1.9362 1.9358 15.9984 145.001 0.00015524 -85.6671 0.95
0.051 0.98801 5.5253e-005 3.8182 0.012049 6.7249e-007 0.001154 0.033486 0.00064709 0.034128 0.030017 0 0.046231 0.0389 0 0.84547 0.22707 0.058816 0.0083387 4.1051 0.052604 6.2739e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99168 2.9812e-006 1.1925e-005 0.13044 0.96347 0.92209 0.0013952 0.9992 0.61981 0.0018798 0.43061 1.9365 1.9361 15.9983 145.001 0.00015519 -85.6671 0.951
0.052 0.98801 5.5253e-005 3.8182 0.012049 6.8567e-007 0.001154 0.033648 0.00064716 0.03429 0.030163 0 0.046215 0.0389 0 0.84547 0.22707 0.058817 0.0083389 4.1051 0.052605 6.274e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99168 2.9811e-006 1.1924e-005 0.13044 0.96354 0.92213 0.0013952 0.99918 0.61994 0.0018798 0.43063 1.9368 1.9364 15.9983 145.0011 0.00015514 -85.6671 0.952
0.053 0.98801 5.5253e-005 3.8182 0.012049 6.9886e-007 0.001154 0.03381 0.00064723 0.034452 0.030309 0 0.046199 0.0389 0 0.84548 0.22707 0.058818 0.008339 4.1051 0.052605 6.274e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99169 2.9811e-006 1.1924e-005 0.13044 0.9636 0.92217 0.0013952 0.99917 0.62007 0.0018798 0.43064 1.9372 1.9367 15.9983 145.0011 0.00015509 -85.6671 0.953
0.054 0.98801 5.5253e-005 3.8182 0.012049 7.1204e-007 0.001154 0.033971 0.00064729 0.034614 0.030455 0 0.046184 0.0389 0 0.84549 0.22708 0.058819 0.0083391 4.1051 0.052605 6.274e-005 0.83746 0.0051031 0.0058411 0.0013828 0.98699 0.99169 2.9811e-006 1.1924e-005 0.13044 0.96366 0.9222 0.0013952 0.99916 0.62021 0.0018798 0.43065 1.9375 1.937 15.9982 145.0011 0.00015504 -85.6672 0.954
0.055 0.98801 5.5253e-005 3.8182 0.012049 7.2523e-007 0.001154 0.034133 0.00064736 0.034776 0.030601 0 0.046168 0.0389 0 0.84549 0.22708 0.058821 0.0083393 4.1051 0.052605 6.2741e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99169 2.9811e-006 1.1924e-005 0.13044 0.96372 0.92224 0.0013952 0.99914 0.62034 0.0018798 0.43066 1.9378 1.9373 15.9982 145.0011 0.00015499 -85.6672 0.955
0.056 0.98801 5.5253e-005 3.8182 0.012049 7.3841e-007 0.001154 0.034294 0.00064743 0.034937 0.030747 0 0.046152 0.0389 0 0.8455 0.22708 0.058822 0.0083394 4.1051 0.052606 6.2741e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99169 2.9811e-006 1.1924e-005 0.13044 0.96379 0.92228 0.0013952 0.99913 0.62047 0.0018798 0.43067 1.9381 1.9376 15.9982 145.0011 0.00015494 -85.6672 0.956
0.057 0.98801 5.5253e-005 3.8182 0.012049 7.516e-007 0.001154 0.034456 0.00064749 0.035099 0.030893 0 0.046137 0.0389 0 0.84551 0.22708 0.058823 0.0083395 4.1051 0.052606 6.2741e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.9811e-006 1.1924e-005 0.13044 0.96385 0.92231 0.0013952 0.99912 0.6206 0.0018798 0.43069 1.9384 1.9379 15.9981 145.0012 0.00015489 -85.6673 0.957
0.058 0.98801 5.5253e-005 3.8182 0.012049 7.6478e-007 0.001154 0.034617 0.00064756 0.03526 0.031038 0 0.046121 0.0389 0 0.84552 0.22709 0.058824 0.0083397 4.1051 0.052606 6.2742e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.9811e-006 1.1924e-005 0.13044 0.96391 0.92235 0.0013952 0.9991 0.62073 0.0018798 0.4307 1.9387 1.9382 15.9981 145.0012 0.00015484 -85.6673 0.958
0.059 0.98801 5.5252e-005 3.8182 0.012049 7.7797e-007 0.001154 0.034778 0.00064762 0.035421 0.031184 0 0.046106 0.0389 0 0.84552 0.22709 0.058825 0.0083398 4.1051 0.052607 6.2742e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.981e-006 1.1924e-005 0.13044 0.96397 0.92238 0.0013952 0.99909 0.62087 0.0018798 0.43071 1.939 1.9385 15.9981 145.0012 0.00015479 -85.6673 0.959
0.06 0.98801 5.5252e-005 3.8182 0.012049 7.9115e-007 0.001154 0.034939 0.00064769 0.035582 0.031329 0 0.04609 0.0389 0 0.84553 0.22709 0.058826 0.00834 4.1051 0.052607 6.2743e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.9917 2.981e-006 1.1924e-005 0.13044 0.96403 0.92242 0.0013952 0.99908 0.621 0.0018798 0.43072 1.9393 1.9389 15.998 145.0012 0.00015474 -85.6673 0.96
0.061 0.98801 5.5252e-005 3.8182 0.012049 8.0434e-007 0.001154 0.0351 0.00064775 0.035743 0.031474 0 0.046075 0.0389 0 0.84554 0.2271 0.058828 0.0083401 4.1051 0.052607 6.2743e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-006 1.1924e-005 0.13044 0.96409 0.92245 0.0013952 0.99907 0.62113 0.0018798 0.43073 1.9396 1.9392 15.998 145.0013 0.0001547 -85.6674 0.961
0.062 0.98801 5.5252e-005 3.8182 0.012049 8.1752e-007 0.001154 0.035261 0.00064782 0.035904 0.03162 0 0.046059 0.0389 0 0.84555 0.2271 0.058829 0.0083403 4.1051 0.052608 6.2743e-005 0.83746 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-006 1.1924e-005 0.13044 0.96415 0.92249 0.0013952 0.99905 0.62126 0.0018798 0.43075 1.9399 1.9395 15.998 145.0013 0.00015465 -85.6674 0.962
0.063 0.98801 5.5252e-005 3.8182 0.012049 8.3071e-007 0.001154 0.035421 0.00064788 0.036064 0.031765 0 0.046044 0.0389 0 0.84555 0.2271 0.05883 0.0083405 4.1051 0.052608 6.2744e-005 0.83745 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-006 1.1924e-005 0.13044 0.96421 0.92252 0.0013952 0.99904 0.62139 0.0018797 0.43076 1.9402 1.9398 15.9979 145.0013 0.0001546 -85.6674 0.963
0.064 0.98801 5.5252e-005 3.8182 0.012049 8.4389e-007 0.001154 0.035582 0.00064795 0.036225 0.03191 0 0.046028 0.0389 0 0.84556 0.22711 0.058831 0.0083406 4.1051 0.052608 6.2744e-005 0.83745 0.0051031 0.0058411 0.0013827 0.98699 0.99171 2.981e-006 1.1924e-005 0.13044 0.96427 0.92256 0.0013952 0.99903 0.62153 0.0018797 0.43077 1.9405 1.9401 15.9979 145.0013 0.00015455 -85.6674 0.964
0.065 0.98801 5.5252e-005 3.8182 0.012049 8.5708e-007 0.001154 0.035742 0.00064801 0.036385 0.032055 0 0.046013 0.0389 0 0.84557 0.22711 0.058833 0.0083408 4.1051 0.052609 6.2745e-005 0.83745 0.0051032 0.0058411 0.0013827 0.98699 0.99171 2.981e-006 1.1924e-005 0.13044 0.96433 0.92259 0.0013952 0.99902 0.62166 0.0018797 0.43078 1.9408 1.9404 15.9979 145.0013 0.0001545 -85.6675 0.965
0.066 0.98801 5.5252e-005 3.8182 0.012049 8.7026e-007 0.001154 0.035902 0.00064808 0.036546 0.032199 0 0.045997 0.0389 0 0.84558 0.22712 0.058834 0.0083409 4.1051 0.052609 6.2745e-005 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99171 2.9809e-006 1.1924e-005 0.13044 0.96439 0.92263 0.0013952 0.99901 0.62179 0.0018797 0.43079 1.9411 1.9407 15.9979 145.0014 0.00015445 -85.6675 0.966
0.067 0.98801 5.5252e-005 3.8182 0.012049 8.8344e-007 0.001154 0.036062 0.00064814 0.036706 0.032344 0 0.045982 0.0389 0 0.84559 0.22712 0.058835 0.0083411 4.1051 0.052609 6.2746e-005 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-006 1.1924e-005 0.13044 0.96445 0.92266 0.0013952 0.99899 0.62192 0.0018797 0.4308 1.9414 1.941 15.9978 145.0014 0.0001544 -85.6675 0.967
0.068 0.98801 5.5252e-005 3.8182 0.012049 8.9663e-007 0.001154 0.036222 0.0006482 0.036866 0.032489 0 0.045967 0.0389 0 0.84559 0.22712 0.058837 0.0083413 4.1051 0.05261 6.2746e-005 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-006 1.1924e-005 0.13044 0.96451 0.9227 0.0013952 0.99898 0.62205 0.0018797 0.43082 1.9417 1.9413 15.9978 145.0014 0.00015436 -85.6675 0.968
0.069 0.98801 5.5252e-005 3.8182 0.012049 9.0981e-007 0.001154 0.036382 0.00064827 0.037025 0.032633 0 0.045951 0.0389 0 0.8456 0.22713 0.058838 0.0083415 4.1051 0.05261 6.2747e-005 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-006 1.1924e-005 0.13044 0.96457 0.92273 0.0013952 0.99897 0.62218 0.0018797 0.43083 1.942 1.9416 15.9978 145.0014 0.00015431 -85.6676 0.969
0.07 0.98801 5.5252e-005 3.8182 0.012049 9.23e-007 0.001154 0.036541 0.00064833 0.037185 0.032777 0 0.045936 0.0389 0 0.84561 0.22713 0.058839 0.0083416 4.1051 0.052611 6.2747e-005 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-006 1.1923e-005 0.13044 0.96463 0.92276 0.0013952 0.99896 0.62231 0.0018797 0.43084 1.9423 1.9419 15.9977 145.0014 0.00015426 -85.6676 0.97
0.071 0.98801 5.5252e-005 3.8182 0.012049 9.3618e-007 0.001154 0.036701 0.00064839 0.037345 0.032922 0 0.045921 0.0389 0 0.84562 0.22713 0.058841 0.0083418 4.1051 0.052611 6.2748e-005 0.83745 0.0051032 0.0058412 0.0013827 0.98699 0.99172 2.9809e-006 1.1923e-005 0.13044 0.96469 0.9228 0.0013952 0.99895 0.62245 0.0018797 0.43085 1.9426 1.9422 15.9977 145.0015 0.00015421 -85.6676 0.971
0.072 0.98801 5.5252e-005 3.8182 0.012049 9.4936e-007 0.001154 0.03686 0.00064845 0.037504 0.033066 0 0.045905 0.0389 0 0.84563 0.22714 0.058842 0.008342 4.1051 0.052612 6.2748e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9809e-006 1.1923e-005 0.13044 0.96475 0.92283 0.0013952 0.99893 0.62258 0.0018797 0.43086 1.9429 1.9425 15.9977 145.0015 0.00015417 -85.6676 0.972
0.073 0.98801 5.5252e-005 3.8182 0.012049 9.6255e-007 0.001154 0.03702 0.00064851 0.037664 0.03321 0 0.04589 0.0389 0 0.84564 0.22714 0.058844 0.0083422 4.1051 0.052612 6.2749e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9809e-006 1.1923e-005 0.13044 0.96481 0.92287 0.0013952 0.99892 0.62271 0.0018797 0.43088 1.9432 1.9428 15.9976 145.0015 0.00015412 -85.6677 0.973
0.074 0.98801 5.5252e-005 3.8182 0.012049 9.7573e-007 0.001154 0.037179 0.00064857 0.037823 0.033354 0 0.045875 0.0389 0 0.84565 0.22715 0.058845 0.0083424 4.1051 0.052612 6.275e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-006 1.1923e-005 0.13044 0.96487 0.9229 0.0013952 0.99891 0.62284 0.0018797 0.43089 1.9435 1.9431 15.9976 145.0015 0.00015407 -85.6677 0.974
0.075 0.98801 5.5251e-005 3.8182 0.012049 9.8892e-007 0.001154 0.037338 0.00064863 0.037982 0.033497 0 0.04586 0.0389 0 0.84566 0.22715 0.058846 0.0083425 4.1051 0.052613 6.275e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-006 1.1923e-005 0.13044 0.96493 0.92293 0.0013952 0.9989 0.62297 0.0018797 0.4309 1.9438 1.9434 15.9976 145.0015 0.00015403 -85.6677 0.975
0.076 0.98801 5.5251e-005 3.8182 0.012049 1.0021e-006 0.001154 0.037497 0.00064869 0.038141 0.033641 0 0.045844 0.0389 0 0.84567 0.22715 0.058848 0.0083427 4.1051 0.052613 6.2751e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-006 1.1923e-005 0.13044 0.96498 0.92297 0.0013952 0.99889 0.6231 0.0018797 0.43091 1.9441 1.9437 15.9975 145.0016 0.00015398 -85.6677 0.976
0.077 0.98801 5.5251e-005 3.8182 0.012049 1.0153e-006 0.001154 0.037656 0.00064875 0.0383 0.033785 0 0.045829 0.0389 0 0.84568 0.22716 0.058849 0.0083429 4.1051 0.052614 6.2751e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99172 2.9808e-006 1.1923e-005 0.13044 0.96504 0.923 0.0013951 0.99888 0.62323 0.0018797 0.43092 1.9444 1.944 15.9975 145.0016 0.00015393 -85.6677 0.977
0.078 0.98801 5.5251e-005 3.8182 0.012049 1.0285e-006 0.001154 0.037814 0.00064881 0.038458 0.033928 0 0.045814 0.0389 0 0.84569 0.22716 0.058851 0.0083431 4.1051 0.052614 6.2752e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13044 0.9651 0.92303 0.0013951 0.99887 0.62337 0.0018797 0.43093 1.9447 1.9443 15.9975 145.0016 0.00015389 -85.6678 0.978
0.079 0.98801 5.5251e-005 3.8182 0.012049 1.0417e-006 0.001154 0.037973 0.00064887 0.038617 0.034072 0 0.045799 0.0389 0 0.8457 0.22717 0.058853 0.0083433 4.1051 0.052615 6.2753e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13044 0.96516 0.92306 0.0013951 0.99886 0.6235 0.0018797 0.43095 1.945 1.9446 15.9974 145.0016 0.00015384 -85.6678 0.979
0.08 0.98801 5.5251e-005 3.8182 0.012049 1.0548e-006 0.001154 0.038131 0.00064893 0.038775 0.034215 0 0.045784 0.0389 0 0.84571 0.22717 0.058854 0.0083435 4.1051 0.052615 6.2753e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13044 0.96521 0.9231 0.0013951 0.99884 0.62363 0.0018797 0.43096 1.9453 1.9449 15.9974 145.0016 0.00015379 -85.6678 0.98
0.081 0.98801 5.5251e-005 3.8182 0.012049 1.068e-006 0.001154 0.038289 0.00064899 0.038934 0.034358 0 0.045769 0.0389 0 0.84572 0.22718 0.058856 0.0083437 4.1051 0.052616 6.2754e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13044 0.96527 0.92313 0.0013951 0.99883 0.62376 0.0018797 0.43097 1.9456 1.9452 15.9973 145.0017 0.00015375 -85.6678 0.981
0.082 0.98801 5.5251e-005 3.8182 0.012049 1.0812e-006 0.001154 0.038448 0.00064905 0.039092 0.034501 0 0.045754 0.0389 0 0.84573 0.22718 0.058857 0.0083439 4.1051 0.052616 6.2755e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96533 0.92316 0.0013951 0.99882 0.62389 0.0018797 0.43098 1.9459 1.9455 15.9973 145.0017 0.0001537 -85.6679 0.982
0.083 0.98801 5.5251e-005 3.8182 0.012049 1.0944e-006 0.001154 0.038606 0.0006491 0.03925 0.034644 0 0.045739 0.0389 0 0.84574 0.22719 0.058859 0.0083441 4.1052 0.052617 6.2755e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96539 0.92319 0.0013951 0.99881 0.62402 0.0018797 0.43099 1.9462 1.9458 15.9973 145.0017 0.00015366 -85.6679 0.983
0.084 0.98801 5.5251e-005 3.8182 0.012049 1.1076e-006 0.001154 0.038763 0.00064916 0.039408 0.034787 0 0.045724 0.0389 0 0.84575 0.22719 0.058861 0.0083443 4.1052 0.052618 6.2756e-005 0.83745 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96544 0.92323 0.0013951 0.9988 0.62415 0.0018797 0.43101 1.9465 1.9461 15.9972 145.0017 0.00015361 -85.6679 0.984
0.085 0.98801 5.5251e-005 3.8182 0.012049 1.1208e-006 0.001154 0.038921 0.00064922 0.039566 0.03493 0 0.045709 0.0389 0 0.84576 0.22719 0.058862 0.0083445 4.1052 0.052618 6.2757e-005 0.83744 0.0051032 0.0058412 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.9655 0.92326 0.0013951 0.99879 0.62428 0.0018797 0.43102 1.9468 1.9464 15.9972 145.0017 0.00015357 -85.6679 0.985
0.086 0.98801 5.5251e-005 3.8182 0.012049 1.1339e-006 0.001154 0.039079 0.00064927 0.039724 0.035072 0 0.045694 0.0389 0 0.84577 0.2272 0.058864 0.0083448 4.1052 0.052619 6.2758e-005 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96556 0.92329 0.0013951 0.99878 0.62441 0.0018797 0.43103 1.9471 1.9467 15.9972 145.0018 0.00015352 -85.6679 0.986
0.087 0.98801 5.5251e-005 3.8182 0.012049 1.1471e-006 0.001154 0.039236 0.00064933 0.039881 0.035215 0 0.045679 0.0389 0 0.84578 0.2272 0.058866 0.008345 4.1052 0.052619 6.2758e-005 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96561 0.92332 0.0013951 0.99877 0.62454 0.0018797 0.43104 1.9474 1.9469 15.9971 145.0018 0.00015348 -85.668 0.987
0.088 0.98801 5.5251e-005 3.8182 0.012049 1.1603e-006 0.001154 0.039394 0.00064938 0.040039 0.035357 0 0.045664 0.0389 0 0.84579 0.22721 0.058867 0.0083452 4.1052 0.05262 6.2759e-005 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96567 0.92335 0.0013951 0.99876 0.62467 0.0018797 0.43105 1.9477 1.9472 15.9971 145.0018 0.00015343 -85.668 0.988
0.089 0.98801 5.5251e-005 3.8182 0.012049 1.1735e-006 0.001154 0.039551 0.00064944 0.040196 0.0355 0 0.045649 0.0389 0 0.8458 0.22721 0.058869 0.0083454 4.1052 0.052621 6.276e-005 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96572 0.92338 0.0013951 0.99875 0.6248 0.0018797 0.43106 1.948 1.9475 15.9971 145.0018 0.00015339 -85.668 0.989
0.09 0.98801 5.5251e-005 3.8182 0.012049 1.1867e-006 0.001154 0.039708 0.00064949 0.040353 0.035642 0 0.045634 0.0389 0 0.84581 0.22722 0.058871 0.0083456 4.1052 0.052621 6.2761e-005 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9807e-006 1.1923e-005 0.13044 0.96578 0.92342 0.0013951 0.99874 0.62493 0.0018796 0.43108 1.9483 1.9478 15.997 145.0018 0.00015334 -85.668 0.99
0.091 0.98801 5.5251e-005 3.8182 0.012049 1.1999e-006 0.001154 0.039865 0.00064954 0.04051 0.035784 0 0.045619 0.0389 0 0.84582 0.22722 0.058873 0.0083459 4.1052 0.052622 6.2762e-005 0.83744 0.0051033 0.0058413 0.0013826 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96583 0.92345 0.0013951 0.99873 0.62507 0.0018796 0.43109 1.9485 1.9481 15.997 145.0019 0.0001533 -85.668 0.991
0.092 0.98801 5.525e-005 3.8182 0.012049 1.213e-006 0.001154 0.040022 0.0006496 0.040667 0.035926 0 0.045604 0.0389 0 0.84583 0.22723 0.058874 0.0083461 4.1052 0.052623 6.2762e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96589 0.92348 0.0013951 0.99872 0.6252 0.0018796 0.4311 1.9488 1.9484 15.997 145.0019 0.00015325 -85.6681 0.992
0.093 0.98801 5.525e-005 3.8182 0.012049 1.2262e-006 0.001154 0.040179 0.00064965 0.040824 0.036068 0 0.045589 0.0389 0 0.84585 0.22723 0.058876 0.0083463 4.1052 0.052623 6.2763e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96595 0.92351 0.0013951 0.99871 0.62533 0.0018796 0.43111 1.9491 1.9487 15.9969 145.0019 0.00015321 -85.6681 0.993
0.094 0.98801 5.525e-005 3.8182 0.012049 1.2394e-006 0.001154 0.040335 0.0006497 0.04098 0.03621 0 0.045574 0.0389 0 0.84586 0.22724 0.058878 0.0083465 4.1052 0.052624 6.2764e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.966 0.92354 0.0013951 0.9987 0.62546 0.0018796 0.43112 1.9494 1.949 15.9969 145.0019 0.00015317 -85.6681 0.994
0.095 0.98801 5.525e-005 3.8182 0.012049 1.2526e-006 0.001154 0.040492 0.00064975 0.041137 0.036351 0 0.04556 0.0389 0 0.84587 0.22724 0.05888 0.0083468 4.1052 0.052625 6.2765e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96606 0.92357 0.0013951 0.99869 0.62559 0.0018796 0.43113 1.9497 1.9493 15.9969 145.002 0.00015312 -85.6681 0.995
0.096 0.98801 5.525e-005 3.8182 0.012049 1.2658e-006 0.001154 0.040648 0.0006498 0.041293 0.036493 0 0.045545 0.0389 0 0.84588 0.22725 0.058882 0.008347 4.1052 0.052625 6.2766e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96611 0.9236 0.0013951 0.99868 0.62572 0.0018796 0.43115 1.95 1.9496 15.9968 145.002 0.00015308 -85.6681 0.996
0.097 0.98801 5.525e-005 3.8182 0.012049 1.279e-006 0.001154 0.040805 0.00064986 0.04145 0.036635 0 0.04553 0.0389 0 0.84589 0.22725 0.058884 0.0083472 4.1052 0.052626 6.2767e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96616 0.92363 0.0013951 0.99867 0.62585 0.0018796 0.43116 1.9503 1.9499 15.9968 145.002 0.00015303 -85.6682 0.997
0.098 0.98801 5.525e-005 3.8182 0.012049 1.2921e-006 0.001154 0.040961 0.00064991 0.041606 0.036776 0 0.045515 0.0389 0 0.8459 0.22726 0.058886 0.0083475 4.1052 0.052627 6.2768e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96622 0.92366 0.0013951 0.99866 0.62598 0.0018796 0.43117 1.9506 1.9502 15.9968 145.002 0.00015299 -85.6682 0.998
0.099 0.98801 5.525e-005 3.8182 0.012049 1.3053e-006 0.001154 0.041117 0.00064996 0.041762 0.036917 0 0.045501 0.0389 0 0.84592 0.22726 0.058888 0.0083477 4.1052 0.052628 6.2769e-005 0.83744 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96627 0.92369 0.0013951 0.99865 0.62611 0.0018796 0.43118 1.9509 1.9504 15.9967 145.002 0.00015295 -85.6682 0.999
0.1 0.98801 5.525e-005 3.8182 0.012049 1.3185e-006 0.001154 0.041273 0.00065001 0.041918 0.037058 0 0.045486 0.0389 0 0.84593 0.22727 0.058889 0.008348 4.1052 0.052628 6.277e-005 0.83743 0.0051033 0.0058413 0.0013825 0.98699 0.99173 2.9806e-006 1.1922e-005 0.13044 0.96633 0.92372 0.0013951 0.99864 0.62624 0.0018796 0.43119 1.9512 1.9507 15.9967 145.0021 0.0001529 -85.6677 1
0.101 0.98801 5.525e-005 3.8182 0.012049 1.3317e-006 0.001154 0.041428 0.00065005 0.042074 0.037199 0 0.045471 0.0389 0 0.84594 0.22728 0.058891 0.0083482 4.1052 0.052629 6.2771e-005 0.83743 0.0051034 0.0058414 0.0064682 0.98325 0.991 1.4506e-005 5.329e-005 0.13044 0.96633 0.92375 0.0027721 0.99862 0.62635 0.0023946 0.43115 1.9514 1.951 15.9967 145.002 0.00015287 -76.1658 1.001
0.102 0.98801 5.525e-005 3.8182 0.012049 1.3449e-006 0.001154 0.041584 0.0006501 0.042229 0.03734 0 0.045457 0.0389 0 0.84595 0.22728 0.058893 0.0083485 4.1052 0.05263 6.2772e-005 0.83743 0.0051034 0.0058414 0.026201 0.97173 0.98768 6.5927e-005 0.00022933 0.13044 0.96611 0.92378 0.0052988 0.99856 0.62645 0.0033354 0.43103 1.9517 1.9513 15.9966 145.002 0.00015286 -67.152 1.002
0.103 0.98801 5.525e-005 3.8182 0.012049 1.358e-006 0.001154 0.041739 0.00065015 0.042385 0.037481 0 0.045442 0.0389 0 0.84597 0.22729 0.058895 0.0083487 4.1052 0.052631 6.2773e-005 0.83743 0.0051034 0.0058414 0.094799 0.94725 0.97734 0.00028414 0.00091235 0.13044 0.96535 0.92381 0.0092447 0.99829 0.62653 0.0044241 0.43087 1.952 1.9516 15.9965 145.002 0.00015287 -58.0214 1.003
0.104 0.98801 5.525e-005 3.8182 0.012049 1.3712e-006 0.001154 0.041895 0.0006502 0.04254 0.037622 0 0.045427 0.0389 0 0.84598 0.22729 0.058897 0.008349 4.1053 0.052631 6.2774e-005 0.83743 0.0051034 0.0058414 0.48704 0.85667 0.93881 0.0021722 0.0054608 0.13044 0.96332 0.92383 0.015745 0.99417 0.62654 0.0056227 0.43068 1.9523 1.9519 15.9973 145.002 0.00015291 -37.2735 0.15765
0.105 0.98801 5.525e-005 3.8182 0.012049 1.3844e-006 0.001154 0.04205 0.00065025 0.042696 0.037763 0 0.045413 0.0389 0 0.84599 0.2273 0.058899 0.0083492 4.1053 0.052632 6.2775e-005 0.83743 0.0051034 0.0058414 0.99958 0.0021914 0.71228 0.93538 0.99563 0.13044 0.92972 0.9209 0.3314 0.96668 0.61279 0.043903 0.43047 1.9123 0.97381 16.0012 145.0017 0.00023146 23.7554 0.0019576
0.106 0.98801 5.525e-005 3.8182 0.012049 1.3976e-006 0.001154 0.042205 0.00065029 0.042851 0.037903 0 0.045398 0.0389 0 0.846 0.2273 0.058901 0.0083495 4.1053 0.052633 6.2776e-005 0.83743 0.0051034 0.0058414 0.99922 1.492e-006 0.5285 0.99578 0.99914 0.13044 0.88962 0.90303 0.59387 0.93946 0.59574 0.093221 0.43027 1.7303 0.59026 16.0008 145.0004 0.00034031 17.2282 0.0029576
0.107 0.98801 5.525e-005 3.8182 0.012049 1.4108e-006 0.001154 0.04236 0.00065034 0.043006 0.038044 0 0.045384 0.0389 0 0.84602 0.22731 0.058904 0.0083498 4.1053 0.052634 6.2777e-005 0.83743 0.0051034 0.0058414 0.99847 1.4033e-008 0.39272 0.99193 0.99759 0.13044 0.85272 0.8799 0.7018 0.913 0.57966 0.12824 0.43006 1.5553 0.56157 16.0004 144.9988 0.00040783 11.0054 0.0039576
0.108 0.98801 5.5249e-005 3.8182 0.012049 1.424e-006 0.001154 0.042515 0.00065039 0.043161 0.038184 0 0.045369 0.0389 0 0.84603 0.22731 0.058906 0.00835 4.1053 0.052635 6.2778e-005 0.83743 0.0051034 0.0058414 0.99759 -2.3924e-009 0.2924 0.98398 0.99505 0.13044 0.81974 0.8545 0.74587 0.8873 0.56492 0.15446 0.42986 1.4089 0.5972 16.0001 144.9971 0.00045761 6.8817 0.0049576
0.109 0.98801 5.5249e-005 3.8182 0.012049 1.4371e-006 0.001154 0.04267 0.00065043 0.043316 0.038324 0 0.045355 0.0389 0 0.84604 0.22732 0.058908 0.0083503 4.1053 0.052636 6.2779e-005 0.83743 0.0051034 0.0058414 0.99672 -5.2015e-010 0.21813 0.97374 0.99183 0.13044 0.79026 0.82824 0.7615 0.86232 0.55155 0.17559 0.42965 1.2923 0.65323 15.9998 144.9956 0.00049538 4.1034 0.0059576
0.11 0.98801 5.5249e-005 3.8182 0.012049 1.4503e-006 0.001154 0.042824 0.00065048 0.04347 0.038464 0 0.04534 0.0389 0 0.84606 0.22733 0.05891 0.0083506 4.1053 0.052636 6.278e-005 0.83743 0.0051034 0.0058414 0.99585 -1.978e-010 0.16302 0.96183 0.98809 0.13044 0.76368 0.80209 0.76272 0.83806 0.53943 0.1934 0.42945 1.2027 0.71416 15.9995 144.9941 0.00052392 1.9696 0.0069576
0.111 0.98801 5.5249e-005 3.8182 0.012049 1.4635e-006 0.001154 0.042979 0.00065052 0.043625 0.038604 0 0.045326 0.0389 0 0.84607 0.22733 0.058912 0.0083508 4.1053 0.052637 6.2781e-005 0.83743 0.0051034 0.0058414 0.9949 -6.7808e-011 0.12206 0.94818 0.98371 0.13044 0.73958 0.77672 0.75565 0.81449 0.52848 0.20868 0.42924 1.1359 0.77218 15.9992 144.9926 0.00054531 0.11945 0.0079576
0.112 0.98801 5.5249e-005 3.8182 0.012049 1.4767e-006 0.001154 0.043133 0.00065057 0.043779 0.038744 0 0.045311 0.0389 0 0.84608 0.22734 0.058914 0.0083511 4.1053 0.052638 6.2782e-005 0.83742 0.0051034 0.0058414 0.99381 2.8719e-011 0.091579 0.93231 0.97842 0.13044 0.71774 0.7526 0.74325 0.79159 0.51863 0.22188 0.42904 1.0876 0.82309 15.999 144.9913 0.00056128 -1.631 0.0089576
0.113 0.98801 5.5249e-005 3.8182 0.012049 1.4899e-006 0.001154 0.043288 0.00065061 0.043934 0.038884 0 0.045297 0.0389 0 0.8461 0.22734 0.058916 0.0083514 4.1053 0.052639 6.2783e-005 0.83742 0.0051035 0.0058414 0.99248 1.6752e-011 0.068865 0.91343 0.97182 0.13044 0.69802 0.73009 0.72694 0.76935 0.50986 0.23322 0.42884 1.0538 0.86516 15.9987 144.9901 0.00057325 -3.3954 0.0099576
0.114 0.98801 5.5249e-005 3.8182 0.012048 1.5031e-006 0.001154 0.043442 0.00065065 0.044088 0.039024 0 0.045282 0.0389 0 0.84611 0.22735 0.058918 0.0083517 4.1053 0.05264 6.2785e-005 0.83742 0.0051035 0.0058415 0.99074 -1.3859e-011 0.05193 0.89039 0.96329 0.13044 0.68034 0.70949 0.70739 0.74775 0.50219 0.24284 0.42863 1.0309 0.89838 15.9984 144.9889 0.00058228 -5.2674 0.010958
0.115 0.98801 5.5249e-005 3.8182 0.012048 1.5162e-006 0.001154 0.043596 0.0006507 0.044242 0.039164 0 0.045268 0.0389 0 0.84613 0.22736 0.058921 0.0083519 4.1053 0.052641 6.2786e-005 0.83742 0.0051035 0.0058415 0.98834 1.4487e-013 0.0393 0.86152 0.95186 0.13044 0.6647 0.69105 0.68475 0.72679 0.49564 0.25079 0.42843 1.016 0.92373 15.9982 144.9879 0.00058914 -7.3481 0.011958
0.116 0.98801 5.5249e-005 3.8182 0.012048 1.5294e-006 0.001154 0.04375 0.00065074 0.044396 0.039303 0 0.045253 0.0389 0 0.84614 0.22736 0.058923 0.0083522 4.1053 0.052642 6.2787e-005 0.83742 0.0051035 0.0058415 0.98474 6.8596e-012 0.029887 0.82427 0.93593 0.13044 0.65114 0.67503 0.65888 0.70645 0.49025 0.2571 0.42822 1.0066 0.94266 15.998 144.9869 0.00059432 -9.7662 0.012958
0.117 0.98801 5.5249e-005 3.8182 0.012048 1.5426e-006 0.001154 0.043903 0.00065078 0.04455 0.039442 0 0.045239 0.0389 0 0.84615 0.22737 0.058925 0.0083525 4.1053 0.052643 6.2788e-005 0.83742 0.0051035 0.0058415 0.97885 -1.9991e-011 0.022892 0.77481 0.91282 0.13044 0.63974 0.6617 0.6294 0.68675 0.48602 0.26176 0.42802 1.0012 0.95665 15.9977 144.986 0.00059809 -12.6971 0.013958
0.118 0.98801 5.5249e-005 3.8182 0.012048 1.5558e-006 0.001154 0.044057 0.00065082 0.044703 0.039582 0 0.045225 0.0389 0 0.84617 0.22738 0.058927 0.0083528 4.1053 0.052644 6.2789e-005 0.83742 0.0051035 0.0058415 0.96817 1.323e-011 0.017729 0.70733 0.8779 0.13044 0.63057 0.65132 0.59593 0.66773 0.48296 0.26475 0.42782 0.99846 0.96704 15.9975 144.9853 0.00060057 -16.3726 0.014958
0.119 0.98801 5.5249e-005 3.8182 0.012048 1.569e-006 0.001154 0.044211 0.00065087 0.044857 0.039721 0 0.04521 0.0389 0 0.84618 0.22738 0.05893 0.0083531 4.1053 0.052645 6.2791e-005 0.83742 0.0051035 0.0058415 0.94654 -3.4669e-011 0.013982 0.61373 0.82336 0.13044 0.62363 0.64402 0.55836 0.6495 0.48095 0.26612 0.42761 0.99751 0.97513 15.9973 144.9846 0.00060172 -21.0381 0.015958
0.12 0.98801 5.5249e-005 3.8182 0.012048 1.5821e-006 0.001154 0.044364 0.00065091 0.04501 0.03986 0 0.045196 0.0389 0 0.8462 0.22739 0.058932 0.0083534 4.1054 0.052646 6.2792e-005 0.83742 0.0051035 0.0058415 0.89964 1.617e-011 0.011359 0.48589 0.73742 0.13044 0.61867 0.63962 0.5168 0.63245 0.47978 0.26606 0.42741 0.99782 0.98181 15.9972 144.9841 0.0006015 -26.7582 0.016958
0.121 0.98801 5.5249e-005 3.8182 0.012048 1.5953e-006 0.001154 0.044517 0.00065095 0.045164 0.039999 0 0.045182 0.0389 0 0.84621 0.22739 0.058934 0.0083537 4.1054 0.052647 6.2793e-005 0.83742 0.0051035 0.0058415 0.80372 2.4521e-011 0.009625 0.32704 0.60832 0.13044 0.6152 0.63734 0.4704 0.61756 0.47919 0.26482 0.42721 0.99898 0.98689 15.997 144.9836 0.00060037 -33.0496 0.017958
0.122 0.98801 5.5249e-005 3.8182 0.012048 1.6085e-006 0.001154 0.04467 0.00065099 0.045317 0.040138 0 0.045168 0.0389 0 0.84623 0.2274 0.058937 0.0083539 4.1054 0.052648 6.2795e-005 0.83741 0.0051035 0.0058415 0.65255 9.4876e-012 0.0085352 0.1705 0.44063 0.13044 0.61269 0.63609 0.41604 0.60676 0.47893 0.26242 0.42701 1.0006 0.99089 15.9969 144.9833 0.00059879 -38.9285 0.018958
0.123 0.98801 5.5249e-005 3.8182 0.012048 1.6217e-006 0.001154 0.044823 0.00065103 0.04547 0.040277 0 0.045153 0.0389 0 0.84624 0.22741 0.058939 0.0083542 4.1054 0.052649 6.2796e-005 0.83741 0.0051036 0.0058415 0.48645 0.00037352 0.0079736 0.063908 0.26874 0.13044 0.61082 0.63534 0.35118 0.60133 0.47885 0.25863 0.42681 1.0026 0.99422 15.9968 144.983 0.00059708 -43.8067 0.019958
0.124 0.98801 5.5248e-005 3.8182 0.012048 1.6349e-006 0.001154 0.044976 0.00065107 0.045623 0.040415 0 0.045139 0.0389 0 0.84626 0.22741 0.058941 0.0083545 4.1054 0.05265 6.2797e-005 0.83741 0.0051036 0.0058416 0.34992 0.0011792 0.0079188 0.017184 0.13496 0.13044 0.60941 0.63525 0.2783 0.59993 0.47887 0.25311 0.42662 1.0047 0.99717 15.9968 144.9828 0.00059531 -47.6904 0.020958
0.125 0.98801 5.5248e-005 3.8182 0.012048 1.6481e-006 0.001154 0.045129 0.00065111 0.045776 0.040554 0 0.045125 0.0389 0 0.84627 0.22742 0.058944 0.0083548 4.1054 0.052651 6.2799e-005 0.83741 0.0051036 0.0058416 0.25515 0.0025148 0.0083273 0.0040177 0.056145 0.13044 0.60839 0.63595 0.20516 0.60036 0.47894 0.24569 0.42643 1.0069 0.99988 15.9967 144.9827 0.00059352 -50.7353 0.021958
0.126 0.98801 5.5248e-005 3.8182 0.012048 1.6612e-006 0.001154 0.045282 0.00065115 0.045928 0.040693 0 0.045111 0.0389 0 0.84629 0.22743 0.058946 0.0083551 4.1054 0.052652 6.28e-005 0.83741 0.0051036 0.0058416 0.19339 0.0044938 0.009167 0.0013555 0.0204 0.13044 0.60768 0.63721 0.14096 0.6014 0.47903 0.23641 0.42624 1.0092 1.0025 15.9967 144.9826 0.0005917 -53.1158 0.022958
0.127 0.98801 5.5248e-005 3.8182 0.012048 1.6744e-006 0.001154 0.045434 0.00065119 0.046081 0.040831 0 0.045097 0.0389 0 0.8463 0.22743 0.058949 0.0083555 4.1054 0.052653 6.2801e-005 0.83741 0.0051036 0.0058416 0.15275 0.007182 0.010405 0.00078089 0.0074152 0.13044 0.60722 0.63872 0.091514 0.60261 0.47914 0.22549 0.42605 1.0116 1.005 15.9967 144.9825 0.00058987 -55.0095 0.023958
0.128 0.98801 5.5248e-005 3.8182 0.012048 1.6876e-006 0.001154 0.045587 0.00065123 0.046233 0.040969 0 0.045083 0.0389 0 0.84632 0.22744 0.058951 0.0083558 4.1054 0.052654 6.2803e-005 0.83741 0.0051036 0.0058416 0.12462 0.010617 0.012016 0.00056051 0.0033289 0.13044 0.60696 0.64031 0.057634 0.60383 0.47925 0.21322 0.42587 1.0139 1.0074 15.9966 144.9824 0.00058802 -56.5747 0.024958
0.129 0.98801 5.5248e-005 3.8182 0.012048 1.7008e-006 0.001154 0.045739 0.00065126 0.046386 0.041107 0 0.045068 0.0389 0 0.84633 0.22745 0.058953 0.0083561 4.1054 0.052655 6.2804e-005 0.83741 0.0051036 0.0058416 0.10388 0.014839 0.013982 0.00043125 0.002023 0.13044 0.60685 0.64192 0.036581 0.60503 0.47937 0.19993 0.42569 1.0162 1.0098 15.9966 144.9824 0.00058617 -57.9333 0.025958
0.13 0.98801 5.5248e-005 3.8182 0.012048 1.714e-006 0.001154 0.045891 0.0006513 0.046538 0.041245 0 0.045054 0.0389 0 0.84635 0.22745 0.058956 0.0083564 4.1054 0.052657 6.2806e-005 0.83741 0.0051036 0.0058416 0.087699 0.019904 0.016304 0.00034242 0.0014845 0.13044 0.60688 0.64352 0.024451 0.60619 0.47949 0.18585 0.42552 1.0186 1.0122 15.9966 144.9824 0.00058431 -59.1682 0.026958
0.131 0.98801 5.5248e-005 3.8182 0.012048 1.7271e-006 0.001154 0.046043 0.00065134 0.04669 0.041383 0 0.04504 0.0389 0 0.84636 0.22746 0.058958 0.0083567 4.1054 0.052658 6.2807e-005 0.83741 0.0051036 0.0058416 0.074548 0.025901 0.018993 0.00027662 0.0011704 0.13044 0.60703 0.64511 0.017775 0.6073 0.47962 0.17123 0.42534 1.0209 1.0146 15.9966 144.9824 0.00058244 -60.3296 0.027958
0.132 0.98801 5.5248e-005 3.8182 0.012048 1.7403e-006 0.001154 0.046195 0.00065138 0.046842 0.041521 0 0.045026 0.0389 0 0.84638 0.22747 0.058961 0.008357 4.1054 0.052659 6.2808e-005 0.8374 0.0051037 0.0058416 0.063605 0.032943 0.022071 0.00022579 0.00094615 0.13044 0.60729 0.64669 0.014099 0.60838 0.47974 0.15628 0.42517 1.0233 1.017 15.9966 144.9823 0.00058057 -61.4451 0.028958
0.133 0.98801 5.5248e-005 3.8182 0.012048 1.7535e-006 0.001154 0.046347 0.00065141 0.046994 0.041659 0 0.045012 0.0389 0 0.8464 0.22748 0.058963 0.0083573 4.1055 0.05266 6.281e-005 0.8374 0.0051037 0.0058417 0.054386 0.041164 0.025565 0.00018555 0.00077282 0.13044 0.60764 0.64826 0.011937 0.60942 0.47987 0.14119 0.42501 1.0256 1.0194 15.9966 144.9823 0.0005787 -62.5285 0.029958
0.134 0.98801 5.5248e-005 3.8182 0.012048 1.7667e-006 0.001154 0.046499 0.00065145 0.047145 0.041797 0 0.044998 0.0389 0 0.84641 0.22748 0.058966 0.0083577 4.1055 0.052661 6.2811e-005 0.8374 0.0051037 0.0058417 0.046578 0.050717 0.029511 0.00015326 0.00063562 0.13044 0.60809 0.64982 0.010502 0.61043 0.47999 0.12618 0.42485 1.028 1.0217 15.9967 144.9823 0.00057683 -63.5863 0.030958
0.135 0.98801 5.5248e-005 3.8182 0.012048 1.7799e-006 0.001154 0.04665 0.00065149 0.047297 0.041934 0 0.044984 0.0389 0 0.84643 0.22749 0.058969 0.008358 4.1055 0.052662 6.2813e-005 0.8374 0.0051037 0.0058417 0.039951 0.06177 0.033947 0.00012723 0.00052544 0.13044 0.60861 0.65136 0.0094189 0.61141 0.48012 0.11146 0.42469 1.0303 1.0241 15.9967 144.9823 0.00057495 -64.6213 0.031958
0.136 0.98801 5.5248e-005 3.8182 0.012048 1.7931e-006 0.001154 0.046802 0.00065152 0.047449 0.042072 0 0.04497 0.0389 0 0.84644 0.2275 0.058971 0.0083583 4.1055 0.052664 6.2814e-005 0.8374 0.0051037 0.0058417 0.034321 0.074496 0.038914 0.00010603 0.00043652 0.13044 0.6092 0.65289 0.0085263 0.61236 0.48025 0.097257 0.42454 1.0327 1.0265 15.9967 144.9822 0.00057307 -65.6345 0.032958
0.137 0.98801 5.5248e-005 3.8182 0.012048 1.8062e-006 0.001154 0.046953 0.00065156 0.0476 0.042209 0 0.044956 0.0389 0 0.84646 0.2275 0.058974 0.0083586 4.1055 0.052665 6.2816e-005 0.8374 0.0051037 0.0058417 0.029537 0.089073 0.044461 8.8745e-005 0.00036424 0.13044 0.60986 0.65441 0.0077572 0.6133 0.48038 0.083764 0.42439 1.035 1.0288 15.9967 144.9822 0.00057119 -66.6262 0.033958
0.138 0.98801 5.5248e-005 3.8182 0.012048 1.8194e-006 0.001154 0.047104 0.00065159 0.047751 0.042346 0 0.044942 0.0389 0 0.84648 0.22751 0.058976 0.008359 4.1055 0.052666 6.2817e-005 0.8374 0.0051037 0.0058417 0.025472 0.10568 0.050637 7.4566e-005 0.00030533 0.13044 0.61057 0.65592 0.007082 0.61423 0.48051 0.071172 0.42424 1.0374 1.0312 15.9968 144.9822 0.00056931 -67.596 0.034958
0.139 0.98801 5.5248e-005 3.8182 0.012048 1.8326e-006 0.001154 0.047255 0.00065163 0.047902 0.042483 0 0.044928 0.0389 0 0.84649 0.22752 0.058979 0.0083593 4.1055 0.052667 6.2819e-005 0.8374 0.0051037 0.0058417 0.022017 0.12448 0.057502 6.2947e-005 0.00025708 0.13045 0.61133 0.65741 0.0064846 0.61516 0.48064 0.059639 0.4241 1.0397 1.0336 15.9968 144.9821 0.00056743 -68.5434 0.035958
0.14 0.98801 5.5247e-005 3.8182 0.012048 1.8458e-006 0.001154 0.047406 0.00065166 0.048053 0.04262 0 0.044914 0.0389 0 0.84651 0.22753 0.058982 0.0083596 4.1055 0.052668 6.2821e-005 0.83739 0.0051038 0.0058417 0.01908 0.14562 0.06512 5.3321e-005 0.00021746 0.13045 0.61214 0.65889 0.005954 0.61608 0.48077 0.049284 0.42397 1.042 1.0359 15.9968 144.9821 0.00056554 -69.4673 0.036958
0.141 0.98801 5.5247e-005 3.8182 0.012048 1.859e-006 0.001154 0.047557 0.0006517 0.048204 0.042757 0 0.0449 0.0389 0 0.84653 0.22753 0.058984 0.00836 4.1055 0.05267 6.2822e-005 0.83739 0.0051038 0.0058418 0.016583 0.16924 0.073562 4.5404e-005 0.00018482 0.13045 0.61299 0.66036 0.0054819 0.617 0.4809 0.040179 0.42384 1.0444 1.0383 15.9969 144.9821 0.00056366 -70.3665 0.037958
0.142 0.98801 5.5247e-005 3.8182 0.012048 1.8721e-006 0.001154 0.047708 0.00065173 0.048355 0.042894 0 0.044887 0.0389 0 0.84654 0.22754 0.058987 0.0083603 4.1055 0.052671 6.2824e-005 0.83739 0.0051038 0.0058418 0.01446 0.1954 0.082904 3.8821e-005 0.00015785 0.13045 0.61387 0.66182 0.0050613 0.61794 0.48103 0.032349 0.42372 1.0467 1.0406 15.9969 144.9821 0.00056178 -71.2398 0.038958
0.143 0.98801 5.5247e-005 3.8182 0.012048 1.8853e-006 0.001154 0.047858 0.00065176 0.048505 0.043031 0 0.044873 0.0389 0 0.84656 0.22755 0.05899 0.0083606 4.1055 0.052672 6.2825e-005 0.83739 0.0051038 0.0058418 0.012655 0.22414 0.09323 3.3412e-005 0.00013552 0.13045 0.61478 0.66327 0.0046861 0.61888 0.48117 0.025768 0.4236 1.049 1.043 15.997 144.982 0.00055989 -72.0854 0.039958
0.144 0.98801 5.5247e-005 3.8182 0.012048 1.8985e-006 0.001154 0.048009 0.0006518 0.048656 0.043168 0 0.044859 0.0389 0 0.84658 0.22756 0.058992 0.008361 4.1056 0.052674 6.2827e-005 0.83739 0.0051038 0.0058418 0.011119 0.25542 0.10462 2.8879e-005 0.00011698 0.13045 0.61571 0.6647 0.0043514 0.61985 0.4813 0.020366 0.42349 1.0513 1.0453 15.997 144.982 0.00055801 -72.9017 0.040958
0.145 0.98801 5.5247e-005 3.8182 0.012048 1.9117e-006 0.001154 0.048159 0.00065183 0.048806 0.043304 0 0.044845 0.0389 0 0.8466 0.22756 0.058995 0.0083613 4.1056 0.052675 6.2829e-005 0.83739 0.0051038 0.0058418 0.0098125 0.28913 0.11717 2.5103e-005 0.00010156 0.13045 0.61667 0.66612 0.0040529 0.62083 0.48144 0.016036 0.42338 1.0536 1.0476 15.9971 144.982 0.00055613 -73.6871 0.041958
0.146 0.98801 5.5247e-005 3.8182 0.012048 1.9249e-006 0.001154 0.048309 0.00065186 0.048957 0.043441 0 0.044831 0.0389 0 0.84661 0.22757 0.058998 0.0083617 4.1056 0.052676 6.283e-005 0.83739 0.0051038 0.0058418 0.0087004 0.32509 0.13094 2.1953e-005 8.8694e-005 0.13045 0.61765 0.66753 0.0037865 0.62184 0.48158 0.012648 0.42328 1.056 1.05 15.9972 144.9819 0.00055426 -74.4399 0.042958
0.147 0.98801 5.5247e-005 3.8182 0.012048 1.938e-006 0.001154 0.048459 0.0006519 0.049107 0.043577 0 0.044817 0.0389 0 0.84663 0.22758 0.059001 0.008362 4.1056 0.052678 6.2832e-005 0.83739 0.0051038 0.0058418 0.007753 0.36301 0.14599 1.931e-005 7.7944e-005 0.13045 0.61864 0.66893 0.0035491 0.62288 0.48171 0.010055 0.42319 1.0583 1.0523 15.9972 144.9819 0.00055238 -75.1588 0.043958
0.148 0.98801 5.5247e-005 3.8182 0.012048 1.9512e-006 0.001154 0.048609 0.00065193 0.049257 0.043713 0 0.044804 0.0389 0 0.84665 0.22759 0.059003 0.0083624 4.1056 0.052679 6.2834e-005 0.83738 0.0051039 0.0058418 0.0069452 0.40253 0.16235 1.7095e-005 6.8938e-005 0.13045 0.61965 0.67032 0.0033376 0.62395 0.48185 0.0081132 0.4231 1.0606 1.0546 15.9973 144.9819 0.00055051 -75.8424 0.044958
0.149 0.98801 5.5247e-005 3.8182 0.012048 1.9644e-006 0.001154 0.048759 0.00065196 0.049407 0.043849 0 0.04479 0.0389 0 0.84667 0.22759 0.059006 0.0083627 4.1056 0.05268 6.2836e-005 0.83738 0.0051039 0.0058419 0.0062562 0.44322 0.18003 1.5234e-005 6.1375e-005 0.13045 0.62067 0.67169 0.0031492 0.62505 0.482 0.0066837 0.42302 1.0629 1.057 15.9974 144.9819 0.00054864 -76.4897 0.045958
0.15 0.98801 5.5247e-005 3.8182 0.012048 1.9776e-006 0.001154 0.048909 0.00065199 0.049557 0.043985 0 0.044776 0.0389 0 0.84668 0.2276 0.059009 0.0083631 4.1056 0.052682 6.2837e-005 0.83738 0.0051039 0.0058419 0.0056676 0.48458 0.199 1.366e-005 5.5007e-005 0.13045 0.6217 0.67306 0.0029815 0.62619 0.48214 0.0056454 0.42294 1.0652 1.0593 15.9974 144.9818 0.00054678 -77.1003 0.046958
0.151 0.98801 5.5247e-005 3.8182 0.012048 1.9908e-006 0.001154 0.049059 0.00065202 0.049706 0.044121 0 0.044763 0.0389 0 0.8467 0.22761 0.059012 0.0083635 4.1056 0.052683 6.2839e-005 0.83738 0.0051039 0.0058419 0.0051637 0.52608 0.21918 1.2331e-005 4.9632e-005 0.13045 0.62273 0.67441 0.0028323 0.62736 0.48228 0.0048964 0.42287 1.0675 1.0616 15.9975 144.9818 0.00054491 -77.6737 0.047958
0.152 0.98801 5.5247e-005 3.8182 0.012048 2.004e-006 0.001154 0.049208 0.00065205 0.049856 0.044257 0 0.044749 0.0389 0 0.84672 0.22762 0.059015 0.0083638 4.1056 0.052684 6.2841e-005 0.83738 0.0051039 0.0058419 0.0047324 0.56718 0.24048 1.1212e-005 4.5083e-005 0.13045 0.62378 0.67576 0.0026997 0.62858 0.48243 0.0043556 0.4228 1.0698 1.0639 15.9976 144.9818 0.00054306 -78.2101 0.048958
0.153 0.98801 5.5247e-005 3.8182 0.012048 2.0171e-006 0.001154 0.049358 0.00065209 0.050005 0.044393 0 0.044735 0.0389 0 0.84674 0.22763 0.059018 0.0083642 4.1057 0.052686 6.2843e-005 0.83738 0.0051039 0.0058419 0.0043622 0.60735 0.26276 1.0257e-005 4.1221e-005 0.13045 0.62482 0.67709 0.0025819 0.62983 0.48258 0.0039612 0.42274 1.0721 1.0662 15.9977 144.9818 0.00054121 -78.7099 0.049958
0.154 0.98801 5.5247e-005 3.8182 0.012048 2.0303e-006 0.001154 0.049507 0.00065212 0.050154 0.044528 0 0.044722 0.0389 0 0.84676 0.22763 0.05902 0.0083645 4.1057 0.052687 6.2845e-005 0.83738 0.005104 0.0058419 0.0040438 0.6461 0.28585 9.4426e-006 3.7934e-005 0.13045 0.62588 0.67841 0.0024772 0.63112 0.48273 0.0036682 0.42268 1.0744 1.0685 15.9977 144.9818 0.00053936 -79.1739 0.050958
0.155 0.98801 5.5247e-005 3.8182 0.012048 2.0435e-006 0.001154 0.049656 0.00065215 0.050304 0.044664 0 0.044708 0.0389 0 0.84677 0.22764 0.059023 0.0083649 4.1057 0.052689 6.2846e-005 0.83737 0.005104 0.0058419 0.0037696 0.683 0.3096 8.7492e-006 3.5128e-005 0.13045 0.62693 0.67973 0.0023842 0.63245 0.48288 0.0034449 0.42263 1.0767 1.0708 15.9978 144.9817 0.00053752 -79.6032 0.051958
0.156 0.98801 5.5247e-005 3.8182 0.012048 2.0567e-006 0.001154 0.049805 0.00065218 0.050453 0.044799 0 0.044694 0.0389 0 0.84679 0.22765 0.059026 0.0083653 4.1057 0.05269 6.2848e-005 0.83737 0.005104 0.005842 0.0035329 0.7177 0.33383 8.1541e-006 3.2725e-005 0.13045 0.62799 0.68103 0.0023016 0.63382 0.48303 0.0032697 0.42258 1.0789 1.0732 15.9979 144.9817 0.00053569 -79.9991 0.052958
0.157 0.98801 5.5246e-005 3.8182 0.012048 2.0699e-006 0.001154 0.049954 0.00065221 0.050602 0.044935 0 0.044681 0.0389 0 0.84681 0.22766 0.059029 0.0083656 4.1057 0.052692 6.285e-005 0.83737 0.005104 0.005842 0.0033281 0.74994 0.35836 7.6414e-006 3.0661e-005 0.13045 0.62905 0.68232 0.0022282 0.63523 0.48318 0.0031283 0.42254 1.0812 1.0755 15.998 144.9817 0.00053386 -80.3632 0.053958
0.158 0.98801 5.5246e-005 3.8182 0.012048 2.083e-006 0.001154 0.050103 0.00065224 0.05075 0.04507 0 0.044667 0.0389 0 0.84683 0.22767 0.059032 0.008366 4.1057 0.052693 6.2852e-005 0.83737 0.005104 0.005842 0.0031503 0.77954 0.38302 7.2005e-006 2.8884e-005 0.13045 0.63012 0.6836 0.0021631 0.63667 0.48334 0.0030112 0.4225 1.0835 1.0777 15.9981 144.9817 0.00053204 -80.697 0.054958
0.159 0.98801 5.5246e-005 3.8182 0.012048 2.0962e-006 0.001154 0.050251 0.00065227 0.050899 0.045205 0 0.044654 0.0389 0 0.84685 0.22767 0.059035 0.0083664 4.1057 0.052695 6.2854e-005 0.83737 0.005104 0.005842 0.0029961 0.80641 0.40766 6.8221e-006 2.7349e-005 0.13045 0.63118 0.68487 0.0021051 0.63814 0.48349 0.0029122 0.42246 1.0858 1.08 15.9982 144.9817 0.00053023 -81.0024 0.055958
0.16 0.98801 5.5246e-005 3.8182 0.012048 2.1094e-006 0.001154 0.0504 0.0006523 0.051048 0.04534 0 0.04464 0.0389 0 0.84687 0.22768 0.059038 0.0083668 4.1057 0.052696 6.2856e-005 0.83737 0.005104 0.005842 0.0028619 0.83056 0.43213 6.4916e-006 2.6019e-005 0.13045 0.63224 0.68614 0.0020536 0.63964 0.48365 0.0028273 0.42243 1.0881 1.0823 15.9983 144.9817 0.00052842 -81.2812 0.056958
0.161 0.98801 5.5246e-005 3.8182 0.012048 2.1226e-006 0.001154 0.050548 0.00065232 0.051196 0.045475 0 0.044627 0.0389 0 0.84689 0.22769 0.059041 0.0083671 4.1057 0.052698 6.2858e-005 0.83737 0.0051041 0.005842 0.0027445 0.85205 0.45631 6.2026e-006 2.4864e-005 0.13045 0.6333 0.68739 0.0020078 0.64118 0.48381 0.0027536 0.4224 1.0903 1.0846 15.9983 144.9817 0.00052662 -81.5352 0.057958
0.162 0.98801 5.5246e-005 3.8182 0.012048 2.1358e-006 0.001154 0.050697 0.00065235 0.051345 0.04561 0 0.044613 0.0389 0 0.8469 0.2277 0.059044 0.0083675 4.1058 0.052699 6.286e-005 0.83736 0.0051041 0.0058421 0.002642 0.871 0.48009 5.9545e-006 2.3859e-005 0.13045 0.63436 0.68863 0.0019671 0.64273 0.48397 0.0026893 0.42237 1.0926 1.0869 15.9984 144.9817 0.00052483 -81.7662 0.058958
0.163 0.98801 5.5246e-005 3.8182 0.012048 2.1489e-006 0.001154 0.050845 0.00065238 0.051493 0.045745 0 0.0446 0.0389 0 0.84692 0.22771 0.059047 0.0083679 4.1058 0.052701 6.2862e-005 0.83736 0.0051041 0.0058421 0.002552 0.88756 0.50338 5.7376e-006 2.2981e-005 0.13045 0.63543 0.68987 0.0019308 0.64432 0.48413 0.0026328 0.42234 1.0948 1.0892 15.9985 144.9817 0.00052305 -81.9761 0.059958
0.164 0.98801 5.5246e-005 3.8182 0.012048 2.1621e-006 0.001154 0.050993 0.00065241 0.051641 0.045879 0 0.044586 0.0389 0 0.84694 0.22772 0.05905 0.0083683 4.1058 0.052702 6.2864e-005 0.83736 0.0051041 0.0058421 0.0024728 0.90193 0.52609 5.5451e-006 2.2212e-005 0.13045 0.63649 0.69109 0.0018985 0.64592 0.48429 0.0025831 0.42232 1.0971 1.0915 15.9986 144.9817 0.00052127 -82.1666 0.060958
0.165 0.98801 5.5246e-005 3.8182 0.012048 2.1753e-006 0.001154 0.051141 0.00065244 0.051789 0.046014 0 0.044573 0.0389 0 0.84696 0.22772 0.059053 0.0083687 4.1058 0.052704 6.2866e-005 0.83736 0.0051041 0.0058421 0.0024032 0.91431 0.54817 5.3773e-006 2.1537e-005 0.13045 0.63754 0.69231 0.0018696 0.64755 0.48445 0.0025391 0.42229 1.0994 1.0937 15.9987 144.9817 0.00051951 -82.3393 0.061958
0.166 0.98801 5.5246e-005 3.8182 0.012048 2.1885e-006 0.001154 0.051289 0.00065247 0.051937 0.046148 0 0.044559 0.0389 0 0.84698 0.22773 0.059056 0.0083691 4.1058 0.052705 6.2868e-005 0.83736 0.0051041 0.0058421 0.0023421 0.9249 0.56956 5.2318e-006 2.0944e-005 0.13045 0.6386 0.69351 0.0018439 0.64919 0.48461 0.0025001 0.42227 1.1016 1.096 15.9988 144.9816 0.00051775 -82.4958 0.062958
0.167 0.98801 5.5246e-005 3.8182 0.012048 2.2017e-006 0.001154 0.051437 0.00065249 0.052085 0.046282 0 0.044546 0.0389 0 0.847 0.22774 0.059059 0.0083695 4.1058 0.052707 6.287e-005 0.83736 0.0051042 0.0058421 0.0022877 0.93391 0.59024 5.1006e-006 2.042e-005 0.13045 0.63965 0.69471 0.0018209 0.65085 0.48477 0.0024655 0.42225 1.1038 1.0983 15.9989 144.9816 0.000516 -82.6376 0.063958
0.168 0.98801 5.5246e-005 3.8182 0.012048 2.2148e-006 0.001154 0.051584 0.00065252 0.052232 0.046417 0 0.044532 0.0389 0 0.84702 0.22775 0.059062 0.0083699 4.1058 0.052709 6.2872e-005 0.83735 0.0051042 0.0058422 0.0022394 0.94155 0.61018 4.9844e-006 1.9958e-005 0.13045 0.64071 0.6959 0.0018003 0.65252 0.48494 0.0024348 0.42224 1.1061 1.1005 15.999 144.9816 0.00051426 -82.766 0.064958
0.169 0.98801 5.5246e-005 3.8182 0.012048 2.228e-006 0.001154 0.051732 0.00065255 0.05238 0.046551 0 0.044519 0.0389 0 0.84704 0.22776 0.059066 0.0083703 4.1058 0.05271 6.2874e-005 0.83735 0.0051042 0.0058422 0.0021968 0.94798 0.62936 4.8832e-006 1.9548e-005 0.13045 0.64176 0.69708 0.0017818 0.6542 0.4851 0.0024074 0.42222 1.1083 1.1028 15.9991 144.9816 0.00051253 -82.8823 0.065958
0.17 0.98801 5.5246e-005 3.8182 0.012048 2.2412e-006 0.001154 0.051879 0.00065258 0.052527 0.046685 0 0.044506 0.0389 0 0.84706 0.22777 0.059069 0.0083707 4.1059 0.052712 6.2876e-005 0.83735 0.0051042 0.0058422 0.0021589 0.95339 0.64777 4.7928e-006 1.9184e-005 0.13045 0.6428 0.69825 0.0017653 0.65589 0.48526 0.0023829 0.42221 1.1106 1.105 15.9992 144.9816 0.00051081 -82.9877 0.066958
0.171 0.98801 5.5246e-005 3.8182 0.012048 2.2544e-006 0.001154 0.052026 0.0006526 0.052674 0.046819 0 0.044492 0.0389 0 0.84708 0.22778 0.059072 0.0083711 4.1059 0.052714 6.2878e-005 0.83735 0.0051042 0.0058422 0.0021249 0.95792 0.66542 4.712e-006 1.8859e-005 0.13045 0.64385 0.69941 0.0017504 0.65759 0.48543 0.0023611 0.42219 1.1128 1.1073 15.9992 144.9817 0.0005091 -83.0832 0.067958
0.172 0.98801 5.5246e-005 3.8182 0.012048 2.2676e-006 0.001154 0.052173 0.00065263 0.052822 0.046952 0 0.044479 0.0389 0 0.8471 0.22779 0.059075 0.0083715 4.1059 0.052715 6.288e-005 0.83735 0.0051043 0.0058422 0.0020946 0.9617 0.6823 4.6398e-006 1.857e-005 0.13045 0.64489 0.70057 0.0017371 0.6593 0.48559 0.0023414 0.42218 1.115 1.1095 15.9993 144.9817 0.00050739 -83.1699 0.068958
0.173 0.98801 5.5245e-005 3.8182 0.012048 2.2807e-006 0.001154 0.052321 0.00065266 0.052969 0.047086 0 0.044466 0.0389 0 0.84712 0.22779 0.059078 0.0083719 4.1059 0.052717 6.2882e-005 0.83735 0.0051043 0.0058422 0.0020674 0.96485 0.69844 4.5753e-006 1.8311e-005 0.13045 0.64593 0.70171 0.001725 0.66101 0.48576 0.0023238 0.42217 1.1172 1.1118 15.9994 144.9817 0.00050569 -83.2486 0.069958
0.174 0.98801 5.5245e-005 3.8182 0.012048 2.2939e-006 0.001154 0.052467 0.00065268 0.053115 0.04722 0 0.044452 0.0389 0 0.84714 0.2278 0.059082 0.0083723 4.1059 0.052719 6.2884e-005 0.83734 0.0051043 0.0058423 0.0020431 0.96747 0.71384 4.5176e-006 1.8079e-005 0.13045 0.64697 0.70285 0.0017141 0.66273 0.48593 0.002308 0.42216 1.1195 1.114 15.9995 144.9817 0.00050401 -83.3202 0.070958
0.175 0.98801 5.5245e-005 3.8182 0.012048 2.3071e-006 0.001154 0.052614 0.00065271 0.053262 0.047353 0 0.044439 0.0389 0 0.84716 0.22781 0.059085 0.0083727 4.1059 0.05272 6.2886e-005 0.83734 0.0051043 0.0058423 0.0020211 0.96965 0.72852 4.4653e-006 1.787e-005 0.13045 0.64801 0.70398 0.0017043 0.66445 0.48609 0.0022938 0.42215 1.1217 1.1163 15.9996 144.9817 0.00050233 -83.3854 0.071958
0.176 0.98801 5.5245e-005 3.8182 0.012048 2.3203e-006 0.001154 0.052761 0.00065273 0.053409 0.047487 0 0.044426 0.0389 0 0.84718 0.22782 0.059088 0.0083731 4.1059 0.052722 6.2889e-005 0.83734 0.0051043 0.0058423 0.0020013 0.97146 0.7425 4.4186e-006 1.7681e-005 0.13045 0.64904 0.7051 0.0016953 0.66617 0.48626 0.0022809 0.42214 1.1239 1.1185 15.9997 144.9817 0.00050066 -83.4449 0.072958
0.177 0.98801 5.5245e-005 3.8182 0.012048 2.3335e-006 0.001154 0.052907 0.00065276 0.053556 0.04762 0 0.044413 0.0389 0 0.8472 0.22783 0.059091 0.0083735 4.106 0.052724 6.2891e-005 0.83734 0.0051043 0.0058423 0.0019834 0.97297 0.7558 4.3767e-006 1.7511e-005 0.13045 0.65007 0.70622 0.0016872 0.66789 0.48642 0.0022692 0.42213 1.1261 1.1207 15.9998 144.9817 0.000499 -83.4992 0.073958
0.178 0.98801 5.5245e-005 3.8182 0.012048 2.3466e-006 0.001154 0.053054 0.00065279 0.053702 0.047753 0 0.044399 0.0389 0 0.84722 0.22784 0.059095 0.0083739 4.106 0.052726 6.2893e-005 0.83734 0.0051044 0.0058423 0.0019671 0.97423 0.76845 4.3382e-006 1.7357e-005 0.13045 0.6511 0.70732 0.0016798 0.66961 0.48659 0.0022586 0.42212 1.1283 1.1229 15.9999 144.9817 0.00049735 -83.549 0.074958
0.179 0.98801 5.5245e-005 3.8182 0.012048 2.3598e-006 0.001154 0.0532 0.00065281 0.053848 0.047886 0 0.044386 0.0389 0 0.84724 0.22785 0.059098 0.0083743 4.106 0.052727 6.2895e-005 0.83734 0.0051044 0.0058424 0.0019521 0.97528 0.78047 4.3027e-006 1.7216e-005 0.13045 0.65212 0.70842 0.0016731 0.67133 0.48676 0.002249 0.42211 1.1305 1.1252 16 144.9817 0.00049571 -83.5946 0.075958
0.18 0.98801 5.5245e-005 3.8182 0.012048 2.373e-006 0.001154 0.053346 0.00065284 0.053995 0.048019 0 0.044373 0.0389 0 0.84727 0.22786 0.059101 0.0083747 4.106 0.052729 6.2897e-005 0.83733 0.0051044 0.0058424 0.0019386 0.97616 0.79188 4.2707e-006 1.7088e-005 0.13045 0.65314 0.70951 0.0016669 0.67305 0.48693 0.0022402 0.4221 1.1327 1.1274 16 144.9817 0.00049407 -83.6366 0.076958
0.181 0.98801 5.5245e-005 3.8182 0.012048 2.3862e-006 0.001154 0.053492 0.00065286 0.054141 0.048152 0 0.04436 0.0389 0 0.84729 0.22787 0.059104 0.0083752 4.106 0.052731 6.29e-005 0.83733 0.0051044 0.0058424 0.0019262 0.97689 0.8027 4.2416e-006 1.6971e-005 0.13045 0.65416 0.71059 0.0016612 0.67476 0.48709 0.0022321 0.4221 1.1349 1.1296 16.0001 144.9817 0.00049245 -83.6753 0.077958
0.182 0.98801 5.5245e-005 3.8182 0.012048 2.3993e-006 0.001154 0.053638 0.00065289 0.054287 0.048285 0 0.044347 0.0389 0 0.84731 0.22788 0.059108 0.0083756 4.106 0.052733 6.2902e-005 0.83733 0.0051044 0.0058424 0.0019148 0.97751 0.81297 4.2149e-006 1.6863e-005 0.13045 0.65518 0.71167 0.001656 0.67648 0.48726 0.0022247 0.42209 1.1371 1.1318 16.0002 144.9817 0.00049083 -83.7111 0.078958
0.183 0.98801 5.5245e-005 3.8182 0.012048 2.4125e-006 0.001154 0.053784 0.00065291 0.054433 0.048418 0 0.044334 0.0389 0 0.84733 0.22789 0.059111 0.008376 4.106 0.052734 6.2904e-005 0.83733 0.0051045 0.0058424 0.0019043 0.97803 0.8227 4.1902e-006 1.6764e-005 0.13045 0.65619 0.71273 0.0016511 0.67819 0.48743 0.0022179 0.42209 1.1393 1.134 16.0003 144.9817 0.00048923 -83.7442 0.079958
0.184 0.98801 5.5245e-005 3.8182 0.012048 2.4257e-006 0.001154 0.05393 0.00065293 0.054578 0.04855 0 0.044321 0.0389 0 0.84735 0.2279 0.059115 0.0083764 4.1061 0.052736 6.2907e-005 0.83733 0.0051045 0.0058425 0.0018946 0.97848 0.83192 4.1673e-006 1.6672e-005 0.13045 0.6572 0.71379 0.0016467 0.67989 0.4876 0.0022117 0.42208 1.1415 1.1362 16.0004 144.9817 0.00048763 -83.7751 0.080958
0.185 0.98801 5.5245e-005 3.8182 0.012048 2.4389e-006 0.001154 0.054076 0.00065296 0.054724 0.048683 0 0.044307 0.0389 0 0.84737 0.2279 0.059118 0.0083769 4.1061 0.052738 6.2909e-005 0.83732 0.0051045 0.0058425 0.0018855 0.97885 0.84065 4.1459e-006 1.6587e-005 0.13045 0.65821 0.71485 0.0016425 0.6816 0.48776 0.0022058 0.42207 1.1437 1.1384 16.0005 144.9817 0.00048604 -83.8038 0.081958
0.186 0.98801 5.5245e-005 3.8182 0.012048 2.4521e-006 0.001154 0.054221 0.00065298 0.054869 0.048815 0 0.044294 0.0389 0 0.84739 0.22791 0.059121 0.0083773 4.1061 0.05274 6.2911e-005 0.83732 0.0051045 0.0058425 0.0018771 0.97918 0.84892 4.1262e-006 1.6508e-005 0.13045 0.65921 0.71589 0.0016386 0.68329 0.48793 0.0022004 0.42207 1.1458 1.1406 16.0006 144.9817 0.00048446 -83.8307 0.082958
0.187 0.98801 5.5245e-005 3.8182 0.012048 2.4652e-006 0.001154 0.054366 0.00065301 0.055015 0.048948 0 0.044281 0.0389 0 0.84741 0.22792 0.059125 0.0083777 4.1061 0.052742 6.2914e-005 0.83732 0.0051046 0.0058425 0.0018693 0.97946 0.85674 4.1079e-006 1.6434e-005 0.13045 0.66021 0.71693 0.001635 0.68499 0.4881 0.0021954 0.42206 1.148 1.1428 16.0007 144.9817 0.00048288 -83.8559 0.083958
0.188 0.98801 5.5245e-005 3.8182 0.012048 2.4784e-006 0.001154 0.054512 0.00065303 0.05516 0.04908 0 0.044268 0.0389 0 0.84744 0.22793 0.059128 0.0083782 4.1061 0.052744 6.2916e-005 0.83732 0.0051046 0.0058425 0.001862 0.9797 0.86414 4.0906e-006 1.6365e-005 0.13045 0.66121 0.71796 0.0016316 0.68668 0.48827 0.0021907 0.42206 1.1502 1.145 16.0007 144.9817 0.00048132 -83.8797 0.084958
0.189 0.98801 5.5244e-005 3.8182 0.012048 2.4916e-006 0.001154 0.054657 0.00065305 0.055305 0.049212 0 0.044255 0.0389 0 0.84746 0.22794 0.059132 0.0083786 4.1061 0.052746 6.2918e-005 0.83732 0.0051046 0.0058426 0.001855 0.97991 0.87115 4.0744e-006 1.63e-005 0.13045 0.66221 0.71899 0.0016284 0.68836 0.48844 0.0021863 0.42206 1.1523 1.1472 16.0008 144.9817 0.00047976 -83.9021 0.085958
0.19 0.98801 5.5244e-005 3.8182 0.012047 2.5048e-006 0.001154 0.054802 0.00065308 0.05545 0.049344 0 0.044242 0.0389 0 0.84748 0.22795 0.059135 0.008379 4.1062 0.052747 6.2921e-005 0.83732 0.0051046 0.0058426 0.0018485 0.9801 0.87777 4.0591e-006 1.6238e-005 0.13045 0.6632 0.72 0.0016253 0.69004 0.4886 0.0021821 0.42205 1.1545 1.1493 16.0009 144.9818 0.00047822 -83.9233 0.086958
0.191 0.98801 5.5244e-005 3.8182 0.012047 2.518e-006 0.001154 0.054947 0.0006531 0.055595 0.049476 0 0.044229 0.0389 0 0.8475 0.22796 0.059139 0.0083795 4.1062 0.052749 6.2923e-005 0.83731 0.0051046 0.0058426 0.0018423 0.98027 0.88404 4.0446e-006 1.618e-005 0.13045 0.66419 0.72101 0.0016224 0.69171 0.48877 0.0021782 0.42205 1.1567 1.1515 16.001 144.9818 0.00047668 -83.9435 0.087958
0.192 0.98801 5.5244e-005 3.8182 0.012047 2.5311e-006 0.001154 0.055092 0.00065312 0.05574 0.049608 0 0.044216 0.0389 0 0.84752 0.22797 0.059142 0.0083799 4.1062 0.052751 6.2926e-005 0.83731 0.0051047 0.0058426 0.0018364 0.98042 0.88996 4.0308e-006 1.6125e-005 0.13045 0.66518 0.72202 0.0016197 0.69338 0.48894 0.0021744 0.42205 1.1588 1.1537 16.0011 144.9818 0.00047515 -83.9627 0.088958
0.193 0.98801 5.5244e-005 3.8182 0.012047 2.5443e-006 0.001154 0.055236 0.00065315 0.055885 0.04974 0 0.044203 0.0389 0 0.84755 0.22798 0.059146 0.0083804 4.1062 0.052753 6.2928e-005 0.83731 0.0051047 0.0058426 0.0018309 0.98055 0.89555 4.0177e-006 1.6073e-005 0.13045 0.66616 0.72301 0.0016171 0.69504 0.48911 0.0021709 0.42204 1.161 1.1559 16.0011 144.9818 0.00047363 -83.9811 0.089958
0.194 0.98801 5.5244e-005 3.8182 0.012047 2.5575e-006 0.001154 0.055381 0.00065317 0.056029 0.049871 0 0.04419 0.0389 0 0.84757 0.22799 0.059149 0.0083808 4.1062 0.052755 6.2931e-005 0.83731 0.0051047 0.0058427 0.0018255 0.98067 0.90084 4.0052e-006 1.6023e-005 0.13045 0.66714 0.724 0.0016146 0.69669 0.48928 0.0021675 0.42204 1.1631 1.158 16.0012 144.9818 0.00047211 -83.9986 0.090958
0.195 0.98801 5.5244e-005 3.8182 0.012047 2.5707e-006 0.001154 0.055525 0.00065319 0.056174 0.050003 0 0.044178 0.0389 0 0.84759 0.228 0.059153 0.0083813 4.1062 0.052757 6.2933e-005 0.83731 0.0051047 0.0058427 0.0018204 0.98078 0.90584 3.9933e-006 1.5975e-005 0.13045 0.66812 0.72499 0.0016122 0.69834 0.48945 0.0021643 0.42204 1.1652 1.1602 16.0013 144.9818 0.00047061 -84.0155 0.091958
0.196 0.98801 5.5244e-005 3.8182 0.012047 2.5839e-006 0.001154 0.05567 0.00065321 0.056318 0.050134 0 0.044165 0.0389 0 0.84761 0.22801 0.059156 0.0083817 4.1063 0.052759 6.2936e-005 0.8373 0.0051048 0.0058427 0.0018155 0.98088 0.91056 3.9818e-006 1.5929e-005 0.13045 0.66909 0.72596 0.0016099 0.69998 0.48961 0.0021612 0.42203 1.1674 1.1623 16.0014 144.9818 0.00046911 -84.0318 0.092958
0.197 0.98801 5.5244e-005 3.8182 0.012047 2.597e-006 0.001154 0.055814 0.00065324 0.056462 0.050266 0 0.044152 0.0389 0 0.84764 0.22802 0.05916 0.0083822 4.1063 0.052761 6.2938e-005 0.8373 0.0051048 0.0058427 0.0018108 0.98098 0.91501 3.9708e-006 1.5884e-005 0.13045 0.67006 0.72693 0.0016077 0.70162 0.48978 0.0021582 0.42203 1.1695 1.1645 16.0015 144.9818 0.00046762 -84.0475 0.093958
0.198 0.98801 5.5244e-005 3.8182 0.012047 2.6102e-006 0.001154 0.055958 0.00065326 0.056607 0.050397 0 0.044139 0.0389 0 0.84766 0.22803 0.059163 0.0083826 4.1063 0.052763 6.2941e-005 0.8373 0.0051048 0.0058428 0.0018062 0.98106 0.91922 3.9601e-006 1.5842e-005 0.13045 0.67103 0.7279 0.0016056 0.70325 0.48995 0.0021553 0.42203 1.1716 1.1666 16.0015 144.9818 0.00046614 -84.0627 0.094958
0.199 0.98801 5.5244e-005 3.8182 0.012047 2.6234e-006 0.001154 0.056102 0.00065328 0.056751 0.050528 0 0.044126 0.0389 0 0.84768 0.22804 0.059167 0.0083831 4.1063 0.052765 6.2943e-005 0.8373 0.0051048 0.0058428 0.0018018 0.98115 0.9232 3.9497e-006 1.58e-005 0.13045 0.672 0.72886 0.0016035 0.70487 0.49012 0.0021526 0.42203 1.1738 1.1688 16.0016 144.9818 0.00046467 -84.0774 0.095958
0.2 0.98801 5.5244e-005 3.8182 0.012047 2.6366e-006 0.001154 0.056246 0.0006533 0.056894 0.050659 0 0.044113 0.0389 0 0.8477 0.22805 0.059171 0.0083835 4.1063 0.052767 6.2946e-005 0.8373 0.0051048 0.0058428 0.0017975 0.98122 0.92696 3.9398e-006 1.576e-005 0.13045 0.67296 0.72981 0.0016015 0.70648 0.49029 0.0021499 0.42202 1.1759 1.1709 16.0017 144.9818 0.0004632 -84.0917 0.096958
0.201 0.98801 5.5244e-005 3.8182 0.012047 2.6497e-006 0.001154 0.05639 0.00065332 0.057038 0.05079 0 0.0441 0.0389 0 0.84773 0.22806 0.059174 0.008384 4.1063 0.052769 6.2948e-005 0.83729 0.0051049 0.0058428 0.0017934 0.9813 0.9305 3.93e-006 1.5721e-005 0.13045 0.67392 0.73075 0.0015995 0.70809 0.49046 0.0021473 0.42202 1.178 1.173 16.0018 144.9818 0.00046175 -84.1056 0.097958
0.202 0.98801 5.5244e-005 3.8182 0.012047 2.6629e-006 0.001154 0.056533 0.00065335 0.057182 0.050921 0 0.044088 0.0389 0 0.84775 0.22807 0.059178 0.0083845 4.1064 0.052771 6.2951e-005 0.83729 0.0051049 0.0058429 0.0017893 0.98137 0.93385 3.9206e-006 1.5684e-005 0.13045 0.67488 0.73169 0.0015976 0.7097 0.49063 0.0021447 0.42202 1.1801 1.1752 16.0019 144.9819 0.0004603 -84.1192 0.098958
0.203 0.98801 5.5244e-005 3.8182 0.012047 2.6761e-006 0.001154 0.056677 0.00065337 0.057325 0.051051 0 0.044075 0.0389 0 0.84777 0.22808 0.059182 0.0083849 4.1064 0.052773 6.2954e-005 0.83729 0.0051049 0.0058429 0.0017853 0.98143 0.93701 3.9114e-006 1.5647e-005 0.13045 0.67583 0.73262 0.0015958 0.71129 0.49079 0.0021423 0.42202 1.1822 1.1773 16.0019 144.9819 0.00045886 -84.1325 0.099958
0.204 0.98801 5.5244e-005 3.8182 0.012047 2.6893e-006 0.001154 0.05682 0.00065339 0.057469 0.051182 0 0.044062 0.0389 0 0.8478 0.22809 0.059185 0.0083854 4.1064 0.052775 6.2956e-005 0.83729 0.0051049 0.0058429 0.0017815 0.9815 0.93999 3.9024e-006 1.5611e-005 0.13046 0.67679 0.73355 0.001594 0.71288 0.49096 0.0021399 0.42202 1.1843 1.1794 16.002 144.9819 0.00045742 -84.1455 0.10096
0.205 0.98801 5.5243e-005 3.8182 0.012047 2.7025e-006 0.001154 0.056963 0.00065341 0.057612 0.051313 0 0.044049 0.0389 0 0.84782 0.2281 0.059189 0.0083859 4.1064 0.052777 6.2959e-005 0.83729 0.005105 0.0058429 0.0017778 0.98156 0.9428 3.8937e-006 1.5576e-005 0.13046 0.67773 0.73447 0.0015922 0.71446 0.49113 0.0021375 0.42202 1.1864 1.1815 16.0021 144.9819 0.000456 -84.1582 0.10196
0.206 0.98801 5.5243e-005 3.8182 0.012047 2.7156e-006 0.001154 0.057107 0.00065343 0.057755 0.051443 0 0.044037 0.0389 0 0.84784 0.22811 0.059193 0.0083863 4.1064 0.05278 6.2962e-005 0.83728 0.005105 0.0058429 0.0017742 0.98162 0.94546 3.8852e-006 1.5541e-005 0.13046 0.67868 0.73539 0.0015904 0.71604 0.4913 0.0021352 0.42202 1.1885 1.1837 16.0022 144.9819 0.00045458 -84.1706 0.10296
0.207 0.98801 5.5243e-005 3.8182 0.012047 2.7288e-006 0.001154 0.05725 0.00065345 0.057898 0.051573 0 0.044024 0.0389 0 0.84787 0.22812 0.059197 0.0083868 4.1065 0.052782 6.2964e-005 0.83728 0.005105 0.005843 0.0017706 0.98167 0.94796 3.8768e-006 1.5508e-005 0.13046 0.67962 0.73629 0.0015887 0.71761 0.49147 0.002133 0.42201 1.1906 1.1858 16.0022 144.9819 0.00045317 -84.1829 0.10396
0.208 0.98801 5.5243e-005 3.8182 0.012047 2.742e-006 0.001154 0.057393 0.00065347 0.058041 0.051704 0 0.044011 0.0389 0 0.84789 0.22813 0.0592 0.0083873 4.1065 0.052784 6.2967e-005 0.83728 0.005105 0.005843 0.001767 0.98173 0.95033 3.8685e-006 1.5475e-005 0.13046 0.68056 0.7372 0.0015871 0.71917 0.49164 0.0021308 0.42201 1.1927 1.1879 16.0023 144.9819 0.00045177 -84.1949 0.10496
0.209 0.98801 5.5243e-005 3.8182 0.012047 2.7552e-006 0.001154 0.057535 0.00065349 0.058184 0.051834 0 0.043998 0.0389 0 0.84791 0.22814 0.059204 0.0083878 4.1065 0.052786 6.297e-005 0.83728 0.0051051 0.005843 0.0017635 0.98178 0.95256 3.8604e-006 1.5442e-005 0.13046 0.6815 0.73809 0.0015854 0.72073 0.49181 0.0021286 0.42201 1.1948 1.19 16.0024 144.9819 0.00045037 -84.2067 0.10596
0.21 0.98801 5.5243e-005 3.8182 0.012047 2.7684e-006 0.001154 0.057678 0.00065351 0.058327 0.051964 0 0.043986 0.0389 0 0.84794 0.22815 0.059208 0.0083882 4.1065 0.052788 6.2972e-005 0.83727 0.0051051 0.005843 0.0017601 0.98184 0.95467 3.8524e-006 1.5411e-005 0.13046 0.68244 0.73899 0.0015838 0.72227 0.49197 0.0021265 0.42201 1.1969 1.1921 16.0025 144.9819 0.00044898 -84.2184 0.10696
0.211 0.98801 5.5243e-005 3.8182 0.012047 2.7815e-006 0.001154 0.057821 0.00065353 0.05847 0.052094 0 0.043973 0.0389 0 0.84796 0.22816 0.059212 0.0083887 4.1065 0.05279 6.2975e-005 0.83727 0.0051051 0.0058431 0.0017567 0.98189 0.95666 3.8445e-006 1.5379e-005 0.13046 0.68337 0.73987 0.0015822 0.72382 0.49214 0.0021244 0.42201 1.199 1.1942 16.0025 144.9819 0.0004476 -84.2298 0.10796
0.212 0.98801 5.5243e-005 3.8182 0.012047 2.7947e-006 0.001154 0.057963 0.00065355 0.058612 0.052224 0 0.043961 0.0389 0 0.84799 0.22818 0.059216 0.0083892 4.1066 0.052793 6.2978e-005 0.83727 0.0051052 0.0058431 0.0017534 0.98194 0.95853 3.8368e-006 1.5348e-005 0.13046 0.6843 0.74075 0.0015806 0.72535 0.49231 0.0021223 0.42201 1.201 1.1963 16.0026 144.9819 0.00044623 -84.2412 0.10896
0.213 0.98801 5.5243e-005 3.8182 0.012047 2.8079e-006 0.001154 0.058106 0.00065357 0.058755 0.052354 0 0.043948 0.0389 0 0.84801 0.22819 0.059219 0.0083897 4.1066 0.052795 6.2981e-005 0.83727 0.0051052 0.0058431 0.0017501 0.98199 0.9603 3.8293e-006 1.5318e-005 0.13046 0.68522 0.74163 0.0015791 0.72688 0.49248 0.0021203 0.42201 1.2031 1.1984 16.0027 144.982 0.00044486 -84.2523 0.10996
0.214 0.98801 5.5243e-005 3.8182 0.012047 2.8211e-006 0.001154 0.058248 0.00065359 0.058897 0.052483 0 0.043935 0.0389 0 0.84804 0.2282 0.059223 0.0083902 4.1066 0.052797 6.2983e-005 0.83727 0.0051052 0.0058432 0.0017469 0.98203 0.96197 3.8218e-006 1.5288e-005 0.13046 0.68615 0.7425 0.0015776 0.7284 0.49265 0.0021183 0.42201 1.2052 1.2004 16.0027 144.982 0.00044351 -84.2634 0.11096
0.215 0.98801 5.5243e-005 3.8182 0.012047 2.8342e-006 0.001154 0.05839 0.00065361 0.059039 0.052613 0 0.043923 0.0389 0 0.84806 0.22821 0.059227 0.0083907 4.1066 0.052799 6.2986e-005 0.83726 0.0051052 0.0058432 0.0017438 0.98208 0.96354 3.8145e-006 1.5259e-005 0.13046 0.68707 0.74336 0.0015761 0.72991 0.49282 0.0021163 0.42201 1.2072 1.2025 16.0028 144.982 0.00044215 -84.2742 0.11196
0.216 0.98801 5.5243e-005 3.8182 0.012047 2.8474e-006 0.001154 0.058532 0.00065363 0.059181 0.052742 0 0.04391 0.0389 0 0.84808 0.22822 0.059231 0.0083911 4.1066 0.052801 6.2989e-005 0.83726 0.0051053 0.0058432 0.0017407 0.98213 0.96503 3.8073e-006 1.523e-005 0.13046 0.68798 0.74422 0.0015746 0.73142 0.49299 0.0021144 0.42201 1.2093 1.2046 16.0029 144.982 0.00044081 -84.285 0.11296
0.217 0.98801 5.5243e-005 3.8182 0.012047 2.8606e-006 0.001154 0.058674 0.00065365 0.059323 0.052872 0 0.043898 0.0389 0 0.84811 0.22823 0.059235 0.0083916 4.1067 0.052804 6.2992e-005 0.83726 0.0051053 0.0058432 0.0017377 0.98217 0.96643 3.8001e-006 1.5201e-005 0.13046 0.6889 0.74507 0.0015731 0.73292 0.49316 0.0021125 0.42201 1.2114 1.2067 16.003 144.982 0.00043947 -84.2956 0.11396
0.218 0.98801 5.5243e-005 3.8182 0.012047 2.8738e-006 0.001154 0.058816 0.00065367 0.059465 0.053001 0 0.043885 0.0389 0 0.84813 0.22824 0.059239 0.0083921 4.1067 0.052806 6.2995e-005 0.83726 0.0051053 0.0058433 0.0017346 0.98221 0.96775 3.793e-006 1.5173e-005 0.13046 0.68981 0.74592 0.0015717 0.73441 0.49332 0.0021106 0.42201 1.2134 1.2087 16.003 144.982 0.00043814 -84.3061 0.11496
0.219 0.98801 5.5243e-005 3.8182 0.012047 2.887e-006 0.001154 0.058958 0.00065369 0.059607 0.05313 0 0.043873 0.0389 0 0.84816 0.22825 0.059243 0.0083926 4.1067 0.052808 6.2998e-005 0.83725 0.0051053 0.0058433 0.0017316 0.98226 0.969 3.786e-006 1.5145e-005 0.13046 0.69072 0.74676 0.0015703 0.7359 0.49349 0.0021087 0.42201 1.2155 1.2108 16.0031 144.982 0.00043682 -84.3165 0.11596
0.22 0.98801 5.5243e-005 3.8182 0.012047 2.9001e-006 0.001154 0.059099 0.00065371 0.059748 0.053259 0 0.04386 0.0389 0 0.84818 0.22826 0.059247 0.0083931 4.1067 0.05281 6.3001e-005 0.83725 0.0051054 0.0058433 0.0017286 0.9823 0.97017 3.7791e-006 1.5117e-005 0.13046 0.69163 0.7476 0.0015688 0.73738 0.49366 0.0021068 0.42201 1.2175 1.2128 16.0032 144.982 0.00043551 -84.3268 0.11696
0.221 0.98801 5.5243e-005 3.8182 0.012047 2.9133e-006 0.001154 0.059241 0.00065373 0.05989 0.053388 0 0.043848 0.0389 0 0.84821 0.22827 0.059251 0.0083936 4.1067 0.052813 6.3004e-005 0.83725 0.0051054 0.0058433 0.0017257 0.98234 0.97128 3.7723e-006 1.509e-005 0.13046 0.69253 0.74843 0.0015674 0.73885 0.49383 0.002105 0.42201 1.2195 1.2149 16.0032 144.982 0.0004342 -84.337 0.11796
0.222 0.98801 5.5242e-005 3.8182 0.012047 2.9265e-006 0.001154 0.059382 0.00065375 0.060031 0.053517 0 0.043835 0.0389 0 0.84823 0.22828 0.059255 0.0083941 4.1068 0.052815 6.3006e-005 0.83725 0.0051054 0.0058434 0.0017228 0.98238 0.97233 3.7656e-006 1.5063e-005 0.13046 0.69343 0.74926 0.0015661 0.74032 0.494 0.0021032 0.42202 1.2216 1.217 16.0033 144.982 0.0004329 -84.3471 0.11896
0.223 0.98801 5.5242e-005 3.8182 0.012047 2.9397e-006 0.001154 0.059523 0.00065377 0.060172 0.053646 0 0.043823 0.0389 0 0.84826 0.2283 0.059259 0.0083946 4.1068 0.052817 6.3009e-005 0.83725 0.0051055 0.0058434 0.0017199 0.98243 0.97332 3.7589e-006 1.5037e-005 0.13046 0.69433 0.75008 0.0015647 0.74178 0.49417 0.0021014 0.42202 1.2236 1.219 16.0034 144.9821 0.0004316 -84.3571 0.11996
0.224 0.98801 5.5242e-005 3.8182 0.012047 2.9528e-006 0.001154 0.059664 0.00065379 0.060313 0.053775 0 0.04381 0.0389 0 0.84828 0.22831 0.059263 0.0083951 4.1068 0.05282 6.3012e-005 0.83724 0.0051055 0.0058434 0.0017171 0.98247 0.97425 3.7524e-006 1.501e-005 0.13046 0.69522 0.7509 0.0015633 0.74323 0.49434 0.0020996 0.42202 1.2256 1.221 16.0034 144.9821 0.00043031 -84.367 0.12096
0.225 0.98801 5.5242e-005 3.8182 0.012047 2.966e-006 0.001154 0.059805 0.0006538 0.060455 0.053903 0 0.043798 0.0389 0 0.84831 0.22832 0.059267 0.0083956 4.1068 0.052822 6.3015e-005 0.83724 0.0051055 0.0058435 0.0017143 0.98251 0.97513 3.7459e-006 1.4984e-005 0.13046 0.69612 0.75171 0.001562 0.74468 0.49451 0.0020979 0.42202 1.2276 1.2231 16.0035 144.9821 0.00042903 -84.3768 0.12196
0.226 0.98801 5.5242e-005 3.8182 0.012047 2.9792e-006 0.001154 0.059946 0.00065382 0.060595 0.054032 0 0.043785 0.0389 0 0.84833 0.22833 0.059271 0.0083962 4.1068 0.052824 6.3018e-005 0.83724 0.0051055 0.0058435 0.0017116 0.98255 0.97595 3.7395e-006 1.4959e-005 0.13046 0.69701 0.75252 0.0015607 0.74611 0.49467 0.0020961 0.42202 1.2297 1.2251 16.0036 144.9821 0.00042776 -84.3865 0.12296
0.227 0.98801 5.5242e-005 3.8182 0.012047 2.9924e-006 0.001154 0.060087 0.00065384 0.060736 0.05416 0 0.043773 0.0389 0 0.84836 0.22834 0.059275 0.0083967 4.1069 0.052827 6.3021e-005 0.83724 0.0051056 0.0058435 0.0017089 0.98258 0.97673 3.7331e-006 1.4933e-005 0.13046 0.69789 0.75332 0.0015594 0.74755 0.49484 0.0020944 0.42202 1.2317 1.2271 16.0036 144.9821 0.00042649 -84.3961 0.12396
0.228 0.98801 5.5242e-005 3.8182 0.012047 3.0055e-006 0.001154 0.060228 0.00065386 0.060877 0.054288 0 0.043761 0.0389 0 0.84839 0.22835 0.059279 0.0083972 4.1069 0.052829 6.3024e-005 0.83723 0.0051056 0.0058435 0.0017062 0.98262 0.97747 3.7268e-006 1.4908e-005 0.13046 0.69878 0.75412 0.0015581 0.74897 0.49501 0.0020927 0.42202 1.2337 1.2292 16.0037 144.9821 0.00042523 -84.4056 0.12496
0.229 0.98801 5.5242e-005 3.8182 0.012047 3.0187e-006 0.001154 0.060368 0.00065388 0.061018 0.054417 0 0.043748 0.0389 0 0.84841 0.22836 0.059283 0.0083977 4.1069 0.052832 6.3027e-005 0.83723 0.0051056 0.0058436 0.0017035 0.98266 0.97817 3.7206e-006 1.4883e-005 0.13046 0.69966 0.75491 0.0015568 0.75039 0.49518 0.002091 0.42203 1.2357 1.2312 16.0038 144.9821 0.00042398 -84.4151 0.12596
0.23 0.98801 5.5242e-005 3.8182 0.012047 3.0319e-006 0.001154 0.060509 0.0006539 0.061158 0.054545 0 0.043736 0.0389 0 0.84844 0.22837 0.059287 0.0083982 4.1069 0.052834 6.303e-005 0.83723 0.0051057 0.0058436 0.0017008 0.9827 0.97882 3.7144e-006 1.4858e-005 0.13046 0.70054 0.7557 0.0015555 0.7518 0.49535 0.0020894 0.42203 1.2377 1.2332 16.0038 144.9821 0.00042273 -84.4245 0.12696
0.231 0.98801 5.5242e-005 3.8182 0.012047 3.0451e-006 0.001154 0.060649 0.00065391 0.061298 0.054673 0 0.043724 0.0389 0 0.84846 0.22839 0.059291 0.0083987 4.107 0.052836 6.3034e-005 0.83723 0.0051057 0.0058436 0.0016982 0.98274 0.97944 3.7083e-006 1.4834e-005 0.13046 0.70142 0.75648 0.0015542 0.75321 0.49552 0.0020877 0.42203 1.2397 1.2352 16.0039 144.9821 0.00042149 -84.4338 0.12796
0.232 0.98801 5.5242e-005 3.8182 0.012047 3.0583e-006 0.001154 0.060789 0.00065393 0.061439 0.054801 0 0.043711 0.0389 0 0.84849 0.2284 0.059295 0.0083992 4.107 0.052839 6.3037e-005 0.83722 0.0051057 0.0058437 0.0016956 0.98277 0.98003 3.7023e-006 1.481e-005 0.13046 0.70229 0.75726 0.001553 0.7546 0.49569 0.0020861 0.42203 1.2417 1.2372 16.004 144.9822 0.00042025 -84.443 0.12896
0.233 0.98801 5.5242e-005 3.8182 0.012047 3.0714e-006 0.001154 0.060929 0.00065395 0.061579 0.054929 0 0.043699 0.0389 0 0.84852 0.22841 0.059299 0.0083998 4.107 0.052841 6.304e-005 0.83722 0.0051058 0.0058437 0.001693 0.98281 0.98058 3.6963e-006 1.4786e-005 0.13046 0.70316 0.75804 0.0015517 0.756 0.49586 0.0020844 0.42203 1.2437 1.2392 16.004 144.9822 0.00041903 -84.4521 0.12996
0.234 0.98801 5.5242e-005 3.8182 0.012047 3.0846e-006 0.001154 0.061069 0.00065397 0.061719 0.055056 0 0.043687 0.0389 0 0.84854 0.22842 0.059303 0.0084003 4.107 0.052844 6.3043e-005 0.83722 0.0051058 0.0058437 0.0016904 0.98285 0.9811 3.6903e-006 1.4762e-005 0.13046 0.70403 0.75881 0.0015505 0.75738 0.49602 0.0020828 0.42204 1.2456 1.2412 16.0041 144.9822 0.0004178 -84.4612 0.13096
0.235 0.98801 5.5242e-005 3.8182 0.012047 3.0978e-006 0.001154 0.061209 0.00065398 0.061859 0.055184 0 0.043675 0.0389 0 0.84857 0.22843 0.059308 0.0084008 4.1071 0.052846 6.3046e-005 0.83722 0.0051058 0.0058438 0.0016879 0.98288 0.98159 3.6845e-006 1.4739e-005 0.13046 0.7049 0.75957 0.0015493 0.75876 0.49619 0.0020812 0.42204 1.2476 1.2432 16.0041 144.9822 0.00041659 -84.4701 0.13196
0.236 0.98801 5.5242e-005 3.8182 0.012047 3.111e-006 0.001154 0.061349 0.000654 0.061998 0.055311 0 0.043662 0.0389 0 0.84859 0.22844 0.059312 0.0084014 4.1071 0.052849 6.3049e-005 0.83721 0.0051059 0.0058438 0.0016854 0.98292 0.98205 3.6787e-006 1.4715e-005 0.13046 0.70576 0.76033 0.0015481 0.76013 0.49636 0.0020797 0.42204 1.2496 1.2452 16.0042 144.9822 0.00041538 -84.479 0.13296
0.237 0.98801 5.5242e-005 3.8182 0.012047 3.1241e-006 0.001154 0.061489 0.00065402 0.062138 0.055439 0 0.04365 0.0389 0 0.84862 0.22845 0.059316 0.0084019 4.1071 0.052851 6.3052e-005 0.83721 0.0051059 0.0058438 0.0016829 0.98295 0.98249 3.6729e-006 1.4692e-005 0.13046 0.70662 0.76109 0.0015469 0.7615 0.49653 0.0020781 0.42204 1.2516 1.2472 16.0043 144.9822 0.00041418 -84.4879 0.13396
0.238 0.98801 5.5241e-005 3.8182 0.012047 3.1373e-006 0.001154 0.061628 0.00065404 0.062278 0.055566 0 0.043638 0.0389 0 0.84865 0.22847 0.05932 0.0084024 4.1071 0.052854 6.3056e-005 0.83721 0.0051059 0.0058438 0.0016805 0.98299 0.9829 3.6673e-006 1.467e-005 0.13046 0.70748 0.76184 0.0015457 0.76285 0.4967 0.0020766 0.42205 1.2535 1.2492 16.0043 144.9822 0.00041298 -84.4966 0.13496
0.239 0.98801 5.5241e-005 3.8182 0.012047 3.1505e-006 0.001154 0.061768 0.00065405 0.062417 0.055694 0 0.043626 0.0389 0 0.84867 0.22848 0.059324 0.0084029 4.1072 0.052856 6.3059e-005 0.83721 0.0051059 0.0058439 0.0016781 0.98302 0.98329 3.6616e-006 1.4647e-005 0.13046 0.70833 0.76259 0.0015445 0.76421 0.49687 0.002075 0.42205 1.2555 1.2512 16.0044 144.9822 0.00041179 -84.5053 0.13596
0.24 0.98801 5.5241e-005 3.8182 0.012047 3.1637e-006 0.001154 0.061907 0.00065407 0.062557 0.055821 0 0.043614 0.0389 0 0.8487 0.22849 0.059329 0.0084035 4.1072 0.052859 6.3062e-005 0.8372 0.005106 0.0058439 0.0016757 0.98305 0.98366 3.656e-006 1.4625e-005 0.13046 0.70919 0.76333 0.0015434 0.76555 0.49704 0.0020735 0.42205 1.2575 1.2531 16.0044 144.9822 0.00041061 -84.5139 0.13696
0.241 0.98801 5.5241e-005 3.8182 0.012047 3.1769e-006 0.001154 0.062046 0.00065409 0.062696 0.055948 0 0.043601 0.0389 0 0.84873 0.2285 0.059333 0.008404 4.1072 0.052861 6.3065e-005 0.8372 0.005106 0.0058439 0.0016733 0.98309 0.98401 3.6505e-006 1.4603e-005 0.13046 0.71004 0.76407 0.0015422 0.76689 0.4972 0.002072 0.42205 1.2594 1.2551 16.0045 144.9823 0.00040943 -84.5225 0.13796
0.242 0.98801 5.5241e-005 3.8182 0.012047 3.19e-006 0.001154 0.062185 0.0006541 0.062835 0.056075 0 0.043589 0.0389 0 0.84875 0.22851 0.059337 0.0084046 4.1072 0.052864 6.3068e-005 0.8372 0.005106 0.005844 0.001671 0.98312 0.98433 3.6451e-006 1.4581e-005 0.13046 0.71088 0.7648 0.0015411 0.76822 0.49737 0.0020705 0.42206 1.2614 1.2571 16.0046 144.9823 0.00040826 -84.531 0.13896
0.243 0.98801 5.5241e-005 3.8182 0.012047 3.2032e-006 0.001154 0.062324 0.00065412 0.062974 0.056202 0 0.043577 0.0389 0 0.84878 0.22853 0.059341 0.0084051 4.1073 0.052867 6.3072e-005 0.8372 0.0051061 0.005844 0.0016686 0.98315 0.98464 3.6396e-006 1.4559e-005 0.13046 0.71173 0.76553 0.0015399 0.76955 0.49754 0.002069 0.42206 1.2633 1.259 16.0046 144.9823 0.00040709 -84.5394 0.13996
0.244 0.98801 5.5241e-005 3.8182 0.012047 3.2164e-006 0.001154 0.062463 0.00065414 0.063113 0.056328 0 0.043565 0.0389 0 0.84881 0.22854 0.059346 0.0084056 4.1073 0.052869 6.3075e-005 0.83719 0.0051061 0.005844 0.0016663 0.98318 0.98494 3.6343e-006 1.4538e-005 0.13046 0.71257 0.76626 0.0015388 0.77087 0.49771 0.0020675 0.42206 1.2652 1.261 16.0047 144.9823 0.00040593 -84.5477 0.14096
0.245 0.98801 5.5241e-005 3.8182 0.012047 3.2296e-006 0.001154 0.062602 0.00065415 0.063252 0.056455 0 0.043553 0.0389 0 0.84884 0.22855 0.05935 0.0084062 4.1073 0.052872 6.3078e-005 0.83719 0.0051062 0.0058441 0.001664 0.98322 0.98521 3.629e-006 1.4516e-005 0.13047 0.71341 0.76698 0.0015377 0.77218 0.49788 0.0020661 0.42207 1.2672 1.2629 16.0047 144.9823 0.00040478 -84.556 0.14196
0.246 0.98801 5.5241e-005 3.8182 0.012047 3.2427e-006 0.001154 0.062741 0.00065417 0.06339 0.056582 0 0.043541 0.0389 0 0.84886 0.22856 0.059354 0.0084067 4.1073 0.052874 6.3082e-005 0.83719 0.0051062 0.0058441 0.0016618 0.98325 0.98547 3.6237e-006 1.4495e-005 0.13047 0.71425 0.7677 0.0015366 0.77348 0.49805 0.0020646 0.42207 1.2691 1.2649 16.0048 144.9823 0.00040363 -84.5642 0.14296
0.247 0.98801 5.5241e-005 3.8182 0.012047 3.2559e-006 0.001154 0.062879 0.00065419 0.063529 0.056708 0 0.043529 0.0389 0 0.84889 0.22857 0.059359 0.0084073 4.1074 0.052877 6.3085e-005 0.83719 0.0051062 0.0058441 0.0016595 0.98328 0.98572 3.6185e-006 1.4474e-005 0.13047 0.71508 0.76841 0.0015355 0.77478 0.49822 0.0020632 0.42207 1.271 1.2668 16.0049 144.9823 0.00040249 -84.5723 0.14396
0.248 0.98801 5.5241e-005 3.8182 0.012047 3.2691e-006 0.001154 0.063018 0.0006542 0.063667 0.056835 0 0.043517 0.0389 0 0.84892 0.22859 0.059363 0.0084078 4.1074 0.05288 6.3088e-005 0.83718 0.0051063 0.0058442 0.0016573 0.98331 0.98595 3.6133e-006 1.4454e-005 0.13047 0.71591 0.76912 0.0015344 0.77608 0.49838 0.0020618 0.42208 1.273 1.2688 16.0049 144.9823 0.00040135 -84.5804 0.14496
0.249 0.98801 5.5241e-005 3.8182 0.012047 3.2823e-006 0.001154 0.063156 0.00065422 0.063806 0.056961 0 0.043505 0.0389 0 0.84895 0.2286 0.059368 0.0084084 4.1074 0.052882 6.3092e-005 0.83718 0.0051063 0.0058442 0.001655 0.98334 0.98617 3.6082e-006 1.4433e-005 0.13047 0.71674 0.76983 0.0015333 0.77736 0.49855 0.0020604 0.42208 1.2749 1.2707 16.005 144.9824 0.00040022 -84.5884 0.14596
0.25 0.98801 5.5241e-005 3.8182 0.012047 3.2954e-006 0.001154 0.063294 0.00065423 0.063944 0.057087 0 0.043493 0.0389 0 0.84897 0.22861 0.059372 0.0084089 4.1074 0.052885 6.3095e-005 0.83718 0.0051063 0.0058442 0.0016529 0.98337 0.98638 3.6031e-006 1.4413e-005 0.13047 0.71757 0.77053 0.0015323 0.77864 0.49872 0.002059 0.42208 1.2768 1.2726 16.005 144.9824 0.0003991 -84.5964 0.14696
0.251 0.98801 5.5241e-005 3.8182 0.012047 3.3086e-006 0.001154 0.063432 0.00065425 0.064082 0.057213 0 0.043481 0.0389 0 0.849 0.22862 0.059376 0.0084095 4.1075 0.052888 6.3098e-005 0.83718 0.0051064 0.0058443 0.0016507 0.9834 0.98658 3.5981e-006 1.4393e-005 0.13047 0.7184 0.77122 0.0015312 0.77992 0.49889 0.0020576 0.42209 1.2787 1.2746 16.0051 144.9824 0.00039798 -84.6043 0.14796
0.252 0.98801 5.5241e-005 3.8182 0.012047 3.3218e-006 0.001154 0.06357 0.00065427 0.06422 0.057339 0 0.043469 0.0389 0 0.84903 0.22863 0.059381 0.0084101 4.1075 0.05289 6.3102e-005 0.83717 0.0051064 0.0058443 0.0016485 0.98343 0.98676 3.5931e-006 1.4373e-005 0.13047 0.71922 0.77192 0.0015302 0.78118 0.49906 0.0020562 0.42209 1.2806 1.2765 16.0051 144.9824 0.00039687 -84.6121 0.14896
0.253 0.98801 5.5241e-005 3.8182 0.012047 3.335e-006 0.001154 0.063708 0.00065428 0.064358 0.057465 0 0.043457 0.0389 0 0.84906 0.22865 0.059385 0.0084106 4.1075 0.052893 6.3105e-005 0.83717 0.0051064 0.0058443 0.0016464 0.98346 0.98694 3.5881e-006 1.4353e-005 0.13047 0.72004 0.77261 0.0015291 0.78244 0.49923 0.0020549 0.4221 1.2825 1.2784 16.0052 144.9824 0.00039576 -84.6199 0.14996
0.254 0.98801 5.524e-005 3.8182 0.012047 3.3481e-006 0.001154 0.063846 0.0006543 0.064496 0.057591 0 0.043445 0.0389 0 0.84909 0.22866 0.05939 0.0084112 4.1075 0.052896 6.3109e-005 0.83717 0.0051065 0.0058444 0.0016443 0.98349 0.9871 3.5832e-006 1.4334e-005 0.13047 0.72085 0.77329 0.0015281 0.7837 0.4994 0.0020535 0.4221 1.2844 1.2803 16.0052 144.9824 0.00039466 -84.6276 0.15096
0.255 0.98801 5.524e-005 3.8182 0.012047 3.3613e-006 0.001154 0.063984 0.00065431 0.064633 0.057717 0 0.043433 0.0389 0 0.84911 0.22867 0.059394 0.0084117 4.1076 0.052898 6.3112e-005 0.83716 0.0051065 0.0058444 0.0016422 0.98352 0.98726 3.5784e-006 1.4314e-005 0.13047 0.72167 0.77397 0.0015271 0.78495 0.49956 0.0020522 0.4221 1.2863 1.2822 16.0053 144.9824 0.00039357 -84.6352 0.15196
0.256 0.98802 5.524e-005 3.8182 0.012047 3.3745e-006 0.001154 0.064121 0.00065433 0.064771 0.057842 0 0.043421 0.0389 0 0.84914 0.22868 0.059399 0.0084123 4.1076 0.052901 6.3116e-005 0.83716 0.0051065 0.0058445 0.0016401 0.98355 0.98741 3.5736e-006 1.4295e-005 0.13047 0.72248 0.77465 0.001526 0.78619 0.49973 0.0020509 0.42211 1.2882 1.2841 16.0054 144.9824 0.00039248 -84.6428 0.15296
0.257 0.98802 5.524e-005 3.8182 0.012047 3.3877e-006 0.001154 0.064259 0.00065434 0.064908 0.057968 0 0.043409 0.0389 0 0.84917 0.2287 0.059403 0.0084129 4.1076 0.052904 6.3119e-005 0.83716 0.0051066 0.0058445 0.0016381 0.98358 0.98755 3.5688e-006 1.4276e-005 0.13047 0.72329 0.77533 0.001525 0.78742 0.4999 0.0020496 0.42211 1.2901 1.286 16.0054 144.9825 0.00039139 -84.6503 0.15396
0.258 0.98802 5.524e-005 3.8182 0.012047 3.4008e-006 0.001154 0.064396 0.00065436 0.065046 0.058093 0 0.043397 0.0389 0 0.8492 0.22871 0.059408 0.0084134 4.1077 0.052907 6.3123e-005 0.83716 0.0051066 0.0058445 0.001636 0.98361 0.98769 3.5641e-006 1.4257e-005 0.13047 0.7241 0.776 0.001524 0.78865 0.50007 0.0020482 0.42212 1.292 1.2879 16.0055 144.9825 0.00039031 -84.6578 0.15496
0.259 0.98802 5.524e-005 3.8182 0.012047 3.414e-006 0.001154 0.064533 0.00065437 0.065183 0.058219 0 0.043385 0.0389 0 0.84923 0.22872 0.059412 0.008414 4.1077 0.052909 6.3126e-005 0.83715 0.0051067 0.0058446 0.001634 0.98363 0.98781 3.5595e-006 1.4238e-005 0.13047 0.7249 0.77666 0.0015231 0.78988 0.50024 0.002047 0.42212 1.2939 1.2898 16.0055 144.9825 0.00038924 -84.6652 0.15596
0.26 0.98802 5.524e-005 3.8182 0.012047 3.4272e-006 0.001154 0.06467 0.00065439 0.06532 0.058344 0 0.043374 0.0389 0 0.84926 0.22873 0.059417 0.0084146 4.1077 0.052912 6.313e-005 0.83715 0.0051067 0.0058446 0.001632 0.98366 0.98793 3.5548e-006 1.422e-005 0.13047 0.7257 0.77733 0.0015221 0.79109 0.50041 0.0020457 0.42213 1.2957 1.2917 16.0056 144.9825 0.00038817 -84.6726 0.15696
0.261 0.98802 5.524e-005 3.8182 0.012047 3.4404e-006 0.001154 0.064807 0.0006544 0.065457 0.058469 0 0.043362 0.0389 0 0.84928 0.22875 0.059421 0.0084152 4.1077 0.052915 6.3133e-005 0.83715 0.0051067 0.0058446 0.00163 0.98369 0.98805 3.5502e-006 1.4201e-005 0.13047 0.7265 0.77799 0.0015211 0.7923 0.50057 0.0020444 0.42213 1.2976 1.2936 16.0056 144.9825 0.00038711 -84.6799 0.15796
0.262 0.98802 5.524e-005 3.8182 0.012047 3.4536e-006 0.001154 0.064944 0.00065442 0.065594 0.058594 0 0.04335 0.0389 0 0.84931 0.22876 0.059426 0.0084157 4.1078 0.052918 6.3137e-005 0.83715 0.0051068 0.0058447 0.0016281 0.98372 0.98815 3.5457e-006 1.4183e-005 0.13047 0.7273 0.77864 0.0015201 0.79351 0.50074 0.0020431 0.42214 1.2995 1.2955 16.0057 144.9825 0.00038605 -84.6871 0.15896
0.263 0.98802 5.524e-005 3.8182 0.012047 3.4667e-006 0.001154 0.065081 0.00065443 0.065731 0.058719 0 0.043338 0.0389 0 0.84934 0.22877 0.05943 0.0084163 4.1078 0.052921 6.314e-005 0.83714 0.0051068 0.0058447 0.0016262 0.98374 0.98826 3.5412e-006 1.4165e-005 0.13047 0.7281 0.7793 0.0015192 0.79471 0.50091 0.0020419 0.42214 1.3013 1.2974 16.0057 144.9825 0.000385 -84.6943 0.15996
0.264 0.98802 5.524e-005 3.8182 0.012047 3.4799e-006 0.001154 0.065218 0.00065445 0.065868 0.058844 0 0.043326 0.0389 0 0.84937 0.22879 0.059435 0.0084169 4.1078 0.052924 6.3144e-005 0.83714 0.0051068 0.0058447 0.0016242 0.98377 0.98835 3.5367e-006 1.4147e-005 0.13047 0.72889 0.77994 0.0015182 0.7959 0.50108 0.0020407 0.42214 1.3032 1.2992 16.0058 144.9825 0.00038396 -84.7014 0.16096
0.265 0.98802 5.524e-005 3.8182 0.012047 3.4931e-006 0.001154 0.065354 0.00065446 0.066004 0.058969 0 0.043314 0.0389 0 0.8494 0.2288 0.05944 0.0084175 4.1079 0.052926 6.3148e-005 0.83714 0.0051069 0.0058448 0.0016223 0.9838 0.98845 3.5323e-006 1.413e-005 0.13047 0.72968 0.78059 0.0015173 0.79708 0.50125 0.0020394 0.42215 1.305 1.3011 16.0058 144.9826 0.00038291 -84.7085 0.16196
0.266 0.98802 5.524e-005 3.8182 0.012046 3.5063e-006 0.001154 0.065491 0.00065448 0.066141 0.059093 0 0.043303 0.0389 0 0.84943 0.22881 0.059444 0.0084181 4.1079 0.052929 6.3151e-005 0.83713 0.0051069 0.0058448 0.0016204 0.98382 0.98853 3.5279e-006 1.4112e-005 0.13047 0.73047 0.78123 0.0015164 0.79826 0.50142 0.0020382 0.42215 1.3069 1.303 16.0059 144.9826 0.00038188 -84.7155 0.16296
0.267 0.98802 5.524e-005 3.8182 0.012046 3.5194e-006 0.001154 0.065627 0.00065449 0.066277 0.059218 0 0.043291 0.0389 0 0.84946 0.22882 0.059449 0.0084187 4.1079 0.052932 6.3155e-005 0.83713 0.005107 0.0058449 0.0016185 0.98385 0.98862 3.5236e-006 1.4095e-005 0.13047 0.73125 0.78187 0.0015155 0.79944 0.50158 0.002037 0.42216 1.3087 1.3048 16.0059 144.9826 0.00038085 -84.7224 0.16396
0.268 0.98802 5.524e-005 3.8182 0.012046 3.5326e-006 0.001154 0.065763 0.00065451 0.066413 0.059343 0 0.043279 0.0389 0 0.84949 0.22884 0.059453 0.0084192 4.1079 0.052935 6.3159e-005 0.83713 0.005107 0.0058449 0.0016167 0.98387 0.9887 3.5193e-006 1.4078e-005 0.13047 0.73203 0.7825 0.0015145 0.8006 0.50175 0.0020358 0.42217 1.3106 1.3067 16.006 144.9826 0.00037982 -84.7293 0.16496
0.269 0.98802 5.524e-005 3.8182 0.012046 3.5458e-006 0.001154 0.065899 0.00065452 0.066549 0.059467 0 0.043268 0.0389 0 0.84952 0.22885 0.059458 0.0084198 4.108 0.052938 6.3162e-005 0.83713 0.005107 0.0058449 0.0016148 0.9839 0.98877 3.515e-006 1.4061e-005 0.13047 0.73281 0.78314 0.0015136 0.80177 0.50192 0.0020346 0.42217 1.3124 1.3085 16.006 144.9826 0.0003788 -84.7362 0.16596
0.27 0.98802 5.5239e-005 3.8182 0.012046 3.559e-006 0.001154 0.066035 0.00065454 0.066685 0.059591 0 0.043256 0.0389 0 0.84955 0.22886 0.059463 0.0084204 4.108 0.052941 6.3166e-005 0.83712 0.0051071 0.005845 0.001613 0.98392 0.98884 3.5108e-006 1.4044e-005 0.13047 0.73359 0.78376 0.0015127 0.80292 0.50209 0.0020334 0.42218 1.3142 1.3104 16.0061 144.9826 0.00037779 -84.743 0.16696
0.271 0.98802 5.5239e-005 3.8182 0.012046 3.5721e-006 0.001154 0.066171 0.00065455 0.066821 0.059716 0 0.043244 0.0389 0 0.84958 0.22888 0.059468 0.008421 4.108 0.052944 6.317e-005 0.83712 0.0051071 0.005845 0.0016112 0.98395 0.98891 3.5066e-006 1.4027e-005 0.13047 0.73437 0.78439 0.0015118 0.80407 0.50226 0.0020323 0.42218 1.3161 1.3122 16.0061 144.9826 0.00037678 -84.7497 0.16796
0.272 0.98802 5.5239e-005 3.8182 0.012046 3.5853e-006 0.001154 0.066307 0.00065456 0.066957 0.05984 0 0.043232 0.0389 0 0.84961 0.22889 0.059472 0.0084216 4.1081 0.052947 6.3173e-005 0.83712 0.0051072 0.0058451 0.0016094 0.98397 0.98898 3.5025e-006 1.401e-005 0.13047 0.73514 0.78501 0.001511 0.80521 0.50243 0.0020311 0.42219 1.3179 1.314 16.0062 144.9826 0.00037577 -84.7564 0.16896
0.273 0.98802 5.5239e-005 3.8182 0.012046 3.5985e-006 0.001154 0.066443 0.00065458 0.067093 0.059964 0 0.043221 0.0389 0 0.84964 0.2289 0.059477 0.0084222 4.1081 0.05295 6.3177e-005 0.83711 0.0051072 0.0058451 0.0016077 0.984 0.98904 3.4984e-006 1.3994e-005 0.13047 0.73591 0.78563 0.0015101 0.80635 0.50259 0.00203 0.42219 1.3197 1.3159 16.0062 144.9827 0.00037478 -84.7631 0.16996
0.274 0.98802 5.5239e-005 3.8182 0.012046 3.6117e-006 0.001154 0.066578 0.00065459 0.067228 0.060088 0 0.043209 0.0389 0 0.84967 0.22891 0.059482 0.0084228 4.1081 0.052953 6.3181e-005 0.83711 0.0051072 0.0058451 0.001606 0.98402 0.9891 3.4943e-006 1.3977e-005 0.13047 0.73668 0.78624 0.0015092 0.80748 0.50276 0.0020288 0.4222 1.3215 1.3177 16.0063 144.9827 0.00037378 -84.7697 0.17096
0.275 0.98802 5.5239e-005 3.8182 0.012046 3.6248e-006 0.001154 0.066714 0.00065461 0.067364 0.060212 0 0.043198 0.0389 0 0.8497 0.22893 0.059486 0.0084234 4.1082 0.052956 6.3185e-005 0.83711 0.0051073 0.0058452 0.0016042 0.98405 0.98915 3.4903e-006 1.3961e-005 0.13047 0.73744 0.78685 0.0015083 0.80861 0.50293 0.0020277 0.4222 1.3233 1.3195 16.0063 144.9827 0.00037279 -84.7762 0.17196
0.276 0.98802 5.5239e-005 3.8182 0.012046 3.638e-006 0.001154 0.066849 0.00065462 0.067499 0.060335 0 0.043186 0.0389 0 0.84973 0.22894 0.059491 0.008424 4.1082 0.052959 6.3188e-005 0.8371 0.0051073 0.0058452 0.0016024 0.98407 0.98921 3.4862e-006 1.3945e-005 0.13047 0.73821 0.78746 0.0015075 0.80973 0.5031 0.0020266 0.42221 1.3251 1.3213 16.0064 144.9827 0.00037181 -84.7827 0.17296
0.277 0.98802 5.5239e-005 3.8182 0.012046 3.6512e-006 0.001154 0.066985 0.00065463 0.067635 0.060459 0 0.043174 0.0389 0 0.84976 0.22895 0.059496 0.0084246 4.1082 0.052962 6.3192e-005 0.8371 0.0051074 0.0058453 0.0016006 0.98409 0.98926 3.4822e-006 1.3929e-005 0.13048 0.73897 0.78807 0.0015066 0.81084 0.50327 0.0020255 0.42222 1.3269 1.3232 16.0064 144.9827 0.00037083 -84.7892 0.17396
0.278 0.98802 5.5239e-005 3.8182 0.012046 3.6644e-006 0.001154 0.06712 0.00065465 0.06777 0.060582 0 0.043163 0.0389 0 0.84979 0.22897 0.059501 0.0084252 4.1083 0.052965 6.3196e-005 0.8371 0.0051074 0.0058453 0.0015988 0.98412 0.98931 3.4782e-006 1.3914e-005 0.13048 0.73973 0.78867 0.0015058 0.81195 0.50343 0.0020244 0.42222 1.3287 1.325 16.0064 144.9827 0.00036985 -84.7956 0.17496
0.279 0.98802 5.5239e-005 3.8182 0.012046 3.6775e-006 0.001154 0.067255 0.00065466 0.067905 0.060706 0 0.043151 0.0389 0 0.84982 0.22898 0.059506 0.0084258 4.1083 0.052968 6.32e-005 0.8371 0.0051075 0.0058453 0.001597 0.98414 0.98935 3.4743e-006 1.3898e-005 0.13048 0.74049 0.78927 0.0015049 0.81305 0.5036 0.0020233 0.42223 1.3305 1.3268 16.0065 144.9827 0.00036888 -84.8019 0.17596
0.28 0.98802 5.5239e-005 3.8182 0.012046 3.6907e-006 0.001154 0.06739 0.00065468 0.06804 0.060829 0 0.04314 0.0389 0 0.84985 0.22899 0.05951 0.0084264 4.1083 0.052971 6.3204e-005 0.83709 0.0051075 0.0058454 0.0015953 0.98416 0.9894 3.4704e-006 1.3882e-005 0.13048 0.74124 0.78986 0.0015041 0.81415 0.50377 0.0020222 0.42223 1.3323 1.3286 16.0065 144.9828 0.00036792 -84.8082 0.17696
0.281 0.98802 5.5239e-005 3.8182 0.012046 3.7039e-006 0.001154 0.067525 0.00065469 0.068175 0.060953 0 0.043128 0.0389 0 0.84988 0.22901 0.059515 0.008427 4.1084 0.052974 6.3208e-005 0.83709 0.0051075 0.0058454 0.0015936 0.98419 0.98944 3.4666e-006 1.3867e-005 0.13048 0.74199 0.79045 0.0015033 0.81524 0.50394 0.0020211 0.42224 1.3341 1.3304 16.0066 144.9828 0.00036696 -84.8144 0.17796
0.282 0.98802 5.5239e-005 3.8182 0.012046 3.7171e-006 0.001154 0.067659 0.0006547 0.068309 0.061076 0 0.043117 0.0389 0 0.84991 0.22902 0.05952 0.0084277 4.1084 0.052977 6.3211e-005 0.83709 0.0051076 0.0058455 0.001592 0.98421 0.98948 3.4628e-006 1.3852e-005 0.13048 0.74274 0.79104 0.0015025 0.81632 0.50411 0.0020201 0.42225 1.3359 1.3322 16.0066 144.9828 0.000366 -84.8206 0.17896
0.283 0.98802 5.5239e-005 3.8182 0.012046 3.7302e-006 0.001154 0.067794 0.00065472 0.068444 0.061199 0 0.043105 0.0389 0 0.84994 0.22904 0.059525 0.0084283 4.1084 0.05298 6.3215e-005 0.83708 0.0051076 0.0058455 0.0015905 0.98423 0.98952 3.4591e-006 1.3837e-005 0.13048 0.74349 0.79163 0.0015017 0.8174 0.50427 0.002019 0.42225 1.3377 1.334 16.0067 144.9828 0.00036505 -84.8268 0.17996
0.284 0.98802 5.5239e-005 3.8182 0.012046 3.7434e-006 0.001154 0.067928 0.00065473 0.068579 0.061322 0 0.043094 0.0389 0 0.84997 0.22905 0.05953 0.0084289 4.1085 0.052983 6.3219e-005 0.83708 0.0051077 0.0058456 0.001589 0.98425 0.98956 3.4554e-006 1.3822e-005 0.13048 0.74423 0.79221 0.0015009 0.81847 0.50444 0.002018 0.42226 1.3394 1.3358 16.0067 144.9828 0.00036411 -84.8329 0.18096
0.285 0.98802 5.5239e-005 3.8182 0.012046 3.7566e-006 0.001154 0.068063 0.00065474 0.068713 0.061445 0 0.043082 0.0389 0 0.85 0.22906 0.059535 0.0084295 4.1085 0.052986 6.3223e-005 0.83708 0.0051077 0.0058456 0.0015874 0.98427 0.9896 3.4517e-006 1.3807e-005 0.13048 0.74498 0.79279 0.0015001 0.81954 0.50461 0.0020169 0.42226 1.3412 1.3375 16.0068 144.9828 0.00036317 -84.8389 0.18196
0.286 0.98802 5.5239e-005 3.8182 0.012046 3.7698e-006 0.001154 0.068197 0.00065476 0.068847 0.061568 0 0.043071 0.0389 0 0.85003 0.22908 0.05954 0.0084301 4.1085 0.052989 6.3227e-005 0.83707 0.0051078 0.0058456 0.0015859 0.9843 0.98963 3.448e-006 1.3792e-005 0.13048 0.74572 0.79337 0.0014993 0.8206 0.50478 0.0020159 0.42227 1.343 1.3393 16.0068 144.9828 0.00036223 -84.845 0.18296
0.287 0.98802 5.5238e-005 3.8182 0.012046 3.7829e-006 0.001154 0.068331 0.00065477 0.068981 0.06169 0 0.043059 0.0389 0 0.85006 0.22909 0.059545 0.0084307 4.1086 0.052992 6.3231e-005 0.83707 0.0051078 0.0058457 0.0015844 0.98432 0.98966 3.4444e-006 1.3778e-005 0.13048 0.74646 0.79394 0.0014985 0.82166 0.50495 0.0020149 0.42228 1.3447 1.3411 16.0068 144.9829 0.0003613 -84.8509 0.18396
0.288 0.98802 5.5238e-005 3.8182 0.012046 3.7961e-006 0.001154 0.068465 0.00065478 0.069116 0.061813 0 0.043048 0.0389 0 0.85009 0.2291 0.05955 0.0084314 4.1086 0.052995 6.3235e-005 0.83707 0.0051079 0.0058457 0.0015829 0.98434 0.9897 3.4408e-006 1.3763e-005 0.13048 0.74719 0.79451 0.0014977 0.82271 0.50511 0.0020138 0.42228 1.3465 1.3429 16.0069 144.9829 0.00036037 -84.8568 0.18496
0.289 0.98802 5.5238e-005 3.8182 0.012046 3.8093e-006 0.001154 0.068599 0.00065479 0.069249 0.061936 0 0.043036 0.0389 0 0.85013 0.22912 0.059555 0.008432 4.1086 0.052998 6.3239e-005 0.83706 0.0051079 0.0058458 0.0015814 0.98436 0.98973 3.4373e-006 1.3749e-005 0.13048 0.74793 0.79508 0.001497 0.82375 0.50528 0.0020128 0.42229 1.3482 1.3446 16.0069 144.9829 0.00035945 -84.8627 0.18596
0.29 0.98802 5.5238e-005 3.8182 0.012046 3.8225e-006 0.001154 0.068733 0.00065481 0.069383 0.062058 0 0.043025 0.0389 0 0.85016 0.22913 0.05956 0.0084326 4.1087 0.053002 6.3243e-005 0.83706 0.0051079 0.0058458 0.0015799 0.98438 0.98976 3.4337e-006 1.3735e-005 0.13048 0.74866 0.79565 0.0014962 0.82479 0.50545 0.0020118 0.4223 1.35 1.3464 16.007 144.9829 0.00035853 -84.8685 0.18696
0.291 0.98802 5.5238e-005 3.8182 0.012046 3.8356e-006 0.001154 0.068867 0.00065482 0.069517 0.06218 0 0.043014 0.0389 0 0.85019 0.22914 0.059564 0.0084332 4.1087 0.053005 6.3247e-005 0.83706 0.005108 0.0058459 0.0015783 0.9844 0.98979 3.4302e-006 1.3721e-005 0.13048 0.74939 0.79621 0.0014954 0.82583 0.50562 0.0020108 0.4223 1.3517 1.3481 16.007 144.9829 0.00035762 -84.8743 0.18796
0.292 0.98802 5.5238e-005 3.8182 0.012046 3.8488e-006 0.001154 0.069001 0.00065483 0.069651 0.062303 0 0.043002 0.0389 0 0.85022 0.22916 0.059569 0.0084339 4.1087 0.053008 6.3251e-005 0.83706 0.005108 0.0058459 0.0015768 0.98442 0.98981 3.4267e-006 1.3707e-005 0.13048 0.75011 0.79677 0.0014947 0.82685 0.50578 0.0020099 0.42231 1.3535 1.3499 16.0071 144.9829 0.00035671 -84.8801 0.18896
0.293 0.98802 5.5238e-005 3.8182 0.012046 3.862e-006 0.001154 0.069134 0.00065485 0.069784 0.062425 0 0.042991 0.0389 0 0.85025 0.22917 0.059574 0.0084345 4.1088 0.053011 6.3255e-005 0.83705 0.0051081 0.005846 0.0015752 0.98444 0.98984 3.4232e-006 1.3693e-005 0.13048 0.75084 0.79732 0.001494 0.82788 0.50595 0.0020089 0.42232 1.3552 1.3516 16.0071 144.9829 0.0003558 -84.8858 0.18996
0.294 0.98802 5.5238e-005 3.8182 0.012046 3.8752e-006 0.001154 0.069268 0.00065486 0.069918 0.062547 0 0.042979 0.0389 0 0.85028 0.22919 0.05958 0.0084351 4.1088 0.053014 6.3259e-005 0.83705 0.0051081 0.005846 0.0015737 0.98446 0.98987 3.4198e-006 1.3679e-005 0.13048 0.75156 0.79788 0.0014932 0.82889 0.50612 0.0020079 0.42233 1.3569 1.3534 16.0071 144.983 0.0003549 -84.8914 0.19096
0.295 0.98802 5.5238e-005 3.8182 0.012046 3.8883e-006 0.001154 0.069401 0.00065487 0.070051 0.062669 0 0.042968 0.0389 0 0.85031 0.2292 0.059585 0.0084358 4.1088 0.053018 6.3263e-005 0.83705 0.0051082 0.005846 0.0015722 0.98448 0.98989 3.4164e-006 1.3666e-005 0.13048 0.75228 0.79843 0.0014925 0.8299 0.50629 0.002007 0.42233 1.3587 1.3551 16.0072 144.983 0.00035401 -84.897 0.19196
0.296 0.98802 5.5238e-005 3.8182 0.012046 3.9015e-006 0.001154 0.069534 0.00065488 0.070184 0.062791 0 0.042957 0.0389 0 0.85035 0.22921 0.05959 0.0084364 4.1089 0.053021 6.3267e-005 0.83704 0.0051082 0.0058461 0.0015707 0.9845 0.98992 3.413e-006 1.3652e-005 0.13048 0.753 0.79898 0.0014917 0.83091 0.50645 0.002006 0.42234 1.3604 1.3568 16.0072 144.983 0.00035312 -84.9026 0.19296
0.297 0.98802 5.5238e-005 3.8182 0.012046 3.9147e-006 0.001154 0.069667 0.0006549 0.070317 0.062913 0 0.042945 0.0389 0 0.85038 0.22923 0.059595 0.0084371 4.1089 0.053024 6.3271e-005 0.83704 0.0051083 0.0058461 0.0015692 0.98452 0.98994 3.4097e-006 1.3639e-005 0.13048 0.75372 0.79952 0.001491 0.83191 0.50662 0.0020051 0.42235 1.3621 1.3586 16.0073 144.983 0.00035223 -84.9081 0.19396
0.298 0.98802 5.5238e-005 3.8182 0.012046 3.9279e-006 0.001154 0.0698 0.00065491 0.07045 0.063034 0 0.042934 0.0389 0 0.85041 0.22924 0.0596 0.0084377 4.109 0.053027 6.3276e-005 0.83704 0.0051083 0.0058462 0.0015678 0.98454 0.98996 3.4064e-006 1.3626e-005 0.13048 0.75443 0.80006 0.0014903 0.8329 0.50679 0.0020041 0.42235 1.3638 1.3603 16.0073 144.983 0.00035135 -84.9136 0.19496
0.299 0.98802 5.5238e-005 3.8182 0.012046 3.941e-006 0.001154 0.069933 0.00065492 0.070583 0.063156 0 0.042923 0.0389 0 0.85044 0.22926 0.059605 0.0084383 4.109 0.05303 6.328e-005 0.83703 0.0051084 0.0058462 0.0015664 0.98456 0.98998 3.4031e-006 1.3613e-005 0.13048 0.75514 0.8006 0.0014896 0.83389 0.50696 0.0020032 0.42236 1.3655 1.362 16.0073 144.983 0.00035047 -84.9191 0.19596
0.3 0.98802 5.5238e-005 3.8182 0.012046 3.9542e-006 0.001154 0.070066 0.00065493 0.070716 0.063277 0 0.042912 0.0389 0 0.85047 0.22927 0.05961 0.008439 4.109 0.053034 6.3284e-005 0.83703 0.0051084 0.0058463 0.0015649 0.98458 0.99001 3.3998e-006 1.36e-005 0.13048 0.75585 0.80114 0.0014889 0.83488 0.50712 0.0020023 0.42237 1.3672 1.3637 16.0074 144.983 0.0003496 -84.9245 0.19696
0.301 0.98802 5.5238e-005 3.8182 0.012046 3.9674e-006 0.001154 0.070199 0.00065495 0.070849 0.063399 0 0.0429 0.0389 0 0.85051 0.22929 0.059615 0.0084396 4.1091 0.053037 6.3288e-005 0.83703 0.0051085 0.0058463 0.0015636 0.9846 0.99003 3.3966e-006 1.3587e-005 0.13048 0.75656 0.80168 0.0014882 0.83586 0.50729 0.0020014 0.42238 1.3689 1.3655 16.0074 144.9831 0.00034873 -84.9298 0.19796
0.302 0.98802 5.5238e-005 3.8182 0.012046 3.9805e-006 0.001154 0.070331 0.00065496 0.070981 0.06352 0 0.042889 0.0389 0 0.85054 0.2293 0.05962 0.0084403 4.1091 0.05304 6.3292e-005 0.83702 0.0051085 0.0058464 0.0015622 0.98462 0.99005 3.3934e-006 1.3574e-005 0.13048 0.75726 0.80221 0.0014875 0.83683 0.50746 0.0020005 0.42238 1.3706 1.3672 16.0074 144.9831 0.00034786 -84.9351 0.19896
0.303 0.98802 5.5237e-005 3.8182 0.012046 3.9937e-006 0.001154 0.070464 0.00065497 0.071114 0.063642 0 0.042878 0.0389 0 0.85057 0.22931 0.059625 0.0084409 4.1091 0.053044 6.3296e-005 0.83702 0.0051086 0.0058464 0.0015609 0.98464 0.99007 3.3903e-006 1.3561e-005 0.13049 0.75796 0.80274 0.0014868 0.8378 0.50763 0.0019996 0.42239 1.3723 1.3689 16.0075 144.9831 0.000347 -84.9404 0.19996
0.304 0.98802 5.5237e-005 3.8182 0.012046 4.0069e-006 0.001154 0.070596 0.00065498 0.071246 0.063763 0 0.042867 0.0389 0 0.8506 0.22933 0.05963 0.0084416 4.1092 0.053047 6.3301e-005 0.83702 0.0051086 0.0058465 0.0015595 0.98465 0.99008 3.3871e-006 1.3549e-005 0.13049 0.75867 0.80326 0.0014861 0.83876 0.50779 0.0019987 0.4224 1.374 1.3706 16.0075 144.9831 0.00034614 -84.9457 0.20096
0.305 0.98802 5.5237e-005 3.8182 0.012046 4.0201e-006 0.001154 0.070728 0.00065499 0.071379 0.063884 0 0.042856 0.0389 0 0.85064 0.22934 0.059636 0.0084422 4.1092 0.05305 6.3305e-005 0.83701 0.0051087 0.0058465 0.0015582 0.98467 0.9901 3.384e-006 1.3536e-005 0.13049 0.75936 0.80379 0.0014855 0.83972 0.50796 0.0019978 0.42241 1.3757 1.3723 16.0076 144.9831 0.00034529 -84.9509 0.20196
0.306 0.98802 5.5237e-005 3.8182 0.012046 4.0332e-006 0.001154 0.07086 0.00065501 0.071511 0.064005 0 0.042844 0.0389 0 0.85067 0.22936 0.059641 0.0084429 4.1093 0.053054 6.3309e-005 0.83701 0.0051087 0.0058466 0.0015569 0.98469 0.99012 3.3809e-006 1.3524e-005 0.13049 0.76006 0.80431 0.0014848 0.84067 0.50813 0.0019969 0.42241 1.3774 1.374 16.0076 144.9831 0.00034444 -84.956 0.20296
0.307 0.98802 5.5237e-005 3.8182 0.012046 4.0464e-006 0.001154 0.070992 0.00065502 0.071643 0.064126 0 0.042833 0.0389 0 0.8507 0.22937 0.059646 0.0084435 4.1093 0.053057 6.3313e-005 0.83701 0.0051088 0.0058466 0.0015555 0.98471 0.99014 3.3779e-006 1.3512e-005 0.13049 0.76075 0.80483 0.0014841 0.84162 0.5083 0.0019961 0.42242 1.379 1.3757 16.0076 144.9831 0.0003436 -84.9611 0.20396
0.308 0.98802 5.5237e-005 3.8182 0.012046 4.0596e-006 0.001154 0.071124 0.00065503 0.071775 0.064246 0 0.042822 0.0389 0 0.85074 0.22939 0.059651 0.0084442 4.1093 0.05306 6.3318e-005 0.837 0.0051088 0.0058467 0.0015542 0.98473 0.99016 3.3748e-006 1.35e-005 0.13049 0.76145 0.80534 0.0014835 0.84256 0.50846 0.0019952 0.42243 1.3807 1.3773 16.0077 144.9832 0.00034276 -84.9662 0.20496
0.309 0.98802 5.5237e-005 3.8182 0.012046 4.0728e-006 0.001154 0.071256 0.00065504 0.071907 0.064367 0 0.042811 0.0389 0 0.85077 0.2294 0.059657 0.0084449 4.1094 0.053064 6.3322e-005 0.837 0.0051089 0.0058467 0.0015529 0.98474 0.99017 3.3718e-006 1.3487e-005 0.13049 0.76214 0.80585 0.0014828 0.84349 0.50863 0.0019943 0.42244 1.3824 1.379 16.0077 144.9832 0.00034192 -84.9713 0.20596
0.31 0.98802 5.5237e-005 3.8182 0.012046 4.0859e-006 0.001154 0.071388 0.00065505 0.072038 0.064488 0 0.0428 0.0389 0 0.8508 0.22941 0.059662 0.0084455 4.1094 0.053067 6.3326e-005 0.837 0.0051089 0.0058468 0.0015516 0.98476 0.99019 3.3688e-006 1.3476e-005 0.13049 0.76282 0.80637 0.0014822 0.84443 0.5088 0.0019935 0.42244 1.3841 1.3807 16.0077 144.9832 0.00034109 -84.9763 0.20696
0.311 0.98802 5.5237e-005 3.8182 0.012046 4.0991e-006 0.001154 0.07152 0.00065506 0.07217 0.064608 0 0.042789 0.0389 0 0.85083 0.22943 0.059667 0.0084462 4.1095 0.053071 6.3331e-005 0.83699 0.005109 0.0058468 0.0015503 0.98478 0.9902 3.3658e-006 1.3464e-005 0.13049 0.76351 0.80687 0.0014815 0.84535 0.50897 0.0019926 0.42245 1.3857 1.3824 16.0078 144.9832 0.00034026 -84.9813 0.20796
0.312 0.98802 5.5237e-005 3.8182 0.012046 4.1123e-006 0.001154 0.071651 0.00065508 0.072302 0.064729 0 0.042778 0.0389 0 0.85087 0.22944 0.059672 0.0084468 4.1095 0.053074 6.3335e-005 0.83699 0.005109 0.0058469 0.001549 0.9848 0.99022 3.3629e-006 1.3452e-005 0.13049 0.76419 0.80738 0.0014809 0.84627 0.50913 0.0019918 0.42246 1.3874 1.384 16.0078 144.9832 0.00033944 -84.9862 0.20896
0.313 0.98802 5.5237e-005 3.8182 0.012046 4.1255e-006 0.001154 0.071782 0.00065509 0.072433 0.064849 0 0.042767 0.0389 0 0.8509 0.22946 0.059678 0.0084475 4.1095 0.053077 6.3339e-005 0.83699 0.0051091 0.0058469 0.0015477 0.98481 0.99024 3.36e-006 1.344e-005 0.13049 0.76488 0.80788 0.0014802 0.84719 0.5093 0.001991 0.42247 1.389 1.3857 16.0078 144.9832 0.00033862 -84.9911 0.20996
0.314 0.98802 5.5237e-005 3.8182 0.012046 4.1386e-006 0.001154 0.071914 0.0006551 0.072564 0.064969 0 0.042756 0.0389 0 0.85093 0.22947 0.059683 0.0084482 4.1096 0.053081 6.3344e-005 0.83698 0.0051091 0.005847 0.0015465 0.98483 0.99025 3.3571e-006 1.3429e-005 0.13049 0.76555 0.80838 0.0014796 0.8481 0.50947 0.0019902 0.42248 1.3907 1.3874 16.0079 144.9833 0.00033781 -84.9959 0.21096
0.315 0.98802 5.5237e-005 3.8182 0.012046 4.1518e-006 0.001154 0.072045 0.00065511 0.072695 0.065089 0 0.042744 0.0389 0 0.85097 0.22949 0.059688 0.0084488 4.1096 0.053084 6.3348e-005 0.83698 0.0051092 0.005847 0.0015452 0.98485 0.99026 3.3542e-006 1.3417e-005 0.13049 0.76623 0.80888 0.001479 0.849 0.50963 0.0019893 0.42248 1.3923 1.389 16.0079 144.9833 0.00033699 -85.0008 0.21196
0.316 0.98802 5.5237e-005 3.8182 0.012046 4.165e-006 0.001154 0.072176 0.00065512 0.072827 0.06521 0 0.042733 0.0389 0 0.851 0.2295 0.059693 0.0084495 4.1097 0.053088 6.3352e-005 0.83698 0.0051092 0.0058471 0.001544 0.98486 0.99028 3.3514e-006 1.3406e-005 0.13049 0.76691 0.80938 0.0014784 0.84991 0.5098 0.0019885 0.42249 1.3939 1.3907 16.0079 144.9833 0.00033619 -85.0055 0.21296
0.317 0.98802 5.5237e-005 3.8182 0.012046 4.1782e-006 0.001154 0.072307 0.00065513 0.072958 0.065329 0 0.042722 0.0389 0 0.85104 0.22952 0.059699 0.0084502 4.1097 0.053091 6.3357e-005 0.83697 0.0051093 0.0058471 0.0015428 0.98488 0.99029 3.3486e-006 1.3395e-005 0.13049 0.76758 0.80987 0.0014778 0.8508 0.50997 0.0019877 0.4225 1.3956 1.3923 16.008 144.9833 0.00033538 -85.0103 0.21396
0.318 0.98802 5.5237e-005 3.8182 0.012046 4.1913e-006 0.001154 0.072438 0.00065514 0.073088 0.065449 0 0.042711 0.0389 0 0.85107 0.22953 0.059704 0.0084509 4.1097 0.053095 6.3361e-005 0.83697 0.0051093 0.0058472 0.0015416 0.9849 0.99031 3.3458e-006 1.3383e-005 0.13049 0.76825 0.81036 0.0014771 0.85169 0.51014 0.0019869 0.42251 1.3972 1.3939 16.008 144.9833 0.00033458 -85.015 0.21496
0.319 0.98802 5.5236e-005 3.8182 0.012046 4.2045e-006 0.001154 0.072569 0.00065516 0.073219 0.065569 0 0.0427 0.0389 0 0.8511 0.22955 0.05971 0.0084515 4.1098 0.053098 6.3366e-005 0.83697 0.0051094 0.0058472 0.0015404 0.98491 0.99032 3.343e-006 1.3372e-005 0.13049 0.76892 0.81085 0.0014765 0.85258 0.5103 0.0019861 0.42252 1.3988 1.3956 16.008 144.9833 0.00033379 -85.0197 0.21596
0.32 0.98802 5.5236e-005 3.8182 0.012046 4.2177e-006 0.001154 0.072699 0.00065517 0.07335 0.065689 0 0.042689 0.0389 0 0.85114 0.22956 0.059715 0.0084522 4.1098 0.053102 6.337e-005 0.83696 0.0051094 0.0058473 0.0015392 0.98493 0.99033 3.3403e-006 1.3361e-005 0.13049 0.76959 0.81134 0.0014759 0.85346 0.51047 0.0019854 0.42253 1.4005 1.3972 16.0081 144.9833 0.00033299 -85.0243 0.21696
0.321 0.98802 5.5236e-005 3.8182 0.012046 4.2308e-006 0.001154 0.07283 0.00065518 0.073481 0.065808 0 0.042678 0.0389 0 0.85117 0.22958 0.05972 0.0084529 4.1099 0.053105 6.3375e-005 0.83696 0.0051095 0.0058473 0.001538 0.98494 0.99035 3.3376e-006 1.335e-005 0.13049 0.77025 0.81182 0.0014754 0.85433 0.51064 0.0019846 0.42253 1.4021 1.3988 16.0081 144.9834 0.0003322 -85.0289 0.21796
0.322 0.98802 5.5236e-005 3.8182 0.012046 4.244e-006 0.001154 0.07296 0.00065519 0.073611 0.065928 0 0.042668 0.0389 0 0.8512 0.22959 0.059726 0.0084536 4.1099 0.053109 6.3379e-005 0.83695 0.0051095 0.0058474 0.0015369 0.98496 0.99036 3.3349e-006 1.334e-005 0.13049 0.77091 0.8123 0.0014748 0.8552 0.5108 0.0019838 0.42254 1.4037 1.4005 16.0081 144.9834 0.00033142 -85.0335 0.21896
0.323 0.98802 5.5236e-005 3.8182 0.012046 4.2572e-006 0.001154 0.073091 0.0006552 0.073741 0.066047 0 0.042657 0.0389 0 0.85124 0.22961 0.059731 0.0084543 4.1099 0.053112 6.3383e-005 0.83695 0.0051096 0.0058474 0.0015357 0.98498 0.99037 3.3322e-006 1.3329e-005 0.13049 0.77158 0.81278 0.0014742 0.85607 0.51097 0.001983 0.42255 1.4053 1.4021 16.0082 144.9834 0.00033064 -85.038 0.21996
0.324 0.98802 5.5236e-005 3.8182 0.012046 4.2704e-006 0.001154 0.073221 0.00065521 0.073872 0.066167 0 0.042646 0.0389 0 0.85127 0.22962 0.059737 0.0084549 4.11 0.053116 6.3388e-005 0.83695 0.0051097 0.0058475 0.0015346 0.98499 0.99038 3.3295e-006 1.3318e-005 0.13049 0.77223 0.81326 0.0014736 0.85693 0.51114 0.0019823 0.42256 1.4069 1.4037 16.0082 144.9834 0.00032986 -85.0426 0.22096
0.325 0.98802 5.5236e-005 3.8182 0.012046 4.2835e-006 0.001154 0.073351 0.00065522 0.074002 0.066286 0 0.042635 0.0389 0 0.85131 0.22964 0.059742 0.0084556 4.11 0.053119 6.3393e-005 0.83694 0.0051097 0.0058476 0.0015334 0.98501 0.9904 3.3269e-006 1.3308e-005 0.13049 0.77289 0.81373 0.001473 0.85779 0.5113 0.0019815 0.42257 1.4085 1.4053 16.0082 144.9834 0.00032909 -85.047 0.22196
0.326 0.98802 5.5236e-005 3.8182 0.012046 4.2967e-006 0.001154 0.073481 0.00065523 0.074132 0.066405 0 0.042624 0.0389 0 0.85134 0.22965 0.059747 0.0084563 4.1101 0.053123 6.3397e-005 0.83694 0.0051098 0.0058476 0.0015323 0.98502 0.99041 3.3243e-006 1.3297e-005 0.1305 0.77355 0.8142 0.0014724 0.85864 0.51147 0.0019808 0.42258 1.4101 1.4069 16.0083 144.9834 0.00032832 -85.0515 0.22296
0.327 0.98802 5.5236e-005 3.8182 0.012046 4.3099e-006 0.001154 0.073611 0.00065524 0.074262 0.066524 0 0.042613 0.0389 0 0.85138 0.22967 0.059753 0.008457 4.1101 0.053127 6.3402e-005 0.83694 0.0051098 0.0058477 0.0015311 0.98504 0.99042 3.3217e-006 1.3287e-005 0.1305 0.7742 0.81467 0.0014719 0.85948 0.51164 0.00198 0.42259 1.4117 1.4085 16.0083 144.9835 0.00032755 -85.0559 0.22396
0.328 0.98802 5.5236e-005 3.8182 0.012046 4.3231e-006 0.001154 0.073741 0.00065525 0.074392 0.066643 0 0.042602 0.0389 0 0.85141 0.22968 0.059758 0.0084577 4.1102 0.05313 6.3406e-005 0.83693 0.0051099 0.0058477 0.00153 0.98505 0.99043 3.3191e-006 1.3277e-005 0.1305 0.77485 0.81514 0.0014713 0.86033 0.5118 0.0019793 0.42259 1.4133 1.4101 16.0083 144.9835 0.00032679 -85.0602 0.22496
0.329 0.98802 5.5236e-005 3.8182 0.012046 4.3362e-006 0.001154 0.073871 0.00065527 0.074521 0.066762 0 0.042591 0.0389 0 0.85145 0.2297 0.059764 0.0084584 4.1102 0.053134 6.3411e-005 0.83693 0.0051099 0.0058478 0.0015289 0.98507 0.99044 3.3166e-006 1.3267e-005 0.1305 0.7755 0.81561 0.0014708 0.86116 0.51197 0.0019786 0.4226 1.4149 1.4117 16.0084 144.9835 0.00032603 -85.0646 0.22596
0.33 0.98802 5.5236e-005 3.8182 0.012046 4.3494e-006 0.001154 0.074 0.00065528 0.074651 0.066881 0 0.04258 0.0389 0 0.85148 0.22971 0.059769 0.0084591 4.1103 0.053137 6.3415e-005 0.83693 0.00511 0.0058478 0.0015278 0.98508 0.99045 3.3141e-006 1.3256e-005 0.1305 0.77614 0.81607 0.0014702 0.862 0.51214 0.0019778 0.42261 1.4165 1.4133 16.0084 144.9835 0.00032528 -85.0689 0.22696
0.331 0.98802 5.5236e-005 3.8182 0.012046 4.3626e-006 0.001154 0.07413 0.00065529 0.074781 0.067 0 0.04257 0.0389 0 0.85152 0.22973 0.059775 0.0084598 4.1103 0.053141 6.342e-005 0.83692 0.00511 0.0058479 0.0015267 0.9851 0.99047 3.3115e-006 1.3246e-005 0.1305 0.77679 0.81653 0.0014697 0.86282 0.5123 0.0019771 0.42262 1.418 1.4149 16.0084 144.9835 0.00032452 -85.0732 0.22796
0.332 0.98802 5.5236e-005 3.8182 0.012046 4.3758e-006 0.001154 0.074259 0.0006553 0.07491 0.067118 0 0.042559 0.0389 0 0.85155 0.22974 0.05978 0.0084605 4.1103 0.053145 6.3425e-005 0.83692 0.0051101 0.0058479 0.0015257 0.98511 0.99048 3.3091e-006 1.3236e-005 0.1305 0.77743 0.81699 0.0014691 0.86365 0.51247 0.0019764 0.42263 1.4196 1.4165 16.0085 144.9835 0.00032378 -85.0774 0.22896
0.333 0.98802 5.5236e-005 3.8182 0.012046 4.3889e-006 0.001154 0.074389 0.00065531 0.075039 0.067237 0 0.042548 0.0389 0 0.85159 0.22976 0.059786 0.0084612 4.1104 0.053148 6.3429e-005 0.83692 0.0051102 0.005848 0.0015246 0.98513 0.99049 3.3066e-006 1.3227e-005 0.1305 0.77807 0.81745 0.0014686 0.86446 0.51264 0.0019757 0.42264 1.4212 1.4181 16.0085 144.9835 0.00032303 -85.0816 0.22996
0.334 0.98802 5.5236e-005 3.8182 0.012046 4.4021e-006 0.001154 0.074518 0.00065532 0.075169 0.067355 0 0.042537 0.0389 0 0.85162 0.22978 0.059792 0.0084619 4.1104 0.053152 6.3434e-005 0.83691 0.0051102 0.0058481 0.0015236 0.98514 0.9905 3.3041e-006 1.3217e-005 0.1305 0.77871 0.8179 0.001468 0.86528 0.5128 0.001975 0.42265 1.4227 1.4197 16.0085 144.9836 0.00032229 -85.0858 0.23096
0.335 0.98802 5.5235e-005 3.8182 0.012046 4.4153e-006 0.001154 0.074647 0.00065533 0.075298 0.067474 0 0.042526 0.0389 0 0.85166 0.22979 0.059797 0.0084626 4.1105 0.053156 6.3439e-005 0.83691 0.0051103 0.0058481 0.0015225 0.98515 0.99051 3.3017e-006 1.3207e-005 0.1305 0.77935 0.81836 0.0014675 0.86609 0.51297 0.0019743 0.42266 1.4243 1.4212 16.0085 144.9836 0.00032155 -85.0899 0.23196
0.336 0.98802 5.5235e-005 3.8182 0.012046 4.4284e-006 0.001154 0.074776 0.00065534 0.075427 0.067592 0 0.042516 0.0389 0 0.85169 0.22981 0.059803 0.0084633 4.1105 0.053159 6.3443e-005 0.8369 0.0051103 0.0058482 0.0015215 0.98517 0.99052 3.2993e-006 1.3197e-005 0.1305 0.77998 0.81881 0.001467 0.86689 0.51314 0.0019736 0.42267 1.4259 1.4228 16.0086 144.9836 0.00032082 -85.0941 0.23296
0.337 0.98802 5.5235e-005 3.8182 0.012046 4.4416e-006 0.001154 0.074905 0.00065535 0.075556 0.06771 0 0.042505 0.0389 0 0.85173 0.22982 0.059808 0.008464 4.1106 0.053163 6.3448e-005 0.8369 0.0051104 0.0058482 0.0015204 0.98518 0.99053 3.2969e-006 1.3188e-005 0.1305 0.78062 0.81925 0.0014664 0.86769 0.5133 0.0019729 0.42268 1.4274 1.4244 16.0086 144.9836 0.00032009 -85.0982 0.23396
0.338 0.98802 5.5235e-005 3.8182 0.012046 4.4548e-006 0.001154 0.075034 0.00065536 0.075685 0.067828 0 0.042494 0.0389 0 0.85176 0.22984 0.059814 0.0084647 4.1106 0.053167 6.3453e-005 0.8369 0.0051105 0.0058483 0.0015194 0.9852 0.99054 3.2946e-006 1.3178e-005 0.1305 0.78125 0.8197 0.0014659 0.86849 0.51347 0.0019722 0.42269 1.429 1.4259 16.0086 144.9836 0.00031936 -85.1022 0.23496
0.339 0.98802 5.5235e-005 3.8182 0.012046 4.468e-006 0.001154 0.075162 0.00065537 0.075813 0.067946 0 0.042484 0.0389 0 0.8518 0.22985 0.05982 0.0084654 4.1107 0.05317 6.3457e-005 0.83689 0.0051105 0.0058483 0.0015184 0.98521 0.99055 3.2922e-006 1.3169e-005 0.1305 0.78188 0.82014 0.0014654 0.86928 0.51363 0.0019716 0.42269 1.4305 1.4275 16.0087 144.9836 0.00031864 -85.1062 0.23596
0.34 0.98802 5.5235e-005 3.8182 0.012046 4.4811e-006 0.001154 0.075291 0.00065538 0.075942 0.068064 0 0.042473 0.0389 0 0.85183 0.22987 0.059825 0.0084661 4.1107 0.053174 6.3462e-005 0.83689 0.0051106 0.0058484 0.0015173 0.98522 0.99056 3.2899e-006 1.316e-005 0.1305 0.7825 0.82059 0.0014649 0.87006 0.5138 0.0019709 0.4227 1.4321 1.429 16.0087 144.9837 0.00031792 -85.1102 0.23696
0.341 0.98802 5.5235e-005 3.8182 0.012045 4.4943e-006 0.001154 0.07542 0.00065539 0.07607 0.068182 0 0.042462 0.0389 0 0.85187 0.22988 0.059831 0.0084668 4.1108 0.053178 6.3467e-005 0.83689 0.0051106 0.0058485 0.0015163 0.98524 0.99057 3.2876e-006 1.315e-005 0.1305 0.78313 0.82102 0.0014644 0.87084 0.51397 0.0019702 0.42271 1.4336 1.4306 16.0087 144.9837 0.0003172 -85.1142 0.23796
0.342 0.98802 5.5235e-005 3.8182 0.012045 4.5075e-006 0.001154 0.075548 0.0006554 0.076199 0.068299 0 0.042451 0.0389 0 0.8519 0.2299 0.059837 0.0084676 4.1108 0.053182 6.3472e-005 0.83688 0.0051107 0.0058485 0.0015153 0.98525 0.99058 3.2853e-006 1.3141e-005 0.1305 0.78375 0.82146 0.0014639 0.87162 0.51413 0.0019696 0.42272 1.4351 1.4321 16.0087 144.9837 0.00031649 -85.1181 0.23896
0.343 0.98802 5.5235e-005 3.8182 0.012045 4.5206e-006 0.001154 0.075676 0.00065541 0.076327 0.068417 0 0.042441 0.0389 0 0.85194 0.22992 0.059842 0.0084683 4.1108 0.053185 6.3476e-005 0.83688 0.0051108 0.0058486 0.0015143 0.98526 0.99059 3.283e-006 1.3132e-005 0.1305 0.78437 0.8219 0.0014634 0.87239 0.5143 0.0019689 0.42273 1.4367 1.4337 16.0088 144.9837 0.00031578 -85.1221 0.23996
0.344 0.98802 5.5235e-005 3.8182 0.012045 4.5338e-006 0.001154 0.075804 0.00065542 0.076455 0.068535 0 0.04243 0.0389 0 0.85198 0.22993 0.059848 0.008469 4.1109 0.053189 6.3481e-005 0.83687 0.0051108 0.0058486 0.0015134 0.98528 0.9906 3.2808e-006 1.3123e-005 0.1305 0.78499 0.82233 0.0014629 0.87316 0.51447 0.0019683 0.42274 1.4382 1.4352 16.0088 144.9837 0.00031507 -85.1259 0.24096
0.345 0.98802 5.5235e-005 3.8182 0.012045 4.547e-006 0.001154 0.075933 0.00065543 0.076583 0.068652 0 0.04242 0.0389 0 0.85201 0.22995 0.059854 0.0084697 4.1109 0.053193 6.3486e-005 0.83687 0.0051109 0.0058487 0.0015124 0.98529 0.9906 3.2785e-006 1.3114e-005 0.1305 0.78561 0.82276 0.0014624 0.87392 0.51463 0.0019676 0.42275 1.4397 1.4367 16.0088 144.9837 0.00031437 -85.1298 0.24196
0.346 0.98802 5.5235e-005 3.8182 0.012045 4.5602e-006 0.001154 0.076061 0.00065544 0.076711 0.068769 0 0.042409 0.0389 0 0.85205 0.22996 0.059859 0.0084704 4.111 0.053197 6.3491e-005 0.83687 0.0051109 0.0058488 0.0015114 0.9853 0.99061 3.2763e-006 1.3105e-005 0.1305 0.78622 0.82319 0.0014619 0.87468 0.5148 0.001967 0.42276 1.4412 1.4383 16.0088 144.9838 0.00031367 -85.1336 0.24296
0.347 0.98802 5.5235e-005 3.8182 0.012045 4.5733e-006 0.001154 0.076188 0.00065545 0.076839 0.068887 0 0.042398 0.0389 0 0.85208 0.22998 0.059865 0.0084711 4.111 0.053201 6.3496e-005 0.83686 0.005111 0.0058488 0.0015105 0.98531 0.99062 3.2741e-006 1.3097e-005 0.13051 0.78684 0.82362 0.0014614 0.87544 0.51496 0.0019664 0.42277 1.4427 1.4398 16.0089 144.9838 0.00031298 -85.1374 0.24396
0.348 0.98802 5.5235e-005 3.8182 0.012045 4.5865e-006 0.001154 0.076316 0.00065546 0.076967 0.069004 0 0.042388 0.0389 0 0.85212 0.23 0.059871 0.0084719 4.1111 0.053204 6.3501e-005 0.83686 0.0051111 0.0058489 0.0015095 0.98533 0.99063 3.2719e-006 1.3088e-005 0.13051 0.78745 0.82405 0.0014609 0.87619 0.51513 0.0019657 0.42278 1.4442 1.4413 16.0089 144.9838 0.00031228 -85.1412 0.24496
0.349 0.98802 5.5235e-005 3.8182 0.012045 4.5997e-006 0.001154 0.076444 0.00065547 0.077095 0.069121 0 0.042377 0.0389 0 0.85216 0.23001 0.059877 0.0084726 4.1111 0.053208 6.3505e-005 0.83686 0.0051111 0.0058489 0.0015086 0.98534 0.99064 3.2698e-006 1.3079e-005 0.13051 0.78806 0.82447 0.0014605 0.87694 0.5153 0.0019651 0.42279 1.4457 1.4428 16.0089 144.9838 0.00031159 -85.1449 0.24596
0.35 0.98802 5.5235e-005 3.8182 0.012045 4.6129e-006 0.001154 0.076571 0.00065548 0.077222 0.069238 0 0.042367 0.0389 0 0.85219 0.23003 0.059882 0.0084733 4.1112 0.053212 6.351e-005 0.83685 0.0051112 0.005849 0.0015077 0.98535 0.99065 3.2676e-006 1.3071e-005 0.13051 0.78867 0.82489 0.00146 0.87768 0.51546 0.0019645 0.4228 1.4472 1.4443 16.0089 144.9838 0.00031091 -85.1486 0.24696
0.351 0.98802 5.5235e-005 3.8182 0.012045 4.626e-006 0.001154 0.076699 0.00065549 0.07735 0.069355 0 0.042356 0.0389 0 0.85223 0.23004 0.059888 0.0084741 4.1112 0.053216 6.3515e-005 0.83685 0.0051113 0.0058491 0.0015067 0.98536 0.99066 3.2655e-006 1.3062e-005 0.13051 0.78927 0.82531 0.0014595 0.87842 0.51563 0.0019639 0.42281 1.4487 1.4458 16.009 144.9838 0.00031022 -85.1523 0.24796
0.352 0.98802 5.5234e-005 3.8182 0.012045 4.6392e-006 0.001154 0.076826 0.0006555 0.077477 0.069472 0 0.042345 0.0389 0 0.85227 0.23006 0.059894 0.0084748 4.1113 0.05322 6.352e-005 0.83684 0.0051113 0.0058491 0.0015058 0.98538 0.99067 3.2634e-006 1.3054e-005 0.13051 0.78988 0.82573 0.001459 0.87915 0.51579 0.0019633 0.42282 1.4502 1.4473 16.009 144.9839 0.00030954 -85.156 0.24896
0.353 0.98802 5.5234e-005 3.8182 0.012045 4.6524e-006 0.001154 0.076954 0.00065551 0.077604 0.069588 0 0.042335 0.0389 0 0.8523 0.23008 0.0599 0.0084755 4.1113 0.053224 6.3525e-005 0.83684 0.0051114 0.0058492 0.0015049 0.98539 0.99068 3.2613e-006 1.3045e-005 0.13051 0.79048 0.82614 0.0014586 0.87988 0.51596 0.0019626 0.42283 1.4517 1.4488 16.009 144.9839 0.00030886 -85.1596 0.24996
0.354 0.98802 5.5234e-005 3.8182 0.012045 4.6655e-006 0.001154 0.077081 0.00065552 0.077732 0.069705 0 0.042324 0.0389 0 0.85234 0.23009 0.059906 0.0084763 4.1114 0.053228 6.353e-005 0.83684 0.0051114 0.0058492 0.001504 0.9854 0.99068 3.2592e-006 1.3037e-005 0.13051 0.79108 0.82656 0.0014581 0.8806 0.51612 0.001962 0.42284 1.4532 1.4503 16.009 144.9839 0.00030819 -85.1632 0.25096
0.355 0.98802 5.5234e-005 3.8182 0.012045 4.6787e-006 0.001154 0.077208 0.00065553 0.077859 0.069822 0 0.042314 0.0389 0 0.85238 0.23011 0.059911 0.008477 4.1114 0.053232 6.3535e-005 0.83683 0.0051115 0.0058493 0.0015031 0.98541 0.99069 3.2571e-006 1.3029e-005 0.13051 0.79168 0.82697 0.0014577 0.88132 0.51629 0.0019614 0.42285 1.4547 1.4518 16.0091 144.9839 0.00030752 -85.1668 0.25196
0.356 0.98802 5.5234e-005 3.8182 0.012045 4.6919e-006 0.001154 0.077335 0.00065554 0.077986 0.069938 0 0.042303 0.0389 0 0.85241 0.23012 0.059917 0.0084777 4.1115 0.053235 6.354e-005 0.83683 0.0051116 0.0058494 0.0015022 0.98542 0.9907 3.2551e-006 1.3021e-005 0.13051 0.79228 0.82738 0.0014572 0.88204 0.51646 0.0019609 0.42286 1.4562 1.4533 16.0091 144.9839 0.00030685 -85.1703 0.25296
0.357 0.98802 5.5234e-005 3.8182 0.012045 4.7051e-006 0.001154 0.077462 0.00065555 0.078113 0.070055 0 0.042293 0.0389 0 0.85245 0.23014 0.059923 0.0084785 4.1115 0.053239 6.3545e-005 0.83682 0.0051116 0.0058494 0.0015013 0.98544 0.99071 3.2531e-006 1.3012e-005 0.13051 0.79287 0.82779 0.0014568 0.88275 0.51662 0.0019603 0.42287 1.4576 1.4548 16.0091 144.9839 0.00030619 -85.1738 0.25396
0.358 0.98802 5.5234e-005 3.8182 0.012045 4.7182e-006 0.001154 0.077588 0.00065556 0.078239 0.070171 0 0.042283 0.0389 0 0.85249 0.23016 0.059929 0.0084792 4.1116 0.053243 6.355e-005 0.83682 0.0051117 0.0058495 0.0015004 0.98545 0.99072 3.2511e-006 1.3004e-005 0.13051 0.79346 0.82819 0.0014563 0.88346 0.51679 0.0019597 0.42288 1.4591 1.4563 16.0091 144.984 0.00030553 -85.1773 0.25496
0.359 0.98802 5.5234e-005 3.8182 0.012045 4.7314e-006 0.001154 0.077715 0.00065557 0.078366 0.070287 0 0.042272 0.0389 0 0.85252 0.23017 0.059935 0.0084799 4.1116 0.053247 6.3555e-005 0.83682 0.0051118 0.0058496 0.0014996 0.98546 0.99072 3.2491e-006 1.2996e-005 0.13051 0.79406 0.8286 0.0014559 0.88416 0.51695 0.0019591 0.42289 1.4606 1.4578 16.0092 144.984 0.00030487 -85.1808 0.25596
0.36 0.98802 5.5234e-005 3.8182 0.012045 4.7446e-006 0.001154 0.077842 0.00065558 0.078493 0.070403 0 0.042262 0.0389 0 0.85256 0.23019 0.059941 0.0084807 4.1117 0.053251 6.356e-005 0.83681 0.0051118 0.0058496 0.0014987 0.98547 0.99073 3.2471e-006 1.2988e-005 0.13051 0.79464 0.829 0.0014554 0.88486 0.51712 0.0019585 0.4229 1.462 1.4592 16.0092 144.984 0.00030421 -85.1843 0.25696
0.361 0.98802 5.5234e-005 3.8182 0.012045 4.7577e-006 0.001154 0.077968 0.00065558 0.078619 0.070519 0 0.042251 0.0389 0 0.8526 0.23021 0.059947 0.0084814 4.1117 0.053255 6.3565e-005 0.83681 0.0051119 0.0058497 0.0014979 0.98548 0.99074 3.2451e-006 1.2981e-005 0.13051 0.79523 0.8294 0.001455 0.88556 0.51728 0.001958 0.42291 1.4635 1.4607 16.0092 144.984 0.00030356 -85.1877 0.25796
0.362 0.98802 5.5234e-005 3.8182 0.012045 4.7709e-006 0.001154 0.078094 0.00065559 0.078745 0.070635 0 0.042241 0.0389 0 0.85264 0.23022 0.059953 0.0084822 4.1118 0.053259 6.357e-005 0.8368 0.005112 0.0058498 0.001497 0.98549 0.99075 3.2432e-006 1.2973e-005 0.13051 0.79582 0.8298 0.0014546 0.88625 0.51745 0.0019574 0.42292 1.465 1.4622 16.0092 144.984 0.00030291 -85.1911 0.25896
0.363 0.98802 5.5234e-005 3.8182 0.012045 4.7841e-006 0.001154 0.078221 0.0006556 0.078872 0.070751 0 0.04223 0.0389 0 0.85267 0.23024 0.059959 0.0084829 4.1118 0.053263 6.3575e-005 0.8368 0.005112 0.0058498 0.0014962 0.9855 0.99076 3.2412e-006 1.2965e-005 0.13051 0.7964 0.8302 0.0014541 0.88694 0.51762 0.0019568 0.42293 1.4664 1.4636 16.0092 144.984 0.00030227 -85.1944 0.25996
0.364 0.98802 5.5234e-005 3.8182 0.012045 4.7973e-006 0.001154 0.078347 0.00065561 0.078998 0.070867 0 0.04222 0.0389 0 0.85271 0.23026 0.059965 0.0084837 4.1119 0.053267 6.358e-005 0.8368 0.0051121 0.0058499 0.0014954 0.98552 0.99076 3.2393e-006 1.2957e-005 0.13051 0.79698 0.83059 0.0014537 0.88762 0.51778 0.0019563 0.42294 1.4679 1.4651 16.0093 144.9841 0.00030162 -85.1978 0.26096
0.365 0.98802 5.5234e-005 3.8182 0.012045 4.8104e-006 0.001154 0.078473 0.00065562 0.079124 0.070982 0 0.04221 0.0389 0 0.85275 0.23027 0.059971 0.0084844 4.112 0.053271 6.3585e-005 0.83679 0.0051122 0.00585 0.0014945 0.98553 0.99077 3.2374e-006 1.295e-005 0.13052 0.79756 0.83099 0.0014533 0.8883 0.51795 0.0019557 0.42295 1.4693 1.4665 16.0093 144.9841 0.00030098 -85.2011 0.26196
0.366 0.98802 5.5234e-005 3.8182 0.012045 4.8236e-006 0.001154 0.078599 0.00065563 0.07925 0.071098 0 0.042199 0.0389 0 0.85279 0.23029 0.059976 0.0084852 4.112 0.053275 6.359e-005 0.83679 0.0051122 0.00585 0.0014937 0.98554 0.99078 3.2355e-006 1.2942e-005 0.13052 0.79814 0.83138 0.0014529 0.88898 0.51811 0.0019552 0.42296 1.4707 1.468 16.0093 144.9841 0.00030035 -85.2044 0.26296
0.367 0.98802 5.5234e-005 3.8182 0.012045 4.8368e-006 0.001154 0.078725 0.00065564 0.079376 0.071214 0 0.042189 0.0389 0 0.85282 0.23031 0.059982 0.0084859 4.1121 0.053279 6.3595e-005 0.83678 0.0051123 0.0058501 0.0014929 0.98555 0.99078 3.2336e-006 1.2935e-005 0.13052 0.79872 0.83177 0.0014525 0.88965 0.51828 0.0019546 0.42297 1.4722 1.4694 16.0093 144.9841 0.00029971 -85.2077 0.26396
0.368 0.98802 5.5233e-005 3.8182 0.012045 4.8499e-006 0.001154 0.07885 0.00065565 0.079501 0.071329 0 0.042179 0.0389 0 0.85286 0.23032 0.059988 0.0084867 4.1121 0.053283 6.3601e-005 0.83678 0.0051124 0.0058502 0.0014921 0.98556 0.99079 3.2318e-006 1.2927e-005 0.13052 0.79929 0.83216 0.001452 0.89032 0.51844 0.0019541 0.42298 1.4736 1.4709 16.0093 144.9841 0.00029908 -85.2109 0.26496
0.369 0.98802 5.5233e-005 3.8182 0.012045 4.8631e-006 0.001154 0.078976 0.00065566 0.079627 0.071444 0 0.042168 0.0389 0 0.8529 0.23034 0.059994 0.0084874 4.1122 0.053287 6.3606e-005 0.83678 0.0051124 0.0058502 0.0014913 0.98557 0.9908 3.2299e-006 1.292e-005 0.13052 0.79987 0.83254 0.0014516 0.89098 0.51861 0.0019536 0.42299 1.475 1.4723 16.0094 144.9841 0.00029845 -85.2142 0.26596
0.37 0.98802 5.5233e-005 3.8182 0.012045 4.8763e-006 0.001154 0.079102 0.00065567 0.079753 0.07156 0 0.042158 0.0389 0 0.85294 0.23036 0.060001 0.0084882 4.1122 0.053291 6.3611e-005 0.83677 0.0051125 0.0058503 0.0014905 0.98558 0.99081 3.2281e-006 1.2913e-005 0.13052 0.80044 0.83293 0.0014512 0.89164 0.51877 0.001953 0.423 1.4765 1.4738 16.0094 144.9842 0.00029783 -85.2174 0.26696
0.371 0.98802 5.5233e-005 3.8182 0.012045 4.8895e-006 0.001154 0.079227 0.00065568 0.079878 0.071675 0 0.042148 0.0389 0 0.85298 0.23037 0.060007 0.008489 4.1123 0.053295 6.3616e-005 0.83677 0.0051126 0.0058504 0.0014897 0.98559 0.99081 3.2263e-006 1.2905e-005 0.13052 0.80101 0.83331 0.0014508 0.8923 0.51894 0.0019525 0.42301 1.4779 1.4752 16.0094 144.9842 0.0002972 -85.2205 0.26796
0.372 0.98802 5.5233e-005 3.8182 0.012045 4.9026e-006 0.001154 0.079352 0.00065568 0.080003 0.07179 0 0.042137 0.0389 0 0.85301 0.23039 0.060013 0.0084897 4.1123 0.0533 6.3621e-005 0.83676 0.0051127 0.0058504 0.0014889 0.9856 0.99082 3.2245e-006 1.2898e-005 0.13052 0.80158 0.83369 0.0014504 0.89295 0.5191 0.001952 0.42302 1.4793 1.4766 16.0094 144.9842 0.00029658 -85.2237 0.26896
0.373 0.98802 5.5233e-005 3.8182 0.012045 4.9158e-006 0.001154 0.079478 0.00065569 0.080129 0.071905 0 0.042127 0.0389 0 0.85305 0.23041 0.060019 0.0084905 4.1124 0.053304 6.3626e-005 0.83676 0.0051127 0.0058505 0.0014881 0.98561 0.99083 3.2227e-006 1.2891e-005 0.13052 0.80214 0.83407 0.00145 0.8936 0.51927 0.0019515 0.42303 1.4807 1.478 16.0094 144.9842 0.00029597 -85.2268 0.26996
0.374 0.98802 5.5233e-005 3.8182 0.012045 4.929e-006 0.001154 0.079603 0.0006557 0.080254 0.07202 0 0.042117 0.0389 0 0.85309 0.23042 0.060025 0.0084913 4.1124 0.053308 6.3632e-005 0.83676 0.0051128 0.0058506 0.0014874 0.98562 0.99083 3.2209e-006 1.2884e-005 0.13052 0.80271 0.83445 0.0014496 0.89424 0.51943 0.0019509 0.42304 1.4821 1.4795 16.0095 144.9842 0.00029535 -85.2299 0.27096
0.375 0.98802 5.5233e-005 3.8182 0.012045 4.9421e-006 0.001154 0.079728 0.00065571 0.080379 0.072134 0 0.042107 0.0389 0 0.85313 0.23044 0.060031 0.008492 4.1125 0.053312 6.3637e-005 0.83675 0.0051129 0.0058506 0.0014866 0.98563 0.99084 3.2192e-006 1.2877e-005 0.13052 0.80327 0.83483 0.0014492 0.89489 0.5196 0.0019504 0.42305 1.4835 1.4809 16.0095 144.9842 0.00029474 -85.233 0.27196
0.376 0.98802 5.5233e-005 3.8182 0.012045 4.9553e-006 0.001154 0.079853 0.00065572 0.080504 0.072249 0 0.042096 0.0389 0 0.85317 0.23046 0.060037 0.0084928 4.1125 0.053316 6.3642e-005 0.83675 0.0051129 0.0058507 0.0014858 0.98564 0.99085 3.2174e-006 1.287e-005 0.13052 0.80383 0.8352 0.0014488 0.89552 0.51976 0.0019499 0.42306 1.4849 1.4823 16.0095 144.9843 0.00029413 -85.2361 0.27296
0.377 0.98802 5.5233e-005 3.8182 0.012045 4.9685e-006 0.001154 0.079978 0.00065573 0.080629 0.072364 0 0.042086 0.0389 0 0.85321 0.23047 0.060043 0.0084936 4.1126 0.05332 6.3647e-005 0.83674 0.005113 0.0058508 0.0014851 0.98565 0.99086 3.2157e-006 1.2863e-005 0.13052 0.80439 0.83557 0.0014485 0.89616 0.51993 0.0019494 0.42307 1.4863 1.4837 16.0095 144.9843 0.00029353 -85.2391 0.27396
0.378 0.98802 5.5233e-005 3.8182 0.012045 4.9817e-006 0.001154 0.080102 0.00065574 0.080753 0.072478 0 0.042076 0.0389 0 0.85324 0.23049 0.060049 0.0084943 4.1127 0.053324 6.3653e-005 0.83674 0.0051131 0.0058508 0.0014843 0.98566 0.99086 3.214e-006 1.2856e-005 0.13052 0.80495 0.83594 0.0014481 0.89679 0.52009 0.0019489 0.42308 1.4877 1.4851 16.0095 144.9843 0.00029293 -85.2422 0.27496
0.379 0.98802 5.5233e-005 3.8182 0.012045 4.9948e-006 0.001154 0.080227 0.00065575 0.080878 0.072593 0 0.042066 0.0389 0 0.85328 0.23051 0.060055 0.0084951 4.1127 0.053328 6.3658e-005 0.83674 0.0051131 0.0058509 0.0014836 0.98567 0.99087 3.2123e-006 1.2849e-005 0.13052 0.8055 0.83631 0.0014477 0.89741 0.52026 0.0019484 0.42309 1.4891 1.4865 16.0096 144.9843 0.00029233 -85.2451 0.27596
0.38 0.98802 5.5233e-005 3.8182 0.012045 5.008e-006 0.001154 0.080351 0.00065575 0.081003 0.072707 0 0.042056 0.0389 0 0.85332 0.23052 0.060061 0.0084959 4.1128 0.053333 6.3663e-005 0.83673 0.0051132 0.005851 0.0014829 0.98568 0.99087 3.2106e-006 1.2842e-005 0.13052 0.80606 0.83668 0.0014473 0.89803 0.52042 0.0019479 0.42311 1.4905 1.4879 16.0096 144.9843 0.00029173 -85.2481 0.27696
0.381 0.98802 5.5233e-005 3.8182 0.012045 5.0212e-006 0.001154 0.080476 0.00065576 0.081127 0.072821 0 0.042045 0.0389 0 0.85336 0.23054 0.060068 0.0084967 4.1128 0.053337 6.3669e-005 0.83673 0.0051133 0.0058511 0.0014821 0.98569 0.99088 3.2089e-006 1.2836e-005 0.13052 0.80661 0.83705 0.0014469 0.89865 0.52059 0.0019474 0.42312 1.4919 1.4893 16.0096 144.9843 0.00029113 -85.2511 0.27796
0.382 0.98802 5.5233e-005 3.8182 0.012045 5.0343e-006 0.001154 0.0806 0.00065577 0.081251 0.072936 0 0.042035 0.0389 0 0.8534 0.23056 0.060074 0.0084974 4.1129 0.053341 6.3674e-005 0.83672 0.0051134 0.0058511 0.0014814 0.9857 0.99089 3.2072e-006 1.2829e-005 0.13053 0.80716 0.83741 0.0014466 0.89927 0.52075 0.001947 0.42313 1.4933 1.4907 16.0096 144.9844 0.00029054 -85.254 0.27896
0.383 0.98802 5.5233e-005 3.8182 0.012045 5.0475e-006 0.001154 0.080724 0.00065578 0.081376 0.07305 0 0.042025 0.0389 0 0.85344 0.23058 0.06008 0.0084982 4.1129 0.053345 6.3679e-005 0.83672 0.0051134 0.0058512 0.0014807 0.98571 0.99089 3.2056e-006 1.2822e-005 0.13053 0.80771 0.83777 0.0014462 0.89988 0.52092 0.0019465 0.42314 1.4946 1.4921 16.0096 144.9844 0.00028995 -85.2569 0.27996
0.384 0.98802 5.5232e-005 3.8182 0.012045 5.0607e-006 0.001154 0.080849 0.00065579 0.0815 0.073164 0 0.042015 0.0389 0 0.85348 0.23059 0.060086 0.008499 4.113 0.053349 6.3685e-005 0.83671 0.0051135 0.0058513 0.00148 0.98572 0.9909 3.2039e-006 1.2816e-005 0.13053 0.80826 0.83814 0.0014458 0.90049 0.52108 0.001946 0.42315 1.496 1.4934 16.0096 144.9844 0.00028937 -85.2598 0.28096
0.385 0.98802 5.5232e-005 3.8182 0.012045 5.0738e-006 0.001154 0.080973 0.0006558 0.081624 0.073278 0 0.042005 0.0389 0 0.85352 0.23061 0.060092 0.0084998 4.1131 0.053354 6.369e-005 0.83671 0.0051136 0.0058513 0.0014793 0.98573 0.99091 3.2023e-006 1.2809e-005 0.13053 0.8088 0.8385 0.0014455 0.90109 0.52124 0.0019455 0.42316 1.4974 1.4948 16.0097 144.9844 0.00028878 -85.2627 0.28196
0.386 0.98802 5.5232e-005 3.8182 0.012045 5.087e-006 0.001154 0.081097 0.00065581 0.081748 0.073391 0 0.041995 0.0389 0 0.85356 0.23063 0.060099 0.0085006 4.1131 0.053358 6.3695e-005 0.83671 0.0051137 0.0058514 0.0014786 0.98574 0.99091 3.2007e-006 1.2803e-005 0.13053 0.80935 0.83885 0.0014451 0.90169 0.52141 0.001945 0.42317 1.4987 1.4962 16.0097 144.9844 0.0002882 -85.2655 0.28296
0.387 0.98802 5.5232e-005 3.8182 0.012045 5.1002e-006 0.001154 0.08122 0.00065581 0.081872 0.073505 0 0.041985 0.0389 0 0.85359 0.23065 0.060105 0.0085013 4.1132 0.053362 6.3701e-005 0.8367 0.0051137 0.0058515 0.0014779 0.98575 0.99092 3.1991e-006 1.2797e-005 0.13053 0.80989 0.83921 0.0014448 0.90229 0.52157 0.0019446 0.42318 1.5001 1.4976 16.0097 144.9845 0.00028762 -85.2684 0.28396
0.388 0.98802 5.5232e-005 3.8182 0.012045 5.1134e-006 0.001154 0.081344 0.00065582 0.081995 0.073619 0 0.041975 0.0389 0 0.85363 0.23066 0.060111 0.0085021 4.1132 0.053366 6.3706e-005 0.8367 0.0051138 0.0058516 0.0014772 0.98576 0.99093 3.1975e-006 1.279e-005 0.13053 0.81043 0.83956 0.0014444 0.90288 0.52174 0.0019441 0.42319 1.5015 1.4989 16.0097 144.9845 0.00028705 -85.2712 0.28496
0.389 0.98802 5.5232e-005 3.8182 0.012045 5.1265e-006 0.001154 0.081468 0.00065583 0.082119 0.073732 0 0.041965 0.0389 0 0.85367 0.23068 0.060117 0.0085029 4.1133 0.053371 6.3712e-005 0.83669 0.0051139 0.0058516 0.0014765 0.98577 0.99093 3.1959e-006 1.2784e-005 0.13053 0.81097 0.83992 0.0014441 0.90347 0.5219 0.0019437 0.4232 1.5028 1.5003 16.0097 144.9845 0.00028647 -85.274 0.28596
0.39 0.98802 5.5232e-005 3.8182 0.012045 5.1397e-006 0.001154 0.081591 0.00065584 0.082243 0.073846 0 0.041955 0.0389 0 0.85371 0.2307 0.060124 0.0085037 4.1134 0.053375 6.3717e-005 0.83669 0.005114 0.0058517 0.0014758 0.98578 0.99094 3.1944e-006 1.2778e-005 0.13053 0.81151 0.84027 0.0014437 0.90406 0.52207 0.0019432 0.42321 1.5042 1.5016 16.0097 144.9845 0.0002859 -85.2767 0.28696
0.391 0.98802 5.5232e-005 3.8182 0.012045 5.1529e-006 0.001154 0.081715 0.00065585 0.082366 0.073959 0 0.041945 0.0389 0 0.85375 0.23072 0.06013 0.0085045 4.1134 0.053379 6.3722e-005 0.83668 0.005114 0.0058518 0.0014751 0.98578 0.99094 3.1928e-006 1.2771e-005 0.13053 0.81204 0.84062 0.0014434 0.90464 0.52223 0.0019427 0.42322 1.5055 1.503 16.0098 144.9845 0.00028534 -85.2795 0.28796
0.392 0.98802 5.5232e-005 3.8182 0.012045 5.166e-006 0.001154 0.081838 0.00065586 0.082489 0.074073 0 0.041934 0.0389 0 0.85379 0.23073 0.060136 0.0085053 4.1135 0.053384 6.3728e-005 0.83668 0.0051141 0.0058519 0.0014744 0.98579 0.99095 3.1913e-006 1.2765e-005 0.13053 0.81257 0.84097 0.001443 0.90522 0.5224 0.0019423 0.42324 1.5069 1.5044 16.0098 144.9845 0.00028477 -85.2822 0.28896
0.393 0.98802 5.5232e-005 3.8182 0.012045 5.1792e-006 0.001154 0.081961 0.00065586 0.082613 0.074186 0 0.041924 0.0389 0 0.85383 0.23075 0.060143 0.0085061 4.1135 0.053388 6.3733e-005 0.83668 0.0051142 0.0058519 0.0014738 0.9858 0.99096 3.1898e-006 1.2759e-005 0.13053 0.81311 0.84132 0.0014427 0.90579 0.52256 0.0019418 0.42325 1.5082 1.5057 16.0098 144.9846 0.00028421 -85.2849 0.28996
0.394 0.98802 5.5232e-005 3.8182 0.012045 5.1924e-006 0.001154 0.082085 0.00065587 0.082736 0.074299 0 0.041914 0.0389 0 0.85387 0.23077 0.060149 0.0085069 4.1136 0.053392 6.3739e-005 0.83667 0.0051143 0.005852 0.0014731 0.98581 0.99096 3.1882e-006 1.2753e-005 0.13053 0.81364 0.84166 0.0014423 0.90637 0.52272 0.0019414 0.42326 1.5095 1.507 16.0098 144.9846 0.00028365 -85.2876 0.29096
0.395 0.98802 5.5232e-005 3.8182 0.012045 5.2055e-006 0.001154 0.082208 0.00065588 0.082859 0.074412 0 0.041904 0.0389 0 0.85391 0.23079 0.060155 0.0085077 4.1137 0.053397 6.3744e-005 0.83667 0.0051143 0.0058521 0.0014725 0.98582 0.99097 3.1867e-006 1.2747e-005 0.13053 0.81417 0.84201 0.001442 0.90693 0.52289 0.001941 0.42327 1.5109 1.5084 16.0098 144.9846 0.00028309 -85.2903 0.29196
0.396 0.98802 5.5232e-005 3.8182 0.012045 5.2187e-006 0.001154 0.082331 0.00065589 0.082982 0.074525 0 0.041895 0.0389 0 0.85395 0.2308 0.060162 0.0085085 4.1137 0.053401 6.375e-005 0.83666 0.0051144 0.0058522 0.0014718 0.98583 0.99097 3.1852e-006 1.2741e-005 0.13053 0.81469 0.84235 0.0014417 0.9075 0.52305 0.0019405 0.42328 1.5122 1.5097 16.0098 144.9846 0.00028253 -85.2929 0.29296
0.397 0.98802 5.5232e-005 3.8182 0.012045 5.2319e-006 0.001154 0.082453 0.0006559 0.083105 0.074638 0 0.041885 0.0389 0 0.85399 0.23082 0.060168 0.0085093 4.1138 0.053405 6.3755e-005 0.83666 0.0051145 0.0058522 0.0014712 0.98584 0.99098 3.1838e-006 1.2735e-005 0.13053 0.81522 0.84269 0.0014413 0.90806 0.52322 0.0019401 0.42329 1.5135 1.5111 16.0098 144.9846 0.00028198 -85.2955 0.29396
0.398 0.98802 5.5232e-005 3.8182 0.012045 5.2451e-006 0.001154 0.082576 0.0006559 0.083227 0.074751 0 0.041875 0.0389 0 0.85403 0.23084 0.060174 0.0085101 4.1138 0.05341 6.3761e-005 0.83665 0.0051146 0.0058523 0.0014706 0.98584 0.99098 3.1823e-006 1.2729e-005 0.13054 0.81574 0.84303 0.001441 0.90862 0.52338 0.0019397 0.4233 1.5148 1.5124 16.0099 144.9846 0.00028143 -85.2981 0.29496
0.399 0.98802 5.5232e-005 3.8182 0.012045 5.2582e-006 0.001154 0.082699 0.00065591 0.08335 0.074864 0 0.041865 0.0389 0 0.85407 0.23086 0.060181 0.0085109 4.1139 0.053414 6.3766e-005 0.83665 0.0051147 0.0058524 0.0014699 0.98585 0.99099 3.1808e-006 1.2723e-005 0.13054 0.81627 0.84337 0.0014407 0.90918 0.52354 0.0019392 0.42331 1.5162 1.5137 16.0099 144.9847 0.00028088 -85.3007 0.29596
0.4 0.98802 5.5231e-005 3.8182 0.012045 5.2714e-006 0.001154 0.082821 0.00065592 0.083473 0.074976 0 0.041855 0.0389 0 0.85411 0.23087 0.060187 0.0085117 4.114 0.053418 6.3772e-005 0.83665 0.0051147 0.0058525 0.0014693 0.98586 0.99099 3.1794e-006 1.2718e-005 0.13054 0.81679 0.8437 0.0014404 0.90973 0.52371 0.0019388 0.42332 1.5175 1.515 16.0099 144.9847 0.00028034 -85.3033 0.29696
0.401 0.98802 5.5231e-005 3.8182 0.012045 5.2846e-006 0.001154 0.082944 0.00065593 0.083595 0.075089 0 0.041845 0.0389 0 0.85415 0.23089 0.060193 0.0085125 4.114 0.053423 6.3778e-005 0.83664 0.0051148 0.0058525 0.0014687 0.98587 0.991 3.1779e-006 1.2712e-005 0.13054 0.81731 0.84404 0.00144 0.91028 0.52387 0.0019384 0.42334 1.5188 1.5164 16.0099 144.9847 0.0002798 -85.3059 0.29796
0.402 0.98802 5.5231e-005 3.8182 0.012045 5.2977e-006 0.001154 0.083066 0.00065594 0.083718 0.075201 0 0.041835 0.0389 0 0.85419 0.23091 0.0602 0.0085133 4.1141 0.053427 6.3783e-005 0.83664 0.0051149 0.0058526 0.001468 0.98588 0.99101 3.1765e-006 1.2706e-005 0.13054 0.81782 0.84437 0.0014397 0.91082 0.52404 0.001938 0.42335 1.5201 1.5177 16.0099 144.9847 0.00027925 -85.3084 0.29896
0.403 0.98802 5.5231e-005 3.8182 0.012045 5.3109e-006 0.001154 0.083188 0.00065594 0.08384 0.075314 0 0.041825 0.0389 0 0.85423 0.23093 0.060206 0.0085141 4.1142 0.053432 6.3789e-005 0.83663 0.005115 0.0058527 0.0014674 0.98589 0.99101 3.1751e-006 1.27e-005 0.13054 0.81834 0.84471 0.0014394 0.91136 0.5242 0.0019376 0.42336 1.5214 1.519 16.0099 144.9847 0.00027872 -85.3109 0.29996
0.404 0.98802 5.5231e-005 3.8182 0.012045 5.3241e-006 0.001154 0.083311 0.00065595 0.083962 0.075426 0 0.041815 0.0389 0 0.85427 0.23095 0.060213 0.0085149 4.1142 0.053436 6.3794e-005 0.83663 0.005115 0.0058528 0.0014668 0.98589 0.99102 3.1737e-006 1.2695e-005 0.13054 0.81885 0.84504 0.0014391 0.9119 0.52436 0.0019371 0.42337 1.5227 1.5203 16.0099 144.9847 0.00027818 -85.3134 0.30096
0.405 0.98802 5.5231e-005 3.8182 0.012045 5.3372e-006 0.001154 0.083433 0.00065596 0.084084 0.075538 0 0.041805 0.0389 0 0.85432 0.23096 0.060219 0.0085157 4.1143 0.05344 6.38e-005 0.83662 0.0051151 0.0058529 0.0014662 0.9859 0.99102 3.1723e-006 1.2689e-005 0.13054 0.81937 0.84537 0.0014388 0.91244 0.52453 0.0019367 0.42338 1.524 1.5216 16.0099 144.9848 0.00027765 -85.3159 0.30196
0.406 0.98802 5.5231e-005 3.8182 0.012045 5.3504e-006 0.001154 0.083555 0.00065597 0.084206 0.07565 0 0.041795 0.0389 0 0.85436 0.23098 0.060226 0.0085166 4.1143 0.053445 6.3806e-005 0.83662 0.0051152 0.0058529 0.0014656 0.98591 0.99103 3.1709e-006 1.2684e-005 0.13054 0.81988 0.84569 0.0014385 0.91297 0.52469 0.0019363 0.42339 1.5253 1.5229 16.01 144.9848 0.00027712 -85.3184 0.30296
0.407 0.98802 5.5231e-005 3.8182 0.012045 5.3636e-006 0.001154 0.083677 0.00065597 0.084328 0.075762 0 0.041786 0.0389 0 0.8544 0.231 0.060232 0.0085174 4.1144 0.053449 6.3811e-005 0.83661 0.0051153 0.005853 0.001465 0.98592 0.99103 3.1696e-006 1.2678e-005 0.13054 0.82039 0.84602 0.0014381 0.9135 0.52486 0.0019359 0.4234 1.5266 1.5242 16.01 144.9848 0.00027659 -85.3208 0.30396
0.408 0.98802 5.5231e-005 3.8182 0.012045 5.3768e-006 0.001154 0.083798 0.00065598 0.08445 0.075874 0 0.041776 0.0389 0 0.85444 0.23102 0.060239 0.0085182 4.1145 0.053454 6.3817e-005 0.83661 0.0051154 0.0058531 0.0014644 0.98593 0.99104 3.1682e-006 1.2673e-005 0.13054 0.82089 0.84635 0.0014378 0.91403 0.52502 0.0019355 0.42342 1.5279 1.5255 16.01 144.9848 0.00027606 -85.3232 0.30496
0.409 0.98802 5.5231e-005 3.8182 0.012045 5.3899e-006 0.001154 0.08392 0.00065599 0.084571 0.075986 0 0.041766 0.0389 0 0.85448 0.23103 0.060245 0.008519 4.1145 0.053458 6.3823e-005 0.83661 0.0051155 0.0058532 0.0014638 0.98593 0.99104 3.1668e-006 1.2667e-005 0.13054 0.8214 0.84667 0.0014375 0.91455 0.52518 0.0019351 0.42343 1.5292 1.5268 16.01 144.9848 0.00027554 -85.3256 0.30596
0.41 0.98802 5.5231e-005 3.8182 0.012045 5.4031e-006 0.001154 0.084042 0.000656 0.084693 0.076098 0 0.041756 0.0389 0 0.85452 0.23105 0.060252 0.0085198 4.1146 0.053463 6.3828e-005 0.8366 0.0051155 0.0058533 0.0014632 0.98594 0.99105 3.1655e-006 1.2662e-005 0.13054 0.82191 0.84699 0.0014372 0.91507 0.52535 0.0019347 0.42344 1.5304 1.5281 16.01 144.9849 0.00027502 -85.328 0.30696
0.411 0.98802 5.5231e-005 3.8182 0.012045 5.4163e-006 0.001154 0.084163 0.00065601 0.084815 0.076209 0 0.041746 0.0389 0 0.85456 0.23107 0.060258 0.0085207 4.1147 0.053467 6.3834e-005 0.8366 0.0051156 0.0058533 0.0014626 0.98595 0.99105 3.1642e-006 1.2657e-005 0.13054 0.82241 0.84731 0.0014369 0.91558 0.52551 0.0019343 0.42345 1.5317 1.5294 16.01 144.9849 0.0002745 -85.3304 0.30796
0.412 0.98802 5.5231e-005 3.8182 0.012045 5.4294e-006 0.001154 0.084284 0.00065601 0.084936 0.076321 0 0.041737 0.0389 0 0.8546 0.23109 0.060265 0.0085215 4.1147 0.053472 6.384e-005 0.83659 0.0051157 0.0058534 0.0014621 0.98596 0.99106 3.1628e-006 1.2651e-005 0.13054 0.82291 0.84763 0.0014366 0.9161 0.52567 0.001934 0.42346 1.533 1.5306 16.01 144.9849 0.00027398 -85.3328 0.30896
0.413 0.98802 5.5231e-005 3.8182 0.012045 5.4426e-006 0.001154 0.084406 0.00065602 0.085057 0.076433 0 0.041727 0.0389 0 0.85464 0.23111 0.060271 0.0085223 4.1148 0.053476 6.3846e-005 0.83659 0.0051158 0.0058535 0.0014615 0.98596 0.99106 3.1615e-006 1.2646e-005 0.13055 0.82341 0.84795 0.0014363 0.91661 0.52584 0.0019336 0.42347 1.5342 1.5319 16.01 144.9849 0.00027347 -85.3351 0.30996
0.414 0.98802 5.5231e-005 3.8182 0.012045 5.4558e-006 0.001154 0.084527 0.00065603 0.085178 0.076544 0 0.041717 0.0389 0 0.85468 0.23113 0.060278 0.0085231 4.1149 0.053481 6.3851e-005 0.83658 0.0051159 0.0058536 0.0014609 0.98597 0.99107 3.1602e-006 1.2641e-005 0.13055 0.82391 0.84827 0.0014361 0.91712 0.526 0.0019332 0.42348 1.5355 1.5332 16.0101 144.9849 0.00027296 -85.3374 0.31096
0.415 0.98802 5.5231e-005 3.8182 0.012045 5.4689e-006 0.001154 0.084648 0.00065604 0.085299 0.076655 0 0.041707 0.0389 0 0.85473 0.23114 0.060284 0.008524 4.1149 0.053485 6.3857e-005 0.83658 0.0051159 0.0058537 0.0014604 0.98598 0.99107 3.1589e-006 1.2636e-005 0.13055 0.82441 0.84858 0.0014358 0.91762 0.52616 0.0019328 0.4235 1.5368 1.5345 16.0101 144.9849 0.00027245 -85.3397 0.31196
0.416 0.98802 5.5231e-005 3.8182 0.012045 5.4821e-006 0.001154 0.084769 0.00065604 0.085421 0.076767 0 0.041698 0.0389 0 0.85477 0.23116 0.060291 0.0085248 4.115 0.05349 6.3863e-005 0.83657 0.005116 0.0058537 0.0014598 0.98599 0.99108 3.1577e-006 1.2631e-005 0.13055 0.8249 0.8489 0.0014355 0.91812 0.52633 0.0019324 0.42351 1.538 1.5357 16.0101 144.985 0.00027194 -85.342 0.31296
0.417 0.98802 5.523e-005 3.8182 0.012044 5.4953e-006 0.001154 0.08489 0.00065605 0.085541 0.076878 0 0.041688 0.0389 0 0.85481 0.23118 0.060298 0.0085256 4.1151 0.053494 6.3869e-005 0.83657 0.0051161 0.0058538 0.0014593 0.98599 0.99108 3.1564e-006 1.2626e-005 0.13055 0.8254 0.84921 0.0014352 0.91862 0.52649 0.0019321 0.42352 1.5393 1.537 16.0101 144.985 0.00027143 -85.3443 0.31396
0.418 0.98802 5.523e-005 3.8182 0.012044 5.5084e-006 0.001154 0.085011 0.00065606 0.085662 0.076989 0 0.041678 0.0389 0 0.85485 0.2312 0.060304 0.0085264 4.1151 0.053499 6.3874e-005 0.83656 0.0051162 0.0058539 0.0014587 0.986 0.99109 3.1551e-006 1.2621e-005 0.13055 0.82589 0.84952 0.0014349 0.91911 0.52665 0.0019317 0.42353 1.5405 1.5383 16.0101 144.985 0.00027093 -85.3466 0.31496
0.419 0.98802 5.523e-005 3.8182 0.012044 5.5216e-006 0.001154 0.085131 0.00065606 0.085783 0.0771 0 0.041668 0.0389 0 0.85489 0.23122 0.060311 0.0085273 4.1152 0.053504 6.388e-005 0.83656 0.0051163 0.005854 0.0014582 0.98601 0.99109 3.1539e-006 1.2616e-005 0.13055 0.82638 0.84983 0.0014346 0.91961 0.52682 0.0019313 0.42354 1.5418 1.5395 16.0101 144.985 0.00027043 -85.3488 0.31596
0.42 0.98802 5.523e-005 3.8182 0.012044 5.5348e-006 0.001154 0.085252 0.00065607 0.085904 0.077211 0 0.041659 0.0389 0 0.85493 0.23124 0.060318 0.0085281 4.1153 0.053508 6.3886e-005 0.83656 0.0051164 0.0058541 0.0014577 0.98602 0.9911 3.1526e-006 1.2611e-005 0.13055 0.82687 0.85014 0.0014344 0.9201 0.52698 0.001931 0.42355 1.543 1.5408 16.0101 144.985 0.00026993 -85.351 0.31696
0.421 0.98802 5.523e-005 3.8182 0.012044 5.548e-006 0.001154 0.085373 0.00065608 0.086024 0.077322 0 0.041649 0.0389 0 0.85498 0.23125 0.060324 0.0085289 4.1153 0.053513 6.3892e-005 0.83655 0.0051165 0.0058542 0.0014571 0.98602 0.9911 3.1514e-006 1.2606e-005 0.13055 0.82736 0.85045 0.0014341 0.92058 0.52714 0.0019306 0.42357 1.5443 1.542 16.0101 144.9851 0.00026943 -85.3533 0.31796
0.422 0.98802 5.523e-005 3.8182 0.012044 5.5611e-006 0.001154 0.085493 0.00065609 0.086145 0.077432 0 0.041639 0.0389 0 0.85502 0.23127 0.060331 0.0085298 4.1154 0.053517 6.3898e-005 0.83655 0.0051165 0.0058542 0.0014566 0.98603 0.99111 3.1502e-006 1.2601e-005 0.13055 0.82784 0.85075 0.0014338 0.92106 0.5273 0.0019302 0.42358 1.5455 1.5433 16.0101 144.9851 0.00026894 -85.3554 0.31896
0.423 0.98802 5.523e-005 3.8182 0.012044 5.5743e-006 0.001154 0.085613 0.00065609 0.086265 0.077543 0 0.04163 0.0389 0 0.85506 0.23129 0.060338 0.0085306 4.1155 0.053522 6.3904e-005 0.83654 0.0051166 0.0058543 0.001456 0.98604 0.99111 3.149e-006 1.2596e-005 0.13055 0.82833 0.85106 0.0014335 0.92154 0.52747 0.0019299 0.42359 1.5468 1.5445 16.0101 144.9851 0.00026845 -85.3576 0.31996
0.424 0.98802 5.523e-005 3.8182 0.012044 5.5875e-006 0.001154 0.085734 0.0006561 0.086385 0.077654 0 0.04162 0.0389 0 0.8551 0.23131 0.060344 0.0085315 4.1155 0.053527 6.391e-005 0.83654 0.0051167 0.0058544 0.0014555 0.98604 0.99112 3.1478e-006 1.2591e-005 0.13055 0.82881 0.85136 0.0014333 0.92202 0.52763 0.0019295 0.4236 1.548 1.5457 16.0102 144.9851 0.00026796 -85.3598 0.32096
0.425 0.98802 5.523e-005 3.8182 0.012044 5.6006e-006 0.001154 0.085854 0.00065611 0.086505 0.077764 0 0.04161 0.0389 0 0.85514 0.23133 0.060351 0.0085323 4.1156 0.053531 6.3915e-005 0.83653 0.0051168 0.0058545 0.001455 0.98605 0.99112 3.1466e-006 1.2586e-005 0.13055 0.82929 0.85166 0.001433 0.9225 0.52779 0.0019292 0.42361 1.5492 1.547 16.0102 144.9851 0.00026747 -85.3619 0.32196
0.426 0.98802 5.523e-005 3.8182 0.012044 5.6138e-006 0.001154 0.085974 0.00065612 0.086625 0.077875 0 0.041601 0.0389 0 0.85519 0.23135 0.060358 0.0085331 4.1157 0.053536 6.3921e-005 0.83653 0.0051169 0.0058546 0.0014545 0.98606 0.99112 3.1454e-006 1.2582e-005 0.13055 0.82977 0.85196 0.0014327 0.92297 0.52796 0.0019288 0.42362 1.5504 1.5482 16.0102 144.9851 0.00026698 -85.3641 0.32296
0.427 0.98802 5.523e-005 3.8182 0.012044 5.627e-006 0.001154 0.086094 0.00065612 0.086745 0.077985 0 0.041591 0.0389 0 0.85523 0.23137 0.060364 0.008534 4.1157 0.053541 6.3927e-005 0.83652 0.005117 0.0058547 0.001454 0.98606 0.99113 3.1442e-006 1.2577e-005 0.13056 0.83025 0.85226 0.0014324 0.92344 0.52812 0.0019285 0.42364 1.5517 1.5494 16.0102 144.9852 0.0002665 -85.3662 0.32396
0.428 0.98802 5.523e-005 3.8182 0.012044 5.6401e-006 0.001154 0.086213 0.00065613 0.086865 0.078095 0 0.041582 0.0389 0 0.85527 0.23138 0.060371 0.0085348 4.1158 0.053545 6.3933e-005 0.83652 0.0051171 0.0058548 0.0014534 0.98607 0.99113 3.143e-006 1.2572e-005 0.13056 0.83073 0.85256 0.0014322 0.9239 0.52828 0.0019281 0.42365 1.5529 1.5507 16.0102 144.9852 0.00026602 -85.3683 0.32496
0.429 0.98802 5.523e-005 3.8182 0.012044 5.6533e-006 0.001154 0.086333 0.00065614 0.086985 0.078205 0 0.041572 0.0389 0 0.85531 0.2314 0.060378 0.0085357 4.1159 0.05355 6.3939e-005 0.83651 0.0051172 0.0058548 0.0014529 0.98608 0.99114 3.1419e-006 1.2568e-005 0.13056 0.83121 0.85286 0.0014319 0.92436 0.52844 0.0019278 0.42366 1.5541 1.5519 16.0102 144.9852 0.00026554 -85.3704 0.32596
0.43 0.98802 5.523e-005 3.8182 0.012044 5.6665e-006 0.001154 0.086453 0.00065614 0.087104 0.078315 0 0.041563 0.0389 0 0.85536 0.23142 0.060385 0.0085365 4.116 0.053555 6.3945e-005 0.83651 0.0051172 0.0058549 0.0014524 0.98608 0.99114 3.1407e-006 1.2563e-005 0.13056 0.83168 0.85316 0.0014317 0.92483 0.52861 0.0019274 0.42367 1.5553 1.5531 16.0102 144.9852 0.00026506 -85.3725 0.32696
0.431 0.98802 5.523e-005 3.8182 0.012044 5.6796e-006 0.001154 0.086572 0.00065615 0.087224 0.078425 0 0.041553 0.0389 0 0.8554 0.23144 0.060391 0.0085374 4.116 0.053559 6.3951e-005 0.8365 0.0051173 0.005855 0.0014519 0.98609 0.99115 3.1396e-006 1.2558e-005 0.13056 0.83215 0.85345 0.0014314 0.92528 0.52877 0.0019271 0.42368 1.5565 1.5543 16.0102 144.9852 0.00026459 -85.3745 0.32796
0.432 0.98802 5.523e-005 3.8182 0.012044 5.6928e-006 0.001154 0.086692 0.00065616 0.087343 0.078535 0 0.041543 0.0389 0 0.85544 0.23146 0.060398 0.0085382 4.1161 0.053564 6.3957e-005 0.8365 0.0051174 0.0058551 0.0014514 0.9861 0.99115 3.1384e-006 1.2554e-005 0.13056 0.83263 0.85374 0.0014312 0.92574 0.52893 0.0019268 0.42369 1.5577 1.5555 16.0102 144.9853 0.00026412 -85.3766 0.32896
0.433 0.98802 5.5229e-005 3.8182 0.012044 5.706e-006 0.001154 0.086811 0.00065617 0.087463 0.078645 0 0.041534 0.0389 0 0.85548 0.23148 0.060405 0.0085391 4.1162 0.053569 6.3963e-005 0.8365 0.0051175 0.0058552 0.001451 0.9861 0.99115 3.1373e-006 1.2549e-005 0.13056 0.8331 0.85404 0.0014309 0.92619 0.52909 0.0019264 0.42371 1.5589 1.5567 16.0102 144.9853 0.00026364 -85.3786 0.32996
0.434 0.98802 5.5229e-005 3.8182 0.012044 5.7191e-006 0.001154 0.086931 0.00065617 0.087582 0.078755 0 0.041524 0.0389 0 0.85553 0.2315 0.060412 0.0085399 4.1162 0.053574 6.3969e-005 0.83649 0.0051176 0.0058553 0.0014505 0.98611 0.99116 3.1362e-006 1.2545e-005 0.13056 0.83357 0.85433 0.0014307 0.92664 0.52926 0.0019261 0.42372 1.5601 1.558 16.0102 144.9853 0.00026318 -85.3806 0.33096
0.435 0.98802 5.5229e-005 3.8182 0.012044 5.7323e-006 0.001154 0.08705 0.00065618 0.087701 0.078865 0 0.041515 0.0389 0 0.85557 0.23152 0.060418 0.0085408 4.1163 0.053578 6.3975e-005 0.83649 0.0051177 0.0058554 0.00145 0.98612 0.99116 3.1351e-006 1.254e-005 0.13056 0.83403 0.85462 0.0014304 0.92708 0.52942 0.0019258 0.42373 1.5613 1.5592 16.0102 144.9853 0.00026271 -85.3826 0.33196
0.436 0.98802 5.5229e-005 3.8182 0.012044 5.7455e-006 0.001154 0.087169 0.00065619 0.08782 0.078974 0 0.041505 0.0389 0 0.85561 0.23153 0.060425 0.0085417 4.1164 0.053583 6.3981e-005 0.83648 0.0051178 0.0058555 0.0014495 0.98612 0.99117 3.134e-006 1.2536e-005 0.13056 0.8345 0.85491 0.0014302 0.92753 0.52958 0.0019255 0.42374 1.5625 1.5604 16.0103 144.9853 0.00026224 -85.3846 0.33296
0.437 0.98802 5.5229e-005 3.8182 0.012044 5.7587e-006 0.001154 0.087288 0.00065619 0.087939 0.079084 0 0.041496 0.0389 0 0.85566 0.23155 0.060432 0.0085425 4.1165 0.053588 6.3987e-005 0.83648 0.0051179 0.0058556 0.001449 0.98613 0.99117 3.1329e-006 1.2532e-005 0.13056 0.83496 0.85519 0.0014299 0.92797 0.52974 0.0019251 0.42375 1.5637 1.5616 16.0103 144.9853 0.00026178 -85.3866 0.33396
0.438 0.98802 5.5229e-005 3.8182 0.012044 5.7718e-006 0.001154 0.087407 0.0006562 0.088058 0.079193 0 0.041486 0.0389 0 0.8557 0.23157 0.060439 0.0085434 4.1165 0.053593 6.3993e-005 0.83647 0.005118 0.0058556 0.0014486 0.98613 0.99118 3.1318e-006 1.2527e-005 0.13056 0.83543 0.85548 0.0014297 0.92841 0.52991 0.0019248 0.42377 1.5649 1.5627 16.0103 144.9854 0.00026132 -85.3885 0.33496
0.439 0.98802 5.5229e-005 3.8182 0.012044 5.785e-006 0.001154 0.087525 0.00065621 0.088177 0.079302 0 0.041477 0.0389 0 0.85574 0.23159 0.060446 0.0085442 4.1166 0.053597 6.3999e-005 0.83647 0.0051181 0.0058557 0.0014481 0.98614 0.99118 3.1307e-006 1.2523e-005 0.13056 0.83589 0.85576 0.0014294 0.92884 0.53007 0.0019245 0.42378 1.5661 1.5639 16.0103 144.9854 0.00026086 -85.3905 0.33596
0.44 0.98802 5.5229e-005 3.8182 0.012044 5.7982e-006 0.001154 0.087644 0.00065621 0.088296 0.079412 0 0.041467 0.0389 0 0.85579 0.23161 0.060453 0.0085451 4.1167 0.053602 6.4005e-005 0.83646 0.0051181 0.0058558 0.0014476 0.98615 0.99118 3.1297e-006 1.2519e-005 0.13056 0.83635 0.85605 0.0014292 0.92927 0.53023 0.0019242 0.42379 1.5672 1.5651 16.0103 144.9854 0.00026041 -85.3924 0.33696
0.441 0.98802 5.5229e-005 3.8182 0.012044 5.8113e-006 0.001154 0.087763 0.00065622 0.088414 0.079521 0 0.041458 0.0389 0 0.85583 0.23163 0.06046 0.008546 4.1168 0.053607 6.4012e-005 0.83646 0.0051182 0.0058559 0.0014472 0.98615 0.99119 3.1286e-006 1.2514e-005 0.13057 0.83681 0.85633 0.0014289 0.9297 0.53039 0.0019239 0.4238 1.5684 1.5663 16.0103 144.9854 0.00025995 -85.3943 0.33796
0.442 0.98802 5.5229e-005 3.8182 0.012044 5.8245e-006 0.001154 0.087881 0.00065623 0.088533 0.07963 0 0.041449 0.0389 0 0.85587 0.23165 0.060466 0.0085468 4.1168 0.053612 6.4018e-005 0.83645 0.0051183 0.005856 0.0014467 0.98616 0.99119 3.1275e-006 1.251e-005 0.13057 0.83726 0.85661 0.0014287 0.93013 0.53056 0.0019236 0.42381 1.5696 1.5675 16.0103 144.9854 0.0002595 -85.3962 0.33896
0.443 0.98802 5.5229e-005 3.8182 0.012044 5.8377e-006 0.001154 0.088 0.00065623 0.088651 0.079739 0 0.041439 0.0389 0 0.85592 0.23167 0.060473 0.0085477 4.1169 0.053617 6.4024e-005 0.83645 0.0051184 0.0058561 0.0014463 0.98616 0.9912 3.1265e-006 1.2506e-005 0.13057 0.83772 0.85689 0.0014285 0.93056 0.53072 0.0019233 0.42383 1.5708 1.5687 16.0103 144.9855 0.00025905 -85.3981 0.33996
0.444 0.98802 5.5229e-005 3.8182 0.012044 5.8508e-006 0.001154 0.088118 0.00065624 0.08877 0.079848 0 0.04143 0.0389 0 0.85596 0.23169 0.06048 0.0085486 4.117 0.053621 6.403e-005 0.83644 0.0051185 0.0058562 0.0014458 0.98617 0.9912 3.1255e-006 1.2502e-005 0.13057 0.83817 0.85717 0.0014282 0.93098 0.53088 0.0019229 0.42384 1.5719 1.5698 16.0103 144.9855 0.0002586 -85.4 0.34096
0.445 0.98802 5.5229e-005 3.8182 0.012044 5.864e-006 0.001154 0.088236 0.00065625 0.088888 0.079957 0 0.04142 0.0389 0 0.856 0.23171 0.060487 0.0085494 4.1171 0.053626 6.4036e-005 0.83644 0.0051186 0.0058563 0.0014454 0.98618 0.9912 3.1244e-006 1.2498e-005 0.13057 0.83863 0.85745 0.001428 0.9314 0.53104 0.0019226 0.42385 1.5731 1.571 16.0103 144.9855 0.00025815 -85.4018 0.34196
0.446 0.98802 5.5229e-005 3.8182 0.012044 5.8772e-006 0.001154 0.088354 0.00065625 0.089006 0.080065 0 0.041411 0.0389 0 0.85605 0.23173 0.060494 0.0085503 4.1171 0.053631 6.4042e-005 0.83643 0.0051187 0.0058564 0.0014449 0.98618 0.99121 3.1234e-006 1.2494e-005 0.13057 0.83908 0.85772 0.0014278 0.93182 0.5312 0.0019223 0.42386 1.5743 1.5722 16.0103 144.9855 0.00025771 -85.4037 0.34296
0.447 0.98802 5.5229e-005 3.8182 0.012044 5.8903e-006 0.001154 0.088472 0.00065626 0.089124 0.080174 0 0.041402 0.0389 0 0.85609 0.23175 0.060501 0.0085512 4.1172 0.053636 6.4048e-005 0.83643 0.0051188 0.0058565 0.0014444 0.98619 0.99121 3.1224e-006 1.249e-005 0.13057 0.83953 0.858 0.0014275 0.93223 0.53136 0.001922 0.42387 1.5754 1.5733 16.0103 144.9855 0.00025726 -85.4055 0.34396
0.448 0.98802 5.5229e-005 3.8182 0.012044 5.9035e-006 0.001154 0.08859 0.00065627 0.089242 0.080283 0 0.041392 0.0389 0 0.85613 0.23176 0.060508 0.0085521 4.1173 0.053641 6.4055e-005 0.83642 0.0051189 0.0058566 0.001444 0.98619 0.99121 3.1214e-006 1.2486e-005 0.13057 0.83998 0.85827 0.0014273 0.93264 0.53153 0.0019217 0.42389 1.5766 1.5745 16.0103 144.9855 0.00025682 -85.4073 0.34496
0.449 0.98802 5.5228e-005 3.8182 0.012044 5.9167e-006 0.001154 0.088708 0.00065627 0.08936 0.080391 0 0.041383 0.0389 0 0.85618 0.23178 0.060515 0.0085529 4.1174 0.053646 6.4061e-005 0.83642 0.005119 0.0058566 0.0014436 0.9862 0.99122 3.1204e-006 1.2482e-005 0.13057 0.84042 0.85855 0.0014271 0.93305 0.53169 0.0019214 0.4239 1.5777 1.5757 16.0103 144.9856 0.00025638 -85.4092 0.34596
0.45 0.98802 5.5228e-005 3.8182 0.012044 5.9298e-006 0.001154 0.088826 0.00065628 0.089477 0.080499 0 0.041374 0.0389 0 0.85622 0.2318 0.060522 0.0085538 4.1174 0.053651 6.4067e-005 0.83641 0.0051191 0.0058567 0.0014431 0.98621 0.99122 3.1194e-006 1.2478e-005 0.13057 0.84087 0.85882 0.0014268 0.93346 0.53185 0.0019212 0.42391 1.5789 1.5768 16.0103 144.9856 0.00025595 -85.4109 0.34696
0.451 0.98802 5.5228e-005 3.8182 0.012044 5.943e-006 0.001154 0.088943 0.00065629 0.089595 0.080608 0 0.041364 0.0389 0 0.85627 0.23182 0.060529 0.0085547 4.1175 0.053655 6.4073e-005 0.83641 0.0051192 0.0058568 0.0014427 0.98621 0.99123 3.1184e-006 1.2474e-005 0.13057 0.84131 0.85909 0.0014266 0.93386 0.53201 0.0019209 0.42392 1.58 1.578 16.0103 144.9856 0.00025551 -85.4127 0.34796
0.452 0.98802 5.5228e-005 3.8182 0.012044 5.9562e-006 0.001154 0.089061 0.00065629 0.089713 0.080716 0 0.041355 0.0389 0 0.85631 0.23184 0.060536 0.0085556 4.1176 0.05366 6.4079e-005 0.8364 0.0051193 0.0058569 0.0014423 0.98622 0.99123 3.1174e-006 1.247e-005 0.13057 0.84176 0.85936 0.0014264 0.93426 0.53217 0.0019206 0.42394 1.5812 1.5791 16.0103 144.9856 0.00025508 -85.4145 0.34896
0.453 0.98802 5.5228e-005 3.8182 0.012044 5.9693e-006 0.001154 0.089178 0.0006563 0.08983 0.080824 0 0.041346 0.0389 0 0.85635 0.23186 0.060543 0.0085565 4.1177 0.053665 6.4086e-005 0.8364 0.0051194 0.005857 0.0014418 0.98622 0.99123 3.1165e-006 1.2466e-005 0.13058 0.8422 0.85963 0.0014262 0.93466 0.53234 0.0019203 0.42395 1.5823 1.5803 16.0103 144.9856 0.00025465 -85.4163 0.34996
0.454 0.98802 5.5228e-005 3.8182 0.012044 5.9825e-006 0.001154 0.089296 0.00065631 0.089948 0.080932 0 0.041336 0.0389 0 0.8564 0.23188 0.06055 0.0085573 4.1177 0.05367 6.4092e-005 0.83639 0.0051195 0.0058571 0.0014414 0.98623 0.99124 3.1155e-006 1.2462e-005 0.13058 0.84264 0.8599 0.001426 0.93506 0.5325 0.00192 0.42396 1.5834 1.5814 16.0103 144.9857 0.00025422 -85.418 0.35096
0.455 0.98802 5.5228e-005 3.8182 0.012044 5.9957e-006 0.001154 0.089413 0.00065631 0.090065 0.08104 0 0.041327 0.0389 0 0.85644 0.2319 0.060557 0.0085582 4.1178 0.053675 6.4098e-005 0.83639 0.0051196 0.0058572 0.001441 0.98623 0.99124 3.1145e-006 1.2458e-005 0.13058 0.84308 0.86016 0.0014258 0.93546 0.53266 0.0019197 0.42397 1.5846 1.5825 16.0104 144.9857 0.00025379 -85.4197 0.35196
0.456 0.98802 5.5228e-005 3.8182 0.012044 6.0088e-006 0.001154 0.08953 0.00065632 0.090182 0.081148 0 0.041318 0.0389 0 0.85649 0.23192 0.060564 0.0085591 4.1179 0.05368 6.4105e-005 0.83638 0.0051197 0.0058573 0.0014406 0.98624 0.99124 3.1136e-006 1.2454e-005 0.13058 0.84352 0.86043 0.0014255 0.93585 0.53282 0.0019194 0.42398 1.5857 1.5837 16.0104 144.9857 0.00025336 -85.4215 0.35296
0.457 0.98802 5.5228e-005 3.8182 0.012044 6.022e-006 0.001154 0.089647 0.00065633 0.090299 0.081256 0 0.041309 0.0389 0 0.85653 0.23194 0.060571 0.00856 4.118 0.053685 6.4111e-005 0.83638 0.0051198 0.0058574 0.0014402 0.98624 0.99125 3.1126e-006 1.2451e-005 0.13058 0.84395 0.86069 0.0014253 0.93624 0.53298 0.0019192 0.424 1.5868 1.5848 16.0104 144.9857 0.00025294 -85.4232 0.35396
0.458 0.98802 5.5228e-005 3.8182 0.012044 6.0352e-006 0.001154 0.089764 0.00065633 0.090416 0.081364 0 0.041299 0.0389 0 0.85658 0.23196 0.060578 0.0085609 4.1181 0.05369 6.4117e-005 0.83637 0.0051199 0.0058575 0.0014398 0.98625 0.99125 3.1117e-006 1.2447e-005 0.13058 0.84439 0.86096 0.0014251 0.93662 0.53314 0.0019189 0.42401 1.5879 1.5859 16.0104 144.9857 0.00025252 -85.4249 0.35496
0.459 0.98802 5.5228e-005 3.8182 0.012044 6.0483e-006 0.001154 0.089881 0.00065634 0.090533 0.081471 0 0.04129 0.0389 0 0.85662 0.23198 0.060585 0.0085618 4.1181 0.053695 6.4123e-005 0.83637 0.00512 0.0058576 0.0014394 0.98625 0.99125 3.1108e-006 1.2443e-005 0.13058 0.84482 0.86122 0.0014249 0.93701 0.5333 0.0019186 0.42402 1.5891 1.5871 16.0104 144.9858 0.0002521 -85.4266 0.35596
0.46 0.98802 5.5228e-005 3.8182 0.012044 6.0615e-006 0.001154 0.089998 0.00065635 0.09065 0.081579 0 0.041281 0.0389 0 0.85667 0.232 0.060592 0.0085627 4.1182 0.0537 6.413e-005 0.83636 0.0051201 0.0058577 0.001439 0.98626 0.99126 3.1099e-006 1.2439e-005 0.13058 0.84525 0.86148 0.0014247 0.93739 0.53347 0.0019183 0.42403 1.5902 1.5882 16.0104 144.9858 0.00025168 -85.4282 0.35696
0.461 0.98802 5.5228e-005 3.8182 0.012044 6.0747e-006 0.001154 0.090115 0.00065635 0.090767 0.081686 0 0.041272 0.0389 0 0.85671 0.23202 0.0606 0.0085636 4.1183 0.053705 6.4136e-005 0.83636 0.0051202 0.0058578 0.0014386 0.98626 0.99126 3.1089e-006 1.2436e-005 0.13058 0.84568 0.86174 0.0014245 0.93777 0.53363 0.0019181 0.42405 1.5913 1.5893 16.0104 144.9858 0.00025126 -85.4299 0.35796
0.462 0.98802 5.5228e-005 3.8182 0.012044 6.0878e-006 0.001154 0.090231 0.00065636 0.090883 0.081794 0 0.041262 0.0389 0 0.85676 0.23204 0.060607 0.0085645 4.1184 0.05371 6.4142e-005 0.83635 0.0051203 0.0058579 0.0014382 0.98627 0.99127 3.108e-006 1.2432e-005 0.13058 0.84611 0.862 0.0014243 0.93815 0.53379 0.0019178 0.42406 1.5924 1.5904 16.0104 144.9858 0.00025085 -85.4316 0.35896
0.463 0.98802 5.5228e-005 3.8182 0.012044 6.101e-006 0.001154 0.090348 0.00065636 0.091 0.081901 0 0.041253 0.0389 0 0.8568 0.23206 0.060614 0.0085654 4.1185 0.053715 6.4149e-005 0.83635 0.0051204 0.005858 0.0014378 0.98628 0.99127 3.1071e-006 1.2429e-005 0.13058 0.84654 0.86226 0.0014241 0.93852 0.53395 0.0019175 0.42407 1.5935 1.5915 16.0104 144.9858 0.00025043 -85.4332 0.35996
0.464 0.98802 5.5228e-005 3.8182 0.012044 6.1142e-006 0.001154 0.090464 0.00065637 0.091116 0.082008 0 0.041244 0.0389 0 0.85685 0.23208 0.060621 0.0085663 4.1185 0.05372 6.4155e-005 0.83634 0.0051205 0.0058581 0.0014374 0.98628 0.99127 3.1062e-006 1.2425e-005 0.13058 0.84697 0.86251 0.0014239 0.9389 0.53411 0.0019173 0.42408 1.5946 1.5927 16.0104 144.9858 0.00025002 -85.4348 0.36096
0.465 0.98802 5.5227e-005 3.8182 0.012044 6.1273e-006 0.001154 0.090581 0.00065638 0.091232 0.082116 0 0.041235 0.0389 0 0.85689 0.2321 0.060628 0.0085672 4.1186 0.053725 6.4162e-005 0.83634 0.0051206 0.0058582 0.001437 0.98629 0.99128 3.1054e-006 1.2421e-005 0.13058 0.84739 0.86277 0.0014237 0.93927 0.53427 0.001917 0.4241 1.5957 1.5938 16.0104 144.9859 0.00024961 -85.4364 0.36196
0.466 0.98802 5.5227e-005 3.8182 0.012044 6.1405e-006 0.001154 0.090697 0.00065638 0.091349 0.082223 0 0.041226 0.0389 0 0.85694 0.23212 0.060635 0.0085681 4.1187 0.05373 6.4168e-005 0.83633 0.0051207 0.0058583 0.0014366 0.98629 0.99128 3.1045e-006 1.2418e-005 0.13059 0.84782 0.86302 0.0014235 0.93964 0.53443 0.0019167 0.42411 1.5968 1.5949 16.0104 144.9859 0.0002492 -85.438 0.36296
0.467 0.98802 5.5227e-005 3.8182 0.012044 6.1537e-006 0.001154 0.090813 0.00065639 0.091465 0.08233 0 0.041217 0.0389 0 0.85698 0.23214 0.060642 0.008569 4.1188 0.053735 6.4174e-005 0.83633 0.0051208 0.0058584 0.0014362 0.9863 0.99128 3.1036e-006 1.2414e-005 0.13059 0.84824 0.86328 0.0014233 0.94 0.53459 0.0019165 0.42412 1.5979 1.596 16.0104 144.9859 0.0002488 -85.4396 0.36396
0.468 0.98802 5.5227e-005 3.8182 0.012044 6.1668e-006 0.001154 0.090929 0.0006564 0.091581 0.082437 0 0.041207 0.0389 0 0.85703 0.23216 0.06065 0.0085699 4.1189 0.05374 6.4181e-005 0.83632 0.0051209 0.0058585 0.0014359 0.9863 0.99128 3.1027e-006 1.2411e-005 0.13059 0.84866 0.86353 0.0014231 0.94037 0.53475 0.0019162 0.42413 1.599 1.5971 16.0104 144.9859 0.00024839 -85.4412 0.36496
0.469 0.98802 5.5227e-005 3.8182 0.012044 6.18e-006 0.001154 0.091045 0.0006564 0.091697 0.082543 0 0.041198 0.0389 0 0.85707 0.23218 0.060657 0.0085708 4.1189 0.053745 6.4187e-005 0.83632 0.005121 0.0058586 0.0014355 0.98631 0.99129 3.1019e-006 1.2407e-005 0.13059 0.84908 0.86378 0.0014229 0.94073 0.53491 0.001916 0.42414 1.6001 1.5982 16.0104 144.9859 0.00024799 -85.4428 0.36596
0.47 0.98802 5.5227e-005 3.8182 0.012044 6.1932e-006 0.001154 0.091161 0.00065641 0.091813 0.08265 0 0.041189 0.0389 0 0.85712 0.2322 0.060664 0.0085717 4.119 0.05375 6.4194e-005 0.83631 0.0051211 0.0058587 0.0014351 0.98631 0.99129 3.101e-006 1.2404e-005 0.13059 0.8495 0.86403 0.0014227 0.94109 0.53508 0.0019157 0.42416 1.6012 1.5993 16.0104 144.986 0.00024759 -85.4443 0.36696
0.471 0.98802 5.5227e-005 3.8182 0.012044 6.2063e-006 0.001154 0.091277 0.00065641 0.091929 0.082757 0 0.04118 0.0389 0 0.85716 0.23222 0.060671 0.0085726 4.1191 0.053755 6.42e-005 0.83631 0.0051212 0.0058588 0.0014347 0.98631 0.99129 3.1002e-006 1.2401e-005 0.13059 0.84992 0.86428 0.0014225 0.94145 0.53524 0.0019155 0.42417 1.6023 1.6004 16.0104 144.986 0.00024719 -85.4459 0.36796
0.472 0.98802 5.5227e-005 3.8182 0.012044 6.2195e-006 0.001154 0.091392 0.00065642 0.092044 0.082863 0 0.041171 0.0389 0 0.85721 0.23224 0.060678 0.0085735 4.1192 0.053761 6.4207e-005 0.8363 0.0051213 0.0058589 0.0014344 0.98632 0.9913 3.0993e-006 1.2397e-005 0.13059 0.85034 0.86453 0.0014223 0.9418 0.5354 0.0019152 0.42418 1.6033 1.6014 16.0104 144.986 0.00024679 -85.4474 0.36896
0.473 0.98802 5.5227e-005 3.8182 0.012044 6.2327e-006 0.001154 0.091508 0.00065643 0.09216 0.08297 0 0.041162 0.0389 0 0.85725 0.23226 0.060686 0.0085744 4.1193 0.053766 6.4213e-005 0.8363 0.0051214 0.005859 0.001434 0.98632 0.9913 3.0985e-006 1.2394e-005 0.13059 0.85075 0.86478 0.0014221 0.94215 0.53556 0.001915 0.42419 1.6044 1.6025 16.0104 144.986 0.00024639 -85.449 0.36996
0.474 0.98802 5.5227e-005 3.8182 0.012044 6.2458e-006 0.001154 0.091624 0.00065643 0.092275 0.083076 0 0.041153 0.0389 0 0.8573 0.23228 0.060693 0.0085753 4.1194 0.053771 6.422e-005 0.83629 0.0051215 0.0058591 0.0014337 0.98633 0.9913 3.0976e-006 1.2391e-005 0.13059 0.85117 0.86502 0.0014219 0.9425 0.53572 0.0019147 0.42421 1.6055 1.6036 16.0104 144.986 0.000246 -85.4505 0.37096
0.475 0.98802 5.5227e-005 3.8182 0.012044 6.259e-006 0.001154 0.091739 0.00065644 0.092391 0.083183 0 0.041144 0.0389 0 0.85734 0.2323 0.0607 0.0085762 4.1194 0.053776 6.4226e-005 0.83629 0.0051216 0.0058592 0.0014333 0.98633 0.99131 3.0968e-006 1.2387e-005 0.13059 0.85158 0.86527 0.0014217 0.94285 0.53588 0.0019145 0.42422 1.6066 1.6047 16.0104 144.9861 0.00024561 -85.452 0.37196
0.476 0.98802 5.5227e-005 3.8182 0.012044 6.2722e-006 0.001154 0.091854 0.00065644 0.092506 0.083289 0 0.041135 0.0389 0 0.85739 0.23232 0.060708 0.0085771 4.1195 0.053781 6.4233e-005 0.83628 0.0051217 0.0058593 0.0014329 0.98634 0.99131 3.096e-006 1.2384e-005 0.13059 0.85199 0.86551 0.0014215 0.9432 0.53604 0.0019142 0.42423 1.6076 1.6058 16.0104 144.9861 0.00024521 -85.4535 0.37296
0.477 0.98802 5.5227e-005 3.8182 0.012044 6.2853e-006 0.001154 0.091969 0.00065645 0.092621 0.083395 0 0.041126 0.0389 0 0.85744 0.23234 0.060715 0.008578 4.1196 0.053786 6.4239e-005 0.83628 0.0051218 0.0058594 0.0014326 0.98634 0.99131 3.0952e-006 1.2381e-005 0.1306 0.8524 0.86575 0.0014214 0.94354 0.5362 0.001914 0.42424 1.6087 1.6068 16.0104 144.9861 0.00024483 -85.455 0.37396
0.478 0.98802 5.5227e-005 3.8182 0.012044 6.2985e-006 0.001154 0.092085 0.00065646 0.092736 0.083501 0 0.041117 0.0389 0 0.85748 0.23236 0.060722 0.008579 4.1197 0.053791 6.4246e-005 0.83627 0.0051219 0.0058595 0.0014322 0.98635 0.99132 3.0944e-006 1.2377e-005 0.1306 0.85281 0.866 0.0014212 0.94389 0.53636 0.0019137 0.42426 1.6098 1.6079 16.0104 144.9861 0.00024444 -85.4564 0.37496
0.479 0.98802 5.5227e-005 3.8182 0.012044 6.3117e-006 0.001154 0.0922 0.00065646 0.092852 0.083607 0 0.041108 0.0389 0 0.85753 0.23238 0.060729 0.0085799 4.1198 0.053796 6.4252e-005 0.83627 0.005122 0.0058596 0.0014319 0.98635 0.99132 3.0936e-006 1.2374e-005 0.1306 0.85322 0.86624 0.001421 0.94423 0.53652 0.0019135 0.42427 1.6108 1.609 16.0104 144.9861 0.00024405 -85.4579 0.37596
0.48 0.98802 5.5227e-005 3.8182 0.012044 6.3248e-006 0.001154 0.092315 0.00065647 0.092966 0.083713 0 0.041099 0.0389 0 0.85757 0.2324 0.060737 0.0085808 4.1199 0.053802 6.4259e-005 0.83626 0.0051221 0.0058597 0.0014315 0.98636 0.99132 3.0928e-006 1.2371e-005 0.1306 0.85362 0.86648 0.0014208 0.94456 0.53668 0.0019133 0.42428 1.6119 1.61 16.0104 144.9861 0.00024367 -85.4594 0.37696
0.481 0.98802 5.5226e-005 3.8182 0.012044 6.338e-006 0.001154 0.092429 0.00065647 0.093081 0.083819 0 0.04109 0.0389 0 0.85762 0.23242 0.060744 0.0085817 4.12 0.053807 6.4266e-005 0.83626 0.0051222 0.0058598 0.0014312 0.98636 0.99133 3.092e-006 1.2368e-005 0.1306 0.85403 0.86672 0.0014206 0.9449 0.53684 0.001913 0.42429 1.6129 1.6111 16.0104 144.9862 0.00024328 -85.4608 0.37796
0.482 0.98802 5.5226e-005 3.8182 0.012044 6.3512e-006 0.001154 0.092544 0.00065648 0.093196 0.083925 0 0.041081 0.0389 0 0.85767 0.23244 0.060751 0.0085826 4.12 0.053812 6.4272e-005 0.83625 0.0051223 0.0058599 0.0014309 0.98637 0.99133 3.0912e-006 1.2365e-005 0.1306 0.85443 0.86696 0.0014205 0.94523 0.537 0.0019128 0.42431 1.614 1.6122 16.0104 144.9862 0.0002429 -85.4622 0.37896
0.483 0.98802 5.5226e-005 3.8182 0.012044 6.3643e-006 0.001154 0.092659 0.00065649 0.093311 0.084031 0 0.041072 0.0389 0 0.85771 0.23246 0.060759 0.0085836 4.1201 0.053817 6.4279e-005 0.83625 0.0051224 0.00586 0.0014305 0.98637 0.99133 3.0904e-006 1.2362e-005 0.1306 0.85483 0.86719 0.0014203 0.94556 0.53716 0.0019126 0.42432 1.615 1.6132 16.0104 144.9862 0.00024252 -85.4637 0.37996
0.484 0.98802 5.5226e-005 3.8182 0.012044 6.3775e-006 0.001154 0.092773 0.00065649 0.093425 0.084136 0 0.041063 0.0389 0 0.85776 0.23248 0.060766 0.0085845 4.1202 0.053822 6.4285e-005 0.83624 0.0051225 0.0058601 0.0014302 0.98637 0.99133 3.0897e-006 1.2359e-005 0.1306 0.85524 0.86743 0.0014201 0.94589 0.53732 0.0019123 0.42433 1.6161 1.6143 16.0104 144.9862 0.00024214 -85.4651 0.38096
0.485 0.98802 5.5226e-005 3.8182 0.012044 6.3907e-006 0.001154 0.092888 0.0006565 0.09354 0.084242 0 0.041054 0.0389 0 0.85781 0.2325 0.060773 0.0085854 4.1203 0.053828 6.4292e-005 0.83624 0.0051226 0.0058602 0.0014298 0.98638 0.99134 3.0889e-006 1.2356e-005 0.1306 0.85564 0.86767 0.0014199 0.94622 0.53748 0.0019121 0.42435 1.6171 1.6153 16.0104 144.9862 0.00024177 -85.4665 0.38196
0.486 0.98802 5.5226e-005 3.8182 0.012044 6.4038e-006 0.001154 0.093002 0.0006565 0.093654 0.084347 0 0.041045 0.0389 0 0.85785 0.23252 0.060781 0.0085863 4.1204 0.053833 6.4299e-005 0.83623 0.0051228 0.0058604 0.0014295 0.98638 0.99134 3.0881e-006 1.2352e-005 0.1306 0.85603 0.8679 0.0014198 0.94655 0.53764 0.0019119 0.42436 1.6182 1.6164 16.0104 144.9863 0.00024139 -85.4679 0.38296
0.487 0.98802 5.5226e-005 3.8182 0.012044 6.417e-006 0.001154 0.093117 0.00065651 0.093769 0.084453 0 0.041036 0.0389 0 0.8579 0.23254 0.060788 0.0085873 4.1205 0.053838 6.4305e-005 0.83623 0.0051229 0.0058605 0.0014292 0.98639 0.99134 3.0874e-006 1.2349e-005 0.1306 0.85643 0.86813 0.0014196 0.94687 0.5378 0.0019117 0.42437 1.6192 1.6174 16.0104 144.9863 0.00024102 -85.4693 0.38396
0.488 0.98802 5.5226e-005 3.8182 0.012044 6.4302e-006 0.001154 0.093231 0.00065652 0.093883 0.084558 0 0.041027 0.0389 0 0.85795 0.23256 0.060796 0.0085882 4.1206 0.053843 6.4312e-005 0.83622 0.005123 0.0058606 0.0014288 0.98639 0.99135 3.0866e-006 1.2346e-005 0.13061 0.85683 0.86837 0.0014194 0.94719 0.53796 0.0019114 0.42438 1.6203 1.6184 16.0104 144.9863 0.00024065 -85.4706 0.38496
0.489 0.98802 5.5226e-005 3.8182 0.012044 6.4433e-006 0.001154 0.093345 0.00065652 0.093997 0.084663 0 0.041018 0.0389 0 0.85799 0.23258 0.060803 0.0085891 4.1207 0.053849 6.4319e-005 0.83622 0.0051231 0.0058607 0.0014285 0.9864 0.99135 3.0859e-006 1.2343e-005 0.13061 0.85722 0.8686 0.0014192 0.94751 0.53812 0.0019112 0.4244 1.6213 1.6195 16.0104 144.9863 0.00024028 -85.472 0.38596
0.49 0.98802 5.5226e-005 3.8182 0.012044 6.4565e-006 0.001154 0.093459 0.00065653 0.094111 0.084768 0 0.041009 0.0389 0 0.85804 0.2326 0.06081 0.0085901 4.1207 0.053854 6.4325e-005 0.83621 0.0051232 0.0058608 0.0014282 0.9864 0.99135 3.0851e-006 1.234e-005 0.13061 0.85762 0.86883 0.0014191 0.94783 0.53828 0.001911 0.42441 1.6223 1.6205 16.0104 144.9863 0.00023991 -85.4734 0.38696
0.491 0.98802 5.5226e-005 3.8182 0.012044 6.4697e-006 0.001154 0.093573 0.00065653 0.094225 0.084873 0 0.041 0.0389 0 0.85809 0.23262 0.060818 0.008591 4.1208 0.053859 6.4332e-005 0.83621 0.0051233 0.0058609 0.0014279 0.9864 0.99135 3.0844e-006 1.2338e-005 0.13061 0.85801 0.86906 0.0014189 0.94814 0.53844 0.0019108 0.42442 1.6233 1.6216 16.0104 144.9864 0.00023954 -85.4747 0.38796
0.492 0.98802 5.5226e-005 3.8182 0.012043 6.4828e-006 0.001154 0.093687 0.00065654 0.094339 0.084978 0 0.040992 0.0389 0 0.85813 0.23265 0.060825 0.0085919 4.1209 0.053864 6.4339e-005 0.8362 0.0051234 0.005861 0.0014276 0.98641 0.99136 3.0837e-006 1.2335e-005 0.13061 0.8584 0.86929 0.0014188 0.94846 0.5386 0.0019106 0.42443 1.6244 1.6226 16.0104 144.9864 0.00023918 -85.476 0.38896
0.493 0.98802 5.5226e-005 3.8182 0.012043 6.496e-006 0.001154 0.093801 0.00065654 0.094452 0.085083 0 0.040983 0.0389 0 0.85818 0.23267 0.060833 0.0085929 4.121 0.05387 6.4346e-005 0.83619 0.0051235 0.0058611 0.0014273 0.98641 0.99136 3.0829e-006 1.2332e-005 0.13061 0.85879 0.86952 0.0014186 0.94877 0.53876 0.0019103 0.42445 1.6254 1.6236 16.0104 144.9864 0.00023881 -85.4774 0.38996
0.494 0.98802 5.5226e-005 3.8182 0.012043 6.5092e-006 0.001154 0.093914 0.00065655 0.094566 0.085188 0 0.040974 0.0389 0 0.85823 0.23269 0.06084 0.0085938 4.1211 0.053875 6.4352e-005 0.83619 0.0051236 0.0058612 0.001427 0.98642 0.99136 3.0822e-006 1.2329e-005 0.13061 0.85918 0.86974 0.0014184 0.94908 0.53892 0.0019101 0.42446 1.6264 1.6246 16.0104 144.9864 0.00023845 -85.4787 0.39096
0.495 0.98802 5.5226e-005 3.8182 0.012043 6.5223e-006 0.001154 0.094028 0.00065656 0.09468 0.085293 0 0.040965 0.0389 0 0.85827 0.23271 0.060848 0.0085947 4.1212 0.05388 6.4359e-005 0.83618 0.0051237 0.0058613 0.0014266 0.98642 0.99136 3.0815e-006 1.2326e-005 0.13061 0.85957 0.86997 0.0014183 0.94938 0.53908 0.0019099 0.42447 1.6274 1.6257 16.0104 144.9864 0.00023809 -85.48 0.39196
0.496 0.98802 5.5226e-005 3.8182 0.012043 6.5355e-006 0.001154 0.094141 0.00065656 0.094793 0.085397 0 0.040956 0.0389 0 0.85832 0.23273 0.060855 0.0085957 4.1213 0.053886 6.4366e-005 0.83618 0.0051239 0.0058614 0.0014263 0.98643 0.99137 3.0808e-006 1.2323e-005 0.13061 0.85995 0.8702 0.0014181 0.94969 0.53924 0.0019097 0.42448 1.6284 1.6267 16.0104 144.9864 0.00023773 -85.4813 0.39296
0.497 0.98802 5.5226e-005 3.8182 0.012043 6.5487e-006 0.001154 0.094255 0.00065657 0.094907 0.085502 0 0.040947 0.0389 0 0.85837 0.23275 0.060863 0.0085966 4.1214 0.053891 6.4373e-005 0.83617 0.005124 0.0058615 0.001426 0.98643 0.99137 3.0801e-006 1.232e-005 0.13061 0.86034 0.87042 0.0014179 0.94999 0.5394 0.0019095 0.4245 1.6294 1.6277 16.0104 144.9865 0.00023737 -85.4826 0.39396
0.498 0.98802 5.5225e-005 3.8182 0.012043 6.5618e-006 0.001154 0.094368 0.00065657 0.09502 0.085606 0 0.040939 0.0389 0 0.85841 0.23277 0.06087 0.0085976 4.1215 0.053896 6.4379e-005 0.83617 0.0051241 0.0058617 0.0014256 0.98643 0.99137 3.0794e-006 1.2317e-005 0.13061 0.86072 0.87064 0.0014177 0.9503 0.53956 0.0019093 0.42451 1.6305 1.6287 16.0104 144.9865 0.00023701 -85.4839 0.39496
0.499 0.98802 5.5225e-005 3.8182 0.012043 6.575e-006 0.001154 0.094481 0.00065658 0.095133 0.085711 0 0.04093 0.0389 0 0.85846 0.23279 0.060878 0.0085985 4.1216 0.053902 6.4386e-005 0.83616 0.0051242 0.0058618 0.0014253 0.98644 0.99137 3.0787e-006 1.2315e-005 0.13062 0.86111 0.87087 0.0014176 0.95059 0.53972 0.0019091 0.42452 1.6315 1.6297 16.0104 144.9865 0.00023666 -85.4852 0.39596
0.5 0.98802 5.5225e-005 3.8182 0.012043 6.5882e-006 0.001154 0.094594 0.00065658 0.095246 0.085815 0 0.040921 0.0389 0 0.85851 0.23281 0.060885 0.0085995 4.1216 0.053907 6.4393e-005 0.83616 0.0051243 0.0058619 0.001425 0.98644 0.99138 3.078e-006 1.2312e-005 0.13062 0.86149 0.87109 0.0014174 0.95089 0.53988 0.0019089 0.42454 1.6325 1.6307 16.0104 144.9865 0.0002363 -85.4864 0.39696
0.501 0.98802 5.5225e-005 3.8182 0.012043 6.6013e-006 0.001154 0.094707 0.00065659 0.095359 0.085919 0 0.040912 0.0389 0 0.85856 0.23283 0.060893 0.0086004 4.1217 0.053912 6.44e-005 0.83615 0.0051244 0.005862 0.0014248 0.98644 0.99138 3.0773e-006 1.2309e-005 0.13062 0.86187 0.87131 0.0014173 0.95119 0.54004 0.0019087 0.42455 1.6335 1.6317 16.0104 144.9865 0.00023595 -85.4877 0.39796
0.502 0.98802 5.5225e-005 3.8182 0.012043 6.6145e-006 0.001154 0.09482 0.00065659 0.095472 0.086024 0 0.040903 0.0389 0 0.8586 0.23285 0.0609 0.0086014 4.1218 0.053918 6.4407e-005 0.83615 0.0051245 0.0058621 0.0014246 0.98645 0.99138 3.0767e-006 1.2307e-005 0.13062 0.86225 0.87153 0.0014172 0.95148 0.5402 0.0019085 0.42456 1.6345 1.6327 16.0104 144.9866 0.0002356 -85.4889 0.39896
0.503 0.98802 5.5225e-005 3.8182 0.012043 6.6277e-006 0.001154 0.094933 0.0006566 0.095585 0.086128 0 0.040895 0.0389 0 0.85865 0.23287 0.060908 0.0086023 4.1219 0.053923 6.4414e-005 0.83614 0.0051246 0.0058622 0.0014243 0.98645 0.99138 3.076e-006 1.2304e-005 0.13062 0.86263 0.87175 0.001417 0.95178 0.54035 0.0019083 0.42457 1.6355 1.6337 16.0104 144.9866 0.00023525 -85.4902 0.39996
0.504 0.98802 5.5225e-005 3.8182 0.012043 6.6408e-006 0.001154 0.095046 0.00065661 0.095698 0.086232 0 0.040886 0.0389 0 0.8587 0.2329 0.060916 0.0086033 4.122 0.053929 6.442e-005 0.83614 0.0051248 0.0058623 0.0014241 0.98646 0.99139 3.0753e-006 1.2301e-005 0.13062 0.863 0.87197 0.0014169 0.95207 0.54051 0.0019081 0.42459 1.6364 1.6347 16.0104 144.9866 0.0002349 -85.4914 0.40096
0.505 0.98802 5.5225e-005 3.8182 0.012043 6.654e-006 0.001154 0.095159 0.00065661 0.095811 0.086336 0 0.040877 0.0389 0 0.85875 0.23292 0.060923 0.0086042 4.1221 0.053934 6.4427e-005 0.83613 0.0051249 0.0058624 0.0014238 0.98646 0.99139 3.0747e-006 1.2299e-005 0.13062 0.86338 0.87218 0.0014167 0.95236 0.54067 0.0019079 0.4246 1.6374 1.6357 16.0104 144.9866 0.00023456 -85.4926 0.40196
0.506 0.98802 5.5225e-005 3.8182 0.012043 6.6672e-006 0.001154 0.095271 0.00065662 0.095923 0.086439 0 0.040868 0.0389 0 0.8588 0.23294 0.060931 0.0086052 4.1222 0.053939 6.4434e-005 0.83612 0.005125 0.0058626 0.0014235 0.98646 0.99139 3.074e-006 1.2296e-005 0.13062 0.86375 0.8724 0.0014166 0.95264 0.54083 0.0019077 0.42461 1.6384 1.6367 16.0104 144.9866 0.00023421 -85.4938 0.40296
0.507 0.98802 5.5225e-005 3.8182 0.012043 6.6803e-006 0.001154 0.095384 0.00065662 0.096036 0.086543 0 0.04086 0.0389 0 0.85884 0.23296 0.060938 0.0086061 4.1223 0.053945 6.4441e-005 0.83612 0.0051251 0.0058627 0.0014232 0.98647 0.99139 3.0733e-006 1.2293e-005 0.13062 0.86413 0.87262 0.0014164 0.95293 0.54099 0.0019075 0.42462 1.6394 1.6377 16.0104 144.9867 0.00023387 -85.495 0.40396
0.508 0.98802 5.5225e-005 3.8182 0.012043 6.6935e-006 0.001154 0.095496 0.00065663 0.096148 0.086647 0 0.040851 0.0389 0 0.85889 0.23298 0.060946 0.0086071 4.1224 0.05395 6.4448e-005 0.83611 0.0051252 0.0058628 0.0014228 0.98647 0.9914 3.0727e-006 1.2291e-005 0.13062 0.8645 0.87283 0.0014163 0.95321 0.54115 0.0019073 0.42464 1.6404 1.6387 16.0104 144.9867 0.00023353 -85.4962 0.40496
0.509 0.98802 5.5225e-005 3.8182 0.012043 6.7066e-006 0.001154 0.095608 0.00065663 0.09626 0.086751 0 0.040842 0.0389 0 0.85894 0.233 0.060954 0.008608 4.1225 0.053956 6.4455e-005 0.83611 0.0051253 0.0058629 0.0014225 0.98648 0.9914 3.072e-006 1.2288e-005 0.13062 0.86487 0.87304 0.0014161 0.95349 0.54131 0.0019071 0.42465 1.6414 1.6397 16.0103 144.9867 0.00023319 -85.4974 0.40596
0.51 0.98802 5.5225e-005 3.8182 0.012043 6.7198e-006 0.001154 0.09572 0.00065664 0.096373 0.086854 0 0.040834 0.0389 0 0.85899 0.23302 0.060961 0.008609 4.1226 0.053961 6.4462e-005 0.8361 0.0051255 0.005863 0.0014222 0.98648 0.9914 3.0714e-006 1.2286e-005 0.13063 0.86524 0.87326 0.001416 0.95377 0.54147 0.0019069 0.42466 1.6423 1.6407 16.0103 144.9867 0.00023285 -85.4986 0.40696
0.511 0.98802 5.5225e-005 3.8182 0.012043 6.733e-006 0.001154 0.095833 0.00065664 0.096485 0.086958 0 0.040825 0.0389 0 0.85904 0.23304 0.060969 0.0086099 4.1227 0.053967 6.4469e-005 0.8361 0.0051256 0.0058631 0.0014219 0.98648 0.9914 3.0708e-006 1.2283e-005 0.13063 0.86561 0.87347 0.0014158 0.95405 0.54163 0.0019067 0.42468 1.6433 1.6416 16.0103 144.9867 0.00023251 -85.4998 0.40796
0.512 0.98802 5.5225e-005 3.8182 0.012043 6.7461e-006 0.001154 0.095945 0.00065665 0.096597 0.087061 0 0.040816 0.0389 0 0.85908 0.23306 0.060977 0.0086109 4.1228 0.053972 6.4476e-005 0.83609 0.0051257 0.0058632 0.0014216 0.98649 0.99141 3.0701e-006 1.228e-005 0.13063 0.86598 0.87368 0.0014157 0.95433 0.54179 0.0019065 0.42469 1.6443 1.6426 16.0103 144.9868 0.00023217 -85.5009 0.40896
0.513 0.98802 5.5225e-005 3.8182 0.012043 6.7593e-006 0.001154 0.096057 0.00065665 0.096709 0.087164 0 0.040808 0.0389 0 0.85913 0.23309 0.060984 0.0086119 4.1229 0.053978 6.4483e-005 0.83609 0.0051258 0.0058634 0.0014214 0.98649 0.99141 3.0695e-006 1.2278e-005 0.13063 0.86634 0.87389 0.0014155 0.9546 0.54194 0.0019063 0.4247 1.6453 1.6436 16.0103 144.9868 0.00023184 -85.5021 0.40996
0.514 0.98802 5.5224e-005 3.8182 0.012043 6.7725e-006 0.001154 0.096168 0.00065666 0.09682 0.087267 0 0.040799 0.0389 0 0.85918 0.23311 0.060992 0.0086128 4.123 0.053983 6.449e-005 0.83608 0.0051259 0.0058635 0.0014211 0.98649 0.99141 3.0689e-006 1.2275e-005 0.13063 0.86671 0.8741 0.0014154 0.95487 0.5421 0.0019061 0.42471 1.6462 1.6446 16.0103 144.9868 0.0002315 -85.5032 0.41096
0.515 0.98802 5.5224e-005 3.8182 0.012043 6.7856e-006 0.001154 0.09628 0.00065666 0.096932 0.087371 0 0.04079 0.0389 0 0.85923 0.23313 0.061 0.0086138 4.1231 0.053989 6.4497e-005 0.83608 0.005126 0.0058636 0.0014208 0.9865 0.99141 3.0682e-006 1.2273e-005 0.13063 0.86707 0.87431 0.0014152 0.95515 0.54226 0.001906 0.42473 1.6472 1.6455 16.0103 144.9868 0.00023117 -85.5044 0.41196
0.516 0.98802 5.5224e-005 3.8182 0.012043 6.7988e-006 0.001154 0.096392 0.00065667 0.097044 0.087474 0 0.040782 0.0389 0 0.85928 0.23315 0.061007 0.0086148 4.1232 0.053994 6.4504e-005 0.83607 0.0051262 0.0058637 0.0014205 0.9865 0.99142 3.0676e-006 1.227e-005 0.13063 0.86744 0.87452 0.0014151 0.95541 0.54242 0.0019058 0.42474 1.6481 1.6465 16.0103 144.9868 0.00023084 -85.5055 0.41296
0.517 0.98802 5.5224e-005 3.8182 0.012043 6.812e-006 0.001154 0.096503 0.00065667 0.097156 0.087577 0 0.040773 0.0389 0 0.85933 0.23317 0.061015 0.0086157 4.1233 0.054 6.4511e-005 0.83606 0.0051263 0.0058638 0.0014203 0.9865 0.99142 3.067e-006 1.2268e-005 0.13063 0.8678 0.87472 0.0014149 0.95568 0.54258 0.0019056 0.42475 1.6491 1.6475 16.0103 144.9869 0.00023051 -85.5066 0.41396
0.518 0.98802 5.5224e-005 3.8182 0.012043 6.8251e-006 0.001154 0.096615 0.00065668 0.097267 0.087679 0 0.040764 0.0389 0 0.85937 0.23319 0.061023 0.0086167 4.1234 0.054005 6.4518e-005 0.83606 0.0051264 0.0058639 0.00142 0.98651 0.99142 3.0664e-006 1.2266e-005 0.13063 0.86816 0.87493 0.0014148 0.95595 0.54274 0.0019054 0.42477 1.6501 1.6484 16.0103 144.9869 0.00023018 -85.5077 0.41496
0.519 0.98802 5.5224e-005 3.8182 0.012043 6.8383e-006 0.001154 0.096726 0.00065669 0.097378 0.087782 0 0.040756 0.0389 0 0.85942 0.23321 0.06103 0.0086177 4.1234 0.054011 6.4525e-005 0.83605 0.0051265 0.0058641 0.0014198 0.98651 0.99142 3.0658e-006 1.2263e-005 0.13063 0.86852 0.87514 0.0014147 0.95621 0.5429 0.0019052 0.42478 1.651 1.6494 16.0103 144.9869 0.00022986 -85.5088 0.41596
0.52 0.98802 5.5224e-005 3.8182 0.012043 6.8515e-006 0.001154 0.096838 0.00065669 0.09749 0.087885 0 0.040747 0.0389 0 0.85947 0.23324 0.061038 0.0086186 4.1235 0.054016 6.4532e-005 0.83605 0.0051266 0.0058642 0.0014195 0.98651 0.99142 3.0652e-006 1.2261e-005 0.13064 0.86888 0.87534 0.0014145 0.95648 0.54305 0.0019051 0.42479 1.652 1.6503 16.0103 144.9869 0.00022953 -85.5099 0.41696
0.521 0.98802 5.5224e-005 3.8182 0.012043 6.8646e-006 0.001154 0.096949 0.0006567 0.097601 0.087988 0 0.040739 0.0389 0 0.85952 0.23326 0.061046 0.0086196 4.1236 0.054022 6.4539e-005 0.83604 0.0051268 0.0058643 0.0014192 0.98652 0.99143 3.0646e-006 1.2258e-005 0.13064 0.86924 0.87555 0.0014144 0.95674 0.54321 0.0019049 0.4248 1.6529 1.6513 16.0103 144.9869 0.00022921 -85.511 0.41796
0.522 0.98802 5.5224e-005 3.8182 0.012043 6.8778e-006 0.001154 0.09706 0.0006567 0.097712 0.08809 0 0.04073 0.0389 0 0.85957 0.23328 0.061054 0.0086206 4.1237 0.054027 6.4546e-005 0.83604 0.0051269 0.0058644 0.001419 0.98652 0.99143 3.064e-006 1.2256e-005 0.13064 0.86959 0.87575 0.0014143 0.957 0.54337 0.0019047 0.42482 1.6539 1.6522 16.0103 144.9869 0.00022888 -85.5121 0.41896
0.523 0.98802 5.5224e-005 3.8182 0.012043 6.891e-006 0.001154 0.097171 0.00065671 0.097823 0.088193 0 0.040722 0.0389 0 0.85962 0.2333 0.061061 0.0086216 4.1238 0.054033 6.4553e-005 0.83603 0.005127 0.0058645 0.0014188 0.98652 0.99143 3.0635e-006 1.2254e-005 0.13064 0.86995 0.87595 0.0014141 0.95725 0.54353 0.0019045 0.42483 1.6548 1.6532 16.0103 144.987 0.00022856 -85.5132 0.41996
0.524 0.98802 5.5224e-005 3.8182 0.012043 6.9041e-006 0.001154 0.097282 0.00065671 0.097934 0.088295 0 0.040713 0.0389 0 0.85967 0.23332 0.061069 0.0086225 4.1239 0.054038 6.456e-005 0.83603 0.0051271 0.0058647 0.0014185 0.98653 0.99143 3.0629e-006 1.2251e-005 0.13064 0.8703 0.87615 0.001414 0.95751 0.54369 0.0019044 0.42484 1.6557 1.6541 16.0103 144.987 0.00022824 -85.5143 0.42096
0.525 0.98802 5.5224e-005 3.8182 0.012043 6.9173e-006 0.001154 0.097393 0.00065672 0.098045 0.088397 0 0.040705 0.0389 0 0.85972 0.23334 0.061077 0.0086235 4.124 0.054044 6.4567e-005 0.83602 0.0051273 0.0058648 0.0014182 0.98653 0.99144 3.0623e-006 1.2249e-005 0.13064 0.87066 0.87635 0.0014139 0.95776 0.54385 0.0019042 0.42486 1.6567 1.6551 16.0103 144.987 0.00022792 -85.5153 0.42196
0.526 0.98802 5.5224e-005 3.8182 0.012043 6.9304e-006 0.001154 0.097504 0.00065672 0.098156 0.0885 0 0.040696 0.0389 0 0.85977 0.23337 0.061085 0.0086245 4.1241 0.05405 6.4574e-005 0.83601 0.0051274 0.0058649 0.001418 0.98653 0.99144 3.0617e-006 1.2247e-005 0.13064 0.87101 0.87655 0.0014138 0.95802 0.544 0.001904 0.42487 1.6576 1.656 16.0103 144.987 0.0002276 -85.5164 0.42296
0.527 0.98802 5.5224e-005 3.8182 0.012043 6.9436e-006 0.001154 0.097614 0.00065673 0.098267 0.088602 0 0.040688 0.0389 0 0.85981 0.23339 0.061093 0.0086255 4.1242 0.054055 6.4581e-005 0.83601 0.0051275 0.005865 0.0014177 0.98654 0.99144 3.0612e-006 1.2245e-005 0.13064 0.87136 0.87675 0.0014136 0.95827 0.54416 0.0019038 0.42488 1.6585 1.6569 16.0103 144.987 0.00022729 -85.5174 0.42396
0.528 0.98802 5.5224e-005 3.8182 0.012043 6.9568e-006 0.001154 0.097725 0.00065673 0.098377 0.088704 0 0.040679 0.0389 0 0.85986 0.23341 0.061101 0.0086265 4.1243 0.054061 6.4588e-005 0.836 0.0051276 0.0058651 0.0014175 0.98654 0.99144 3.0606e-006 1.2242e-005 0.13064 0.87171 0.87695 0.0014135 0.95852 0.54432 0.0019037 0.42489 1.6595 1.6579 16.0103 144.9871 0.00022697 -85.5185 0.42496
0.529 0.98802 5.5224e-005 3.8182 0.012043 6.9699e-006 0.001154 0.097836 0.00065674 0.098488 0.088806 0 0.040671 0.0389 0 0.85991 0.23343 0.061108 0.0086274 4.1244 0.054066 6.4596e-005 0.836 0.0051277 0.0058653 0.0014173 0.98654 0.99144 3.06e-006 1.224e-005 0.13064 0.87206 0.87715 0.0014134 0.95877 0.54448 0.0019035 0.42491 1.6604 1.6588 16.0102 144.9871 0.00022666 -85.5195 0.42596
0.53 0.98802 5.5223e-005 3.8182 0.012043 6.9831e-006 0.001154 0.097946 0.00065674 0.098598 0.088908 0 0.040662 0.0389 0 0.85996 0.23345 0.061116 0.0086284 4.1245 0.054072 6.4603e-005 0.83599 0.0051279 0.0058654 0.001417 0.98655 0.99145 3.0595e-006 1.2238e-005 0.13065 0.87241 0.87734 0.0014132 0.95901 0.54464 0.0019033 0.42492 1.6613 1.6597 16.0102 144.9871 0.00022634 -85.5205 0.42696
0.531 0.98802 5.5223e-005 3.8182 0.012043 6.9963e-006 0.001154 0.098056 0.00065675 0.098708 0.08901 0 0.040654 0.0389 0 0.86001 0.23347 0.061124 0.0086294 4.1246 0.054078 6.461e-005 0.83599 0.005128 0.0058655 0.0014168 0.98655 0.99145 3.0589e-006 1.2236e-005 0.13065 0.87275 0.87754 0.0014131 0.95926 0.54479 0.0019032 0.42493 1.6622 1.6607 16.0102 144.9871 0.00022603 -85.5216 0.42796
0.532 0.98802 5.5223e-005 3.8182 0.012043 7.0094e-006 0.001154 0.098167 0.00065675 0.098819 0.089112 0 0.040645 0.0389 0 0.86006 0.2335 0.061132 0.0086304 4.1248 0.054083 6.4617e-005 0.83598 0.0051281 0.0058656 0.0014165 0.98655 0.99145 3.0584e-006 1.2233e-005 0.13065 0.8731 0.87774 0.001413 0.9595 0.54495 0.001903 0.42495 1.6632 1.6616 16.0102 144.9871 0.00022572 -85.5226 0.42896
0.533 0.98802 5.5223e-005 3.8182 0.012043 7.0226e-006 0.001154 0.098277 0.00065676 0.098929 0.089213 0 0.040637 0.0389 0 0.86011 0.23352 0.06114 0.0086314 4.1249 0.054089 6.4624e-005 0.83598 0.0051282 0.0058658 0.0014163 0.98656 0.99145 3.0578e-006 1.2231e-005 0.13065 0.87344 0.87793 0.0014129 0.95974 0.54511 0.0019029 0.42496 1.6641 1.6625 16.0102 144.9872 0.00022541 -85.5236 0.42996
0.534 0.98802 5.5223e-005 3.8182 0.012043 7.0358e-006 0.001154 0.098387 0.00065676 0.099039 0.089315 0 0.040628 0.0389 0 0.86016 0.23354 0.061148 0.0086324 4.125 0.054095 6.4632e-005 0.83597 0.0051284 0.0058659 0.001416 0.98656 0.99145 3.0573e-006 1.2229e-005 0.13065 0.87379 0.87812 0.0014127 0.95998 0.54527 0.0019027 0.42497 1.665 1.6634 16.0102 144.9872 0.00022511 -85.5246 0.43096
0.535 0.98802 5.5223e-005 3.8182 0.012043 7.0489e-006 0.001154 0.098497 0.00065677 0.099149 0.089417 0 0.04062 0.0389 0 0.86021 0.23356 0.061156 0.0086334 4.1251 0.0541 6.4639e-005 0.83596 0.0051285 0.005866 0.0014158 0.98656 0.99146 3.0568e-006 1.2227e-005 0.13065 0.87413 0.87832 0.0014126 0.96022 0.54542 0.0019025 0.42499 1.6659 1.6644 16.0102 144.9872 0.0002248 -85.5256 0.43196
0.536 0.98802 5.5223e-005 3.8182 0.012043 7.0621e-006 0.001154 0.098607 0.00065677 0.099259 0.089518 0 0.040611 0.0389 0 0.86026 0.23358 0.061164 0.0086344 4.1252 0.054106 6.4646e-005 0.83596 0.0051286 0.0058661 0.0014156 0.98656 0.99146 3.0562e-006 1.2225e-005 0.13065 0.87447 0.87851 0.0014125 0.96046 0.54558 0.0019024 0.425 1.6668 1.6653 16.0102 144.9872 0.0002245 -85.5265 0.43296
0.537 0.98802 5.5223e-005 3.8182 0.012043 7.0753e-006 0.001154 0.098716 0.00065678 0.099369 0.089619 0 0.040603 0.0389 0 0.86031 0.23361 0.061171 0.0086353 4.1253 0.054112 6.4653e-005 0.83595 0.0051288 0.0058663 0.0014154 0.98657 0.99146 3.0557e-006 1.2223e-005 0.13065 0.87481 0.8787 0.0014124 0.9607 0.54574 0.0019022 0.42501 1.6677 1.6662 16.0102 144.9872 0.00022419 -85.5275 0.43396
0.538 0.98802 5.5223e-005 3.8182 0.012043 7.0884e-006 0.001154 0.098826 0.00065678 0.099478 0.089721 0 0.040595 0.0389 0 0.86036 0.23363 0.061179 0.0086363 4.1254 0.054117 6.466e-005 0.83595 0.0051289 0.0058664 0.0014151 0.98657 0.99146 3.0552e-006 1.2221e-005 0.13065 0.87515 0.87889 0.0014123 0.96093 0.5459 0.0019021 0.42502 1.6686 1.6671 16.0102 144.9873 0.00022389 -85.5285 0.43496
0.539 0.98802 5.5223e-005 3.8182 0.012043 7.1016e-006 0.001154 0.098936 0.00065679 0.099588 0.089822 0 0.040586 0.0389 0 0.86041 0.23365 0.061187 0.0086373 4.1255 0.054123 6.4668e-005 0.83594 0.005129 0.0058665 0.0014149 0.98657 0.99146 3.0546e-006 1.2219e-005 0.13066 0.87549 0.87908 0.0014121 0.96116 0.54605 0.0019019 0.42504 1.6695 1.668 16.0102 144.9873 0.00022359 -85.5295 0.43596
0.54 0.98802 5.5223e-005 3.8182 0.012043 7.1147e-006 0.001154 0.099045 0.00065679 0.099698 0.089923 0 0.040578 0.0389 0 0.86046 0.23367 0.061195 0.0086383 4.1256 0.054129 6.4675e-005 0.83594 0.0051291 0.0058666 0.0014147 0.98658 0.99147 3.0541e-006 1.2216e-005 0.13066 0.87582 0.87927 0.001412 0.9614 0.54621 0.0019017 0.42505 1.6704 1.6689 16.0102 144.9873 0.00022329 -85.5304 0.43696
0.541 0.98802 5.5223e-005 3.8182 0.012043 7.1279e-006 0.001154 0.099155 0.0006568 0.099807 0.090024 0 0.040569 0.0389 0 0.86051 0.23369 0.061203 0.0086393 4.1257 0.054135 6.4682e-005 0.83593 0.0051293 0.0058668 0.0014145 0.98658 0.99147 3.0536e-006 1.2214e-005 0.13066 0.87616 0.87946 0.0014119 0.96163 0.54637 0.0019016 0.42506 1.6713 1.6698 16.0102 144.9873 0.00022299 -85.5314 0.43796
0.542 0.98802 5.5223e-005 3.8182 0.012043 7.1411e-006 0.001154 0.099264 0.0006568 0.099916 0.090125 0 0.040561 0.0389 0 0.86056 0.23372 0.061211 0.0086403 4.1258 0.05414 6.469e-005 0.83592 0.0051294 0.0058669 0.0014142 0.98658 0.99147 3.0531e-006 1.2212e-005 0.13066 0.87649 0.87965 0.0014118 0.96185 0.54653 0.0019014 0.42508 1.6722 1.6707 16.0102 144.9873 0.00022269 -85.5323 0.43896
0.543 0.98802 5.5223e-005 3.8182 0.012043 7.1542e-006 0.001154 0.099374 0.00065681 0.10003 0.090226 0 0.040553 0.0389 0 0.86061 0.23374 0.061219 0.0086413 4.1259 0.054146 6.4697e-005 0.83592 0.0051295 0.005867 0.001414 0.98659 0.99147 3.0526e-006 1.221e-005 0.13066 0.87683 0.87983 0.0014117 0.96208 0.54668 0.0019013 0.42509 1.6731 1.6716 16.0102 144.9874 0.00022239 -85.5333 0.43996
0.544 0.98802 5.5223e-005 3.8182 0.012043 7.1674e-006 0.001154 0.099483 0.00065681 0.10013 0.090327 0 0.040544 0.0389 0 0.86066 0.23376 0.061227 0.0086423 4.126 0.054152 6.4704e-005 0.83591 0.0051296 0.0058671 0.0014138 0.98659 0.99147 3.0521e-006 1.2208e-005 0.13066 0.87716 0.88002 0.0014116 0.96231 0.54684 0.0019011 0.4251 1.674 1.6725 16.0101 144.9874 0.0002221 -85.5342 0.44096
0.545 0.98802 5.5223e-005 3.8182 0.012043 7.1806e-006 0.001154 0.099592 0.00065682 0.10024 0.090428 0 0.040536 0.0389 0 0.86071 0.23378 0.061235 0.0086433 4.1261 0.054157 6.4711e-005 0.83591 0.0051298 0.0058673 0.0014136 0.98659 0.99148 3.0516e-006 1.2206e-005 0.13066 0.87749 0.8802 0.0014114 0.96253 0.547 0.001901 0.42512 1.6749 1.6734 16.0101 144.9874 0.0002218 -85.5351 0.44196
0.546 0.98802 5.5222e-005 3.8182 0.012043 7.1937e-006 0.001154 0.099701 0.00065682 0.10035 0.090529 0 0.040528 0.0389 0 0.86076 0.2338 0.061243 0.0086443 4.1262 0.054163 6.4719e-005 0.8359 0.0051299 0.0058674 0.0014133 0.98659 0.99148 3.0511e-006 1.2204e-005 0.13066 0.87782 0.88039 0.0014113 0.96275 0.54715 0.0019008 0.42513 1.6758 1.6743 16.0101 144.9874 0.00022151 -85.536 0.44296
0.547 0.98802 5.5222e-005 3.8182 0.012043 7.2069e-006 0.001154 0.09981 0.00065683 0.10046 0.090629 0 0.040519 0.0389 0 0.86081 0.23383 0.061251 0.0086453 4.1263 0.054169 6.4726e-005 0.8359 0.00513 0.0058675 0.0014131 0.9866 0.99148 3.0506e-006 1.2202e-005 0.13066 0.87815 0.88057 0.0014112 0.96297 0.54731 0.0019007 0.42514 1.6767 1.6752 16.0101 144.9874 0.00022122 -85.5369 0.44396
0.548 0.98802 5.5222e-005 3.8182 0.012043 7.2201e-006 0.001154 0.099919 0.00065683 0.10057 0.09073 0 0.040511 0.0389 0 0.86086 0.23385 0.061259 0.0086463 4.1264 0.054175 6.4734e-005 0.83589 0.0051302 0.0058677 0.0014129 0.9866 0.99148 3.0501e-006 1.22e-005 0.13066 0.87848 0.88076 0.0014111 0.96319 0.54747 0.0019005 0.42515 1.6776 1.6761 16.0101 144.9875 0.00022093 -85.5379 0.44496
0.549 0.98802 5.5222e-005 3.8182 0.012043 7.2332e-006 0.001154 0.10003 0.00065683 0.10068 0.09083 0 0.040503 0.0389 0 0.86091 0.23387 0.061267 0.0086474 4.1265 0.054181 6.4741e-005 0.83588 0.0051303 0.0058678 0.0014127 0.9866 0.99148 3.0496e-006 1.2198e-005 0.13067 0.87881 0.88094 0.001411 0.96341 0.54763 0.0019004 0.42517 1.6784 1.677 16.0101 144.9875 0.00022064 -85.5388 0.44596
0.55 0.98802 5.5222e-005 3.8182 0.012043 7.2464e-006 0.001154 0.10014 0.00065684 0.10079 0.090931 0 0.040495 0.0389 0 0.86096 0.23389 0.061275 0.0086484 4.1266 0.054186 6.4748e-005 0.83588 0.0051304 0.0058679 0.0014125 0.9866 0.99148 3.0491e-006 1.2197e-005 0.13067 0.87914 0.88112 0.0014109 0.96363 0.54778 0.0019003 0.42518 1.6793 1.6778 16.0101 144.9875 0.00022035 -85.5397 0.44696
0.551 0.98802 5.5222e-005 3.8182 0.012043 7.2595e-006 0.001154 0.10024 0.00065684 0.1009 0.091031 0 0.040486 0.0389 0 0.86101 0.23392 0.061283 0.0086494 4.1268 0.054192 6.4756e-005 0.83587 0.0051306 0.005868 0.0014123 0.98661 0.99149 3.0487e-006 1.2195e-005 0.13067 0.87946 0.8813 0.0014108 0.96385 0.54794 0.0019001 0.42519 1.6802 1.6787 16.0101 144.9875 0.00022006 -85.5405 0.44796
0.552 0.98802 5.5222e-005 3.8182 0.012043 7.2727e-006 0.001154 0.10035 0.00065685 0.10101 0.091131 0 0.040478 0.0389 0 0.86106 0.23394 0.061291 0.0086504 4.1269 0.054198 6.4763e-005 0.83587 0.0051307 0.0058682 0.0014121 0.98661 0.99149 3.0482e-006 1.2193e-005 0.13067 0.87979 0.88148 0.0014107 0.96406 0.5481 0.0019 0.42521 1.6811 1.6796 16.0101 144.9875 0.00021978 -85.5414 0.44896
0.553 0.98802 5.5222e-005 3.8182 0.012043 7.2859e-006 0.001154 0.10046 0.00065685 0.10111 0.091231 0 0.04047 0.0389 0 0.86112 0.23396 0.061299 0.0086514 4.127 0.054204 6.477e-005 0.83586 0.0051308 0.0058683 0.0014119 0.98661 0.99149 3.0477e-006 1.2191e-005 0.13067 0.88011 0.88166 0.0014105 0.96427 0.54825 0.0018998 0.42522 1.6819 1.6805 16.0101 144.9876 0.00021949 -85.5423 0.44996
0.554 0.98802 5.5222e-005 3.8182 0.012043 7.299e-006 0.001154 0.10057 0.00065686 0.10122 0.091331 0 0.040461 0.0389 0 0.86117 0.23398 0.061308 0.0086524 4.1271 0.05421 6.4778e-005 0.83586 0.005131 0.0058684 0.0014117 0.98662 0.99149 3.0473e-006 1.2189e-005 0.13067 0.88043 0.88184 0.0014104 0.96449 0.54841 0.0018997 0.42523 1.6828 1.6813 16.0101 144.9876 0.00021921 -85.5432 0.45096
0.555 0.98802 5.5222e-005 3.8182 0.012043 7.3122e-006 0.001154 0.10068 0.00065686 0.10133 0.091431 0 0.040453 0.0389 0 0.86122 0.23401 0.061316 0.0086534 4.1272 0.054216 6.4785e-005 0.83585 0.0051311 0.0058686 0.0014115 0.98662 0.99149 3.0468e-006 1.2187e-005 0.13067 0.88076 0.88202 0.0014103 0.9647 0.54857 0.0018996 0.42525 1.6837 1.6822 16.0101 144.9876 0.00021893 -85.544 0.45196
0.556 0.98802 5.5222e-005 3.8182 0.012043 7.3254e-006 0.001154 0.10079 0.00065687 0.10144 0.091531 0 0.040445 0.0389 0 0.86127 0.23403 0.061324 0.0086544 4.1273 0.054221 6.4793e-005 0.83584 0.0051312 0.0058687 0.0014113 0.98662 0.99149 3.0463e-006 1.2185e-005 0.13067 0.88108 0.8822 0.0014102 0.96491 0.54872 0.0018994 0.42526 1.6845 1.6831 16.01 144.9876 0.00021864 -85.5449 0.45296
0.557 0.98802 5.5222e-005 3.8182 0.012043 7.3385e-006 0.001154 0.10089 0.00065687 0.10155 0.091631 0 0.040437 0.0389 0 0.86132 0.23405 0.061332 0.0086555 4.1274 0.054227 6.48e-005 0.83584 0.0051314 0.0058688 0.0014111 0.98662 0.9915 3.0459e-006 1.2183e-005 0.13067 0.8814 0.88238 0.0014101 0.96511 0.54888 0.0018993 0.42527 1.6854 1.6839 16.01 144.9876 0.00021836 -85.5457 0.45396
0.558 0.98802 5.5222e-005 3.8182 0.012043 7.3517e-006 0.001154 0.101 0.00065688 0.10165 0.091731 0 0.040429 0.0389 0 0.86137 0.23407 0.06134 0.0086565 4.1275 0.054233 6.4808e-005 0.83583 0.0051315 0.005869 0.0014109 0.98663 0.9915 3.0454e-006 1.2182e-005 0.13068 0.88171 0.88255 0.00141 0.96532 0.54904 0.0018991 0.42528 1.6863 1.6848 16.01 144.9876 0.00021808 -85.5466 0.45496
0.559 0.98802 5.5222e-005 3.8182 0.012043 7.3648e-006 0.001154 0.10111 0.00065688 0.10176 0.091831 0 0.04042 0.0389 0 0.86142 0.2341 0.061348 0.0086575 4.1276 0.054239 6.4815e-005 0.83583 0.0051316 0.0058691 0.0014107 0.98663 0.9915 3.0449e-006 1.218e-005 0.13068 0.88203 0.88273 0.0014099 0.96552 0.54919 0.001899 0.4253 1.6871 1.6857 16.01 144.9877 0.00021781 -85.5474 0.45596
0.56 0.98802 5.5222e-005 3.8182 0.012043 7.378e-006 0.001154 0.10122 0.00065689 0.10187 0.09193 0 0.040412 0.0389 0 0.86147 0.23412 0.061356 0.0086585 4.1277 0.054245 6.4823e-005 0.83582 0.0051318 0.0058692 0.0014105 0.98663 0.9915 3.0445e-006 1.2178e-005 0.13068 0.88235 0.8829 0.0014098 0.96573 0.54935 0.0018989 0.42531 1.688 1.6865 16.01 144.9877 0.00021753 -85.5483 0.45696
0.561 0.98802 5.5222e-005 3.8182 0.012043 7.3912e-006 0.001154 0.10133 0.00065689 0.10198 0.09203 0 0.040404 0.0389 0 0.86152 0.23414 0.061364 0.0086595 4.1279 0.054251 6.483e-005 0.83581 0.0051319 0.0058694 0.0014103 0.98663 0.9915 3.044e-006 1.2176e-005 0.13068 0.88266 0.88308 0.0014097 0.96593 0.54951 0.0018987 0.42532 1.6888 1.6874 16.01 144.9877 0.00021725 -85.5491 0.45796
0.562 0.98802 5.5221e-005 3.8182 0.012043 7.4043e-006 0.001154 0.10143 0.0006569 0.10209 0.092129 0 0.040396 0.0389 0 0.86158 0.23416 0.061373 0.0086606 4.128 0.054257 6.4838e-005 0.83581 0.005132 0.0058695 0.0014101 0.98664 0.9915 3.0436e-006 1.2174e-005 0.13068 0.88298 0.88325 0.0014096 0.96613 0.54966 0.0018986 0.42534 1.6897 1.6882 16.01 144.9877 0.00021698 -85.5499 0.45896
0.563 0.98802 5.5221e-005 3.8182 0.012043 7.4175e-006 0.001154 0.10154 0.0006569 0.10219 0.092229 0 0.040388 0.0389 0 0.86163 0.23419 0.061381 0.0086616 4.1281 0.054263 6.4845e-005 0.8358 0.0051322 0.0058696 0.0014099 0.98664 0.99151 3.0432e-006 1.2173e-005 0.13068 0.88329 0.88342 0.0014095 0.96633 0.54982 0.0018985 0.42535 1.6905 1.6891 16.01 144.9877 0.0002167 -85.5507 0.45996
0.564 0.98802 5.5221e-005 3.8182 0.012043 7.4307e-006 0.001154 0.10165 0.0006569 0.1023 0.092328 0 0.04038 0.0389 0 0.86168 0.23421 0.061389 0.0086626 4.1282 0.054268 6.4853e-005 0.8358 0.0051323 0.0058698 0.0014097 0.98664 0.99151 3.0427e-006 1.2171e-005 0.13068 0.88361 0.8836 0.0014094 0.96653 0.54997 0.0018983 0.42536 1.6914 1.6899 16.01 144.9878 0.00021643 -85.5516 0.46096
0.565 0.98802 5.5221e-005 3.8182 0.012043 7.4438e-006 0.001154 0.10176 0.00065691 0.10241 0.092427 0 0.040371 0.0389 0 0.86173 0.23423 0.061397 0.0086636 4.1283 0.054274 6.486e-005 0.83579 0.0051325 0.0058699 0.0014095 0.98664 0.99151 3.0423e-006 1.2169e-005 0.13068 0.88392 0.88377 0.0014093 0.96673 0.55013 0.0018982 0.42538 1.6922 1.6908 16.01 144.9878 0.00021616 -85.5524 0.46196
0.566 0.98802 5.5221e-005 3.8182 0.012043 7.457e-006 0.001154 0.10186 0.00065691 0.10252 0.092526 0 0.040363 0.0389 0 0.86178 0.23426 0.061405 0.0086647 4.1284 0.05428 6.4868e-005 0.83578 0.0051326 0.00587 0.0014093 0.98665 0.99151 3.0419e-006 1.2167e-005 0.13069 0.88423 0.88394 0.0014092 0.96692 0.55029 0.0018981 0.42539 1.693 1.6916 16.0099 144.9878 0.00021589 -85.5532 0.46296
0.567 0.98802 5.5221e-005 3.8182 0.012043 7.4701e-006 0.001154 0.10197 0.00065692 0.10262 0.092625 0 0.040355 0.0389 0 0.86183 0.23428 0.061414 0.0086657 4.1285 0.054286 6.4875e-005 0.83578 0.0051327 0.0058702 0.0014091 0.98665 0.99151 3.0414e-006 1.2166e-005 0.13069 0.88454 0.88411 0.0014091 0.96712 0.55044 0.0018979 0.4254 1.6939 1.6925 16.0099 144.9878 0.00021562 -85.554 0.46396
0.568 0.98802 5.5221e-005 3.8182 0.012042 7.4833e-006 0.001154 0.10208 0.00065692 0.10273 0.092724 0 0.040347 0.0389 0 0.86189 0.2343 0.061422 0.0086667 4.1286 0.054292 6.4883e-005 0.83577 0.0051329 0.0058703 0.0014089 0.98665 0.99151 3.041e-006 1.2164e-005 0.13069 0.88485 0.88428 0.001409 0.96731 0.5506 0.0018978 0.42542 1.6947 1.6933 16.0099 144.9878 0.00021535 -85.5547 0.46496
0.569 0.98802 5.5221e-005 3.8182 0.012042 7.4965e-006 0.001154 0.10218 0.00065693 0.10284 0.092823 0 0.040339 0.0389 0 0.86194 0.23432 0.06143 0.0086678 4.1288 0.054298 6.489e-005 0.83577 0.005133 0.0058705 0.0014088 0.98665 0.99152 3.0406e-006 1.2162e-005 0.13069 0.88516 0.88445 0.0014089 0.96751 0.55075 0.0018977 0.42543 1.6956 1.6942 16.0099 144.9879 0.00021508 -85.5555 0.46596
0.57 0.98802 5.5221e-005 3.8182 0.012042 7.5096e-006 0.001154 0.10229 0.00065693 0.10294 0.092922 0 0.040331 0.0389 0 0.86199 0.23435 0.061438 0.0086688 4.1289 0.054304 6.4898e-005 0.83576 0.0051331 0.0058706 0.0014086 0.98666 0.99152 3.0402e-006 1.2161e-005 0.13069 0.88546 0.88462 0.0014088 0.9677 0.55091 0.0018976 0.42544 1.6964 1.695 16.0099 144.9879 0.00021482 -85.5563 0.46696
0.571 0.98802 5.5221e-005 3.8182 0.012042 7.5228e-006 0.001154 0.1024 0.00065694 0.10305 0.093021 0 0.040323 0.0389 0 0.86204 0.23437 0.061447 0.0086698 4.129 0.05431 6.4906e-005 0.83575 0.0051333 0.0058707 0.0014084 0.98666 0.99152 3.0398e-006 1.2159e-005 0.13069 0.88577 0.88478 0.0014087 0.96789 0.55107 0.0018974 0.42545 1.6972 1.6958 16.0099 144.9879 0.00021455 -85.5571 0.46796
0.572 0.98802 5.5221e-005 3.8182 0.012042 7.536e-006 0.001154 0.1025 0.00065694 0.10316 0.09312 0 0.040315 0.0389 0 0.86209 0.23439 0.061455 0.0086709 4.1291 0.054316 6.4913e-005 0.83575 0.0051334 0.0058709 0.0014082 0.98666 0.99152 3.0393e-006 1.2157e-005 0.13069 0.88607 0.88495 0.0014086 0.96808 0.55122 0.0018973 0.42547 1.698 1.6967 16.0099 144.9879 0.00021429 -85.5579 0.46896
0.573 0.98802 5.5221e-005 3.8182 0.012042 7.5491e-006 0.001154 0.10261 0.00065694 0.10326 0.093218 0 0.040307 0.0389 0 0.86215 0.23442 0.061463 0.0086719 4.1292 0.054322 6.4921e-005 0.83574 0.0051336 0.005871 0.001408 0.98666 0.99152 3.0389e-006 1.2156e-005 0.13069 0.88638 0.88512 0.0014085 0.96826 0.55138 0.0018972 0.42548 1.6989 1.6975 16.0099 144.9879 0.00021402 -85.5586 0.46996
0.574 0.98802 5.5221e-005 3.8182 0.012042 7.5623e-006 0.001154 0.10272 0.00065695 0.10337 0.093317 0 0.040299 0.0389 0 0.8622 0.23444 0.061471 0.0086729 4.1293 0.054328 6.4929e-005 0.83574 0.0051337 0.0058711 0.0014079 0.98666 0.99152 3.0385e-006 1.2154e-005 0.13069 0.88668 0.88528 0.0014084 0.96845 0.55153 0.0018971 0.42549 1.6997 1.6983 16.0099 144.988 0.00021376 -85.5594 0.47096
0.575 0.98802 5.5221e-005 3.8182 0.012042 7.5754e-006 0.001154 0.10282 0.00065695 0.10348 0.093415 0 0.040291 0.0389 0 0.86225 0.23446 0.06148 0.008674 4.1295 0.054334 6.4936e-005 0.83573 0.0051338 0.0058713 0.0014077 0.98667 0.99152 3.0381e-006 1.2152e-005 0.1307 0.88698 0.88545 0.0014083 0.96863 0.55169 0.001897 0.42551 1.7005 1.6991 16.0098 144.988 0.0002135 -85.5601 0.47196
0.576 0.98802 5.5221e-005 3.8182 0.012042 7.5886e-006 0.001154 0.10293 0.00065696 0.10358 0.093514 0 0.040283 0.0389 0 0.8623 0.23448 0.061488 0.008675 4.1296 0.05434 6.4944e-005 0.83572 0.005134 0.0058714 0.0014075 0.98667 0.99153 3.0377e-006 1.2151e-005 0.1307 0.88728 0.88561 0.0014083 0.96882 0.55184 0.0018968 0.42552 1.7013 1.7 16.0098 144.988 0.00021324 -85.5609 0.47296
0.577 0.98802 5.5221e-005 3.8182 0.012042 7.6018e-006 0.001154 0.10304 0.00065696 0.10369 0.093612 0 0.040275 0.0389 0 0.86235 0.23451 0.061496 0.0086761 4.1297 0.054346 6.4952e-005 0.83572 0.0051341 0.0058716 0.0014073 0.98667 0.99153 3.0373e-006 1.2149e-005 0.1307 0.88758 0.88578 0.0014082 0.969 0.552 0.0018967 0.42553 1.7022 1.7008 16.0098 144.988 0.00021298 -85.5616 0.47396
0.578 0.98802 5.5221e-005 3.8182 0.012042 7.6149e-006 0.001154 0.10314 0.00065697 0.1038 0.09371 0 0.040267 0.0389 0 0.86241 0.23453 0.061505 0.0086771 4.1298 0.054352 6.4959e-005 0.83571 0.0051343 0.0058717 0.0014071 0.98667 0.99153 3.0369e-006 1.2148e-005 0.1307 0.88788 0.88594 0.0014081 0.96918 0.55216 0.0018966 0.42555 1.703 1.7016 16.0098 144.988 0.00021272 -85.5624 0.47496
0.579 0.98802 5.522e-005 3.8182 0.012042 7.6281e-006 0.001154 0.10325 0.00065697 0.1039 0.093808 0 0.040259 0.0389 0 0.86246 0.23455 0.061513 0.0086781 4.1299 0.054358 6.4967e-005 0.83571 0.0051344 0.0058718 0.001407 0.98668 0.99153 3.0365e-006 1.2146e-005 0.1307 0.88818 0.8861 0.001408 0.96936 0.55231 0.0018965 0.42556 1.7038 1.7024 16.0098 144.9881 0.00021247 -85.5631 0.47596
0.58 0.98802 5.522e-005 3.8182 0.012042 7.6413e-006 0.001154 0.10336 0.00065698 0.10401 0.093907 0 0.040251 0.0389 0 0.86251 0.23458 0.061521 0.0086792 4.13 0.054364 6.4975e-005 0.8357 0.0051346 0.005872 0.0014068 0.98668 0.99153 3.0361e-006 1.2144e-005 0.1307 0.88848 0.88626 0.0014079 0.96954 0.55247 0.0018964 0.42557 1.7046 1.7032 16.0098 144.9881 0.00021221 -85.5638 0.47696
0.581 0.98802 5.522e-005 3.8182 0.012042 7.6544e-006 0.001154 0.10346 0.00065698 0.10411 0.094005 0 0.040243 0.0389 0 0.86256 0.2346 0.06153 0.0086802 4.1302 0.05437 6.4982e-005 0.83569 0.0051347 0.0058721 0.0014066 0.98668 0.99153 3.0357e-006 1.2143e-005 0.1307 0.88878 0.88643 0.0014078 0.96972 0.55262 0.0018962 0.42559 1.7054 1.7041 16.0098 144.9881 0.00021196 -85.5646 0.47796
0.582 0.98802 5.522e-005 3.8182 0.012042 7.6676e-006 0.001154 0.10357 0.00065698 0.10422 0.094102 0 0.040235 0.0389 0 0.86262 0.23462 0.061538 0.0086813 4.1303 0.054376 6.499e-005 0.83569 0.0051348 0.0058723 0.0014065 0.98668 0.99153 3.0353e-006 1.2141e-005 0.1307 0.88907 0.88659 0.0014077 0.9699 0.55278 0.0018961 0.4256 1.7062 1.7049 16.0098 144.9881 0.0002117 -85.5653 0.47896
0.583 0.98802 5.522e-005 3.8182 0.012042 7.6807e-006 0.001154 0.10367 0.00065699 0.10433 0.0942 0 0.040227 0.0389 0 0.86267 0.23465 0.061546 0.0086823 4.1304 0.054382 6.4998e-005 0.83568 0.005135 0.0058724 0.0014063 0.98669 0.99154 3.035e-006 1.214e-005 0.1307 0.88937 0.88675 0.0014076 0.97007 0.55293 0.001896 0.42561 1.707 1.7057 16.0098 144.9881 0.00021145 -85.566 0.47996
0.584 0.98802 5.522e-005 3.8182 0.012042 7.6939e-006 0.001154 0.10378 0.00065699 0.10443 0.094298 0 0.040219 0.0389 0 0.86272 0.23467 0.061555 0.0086834 4.1305 0.054389 6.5005e-005 0.83568 0.0051351 0.0058726 0.0014062 0.98669 0.99154 3.0346e-006 1.2138e-005 0.13071 0.88966 0.88691 0.0014075 0.97025 0.55309 0.0018959 0.42563 1.7078 1.7065 16.0097 144.9882 0.0002112 -85.5667 0.48096
0.585 0.98802 5.522e-005 3.8182 0.012042 7.7071e-006 0.001154 0.10389 0.000657 0.10454 0.094396 0 0.040211 0.0389 0 0.86277 0.23469 0.061563 0.0086844 4.1306 0.054395 6.5013e-005 0.83567 0.0051353 0.0058727 0.001406 0.98669 0.99154 3.0342e-006 1.2137e-005 0.13071 0.88995 0.88706 0.0014075 0.97042 0.55324 0.0018958 0.42564 1.7086 1.7073 16.0097 144.9882 0.00021094 -85.5674 0.48196
0.586 0.98802 5.522e-005 3.8182 0.012042 7.7202e-006 0.001154 0.10399 0.000657 0.10464 0.094494 0 0.040203 0.0389 0 0.86283 0.23472 0.061572 0.0086855 4.1308 0.054401 6.5021e-005 0.83566 0.0051354 0.0058728 0.0014058 0.98669 0.99154 3.0338e-006 1.2135e-005 0.13071 0.89025 0.88722 0.0014074 0.9706 0.5534 0.0018957 0.42565 1.7094 1.7081 16.0097 144.9882 0.00021069 -85.5681 0.48296
0.587 0.98802 5.522e-005 3.8182 0.012042 7.7334e-006 0.001154 0.1041 0.00065701 0.10475 0.094591 0 0.040195 0.0389 0 0.86288 0.23474 0.06158 0.0086865 4.1309 0.054407 6.5029e-005 0.83566 0.0051356 0.005873 0.0014056 0.98669 0.99154 3.0335e-006 1.2134e-005 0.13071 0.89054 0.88738 0.0014073 0.97077 0.55355 0.0018956 0.42566 1.7102 1.7089 16.0097 144.9882 0.00021045 -85.5688 0.48396
0.588 0.98802 5.522e-005 3.8182 0.012042 7.7466e-006 0.001154 0.1042 0.00065701 0.10485 0.094689 0 0.040187 0.0389 0 0.86293 0.23476 0.061588 0.0086876 4.131 0.054413 6.5037e-005 0.83565 0.0051357 0.0058731 0.0014054 0.9867 0.99154 3.0331e-006 1.2132e-005 0.13071 0.89083 0.88754 0.0014072 0.97094 0.55371 0.0018954 0.42568 1.711 1.7097 16.0097 144.9882 0.0002102 -85.5695 0.48496
0.589 0.98802 5.522e-005 3.8182 0.012042 7.7597e-006 0.001154 0.10431 0.00065701 0.10496 0.094786 0 0.040179 0.0389 0 0.86299 0.23479 0.061597 0.0086887 4.1311 0.054419 6.5044e-005 0.83565 0.0051359 0.0058733 0.0014053 0.9867 0.99154 3.0327e-006 1.2131e-005 0.13071 0.89112 0.88769 0.0014071 0.97111 0.55386 0.0018953 0.42569 1.7118 1.7105 16.0097 144.9883 0.00020995 -85.5702 0.48596
0.59 0.98802 5.522e-005 3.8182 0.012042 7.7729e-006 0.001154 0.10441 0.00065702 0.10506 0.094883 0 0.040171 0.0389 0 0.86304 0.23481 0.061605 0.0086897 4.1312 0.054425 6.5052e-005 0.83564 0.005136 0.0058734 0.0014051 0.9867 0.99155 3.0324e-006 1.2129e-005 0.13071 0.89141 0.88785 0.001407 0.97128 0.55402 0.0018952 0.4257 1.7126 1.7113 16.0097 144.9883 0.0002097 -85.5709 0.48696
0.591 0.98802 5.522e-005 3.8182 0.012042 7.786e-006 0.001154 0.10452 0.00065702 0.10517 0.094981 0 0.040163 0.0389 0 0.86309 0.23483 0.061614 0.0086908 4.1314 0.054431 6.506e-005 0.83563 0.0051362 0.0058736 0.001405 0.9867 0.99155 3.032e-006 1.2128e-005 0.13071 0.89169 0.88801 0.0014069 0.97144 0.55417 0.0018951 0.42572 1.7134 1.7121 16.0097 144.9883 0.00020946 -85.5715 0.48796
0.592 0.98802 5.522e-005 3.8182 0.012042 7.7992e-006 0.001154 0.10462 0.00065703 0.10527 0.095078 0 0.040155 0.0389 0 0.86315 0.23486 0.061622 0.0086918 4.1315 0.054438 6.5068e-005 0.83563 0.0051363 0.0058737 0.0014049 0.9867 0.99155 3.0316e-006 1.2126e-005 0.13072 0.89198 0.88816 0.0014069 0.97161 0.55433 0.001895 0.42573 1.7142 1.7129 16.0096 144.9883 0.00020921 -85.5722 0.48896
0.593 0.98802 5.522e-005 3.8182 0.012042 7.8124e-006 0.001154 0.10473 0.00065703 0.10538 0.095175 0 0.040147 0.0389 0 0.8632 0.23488 0.061631 0.0086929 4.1316 0.054444 6.5076e-005 0.83562 0.0051365 0.0058739 0.0014047 0.98671 0.99155 3.0312e-006 1.2125e-005 0.13072 0.89227 0.88831 0.0014068 0.97177 0.55448 0.0018949 0.42574 1.715 1.7137 16.0096 144.9883 0.00020897 -85.5729 0.48996
0.594 0.98802 5.522e-005 3.8182 0.012042 7.8255e-006 0.001154 0.10483 0.00065704 0.10548 0.095272 0 0.04014 0.0389 0 0.86325 0.2349 0.061639 0.0086939 4.1317 0.05445 6.5083e-005 0.83562 0.0051366 0.005874 0.0014046 0.98671 0.99155 3.0309e-006 1.2124e-005 0.13072 0.89255 0.88847 0.0014067 0.97194 0.55464 0.0018948 0.42576 1.7157 1.7144 16.0096 144.9884 0.00020873 -85.5735 0.49096
0.595 0.98802 5.5219e-005 3.8182 0.012042 7.8387e-006 0.001154 0.10494 0.00065704 0.10559 0.095369 0 0.040132 0.0389 0 0.86331 0.23493 0.061648 0.008695 4.1319 0.054456 6.5091e-005 0.83561 0.0051367 0.0058741 0.0014044 0.98671 0.99155 3.0305e-006 1.2122e-005 0.13072 0.89283 0.88862 0.0014066 0.9721 0.55479 0.0018947 0.42577 1.7165 1.7152 16.0096 144.9884 0.00020849 -85.5742 0.49196
0.596 0.98802 5.5219e-005 3.8182 0.012042 7.8518e-006 0.001154 0.10504 0.00065704 0.10569 0.095466 0 0.040124 0.0389 0 0.86336 0.23495 0.061656 0.0086961 4.132 0.054462 6.5099e-005 0.8356 0.0051369 0.0058743 0.0014042 0.98671 0.99155 3.0302e-006 1.2121e-005 0.13072 0.89312 0.88877 0.0014065 0.97226 0.55495 0.0018946 0.42578 1.7173 1.716 16.0096 144.9884 0.00020825 -85.5748 0.49296
0.597 0.98802 5.5219e-005 3.8182 0.012042 7.865e-006 0.001154 0.10515 0.00065705 0.1058 0.095563 0 0.040116 0.0389 0 0.86341 0.23497 0.061665 0.0086971 4.1321 0.054468 6.5107e-005 0.8356 0.005137 0.0058744 0.001404 0.98671 0.99155 3.0299e-006 1.2119e-005 0.13072 0.8934 0.88893 0.0014064 0.97242 0.5551 0.0018945 0.4258 1.7181 1.7168 16.0096 144.9884 0.00020801 -85.5755 0.49396
0.598 0.98802 5.5219e-005 3.8182 0.012042 7.8782e-006 0.001154 0.10525 0.00065705 0.1059 0.095659 0 0.040108 0.0389 0 0.86347 0.235 0.061673 0.0086982 4.1322 0.054475 6.5115e-005 0.83559 0.0051372 0.0058746 0.0014038 0.98672 0.99156 3.0296e-006 1.2118e-005 0.13072 0.89368 0.88908 0.0014063 0.97258 0.55525 0.0018944 0.42581 1.7189 1.7176 16.0096 144.9884 0.00020777 -85.5761 0.49496
0.599 0.98802 5.5219e-005 3.8182 0.012042 7.8913e-006 0.001154 0.10536 0.00065706 0.10601 0.095756 0 0.0401 0.0389 0 0.86352 0.23502 0.061682 0.0086993 4.1324 0.054481 6.5123e-005 0.83558 0.0051373 0.0058747 0.0014037 0.98672 0.99156 3.0292e-006 1.2117e-005 0.13072 0.89396 0.88923 0.0014062 0.97274 0.55541 0.0018943 0.42582 1.7196 1.7183 16.0096 144.9885 0.00020753 -85.5768 0.49596
0.6 0.98802 5.5219e-005 3.8182 0.012042 7.9045e-006 0.001154 0.10546 0.00065706 0.10611 0.095853 0 0.040093 0.0389 0 0.86357 0.23505 0.06169 0.0087003 4.1325 0.054487 6.5131e-005 0.83558 0.0051375 0.0058749 0.0014036 0.98672 0.99156 3.0289e-006 1.2115e-005 0.13073 0.89424 0.88938 0.0014062 0.9729 0.55556 0.0018942 0.42584 1.7204 1.7191 16.0095 144.9885 0.00020729 -85.5774 0.49696
0.601 0.98802 5.5219e-005 3.8182 0.012042 7.9177e-006 0.001154 0.10556 0.00065706 0.10622 0.095949 0 0.040085 0.0389 0 0.86363 0.23507 0.061699 0.0087014 4.1326 0.054493 6.5139e-005 0.83557 0.0051376 0.005875 0.0014035 0.98672 0.99156 3.0285e-006 1.2114e-005 0.13073 0.89452 0.88953 0.0014061 0.97306 0.55572 0.0018941 0.42585 1.7212 1.7199 16.0095 144.9885 0.00020706 -85.578 0.49796
0.602 0.98802 5.5219e-005 3.8182 0.012042 7.9308e-006 0.001154 0.10567 0.00065707 0.10632 0.096046 0 0.040077 0.0389 0 0.86368 0.23509 0.061707 0.0087025 4.1327 0.054499 6.5147e-005 0.83557 0.0051378 0.0058752 0.0014034 0.98672 0.99156 3.0281e-006 1.2112e-005 0.13073 0.8948 0.88968 0.0014061 0.97321 0.55587 0.001894 0.42586 1.7219 1.7207 16.0095 144.9885 0.00020682 -85.5787 0.49896
0.603 0.98802 5.5219e-005 3.8182 0.012042 7.944e-006 0.001154 0.10577 0.00065707 0.10643 0.096142 0 0.040069 0.0389 0 0.86373 0.23512 0.061716 0.0087035 4.1329 0.054506 6.5155e-005 0.83556 0.005138 0.0058753 0.0014034 0.98673 0.99156 3.0278e-006 1.2111e-005 0.13073 0.89507 0.88982 0.0014061 0.97337 0.55603 0.0018939 0.42588 1.7227 1.7214 16.0095 144.9885 0.00020659 -85.5793 0.49996
0.604 0.98802 5.5219e-005 3.8182 0.012042 7.9571e-006 0.001154 0.10588 0.00065708 0.10653 0.096238 0 0.040061 0.0389 0 0.86379 0.23514 0.061725 0.0087046 4.133 0.054512 6.5162e-005 0.83555 0.0051381 0.0058755 0.0014032 0.98673 0.99156 3.0274e-006 1.211e-005 0.13073 0.89535 0.88997 0.001406 0.97352 0.55618 0.0018938 0.42589 1.7235 1.7222 16.0095 144.9886 0.00020635 -85.5799 0.50096
0.605 0.98802 5.5219e-005 3.8182 0.012042 7.9703e-006 0.001154 0.10598 0.00065708 0.10663 0.096334 0 0.040054 0.0389 0 0.86384 0.23516 0.061733 0.0087057 4.1331 0.054518 6.517e-005 0.83555 0.0051383 0.0058756 0.0014031 0.98673 0.99156 3.0271e-006 1.2108e-005 0.13073 0.89563 0.89012 0.001406 0.97367 0.55633 0.0018937 0.4259 1.7242 1.723 16.0095 144.9886 0.00020612 -85.5805 0.50196
0.606 0.98802 5.5219e-005 3.8182 0.012042 7.9835e-006 0.001154 0.10608 0.00065708 0.10674 0.096431 0 0.040046 0.0389 0 0.8639 0.23519 0.061742 0.0087068 4.1332 0.054524 6.5178e-005 0.83554 0.0051384 0.0058758 0.0014029 0.98673 0.99157 3.0268e-006 1.2107e-005 0.13073 0.8959 0.89027 0.0014059 0.97383 0.55649 0.0018936 0.42591 1.725 1.7237 16.0095 144.9886 0.00020589 -85.5811 0.50296
0.607 0.98802 5.5219e-005 3.8182 0.012042 7.9966e-006 0.001154 0.10619 0.00065709 0.10684 0.096527 0 0.040038 0.0389 0 0.86395 0.23521 0.06175 0.0087078 4.1334 0.054531 6.5186e-005 0.83553 0.0051386 0.0058759 0.0014028 0.98673 0.99157 3.0265e-006 1.2106e-005 0.13073 0.89617 0.89041 0.0014058 0.97398 0.55664 0.0018935 0.42593 1.7257 1.7245 16.0094 144.9886 0.00020566 -85.5818 0.50396
0.608 0.98802 5.5219e-005 3.8182 0.012042 8.0098e-006 0.001154 0.10629 0.00065709 0.10694 0.096623 0 0.04003 0.0389 0 0.864 0.23524 0.061759 0.0087089 4.1335 0.054537 6.5194e-005 0.83553 0.0051387 0.0058761 0.0014026 0.98673 0.99157 3.0262e-006 1.2105e-005 0.13074 0.89645 0.89056 0.0014057 0.97413 0.5568 0.0018934 0.42594 1.7265 1.7252 16.0094 144.9886 0.00020543 -85.5824 0.50496
0.609 0.98802 5.5219e-005 3.8182 0.012042 8.0229e-006 0.001154 0.1064 0.0006571 0.10705 0.096719 0 0.040023 0.0389 0 0.86406 0.23526 0.061768 0.00871 4.1336 0.054543 6.5202e-005 0.83552 0.0051389 0.0058762 0.0014024 0.98674 0.99157 3.0258e-006 1.2103e-005 0.13074 0.89672 0.8907 0.0014056 0.97428 0.55695 0.0018933 0.42595 1.7272 1.726 16.0094 144.9887 0.0002052 -85.583 0.50596
0.61 0.98802 5.5219e-005 3.8182 0.012042 8.0361e-006 0.001154 0.1065 0.0006571 0.10715 0.096814 0 0.040015 0.0389 0 0.86411 0.23528 0.061776 0.0087111 4.1338 0.05455 6.521e-005 0.83552 0.005139 0.0058764 0.0014022 0.98674 0.99157 3.0255e-006 1.2102e-005 0.13074 0.89699 0.89085 0.0014055 0.97442 0.5571 0.0018932 0.42597 1.728 1.7268 16.0094 144.9887 0.00020497 -85.5835 0.50696
0.611 0.98802 5.5218e-005 3.8182 0.012042 8.0493e-006 0.001154 0.1066 0.0006571 0.10726 0.09691 0 0.040007 0.0389 0 0.86417 0.23531 0.061785 0.0087122 4.1339 0.054556 6.5218e-005 0.83551 0.0051392 0.0058766 0.0014021 0.98674 0.99157 3.0252e-006 1.2101e-005 0.13074 0.89726 0.89099 0.0014054 0.97457 0.55726 0.0018931 0.42598 1.7287 1.7275 16.0094 144.9887 0.00020475 -85.5841 0.50796
0.612 0.98802 5.5218e-005 3.8182 0.012042 8.0624e-006 0.001154 0.10671 0.00065711 0.10736 0.097006 0 0.04 0.0389 0 0.86422 0.23533 0.061793 0.0087132 4.134 0.054562 6.5226e-005 0.8355 0.0051393 0.0058767 0.0014019 0.98674 0.99157 3.0249e-006 1.21e-005 0.13074 0.89753 0.89113 0.0014053 0.97472 0.55741 0.001893 0.42599 1.7295 1.7283 16.0094 144.9887 0.00020452 -85.5847 0.50896
0.613 0.98802 5.5218e-005 3.8182 0.012042 8.0756e-006 0.001154 0.10681 0.00065711 0.10746 0.097101 0 0.039992 0.0389 0 0.86428 0.23536 0.061802 0.0087143 4.1341 0.054568 6.5234e-005 0.8355 0.0051395 0.0058769 0.0014017 0.98674 0.99157 3.0246e-006 1.2098e-005 0.13074 0.8978 0.89128 0.0014052 0.97486 0.55757 0.0018929 0.42601 1.7302 1.729 16.0094 144.9887 0.00020429 -85.5853 0.50996
0.614 0.98802 5.5218e-005 3.8182 0.012042 8.0887e-006 0.001154 0.10691 0.00065712 0.10757 0.097197 0 0.039984 0.0389 0 0.86433 0.23538 0.061811 0.0087154 4.1343 0.054575 6.5243e-005 0.83549 0.0051396 0.005877 0.0014016 0.98675 0.99158 3.0243e-006 1.2097e-005 0.13074 0.89806 0.89142 0.0014051 0.97501 0.55772 0.0018928 0.42602 1.731 1.7298 16.0093 144.9888 0.00020407 -85.5859 0.51096
0.615 0.98802 5.5218e-005 3.8182 0.012042 8.1019e-006 0.001154 0.10702 0.00065712 0.10767 0.097292 0 0.039976 0.0389 0 0.86438 0.2354 0.061819 0.0087165 4.1344 0.054581 6.5251e-005 0.83548 0.0051398 0.0058772 0.0014014 0.98675 0.99158 3.024e-006 1.2096e-005 0.13075 0.89833 0.89156 0.0014051 0.97515 0.55787 0.0018927 0.42603 1.7317 1.7305 16.0093 144.9888 0.00020385 -85.5865 0.51196
0.616 0.98802 5.5218e-005 3.8182 0.012042 8.1151e-006 0.001154 0.10712 0.00065712 0.10777 0.097388 0 0.039969 0.0389 0 0.86444 0.23543 0.061828 0.0087176 4.1345 0.054587 6.5259e-005 0.83548 0.00514 0.0058773 0.0014013 0.98675 0.99158 3.0237e-006 1.2095e-005 0.13075 0.8986 0.8917 0.001405 0.97529 0.55803 0.0018926 0.42605 1.7325 1.7312 16.0093 144.9888 0.00020362 -85.587 0.51296
0.617 0.98802 5.5218e-005 3.8182 0.012042 8.1282e-006 0.001154 0.10722 0.00065713 0.10787 0.097483 0 0.039961 0.0389 0 0.86449 0.23545 0.061837 0.0087187 4.1347 0.054594 6.5267e-005 0.83547 0.0051401 0.0058775 0.0014012 0.98675 0.99158 3.0234e-006 1.2094e-005 0.13075 0.89886 0.89184 0.0014049 0.97543 0.55818 0.0018925 0.42606 1.7332 1.732 16.0093 144.9888 0.0002034 -85.5876 0.51396
0.618 0.98802 5.5218e-005 3.8182 0.012042 8.1414e-006 0.001154 0.10732 0.00065713 0.10798 0.097578 0 0.039953 0.0389 0 0.86455 0.23548 0.061846 0.0087198 4.1348 0.0546 6.5275e-005 0.83547 0.0051403 0.0058776 0.0014011 0.98675 0.99158 3.0231e-006 1.2092e-005 0.13075 0.89913 0.89198 0.0014049 0.97557 0.55833 0.0018924 0.42607 1.7339 1.7327 16.0093 144.9888 0.00020318 -85.5882 0.51496
0.619 0.98802 5.5218e-005 3.8182 0.012042 8.1545e-006 0.001154 0.10743 0.00065714 0.10808 0.097674 0 0.039946 0.0389 0 0.8646 0.2355 0.061854 0.0087208 4.1349 0.054606 6.5283e-005 0.83546 0.0051404 0.0058778 0.001401 0.98675 0.99158 3.0228e-006 1.2091e-005 0.13075 0.89939 0.89212 0.0014048 0.97571 0.55849 0.0018924 0.42609 1.7347 1.7335 16.0093 144.9889 0.00020296 -85.5887 0.51596
0.62 0.98802 5.5218e-005 3.8182 0.012042 8.1677e-006 0.001154 0.10753 0.00065714 0.10818 0.097769 0 0.039938 0.0389 0 0.86466 0.23552 0.061863 0.0087219 4.1351 0.054613 6.5291e-005 0.83545 0.0051406 0.0058779 0.0014008 0.98676 0.99158 3.0225e-006 1.209e-005 0.13075 0.89965 0.89226 0.0014047 0.97585 0.55864 0.0018923 0.4261 1.7354 1.7342 16.0093 144.9889 0.00020274 -85.5893 0.51696
0.621 0.98802 5.5218e-005 3.8182 0.012042 8.1809e-006 0.001154 0.10763 0.00065714 0.10829 0.097864 0 0.039931 0.0389 0 0.86471 0.23555 0.061872 0.008723 4.1352 0.054619 6.5299e-005 0.83545 0.0051407 0.0058781 0.0014007 0.98676 0.99158 3.0222e-006 1.2089e-005 0.13075 0.89992 0.8924 0.0014047 0.97599 0.55879 0.0018922 0.42611 1.7361 1.7349 16.0092 144.9889 0.00020252 -85.5898 0.51796
0.622 0.98802 5.5218e-005 3.8182 0.012042 8.194e-006 0.001154 0.10774 0.00065715 0.10839 0.097959 0 0.039923 0.0389 0 0.86477 0.23557 0.06188 0.0087241 4.1353 0.054626 6.5307e-005 0.83544 0.0051409 0.0058783 0.0014006 0.98676 0.99158 3.0219e-006 1.2088e-005 0.13075 0.90018 0.89254 0.0014046 0.97613 0.55895 0.0018921 0.42613 1.7369 1.7357 16.0092 144.9889 0.0002023 -85.5904 0.51896
0.623 0.98802 5.5218e-005 3.8182 0.012042 8.2072e-006 0.001154 0.10784 0.00065715 0.10849 0.098054 0 0.039915 0.0389 0 0.86482 0.2356 0.061889 0.0087252 4.1355 0.054632 6.5315e-005 0.83543 0.0051411 0.0058784 0.0014005 0.98676 0.99159 3.0216e-006 1.2086e-005 0.13076 0.90044 0.89268 0.0014046 0.97626 0.5591 0.001892 0.42614 1.7376 1.7364 16.0092 144.9889 0.00020209 -85.5909 0.51996
0.624 0.98802 5.5218e-005 3.8182 0.012042 8.2203e-006 0.001154 0.10794 0.00065715 0.10859 0.098148 0 0.039908 0.0389 0 0.86488 0.23562 0.061898 0.0087263 4.1356 0.054638 6.5324e-005 0.83543 0.0051412 0.0058786 0.0014004 0.98676 0.99159 3.0213e-006 1.2085e-005 0.13076 0.9007 0.89281 0.0014045 0.9764 0.55925 0.0018919 0.42615 1.7383 1.7371 16.0092 144.989 0.00020187 -85.5915 0.52096
0.625 0.98802 5.5218e-005 3.8182 0.012042 8.2335e-006 0.001154 0.10804 0.00065716 0.1087 0.098243 0 0.0399 0.0389 0 0.86493 0.23565 0.061907 0.0087274 4.1357 0.054645 6.5332e-005 0.83542 0.0051414 0.0058787 0.0014002 0.98676 0.99159 3.021e-006 1.2084e-005 0.13076 0.90095 0.89295 0.0014044 0.97653 0.55941 0.0018918 0.42617 1.739 1.7379 16.0092 144.989 0.00020166 -85.592 0.52196
0.626 0.98802 5.5218e-005 3.8182 0.012042 8.2467e-006 0.001154 0.10815 0.00065716 0.1088 0.098338 0 0.039893 0.0389 0 0.86499 0.23567 0.061915 0.0087285 4.1359 0.054651 6.534e-005 0.83541 0.0051415 0.0058789 0.0014001 0.98677 0.99159 3.0207e-006 1.2083e-005 0.13076 0.90121 0.89309 0.0014044 0.97667 0.55956 0.0018917 0.42618 1.7398 1.7386 16.0092 144.989 0.00020144 -85.5925 0.52296
0.627 0.98802 5.5217e-005 3.8182 0.012042 8.2598e-006 0.001154 0.10825 0.00065717 0.1089 0.098432 0 0.039885 0.0389 0 0.86504 0.23569 0.061924 0.0087296 4.136 0.054658 6.5348e-005 0.83541 0.0051417 0.0058791 0.0014 0.98677 0.99159 3.0205e-006 1.2082e-005 0.13076 0.90147 0.89322 0.0014043 0.9768 0.55971 0.0018917 0.42619 1.7405 1.7393 16.0092 144.989 0.00020123 -85.5931 0.52396
0.628 0.98802 5.5217e-005 3.8182 0.012042 8.273e-006 0.001154 0.10835 0.00065717 0.109 0.098527 0 0.039877 0.0389 0 0.8651 0.23572 0.061933 0.0087307 4.1361 0.054664 6.5356e-005 0.8354 0.0051419 0.0058792 0.0013998 0.98677 0.99159 3.0202e-006 1.2081e-005 0.13076 0.90173 0.89336 0.0014042 0.97693 0.55987 0.0018916 0.4262 1.7412 1.74 16.0091 144.989 0.00020102 -85.5936 0.52496
0.629 0.98802 5.5217e-005 3.8182 0.012042 8.2861e-006 0.001154 0.10845 0.00065717 0.1091 0.098621 0 0.03987 0.0389 0 0.86515 0.23574 0.061942 0.0087318 4.1363 0.05467 6.5364e-005 0.83539 0.005142 0.0058794 0.0013997 0.98677 0.99159 3.0199e-006 1.208e-005 0.13076 0.90198 0.89349 0.0014042 0.97706 0.56002 0.0018915 0.42622 1.7419 1.7407 16.0091 144.9891 0.0002008 -85.5941 0.52596
0.63 0.98802 5.5217e-005 3.8182 0.012042 8.2993e-006 0.001154 0.10855 0.00065718 0.10921 0.098716 0 0.039862 0.0389 0 0.86521 0.23577 0.061951 0.0087329 4.1364 0.054677 6.5373e-005 0.83539 0.0051422 0.0058795 0.0013996 0.98677 0.99159 3.0196e-006 1.2078e-005 0.13076 0.90224 0.89363 0.0014041 0.97719 0.56017 0.0018914 0.42623 1.7426 1.7415 16.0091 144.9891 0.00020059 -85.5946 0.52696
0.631 0.98802 5.5217e-005 3.8182 0.012042 8.3125e-006 0.001154 0.10866 0.00065718 0.10931 0.09881 0 0.039855 0.0389 0 0.86527 0.23579 0.06196 0.008734 4.1365 0.054683 6.5381e-005 0.83538 0.0051424 0.0058797 0.0013995 0.98677 0.99159 3.0193e-006 1.2077e-005 0.13077 0.90249 0.89376 0.001404 0.97732 0.56032 0.0018913 0.42624 1.7433 1.7422 16.0091 144.9891 0.00020038 -85.5951 0.52796
0.632 0.98802 5.5217e-005 3.8182 0.012042 8.3256e-006 0.001154 0.10876 0.00065719 0.10941 0.098904 0 0.039847 0.0389 0 0.86532 0.23582 0.061968 0.0087351 4.1367 0.05469 6.5389e-005 0.83538 0.0051425 0.0058799 0.0013994 0.98677 0.99159 3.0191e-006 1.2076e-005 0.13077 0.90274 0.89389 0.001404 0.97745 0.56048 0.0018912 0.42626 1.7441 1.7429 16.0091 144.9891 0.00020017 -85.5957 0.52896
0.633 0.98802 5.5217e-005 3.8182 0.012042 8.3388e-006 0.001154 0.10886 0.00065719 0.10951 0.098998 0 0.03984 0.0389 0 0.86538 0.23584 0.061977 0.0087362 4.1368 0.054696 6.5397e-005 0.83537 0.0051427 0.00588 0.0013992 0.98678 0.9916 3.0188e-006 1.2075e-005 0.13077 0.90299 0.89403 0.0014039 0.97758 0.56063 0.0018912 0.42627 1.7448 1.7436 16.0091 144.9891 0.00019996 -85.5962 0.52996
0.634 0.98802 5.5217e-005 3.8182 0.012042 8.3519e-006 0.001154 0.10896 0.00065719 0.10961 0.099093 0 0.039832 0.0389 0 0.86543 0.23587 0.061986 0.0087373 4.137 0.054703 6.5406e-005 0.83536 0.0051428 0.0058802 0.0013991 0.98678 0.9916 3.0185e-006 1.2074e-005 0.13077 0.90325 0.89416 0.0014039 0.97771 0.56078 0.0018911 0.42628 1.7455 1.7443 16.009 144.9892 0.00019975 -85.5967 0.53096
0.635 0.98802 5.5217e-005 3.8182 0.012042 8.3651e-006 0.001154 0.10906 0.0006572 0.10971 0.099187 0 0.039825 0.0389 0 0.86549 0.23589 0.061995 0.0087384 4.1371 0.054709 6.5414e-005 0.83536 0.005143 0.0058803 0.001399 0.98678 0.9916 3.0183e-006 1.2073e-005 0.13077 0.9035 0.89429 0.0014038 0.97783 0.56094 0.001891 0.4263 1.7462 1.745 16.009 144.9892 0.00019955 -85.5972 0.53196
0.636 0.98802 5.5217e-005 3.8182 0.012042 8.3783e-006 0.001154 0.10916 0.0006572 0.10982 0.099281 0 0.039817 0.0389 0 0.86554 0.23592 0.062004 0.0087395 4.1372 0.054716 6.5422e-005 0.83535 0.0051432 0.0058805 0.0013989 0.98678 0.9916 3.018e-006 1.2072e-005 0.13077 0.90375 0.89442 0.0014037 0.97796 0.56109 0.0018909 0.42631 1.7469 1.7457 16.009 144.9892 0.00019934 -85.5977 0.53296
0.637 0.98802 5.5217e-005 3.8182 0.012042 8.3914e-006 0.001154 0.10926 0.0006572 0.10992 0.099374 0 0.03981 0.0389 0 0.8656 0.23594 0.062013 0.0087406 4.1374 0.054722 6.543e-005 0.83534 0.0051433 0.0058807 0.0013988 0.98678 0.9916 3.0177e-006 1.2071e-005 0.13077 0.904 0.89455 0.0014037 0.97808 0.56124 0.0018908 0.42632 1.7476 1.7464 16.009 144.9892 0.00019914 -85.5982 0.53396
0.638 0.98802 5.5217e-005 3.8182 0.012042 8.4046e-006 0.001154 0.10937 0.00065721 0.11002 0.099468 0 0.039802 0.0389 0 0.86565 0.23596 0.062022 0.0087418 4.1375 0.054729 6.5439e-005 0.83534 0.0051435 0.0058808 0.0013986 0.98678 0.9916 3.0175e-006 1.207e-005 0.13078 0.90424 0.89468 0.0014036 0.9782 0.56139 0.0018908 0.42634 1.7483 1.7471 16.009 144.9892 0.00019893 -85.5987 0.53496
0.639 0.98802 5.5217e-005 3.8182 0.012042 8.4177e-006 0.001154 0.10947 0.00065721 0.11012 0.099562 0 0.039795 0.0389 0 0.86571 0.23599 0.06203 0.0087429 4.1376 0.054735 6.5447e-005 0.83533 0.0051437 0.005881 0.0013985 0.98679 0.9916 3.0172e-006 1.2069e-005 0.13078 0.90449 0.89481 0.0014035 0.97833 0.56155 0.0018907 0.42635 1.749 1.7478 16.009 144.9893 0.00019873 -85.5992 0.53596
0.64 0.98802 5.5217e-005 3.8182 0.012042 8.4309e-006 0.001154 0.10957 0.00065721 0.11022 0.099656 0 0.039787 0.0389 0 0.86577 0.23601 0.062039 0.008744 4.1378 0.054742 6.5455e-005 0.83532 0.0051438 0.0058812 0.0013984 0.98679 0.9916 3.017e-006 1.2068e-005 0.13078 0.90474 0.89494 0.0014035 0.97845 0.5617 0.0018906 0.42636 1.7497 1.7485 16.0089 144.9893 0.00019852 -85.5996 0.53696
0.641 0.98802 5.5217e-005 3.8182 0.012042 8.4441e-006 0.001154 0.10967 0.00065722 0.11032 0.099749 0 0.03978 0.0389 0 0.86582 0.23604 0.062048 0.0087451 4.1379 0.054748 6.5464e-005 0.83532 0.005144 0.0058813 0.0013983 0.98679 0.9916 3.0167e-006 1.2067e-005 0.13078 0.90498 0.89507 0.0014034 0.97857 0.56185 0.0018905 0.42638 1.7504 1.7492 16.0089 144.9893 0.00019832 -85.6001 0.53796
0.642 0.98802 5.5217e-005 3.8182 0.012042 8.4572e-006 0.001154 0.10977 0.00065722 0.11042 0.099843 0 0.039773 0.0389 0 0.86588 0.23606 0.062057 0.0087462 4.1381 0.054755 6.5472e-005 0.83531 0.0051442 0.0058815 0.0013982 0.98679 0.9916 3.0164e-006 1.2066e-005 0.13078 0.90523 0.8952 0.0014034 0.97869 0.562 0.0018904 0.42639 1.7511 1.7499 16.0089 144.9893 0.00019812 -85.6006 0.53896
0.643 0.98802 5.5216e-005 3.8182 0.012041 8.4704e-006 0.001154 0.10987 0.00065723 0.11052 0.099936 0 0.039765 0.0389 0 0.86593 0.23609 0.062066 0.0087473 4.1382 0.054761 6.548e-005 0.8353 0.0051443 0.0058817 0.0013981 0.98679 0.99161 3.0162e-006 1.2065e-005 0.13078 0.90547 0.89532 0.0014033 0.97881 0.56215 0.0018904 0.4264 1.7518 1.7506 16.0089 144.9893 0.00019792 -85.6011 0.53996
0.644 0.98802 5.5216e-005 3.8182 0.012041 8.4835e-006 0.001154 0.10997 0.00065723 0.11062 0.10003 0 0.039758 0.0389 0 0.86599 0.23611 0.062075 0.0087484 4.1383 0.054768 6.5489e-005 0.8353 0.0051445 0.0058818 0.001398 0.98679 0.99161 3.0159e-006 1.2064e-005 0.13078 0.90572 0.89545 0.0014033 0.97893 0.56231 0.0018903 0.42642 1.7525 1.7513 16.0089 144.9894 0.00019772 -85.6015 0.54096
0.645 0.98802 5.5216e-005 3.8182 0.012041 8.4967e-006 0.001154 0.11007 0.00065723 0.11073 0.10012 0 0.03975 0.0389 0 0.86605 0.23614 0.062084 0.0087496 4.1385 0.054774 6.5497e-005 0.83529 0.0051447 0.005882 0.0013979 0.98679 0.99161 3.0157e-006 1.2063e-005 0.13079 0.90596 0.89558 0.0014032 0.97905 0.56246 0.0018902 0.42643 1.7531 1.752 16.0089 144.9894 0.00019752 -85.602 0.54196
0.646 0.98802 5.5216e-005 3.8182 0.012041 8.5099e-006 0.001154 0.11017 0.00065724 0.11083 0.10022 0 0.039743 0.0389 0 0.8661 0.23616 0.062093 0.0087507 4.1386 0.054781 6.5505e-005 0.83528 0.0051448 0.0058822 0.0013978 0.9868 0.99161 3.0154e-006 1.2062e-005 0.13079 0.9062 0.89571 0.0014031 0.97917 0.56261 0.0018901 0.42644 1.7538 1.7527 16.0088 144.9894 0.00019732 -85.6025 0.54296
0.647 0.98802 5.5216e-005 3.8182 0.012041 8.523e-006 0.001154 0.11027 0.00065724 0.11093 0.10031 0 0.039735 0.0389 0 0.86616 0.23619 0.062102 0.0087518 4.1388 0.054788 6.5514e-005 0.83528 0.005145 0.0058823 0.0013977 0.9868 0.99161 3.0152e-006 1.2061e-005 0.13079 0.90644 0.89583 0.0014031 0.97928 0.56276 0.0018901 0.42645 1.7545 1.7534 16.0088 144.9894 0.00019712 -85.6029 0.54396
0.648 0.98802 5.5216e-005 3.8182 0.012041 8.5362e-006 0.001154 0.11037 0.00065724 0.11103 0.1004 0 0.039728 0.0389 0 0.86622 0.23621 0.062111 0.0087529 4.1389 0.054794 6.5522e-005 0.83527 0.0051452 0.0058825 0.0013976 0.9868 0.99161 3.0149e-006 1.206e-005 0.13079 0.90669 0.89596 0.001403 0.9794 0.56291 0.00189 0.42647 1.7552 1.7541 16.0088 144.9894 0.00019692 -85.6034 0.54496
0.649 0.98802 5.5216e-005 3.8182 0.012041 8.5493e-006 0.001154 0.11047 0.00065725 0.11113 0.1005 0 0.039721 0.0389 0 0.86627 0.23624 0.06212 0.008754 4.1391 0.054801 6.553e-005 0.83526 0.0051454 0.0058827 0.0013975 0.9868 0.99161 3.0147e-006 1.2059e-005 0.13079 0.90693 0.89608 0.001403 0.97951 0.56307 0.0018899 0.42648 1.7559 1.7548 16.0088 144.9895 0.00019673 -85.6039 0.54596
0.65 0.98802 5.5216e-005 3.8182 0.012041 8.5625e-006 0.001154 0.11057 0.00065725 0.11123 0.10059 0 0.039713 0.0389 0 0.86633 0.23626 0.062129 0.0087552 4.1392 0.054807 6.5539e-005 0.83526 0.0051455 0.0058828 0.0013973 0.9868 0.99161 3.0145e-006 1.2058e-005 0.13079 0.90716 0.89621 0.0014029 0.97963 0.56322 0.0018898 0.42649 1.7566 1.7555 16.0088 144.9895 0.00019653 -85.6043 0.54696
0.651 0.98802 5.5216e-005 3.8182 0.012041 8.5757e-006 0.001154 0.11067 0.00065725 0.11133 0.10068 0 0.039706 0.0389 0 0.86639 0.23629 0.062138 0.0087563 4.1393 0.054814 6.5547e-005 0.83525 0.0051457 0.005883 0.0013972 0.9868 0.99161 3.0142e-006 1.2057e-005 0.13079 0.9074 0.89633 0.0014029 0.97974 0.56337 0.0018898 0.42651 1.7572 1.7561 16.0088 144.9895 0.00019634 -85.6048 0.54796
0.652 0.98802 5.5216e-005 3.8182 0.012041 8.5888e-006 0.001154 0.11078 0.00065726 0.11143 0.10077 0 0.039699 0.0389 0 0.86644 0.23631 0.062147 0.0087574 4.1395 0.054821 6.5556e-005 0.83524 0.0051459 0.0058832 0.0013971 0.9868 0.99161 3.014e-006 1.2056e-005 0.1308 0.90764 0.89645 0.0014028 0.97985 0.56352 0.0018897 0.42652 1.7579 1.7568 16.0087 144.9895 0.00019614 -85.6052 0.54896
0.653 0.98802 5.5216e-005 3.8182 0.012041 8.602e-006 0.001154 0.11088 0.00065726 0.11153 0.10087 0 0.039691 0.0389 0 0.8665 0.23634 0.062156 0.0087585 4.1396 0.054827 6.5564e-005 0.83524 0.005146 0.0058833 0.001397 0.9868 0.99161 3.0137e-006 1.2055e-005 0.1308 0.90788 0.89658 0.0014027 0.97997 0.56367 0.0018896 0.42653 1.7586 1.7575 16.0087 144.9895 0.00019595 -85.6057 0.54996
0.654 0.98802 5.5216e-005 3.8182 0.012041 8.6151e-006 0.001154 0.11098 0.00065727 0.11163 0.10096 0 0.039684 0.0389 0 0.86656 0.23636 0.062165 0.0087597 4.1398 0.054834 6.5573e-005 0.83523 0.0051462 0.0058835 0.0013969 0.98681 0.99161 3.0135e-006 1.2054e-005 0.1308 0.90811 0.8967 0.0014027 0.98008 0.56383 0.0018896 0.42655 1.7593 1.7582 16.0087 144.9896 0.00019575 -85.6061 0.55096
0.655 0.98802 5.5216e-005 3.8182 0.012041 8.6283e-006 0.001154 0.11107 0.00065727 0.11173 0.10105 0 0.039677 0.0389 0 0.86661 0.23639 0.062174 0.0087608 4.1399 0.05484 6.5581e-005 0.83523 0.0051464 0.0058837 0.0013968 0.98681 0.99162 3.0133e-006 1.2053e-005 0.1308 0.90835 0.89682 0.0014026 0.98019 0.56398 0.0018895 0.42656 1.7599 1.7588 16.0087 144.9896 0.00019556 -85.6065 0.55196
0.656 0.98802 5.5216e-005 3.8182 0.012041 8.6414e-006 0.001154 0.11117 0.00065727 0.11183 0.10114 0 0.039669 0.0389 0 0.86667 0.23641 0.062183 0.0087619 4.1401 0.054847 6.5589e-005 0.83522 0.0051465 0.0058838 0.0013967 0.98681 0.99162 3.013e-006 1.2052e-005 0.1308 0.90858 0.89694 0.0014026 0.9803 0.56413 0.0018894 0.42657 1.7606 1.7595 16.0087 144.9896 0.00019537 -85.607 0.55296
0.657 0.98802 5.5216e-005 3.8182 0.012041 8.6546e-006 0.001154 0.11127 0.00065728 0.11193 0.10124 0 0.039662 0.0389 0 0.86673 0.23644 0.062192 0.0087631 4.1402 0.054854 6.5598e-005 0.83521 0.0051467 0.005884 0.0013966 0.98681 0.99162 3.0128e-006 1.2051e-005 0.1308 0.90882 0.89706 0.0014025 0.98041 0.56428 0.0018894 0.42659 1.7613 1.7602 16.0086 144.9896 0.00019518 -85.6074 0.55396
0.658 0.98802 5.5216e-005 3.8182 0.012041 8.6678e-006 0.001154 0.11137 0.00065728 0.11203 0.10133 0 0.039655 0.0389 0 0.86678 0.23646 0.062201 0.0087642 4.1404 0.05486 6.5606e-005 0.83521 0.0051469 0.0058842 0.0013965 0.98681 0.99162 3.0126e-006 1.205e-005 0.1308 0.90905 0.89719 0.0014025 0.98052 0.56443 0.0018893 0.4266 1.7619 1.7609 16.0086 144.9896 0.00019499 -85.6078 0.55496
0.659 0.98802 5.5215e-005 3.8182 0.012041 8.6809e-006 0.001154 0.11147 0.00065728 0.11213 0.10142 0 0.039647 0.0389 0 0.86684 0.23649 0.06221 0.0087653 4.1405 0.054867 6.5615e-005 0.8352 0.0051471 0.0058844 0.0013964 0.98681 0.99162 3.0124e-006 1.2049e-005 0.13081 0.90928 0.89731 0.0014024 0.98062 0.56458 0.0018892 0.42661 1.7626 1.7615 16.0086 144.9897 0.0001948 -85.6083 0.55596
0.66 0.98802 5.5215e-005 3.8182 0.012041 8.6941e-006 0.001154 0.11157 0.00065729 0.11223 0.10151 0 0.03964 0.0389 0 0.8669 0.23651 0.062219 0.0087665 4.1407 0.054874 6.5623e-005 0.83519 0.0051472 0.0058845 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.13081 0.90952 0.89743 0.0014024 0.98073 0.56473 0.0018891 0.42663 1.7633 1.7622 16.0086 144.9897 0.00019461 -85.6087 0.55696
0.661 0.98802 5.5215e-005 3.8182 0.012041 8.7072e-006 0.001154 0.11167 0.00065729 0.11233 0.10161 0 0.039633 0.0389 0 0.86695 0.23654 0.062228 0.0087676 4.1408 0.05488 6.5632e-005 0.83519 0.0051474 0.0058847 0.0013962 0.98682 0.99162 3.0119e-006 1.2047e-005 0.13081 0.90975 0.89754 0.0014023 0.98084 0.56489 0.0018891 0.42664 1.7639 1.7629 16.0086 144.9897 0.00019442 -85.6091 0.55796
0.662 0.98802 5.5215e-005 3.8182 0.012041 8.7204e-006 0.001154 0.11177 0.00065729 0.11242 0.1017 0 0.039625 0.0389 0 0.86701 0.23656 0.062237 0.0087687 4.1409 0.054887 6.564e-005 0.83518 0.0051476 0.0058849 0.0013961 0.98682 0.99162 3.0117e-006 1.2047e-005 0.13081 0.90998 0.89766 0.0014023 0.98094 0.56504 0.001889 0.42665 1.7646 1.7635 16.0086 144.9897 0.00019424 -85.6095 0.55896
0.663 0.98802 5.5215e-005 3.8182 0.012041 8.7336e-006 0.001154 0.11187 0.0006573 0.11252 0.10179 0 0.039618 0.0389 0 0.86707 0.23659 0.062247 0.0087699 4.1411 0.054894 6.5649e-005 0.83517 0.0051478 0.0058851 0.001396 0.98682 0.99162 3.0114e-006 1.2046e-005 0.13081 0.91021 0.89778 0.0014022 0.98105 0.56519 0.0018889 0.42667 1.7652 1.7642 16.0085 144.9897 0.00019405 -85.61 0.55996
0.664 0.98802 5.5215e-005 3.8182 0.012041 8.7467e-006 0.001154 0.11197 0.0006573 0.11262 0.10188 0 0.039611 0.0389 0 0.86713 0.23661 0.062256 0.008771 4.1412 0.0549 6.5657e-005 0.83517 0.0051479 0.0058852 0.0013959 0.98682 0.99162 3.0112e-006 1.2045e-005 0.13081 0.91044 0.8979 0.0014022 0.98115 0.56534 0.0018889 0.42668 1.7659 1.7648 16.0085 144.9898 0.00019386 -85.6104 0.56096
0.665 0.98802 5.5215e-005 3.8182 0.012041 8.7599e-006 0.001154 0.11207 0.0006573 0.11272 0.10197 0 0.039604 0.0389 0 0.86718 0.23664 0.062265 0.0087722 4.1414 0.054907 6.5666e-005 0.83516 0.0051481 0.0058854 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.13081 0.91066 0.89802 0.0014021 0.98126 0.56549 0.0018888 0.42669 1.7666 1.7655 16.0085 144.9898 0.00019368 -85.6108 0.56196
0.666 0.98802 5.5215e-005 3.8182 0.012041 8.773e-006 0.001154 0.11217 0.00065731 0.11282 0.10207 0 0.039596 0.0389 0 0.86724 0.23666 0.062274 0.0087733 4.1415 0.054914 6.5675e-005 0.83515 0.0051483 0.0058856 0.0013957 0.98682 0.99162 3.0108e-006 1.2043e-005 0.13082 0.91089 0.89814 0.0014021 0.98136 0.56564 0.0018887 0.4267 1.7672 1.7662 16.0085 144.9898 0.00019349 -85.6112 0.56296
0.667 0.98802 5.5215e-005 3.8182 0.012041 8.7862e-006 0.001154 0.11227 0.00065731 0.11292 0.10216 0 0.039589 0.0389 0 0.8673 0.23669 0.062283 0.0087744 4.1417 0.054921 6.5683e-005 0.83515 0.0051485 0.0058858 0.0013956 0.98682 0.99163 3.0106e-006 1.2042e-005 0.13082 0.91112 0.89825 0.001402 0.98146 0.56579 0.0018887 0.42672 1.7679 1.7668 16.0085 144.9898 0.00019331 -85.6116 0.56396
0.668 0.98802 5.5215e-005 3.8182 0.012041 8.7993e-006 0.001154 0.11237 0.00065731 0.11302 0.10225 0 0.039582 0.0389 0 0.86736 0.23672 0.062292 0.0087756 4.1418 0.054927 6.5692e-005 0.83514 0.0051486 0.0058859 0.0013955 0.98682 0.99163 3.0104e-006 1.2041e-005 0.13082 0.91134 0.89837 0.001402 0.98157 0.56594 0.0018886 0.42673 1.7685 1.7675 16.0084 144.9898 0.00019313 -85.612 0.56496
0.669 0.98802 5.5215e-005 3.8182 0.012041 8.8125e-006 0.001154 0.11247 0.00065732 0.11312 0.10234 0 0.039575 0.0389 0 0.86741 0.23674 0.062301 0.0087767 4.142 0.054934 6.57e-005 0.83513 0.0051488 0.0058861 0.0013954 0.98683 0.99163 3.0102e-006 1.2041e-005 0.13082 0.91157 0.89849 0.0014019 0.98167 0.56609 0.0018886 0.42674 1.7692 1.7681 16.0084 144.9899 0.00019294 -85.6124 0.56596
0.67 0.98802 5.5215e-005 3.8182 0.012041 8.8257e-006 0.001154 0.11256 0.00065732 0.11322 0.10243 0 0.039568 0.0389 0 0.86747 0.23677 0.062311 0.0087779 4.1421 0.054941 6.5709e-005 0.83512 0.005149 0.0058863 0.0013953 0.98683 0.99163 3.01e-006 1.204e-005 0.13082 0.9118 0.8986 0.0014019 0.98177 0.56624 0.0018885 0.42676 1.7698 1.7688 16.0084 144.9899 0.00019276 -85.6128 0.56696
0.671 0.98802 5.5215e-005 3.8182 0.012041 8.8388e-006 0.001154 0.11266 0.00065732 0.11332 0.10252 0 0.03956 0.0389 0 0.86753 0.23679 0.06232 0.008779 4.1423 0.054948 6.5717e-005 0.83512 0.0051492 0.0058865 0.0013952 0.98683 0.99163 3.0097e-006 1.2039e-005 0.13082 0.91202 0.89872 0.0014018 0.98187 0.5664 0.0018884 0.42677 1.7705 1.7694 16.0084 144.9899 0.00019258 -85.6132 0.56796
0.672 0.98802 5.5215e-005 3.8182 0.012041 8.852e-006 0.001154 0.11276 0.00065733 0.11341 0.10261 0 0.039553 0.0389 0 0.86759 0.23682 0.062329 0.0087802 4.1424 0.054954 6.5726e-005 0.83511 0.0051494 0.0058866 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.13082 0.91224 0.89883 0.0014018 0.98197 0.56655 0.0018884 0.42678 1.7711 1.7701 16.0084 144.9899 0.0001924 -85.6136 0.56896
0.673 0.98802 5.5215e-005 3.8182 0.012041 8.8651e-006 0.001154 0.11286 0.00065733 0.11351 0.10271 0 0.039546 0.0389 0 0.86764 0.23684 0.062338 0.0087813 4.1426 0.054961 6.5735e-005 0.8351 0.0051495 0.0058868 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.13083 0.91247 0.89895 0.0014017 0.98207 0.5667 0.0018883 0.4268 1.7717 1.7707 16.0084 144.9899 0.00019222 -85.614 0.56996
0.674 0.98802 5.5215e-005 3.8182 0.012041 8.8783e-006 0.001154 0.11296 0.00065733 0.11361 0.1028 0 0.039539 0.0389 0 0.8677 0.23687 0.062347 0.0087825 4.1427 0.054968 6.5743e-005 0.8351 0.0051497 0.005887 0.001395 0.98683 0.99163 3.0091e-006 1.2036e-005 0.13083 0.91269 0.89906 0.0014017 0.98216 0.56685 0.0018882 0.42681 1.7724 1.7714 16.0083 144.99 0.00019204 -85.6143 0.57096
0.675 0.98802 5.5214e-005 3.8182 0.012041 8.8915e-006 0.001154 0.11306 0.00065734 0.11371 0.10289 0 0.039532 0.0389 0 0.86776 0.23689 0.062357 0.0087836 4.1429 0.054975 6.5752e-005 0.83509 0.0051499 0.0058872 0.0013949 0.98683 0.99163 3.0089e-006 1.2036e-005 0.13083 0.91291 0.89917 0.0014016 0.98226 0.567 0.0018882 0.42682 1.773 1.772 16.0083 144.99 0.00019186 -85.6147 0.57196
0.676 0.98802 5.5214e-005 3.8182 0.012041 8.9046e-006 0.001154 0.11315 0.00065734 0.11381 0.10298 0 0.039525 0.0389 0 0.86782 0.23692 0.062366 0.0087848 4.1431 0.054981 6.5761e-005 0.83508 0.0051501 0.0058873 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.13083 0.91313 0.89929 0.0014016 0.98236 0.56715 0.0018881 0.42684 1.7737 1.7726 16.0083 144.99 0.00019169 -85.6151 0.57296
0.677 0.98802 5.5214e-005 3.8182 0.012041 8.9178e-006 0.001154 0.11325 0.00065734 0.11391 0.10307 0 0.039517 0.0389 0 0.86788 0.23694 0.062375 0.0087859 4.1432 0.054988 6.5769e-005 0.83508 0.0051503 0.0058875 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.13083 0.91335 0.8994 0.0014015 0.98245 0.5673 0.0018881 0.42685 1.7743 1.7733 16.0083 144.99 0.00019151 -85.6155 0.57396
0.678 0.98802 5.5214e-005 3.8182 0.012041 8.9309e-006 0.001154 0.11335 0.00065735 0.114 0.10316 0 0.03951 0.0389 0 0.86793 0.23697 0.062384 0.0087871 4.1434 0.054995 6.5778e-005 0.83507 0.0051504 0.0058877 0.0013946 0.98684 0.99163 3.0083e-006 1.2033e-005 0.13083 0.91357 0.89951 0.0014015 0.98255 0.56745 0.001888 0.42686 1.7749 1.7739 16.0083 144.99 0.00019133 -85.6159 0.57496
0.679 0.98802 5.5214e-005 3.8182 0.012041 8.9441e-006 0.001154 0.11345 0.00065735 0.1141 0.10325 0 0.039503 0.0389 0 0.86799 0.237 0.062393 0.0087882 4.1435 0.055002 6.5787e-005 0.83506 0.0051506 0.0058879 0.0013945 0.98684 0.99163 3.0081e-006 1.2032e-005 0.13084 0.91379 0.89962 0.0014015 0.98264 0.5676 0.0018879 0.42688 1.7756 1.7746 16.0082 144.9901 0.00019116 -85.6162 0.57596
0.68 0.98802 5.5214e-005 3.8182 0.012041 8.9572e-006 0.001154 0.11355 0.00065735 0.1142 0.10334 0 0.039496 0.0389 0 0.86805 0.23702 0.062403 0.0087894 4.1437 0.055009 6.5795e-005 0.83506 0.0051508 0.0058881 0.0013945 0.98684 0.99164 3.0079e-006 1.2032e-005 0.13084 0.914 0.89973 0.0014014 0.98274 0.56775 0.0018879 0.42689 1.7762 1.7752 16.0082 144.9901 0.00019098 -85.6166 0.57696
0.681 0.98802 5.5214e-005 3.8182 0.012041 8.9704e-006 0.001154 0.11364 0.00065736 0.1143 0.10343 0 0.039489 0.0389 0 0.86811 0.23705 0.062412 0.0087905 4.1438 0.055015 6.5804e-005 0.83505 0.005151 0.0058882 0.0013944 0.98684 0.99164 3.0077e-006 1.2031e-005 0.13084 0.91422 0.89985 0.0014014 0.98283 0.5679 0.0018878 0.4269 1.7768 1.7758 16.0082 144.9901 0.00019081 -85.617 0.57796
0.682 0.98802 5.5214e-005 3.8182 0.012041 8.9836e-006 0.001154 0.11374 0.00065736 0.11439 0.10352 0 0.039482 0.0389 0 0.86817 0.23707 0.062421 0.0087917 4.144 0.055022 6.5813e-005 0.83504 0.0051512 0.0058884 0.0013943 0.98684 0.99164 3.0075e-006 1.203e-005 0.13084 0.91444 0.89996 0.0014013 0.98292 0.56805 0.0018878 0.42691 1.7775 1.7765 16.0082 144.9901 0.00019063 -85.6173 0.57896
0.683 0.98802 5.5214e-005 3.8182 0.012041 8.9967e-006 0.001154 0.11384 0.00065736 0.11449 0.10361 0 0.039475 0.0389 0 0.86822 0.2371 0.062431 0.0087928 4.1441 0.055029 6.5821e-005 0.83504 0.0051514 0.0058886 0.0013942 0.98684 0.99164 3.0073e-006 1.2029e-005 0.13084 0.91465 0.90007 0.0014013 0.98302 0.5682 0.0018877 0.42693 1.7781 1.7771 16.0082 144.9901 0.00019046 -85.6177 0.57996
0.684 0.98802 5.5214e-005 3.8182 0.012041 9.0099e-006 0.001154 0.11394 0.00065737 0.11459 0.1037 0 0.039468 0.0389 0 0.86828 0.23712 0.06244 0.008794 4.1443 0.055036 6.583e-005 0.83503 0.0051515 0.0058888 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.13084 0.91487 0.90018 0.0014012 0.98311 0.56835 0.0018876 0.42694 1.7787 1.7777 16.0081 144.9902 0.00019029 -85.6181 0.58096
0.685 0.98802 5.5214e-005 3.8182 0.012041 9.023e-006 0.001154 0.11403 0.00065737 0.11469 0.1038 0 0.03946 0.0389 0 0.86834 0.23715 0.062449 0.0087952 4.1444 0.055043 6.5839e-005 0.83502 0.0051517 0.005889 0.0013941 0.98684 0.99164 3.0069e-006 1.2028e-005 0.13084 0.91508 0.90029 0.0014012 0.9832 0.5685 0.0018876 0.42695 1.7793 1.7783 16.0081 144.9902 0.00019011 -85.6184 0.58196
0.686 0.98802 5.5214e-005 3.8182 0.012041 9.0362e-006 0.001154 0.11413 0.00065737 0.11479 0.10389 0 0.039453 0.0389 0 0.8684 0.23718 0.062458 0.0087963 4.1446 0.05505 6.5848e-005 0.83502 0.0051519 0.0058892 0.001394 0.98684 0.99164 3.0067e-006 1.2027e-005 0.13085 0.9153 0.90039 0.0014011 0.98329 0.56865 0.0018875 0.42697 1.78 1.779 16.0081 144.9902 0.00018994 -85.6188 0.58296
0.687 0.98802 5.5214e-005 3.8182 0.012041 9.0493e-006 0.001154 0.11423 0.00065738 0.11488 0.10398 0 0.039446 0.0389 0 0.86846 0.2372 0.062468 0.0087975 4.1448 0.055057 6.5856e-005 0.83501 0.0051521 0.0058893 0.0013939 0.98685 0.99164 3.0066e-006 1.2026e-005 0.13085 0.91551 0.9005 0.0014011 0.98338 0.5688 0.0018875 0.42698 1.7806 1.7796 16.0081 144.9902 0.00018977 -85.6191 0.58396
0.688 0.98802 5.5214e-005 3.8182 0.012041 9.0625e-006 0.001154 0.11433 0.00065738 0.11498 0.10407 0 0.039439 0.0389 0 0.86852 0.23723 0.062477 0.0087986 4.1449 0.055063 6.5865e-005 0.835 0.0051523 0.0058895 0.0013938 0.98685 0.99164 3.0064e-006 1.2025e-005 0.13085 0.91572 0.90061 0.0014011 0.98347 0.56895 0.0018874 0.42699 1.7812 1.7802 16.0081 144.9902 0.0001896 -85.6195 0.58496
0.689 0.98802 5.5214e-005 3.8182 0.012041 9.0757e-006 0.001154 0.11442 0.00065738 0.11508 0.10416 0 0.039432 0.0389 0 0.86858 0.23725 0.062486 0.0087998 4.1451 0.05507 6.5874e-005 0.835 0.0051525 0.0058897 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.13085 0.91593 0.90072 0.001401 0.98356 0.5691 0.0018874 0.42701 1.7818 1.7808 16.008 144.9903 0.00018943 -85.6198 0.58596
0.69 0.98802 5.5214e-005 3.8182 0.012041 9.0888e-006 0.001154 0.11452 0.00065739 0.11517 0.10425 0 0.039425 0.0389 0 0.86863 0.23728 0.062496 0.008801 4.1452 0.055077 6.5883e-005 0.83499 0.0051526 0.0058899 0.0013936 0.98685 0.99164 3.006e-006 1.2024e-005 0.13085 0.91615 0.90083 0.001401 0.98365 0.56925 0.0018873 0.42702 1.7825 1.7815 16.008 144.9903 0.00018926 -85.6202 0.58696
0.691 0.98802 5.5214e-005 3.8182 0.012041 9.102e-006 0.001154 0.11462 0.00065739 0.11527 0.10434 0 0.039418 0.0389 0 0.86869 0.23731 0.062505 0.0088021 4.1454 0.055084 6.5891e-005 0.83498 0.0051528 0.0058901 0.0013935 0.98685 0.99164 3.0058e-006 1.2023e-005 0.13085 0.91636 0.90093 0.0014009 0.98374 0.5694 0.0018872 0.42703 1.7831 1.7821 16.008 144.9903 0.00018909 -85.6205 0.58796
0.692 0.98802 5.5213e-005 3.8182 0.012041 9.1151e-006 0.001154 0.11472 0.00065739 0.11537 0.10443 0 0.039411 0.0389 0 0.86875 0.23733 0.062514 0.0088033 4.1455 0.055091 6.59e-005 0.83497 0.005153 0.0058903 0.0013935 0.98685 0.99164 3.0056e-006 1.2022e-005 0.13086 0.91657 0.90104 0.0014009 0.98382 0.56955 0.0018872 0.42705 1.7837 1.7827 16.008 144.9903 0.00018893 -85.6209 0.58896
0.693 0.98802 5.5213e-005 3.8182 0.012041 9.1283e-006 0.001154 0.11481 0.0006574 0.11547 0.10452 0 0.039404 0.0389 0 0.86881 0.23736 0.062524 0.0088045 4.1457 0.055098 6.5909e-005 0.83497 0.0051532 0.0058904 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.13086 0.91677 0.90115 0.0014008 0.98391 0.5697 0.0018871 0.42706 1.7843 1.7833 16.008 144.9903 0.00018876 -85.6212 0.58996
0.694 0.98802 5.5213e-005 3.8182 0.012041 9.1414e-006 0.001154 0.11491 0.0006574 0.11556 0.10461 0 0.039397 0.0389 0 0.86887 0.23738 0.062533 0.0088056 4.1459 0.055105 6.5918e-005 0.83496 0.0051534 0.0058906 0.0013933 0.98685 0.99164 3.0053e-006 1.2021e-005 0.13086 0.91698 0.90125 0.0014008 0.984 0.56985 0.0018871 0.42707 1.7849 1.7839 16.0079 144.9904 0.00018859 -85.6216 0.59096
0.695 0.98802 5.5213e-005 3.8182 0.012041 9.1546e-006 0.001154 0.11501 0.0006574 0.11566 0.1047 0 0.03939 0.0389 0 0.86893 0.23741 0.062543 0.0088068 4.146 0.055112 6.5927e-005 0.83495 0.0051536 0.0058908 0.0013932 0.98685 0.99165 3.0051e-006 1.202e-005 0.13086 0.91719 0.90136 0.0014008 0.98408 0.57 0.001887 0.42708 1.7855 1.7845 16.0079 144.9904 0.00018843 -85.6219 0.59196
0.696 0.98802 5.5213e-005 3.8182 0.012041 9.1678e-006 0.001154 0.1151 0.00065741 0.11576 0.10479 0 0.039383 0.0389 0 0.86899 0.23744 0.062552 0.008808 4.1462 0.055119 6.5935e-005 0.83495 0.0051538 0.005891 0.0013932 0.98685 0.99165 3.0049e-006 1.202e-005 0.13086 0.9174 0.90146 0.0014007 0.98417 0.57015 0.001887 0.4271 1.7861 1.7852 16.0079 144.9904 0.00018826 -85.6222 0.59296
0.697 0.98802 5.5213e-005 3.8182 0.012041 9.1809e-006 0.001154 0.1152 0.00065741 0.11585 0.10488 0 0.039376 0.0389 0 0.86905 0.23746 0.062561 0.0088092 4.1463 0.055126 6.5944e-005 0.83494 0.005154 0.0058912 0.0013931 0.98686 0.99165 3.0047e-006 1.2019e-005 0.13086 0.91761 0.90157 0.0014007 0.98425 0.5703 0.0018869 0.42711 1.7867 1.7858 16.0079 144.9904 0.0001881 -85.6226 0.59396
0.698 0.98802 5.5213e-005 3.8182 0.012041 9.1941e-006 0.001154 0.1153 0.00065741 0.11595 0.10496 0 0.039369 0.0389 0 0.8691 0.23749 0.062571 0.0088103 4.1465 0.055132 6.5953e-005 0.83493 0.0051541 0.0058914 0.001393 0.98686 0.99165 3.0046e-006 1.2018e-005 0.13086 0.91781 0.90167 0.0014006 0.98433 0.57045 0.0018869 0.42712 1.7873 1.7864 16.0079 144.9904 0.00018793 -85.6229 0.59496
0.699 0.98802 5.5213e-005 3.8182 0.012041 9.2072e-006 0.001154 0.11539 0.00065742 0.11604 0.10505 0 0.039362 0.0389 0 0.86916 0.23751 0.06258 0.0088115 4.1467 0.055139 6.5962e-005 0.83493 0.0051543 0.0058916 0.0013929 0.98686 0.99165 3.0044e-006 1.2017e-005 0.13087 0.91802 0.90178 0.0014006 0.98442 0.5706 0.0018868 0.42714 1.7879 1.787 16.0078 144.9905 0.00018777 -85.6232 0.59596
0.7 0.98802 5.5213e-005 3.8182 0.012041 9.2204e-006 0.001154 0.11549 0.00065742 0.11614 0.10514 0 0.039355 0.0389 0 0.86922 0.23754 0.06259 0.0088127 4.1468 0.055146 6.5971e-005 0.83492 0.0051545 0.0058918 0.0013929 0.98686 0.99165 3.0042e-006 1.2017e-005 0.13087 0.91822 0.90188 0.0014006 0.9845 0.57075 0.0018868 0.42715 1.7885 1.7876 16.0078 144.9905 0.00018761 -85.6235 0.59696
0.701 0.98802 5.5213e-005 3.8182 0.012041 9.2335e-006 0.001154 0.11558 0.00065742 0.11624 0.10523 0 0.039348 0.0389 0 0.86928 0.23757 0.062599 0.0088139 4.147 0.055153 6.598e-005 0.83491 0.0051547 0.0058919 0.0013928 0.98686 0.99165 3.004e-006 1.2016e-005 0.13087 0.91842 0.90198 0.0014005 0.98458 0.5709 0.0018867 0.42716 1.7891 1.7882 16.0078 144.9905 0.00018745 -85.6239 0.59796
0.702 0.98802 5.5213e-005 3.8182 0.012041 9.2467e-006 0.001154 0.11568 0.00065742 0.11633 0.10532 0 0.039341 0.0389 0 0.86934 0.23759 0.062608 0.008815 4.1472 0.05516 6.5989e-005 0.83491 0.0051549 0.0058921 0.0013927 0.98686 0.99165 3.0039e-006 1.2015e-005 0.13087 0.91863 0.90209 0.0014005 0.98466 0.57105 0.0018867 0.42718 1.7897 1.7888 16.0078 144.9905 0.00018728 -85.6242 0.59896
0.703 0.98802 5.5213e-005 3.8182 0.012041 9.2599e-006 0.001154 0.11578 0.00065743 0.11643 0.10541 0 0.039334 0.0389 0 0.8694 0.23762 0.062618 0.0088162 4.1473 0.055167 6.5998e-005 0.8349 0.0051551 0.0058923 0.0013926 0.98686 0.99165 3.0037e-006 1.2015e-005 0.13087 0.91883 0.90219 0.0014004 0.98475 0.57119 0.0018866 0.42719 1.7903 1.7894 16.0078 144.9905 0.00018712 -85.6245 0.59996
0.704 0.98802 5.5213e-005 3.8182 0.012041 9.273e-006 0.001154 0.11587 0.00065743 0.11653 0.1055 0 0.039327 0.0389 0 0.86946 0.23764 0.062627 0.0088174 4.1475 0.055174 6.6006e-005 0.83489 0.0051553 0.0058925 0.0013926 0.98686 0.99165 3.0035e-006 1.2014e-005 0.13087 0.91903 0.90229 0.0014004 0.98483 0.57134 0.0018866 0.4272 1.7909 1.79 16.0077 144.9906 0.00018696 -85.6248 0.60096
0.705 0.98802 5.5213e-005 3.8182 0.012041 9.2862e-006 0.001154 0.11597 0.00065743 0.11662 0.10559 0 0.03932 0.0389 0 0.86952 0.23767 0.062637 0.0088186 4.1476 0.055181 6.6015e-005 0.83488 0.0051555 0.0058927 0.0013925 0.98686 0.99165 3.0034e-006 1.2013e-005 0.13088 0.91923 0.90239 0.0014004 0.98491 0.57149 0.0018865 0.42722 1.7915 1.7906 16.0077 144.9906 0.0001868 -85.6251 0.60196
0.706 0.98802 5.5213e-005 3.8182 0.012041 9.2993e-006 0.001154 0.11606 0.00065744 0.11672 0.10568 0 0.039314 0.0389 0 0.86958 0.2377 0.062646 0.0088198 4.1478 0.055188 6.6024e-005 0.83488 0.0051557 0.0058929 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.13088 0.91944 0.90249 0.0014003 0.98499 0.57164 0.0018865 0.42723 1.7921 1.7912 16.0077 144.9906 0.00018664 -85.6254 0.60296
0.707 0.98802 5.5213e-005 3.8182 0.012041 9.3125e-006 0.001154 0.11616 0.00065744 0.11681 0.10577 0 0.039307 0.0389 0 0.86964 0.23772 0.062656 0.0088209 4.148 0.055195 6.6033e-005 0.83487 0.0051559 0.0058931 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.13088 0.91964 0.9026 0.0014003 0.98507 0.57179 0.0018864 0.42724 1.7927 1.7918 16.0077 144.9906 0.00018648 -85.6258 0.60396
0.708 0.98802 5.5212e-005 3.8182 0.012041 9.3256e-006 0.0011541 0.11626 0.00065744 0.11691 0.10586 0 0.0393 0.0389 0 0.8697 0.23775 0.062665 0.0088221 4.1481 0.055202 6.6042e-005 0.83486 0.0051561 0.0058933 0.0013923 0.98687 0.99165 3.0029e-006 1.2011e-005 0.13088 0.91984 0.9027 0.0014002 0.98514 0.57194 0.0018864 0.42725 1.7933 1.7924 16.0076 144.9906 0.00018633 -85.6261 0.60496
0.709 0.98802 5.5212e-005 3.8182 0.012041 9.3388e-006 0.0011541 0.11635 0.00065745 0.117 0.10594 0 0.039293 0.0389 0 0.86976 0.23778 0.062675 0.0088233 4.1483 0.055209 6.6051e-005 0.83486 0.0051563 0.0058935 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.13088 0.92003 0.9028 0.0014002 0.98522 0.57209 0.0018863 0.42727 1.7939 1.793 16.0076 144.9907 0.00018617 -85.6264 0.60596
0.71 0.98802 5.5212e-005 3.8182 0.012041 9.3519e-006 0.0011541 0.11645 0.00065745 0.1171 0.10603 0 0.039286 0.0389 0 0.86982 0.2378 0.062684 0.0088245 4.1485 0.055216 6.606e-005 0.83485 0.0051564 0.0058937 0.0013921 0.98687 0.99165 3.0026e-006 1.201e-005 0.13088 0.92023 0.9029 0.0014002 0.9853 0.57224 0.0018863 0.42728 1.7945 1.7936 16.0076 144.9907 0.00018601 -85.6267 0.60696
0.711 0.98802 5.5212e-005 3.8182 0.012041 9.3651e-006 0.0011541 0.11654 0.00065745 0.1172 0.10612 0 0.039279 0.0389 0 0.86988 0.23783 0.062694 0.0088257 4.1486 0.055223 6.6069e-005 0.83484 0.0051566 0.0058939 0.001392 0.98687 0.99166 3.0024e-006 1.2009e-005 0.13089 0.92043 0.903 0.0014001 0.98538 0.57239 0.0018862 0.42729 1.7951 1.7942 16.0076 144.9907 0.00018585 -85.627 0.60796
0.712 0.98802 5.5212e-005 3.8182 0.012041 9.3783e-006 0.0011541 0.11664 0.00065746 0.11729 0.10621 0 0.039272 0.0389 0 0.86994 0.23786 0.062703 0.0088269 4.1488 0.05523 6.6078e-005 0.83484 0.0051568 0.005894 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.13089 0.92063 0.90309 0.0014001 0.98545 0.57253 0.0018862 0.42731 1.7957 1.7947 16.0076 144.9907 0.0001857 -85.6273 0.60896
0.713 0.98802 5.5212e-005 3.8182 0.012041 9.3914e-006 0.0011541 0.11673 0.00065746 0.11739 0.1063 0 0.039265 0.0389 0 0.87 0.23788 0.062713 0.008828 4.149 0.055237 6.6087e-005 0.83483 0.005157 0.0058942 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.13089 0.92082 0.90319 0.0014001 0.98553 0.57268 0.0018861 0.42732 1.7963 1.7953 16.0075 144.9907 0.00018554 -85.6276 0.60996
0.714 0.98802 5.5212e-005 3.8182 0.012041 9.4046e-006 0.0011541 0.11683 0.00065746 0.11748 0.10639 0 0.039258 0.0389 0 0.87006 0.23791 0.062722 0.0088292 4.1491 0.055244 6.6096e-005 0.83482 0.0051572 0.0058944 0.0013918 0.98687 0.99166 3.0019e-006 1.2008e-005 0.13089 0.92102 0.90329 0.0014 0.98561 0.57283 0.0018861 0.42733 1.7968 1.7959 16.0075 144.9908 0.00018539 -85.6279 0.61096
0.715 0.98802 5.5212e-005 3.8182 0.012041 9.4177e-006 0.0011541 0.11692 0.00065746 0.11758 0.10648 0 0.039252 0.0389 0 0.87012 0.23793 0.062732 0.0088304 4.1493 0.055251 6.6105e-005 0.83481 0.0051574 0.0058946 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.13089 0.92122 0.90339 0.0014 0.98568 0.57298 0.001886 0.42735 1.7974 1.7965 16.0075 144.9908 0.00018523 -85.6282 0.61196
0.716 0.98802 5.5212e-005 3.8182 0.012041 9.4309e-006 0.0011541 0.11702 0.00065747 0.11767 0.10656 0 0.039245 0.0389 0 0.87018 0.23796 0.062742 0.0088316 4.1495 0.055259 6.6114e-005 0.83481 0.0051576 0.0058948 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.13089 0.92141 0.90349 0.0014 0.98575 0.57313 0.001886 0.42736 1.798 1.7971 16.0075 144.9908 0.00018508 -85.6284 0.61296
0.717 0.98802 5.5212e-005 3.8182 0.012041 9.444e-006 0.0011541 0.11711 0.00065747 0.11777 0.10665 0 0.039238 0.0389 0 0.87024 0.23799 0.062751 0.0088328 4.1496 0.055266 6.6123e-005 0.8348 0.0051578 0.005895 0.0013916 0.98687 0.99166 3.0015e-006 1.2006e-005 0.13089 0.9216 0.90359 0.0013999 0.98583 0.57328 0.0018859 0.42737 1.7986 1.7977 16.0075 144.9908 0.00018493 -85.6287 0.61396
0.718 0.98802 5.5212e-005 3.8182 0.01204 9.4572e-006 0.0011541 0.11721 0.00065747 0.11786 0.10674 0 0.039231 0.0389 0 0.8703 0.23801 0.062761 0.008834 4.1498 0.055273 6.6132e-005 0.83479 0.005158 0.0058952 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.1309 0.9218 0.90368 0.0013999 0.9859 0.57343 0.0018859 0.42738 1.7992 1.7982 16.0074 144.9908 0.00018477 -85.629 0.61496
0.719 0.98802 5.5212e-005 3.8182 0.01204 9.4704e-006 0.0011541 0.1173 0.00065748 0.11796 0.10683 0 0.039224 0.0389 0 0.87036 0.23804 0.06277 0.0088352 4.15 0.05528 6.6141e-005 0.83479 0.0051582 0.0058954 0.0013915 0.98688 0.99166 3.0011e-006 1.2005e-005 0.1309 0.92199 0.90378 0.0013998 0.98598 0.57357 0.0018858 0.4274 1.7997 1.7988 16.0074 144.9909 0.00018462 -85.6293 0.61596
0.72 0.98802 5.5212e-005 3.8182 0.01204 9.4835e-006 0.0011541 0.1174 0.00065748 0.11805 0.10692 0 0.039217 0.0389 0 0.87042 0.23807 0.06278 0.0088364 4.1501 0.055287 6.615e-005 0.83478 0.0051584 0.0058956 0.0013914 0.98688 0.99166 3.001e-006 1.2004e-005 0.1309 0.92218 0.90388 0.0013998 0.98605 0.57372 0.0018858 0.42741 1.8003 1.7994 16.0074 144.9909 0.00018447 -85.6296 0.61696
0.721 0.98802 5.5212e-005 3.8182 0.01204 9.4967e-006 0.0011541 0.11749 0.00065748 0.11815 0.107 0 0.039211 0.0389 0 0.87048 0.23809 0.062789 0.0088376 4.1503 0.055294 6.6159e-005 0.83477 0.0051586 0.0058958 0.0013914 0.98688 0.99166 3.0008e-006 1.2003e-005 0.1309 0.92237 0.90397 0.0013998 0.98612 0.57387 0.0018857 0.42742 1.8009 1.8 16.0074 144.9909 0.00018432 -85.6299 0.61796
0.722 0.98802 5.5212e-005 3.8182 0.01204 9.5098e-006 0.0011541 0.11759 0.00065749 0.11824 0.10709 0 0.039204 0.0389 0 0.87054 0.23812 0.062799 0.0088388 4.1505 0.055301 6.6168e-005 0.83477 0.0051588 0.005896 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.1309 0.92256 0.90407 0.0013997 0.98619 0.57402 0.0018857 0.42744 1.8015 1.8006 16.0073 144.9909 0.00018417 -85.6302 0.61896
0.723 0.98802 5.5212e-005 3.8182 0.01204 9.523e-006 0.0011541 0.11768 0.00065749 0.11834 0.10718 0 0.039197 0.0389 0 0.8706 0.23815 0.062809 0.00884 4.1507 0.055308 6.6177e-005 0.83476 0.005159 0.0058962 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.1309 0.92276 0.90416 0.0013997 0.98626 0.57417 0.0018857 0.42745 1.802 1.8011 16.0073 144.9909 0.00018402 -85.6304 0.61996
0.724 0.98802 5.5211e-005 3.8182 0.01204 9.5361e-006 0.0011541 0.11778 0.00065749 0.11843 0.10727 0 0.03919 0.0389 0 0.87066 0.23817 0.062818 0.0088412 4.1508 0.055315 6.6186e-005 0.83475 0.0051592 0.0058964 0.0013912 0.98688 0.99166 3.0004e-006 1.2002e-005 0.13091 0.92295 0.90426 0.0013997 0.98633 0.57432 0.0018856 0.42746 1.8026 1.8017 16.0073 144.991 0.00018387 -85.6307 0.62096
0.725 0.98802 5.5211e-005 3.8182 0.01204 9.5493e-006 0.0011541 0.11787 0.00065749 0.11853 0.10736 0 0.039184 0.0389 0 0.87072 0.2382 0.062828 0.0088424 4.151 0.055322 6.6195e-005 0.83474 0.0051594 0.0058966 0.0013911 0.98688 0.99166 3.0003e-006 1.2001e-005 0.13091 0.92313 0.90435 0.0013996 0.98641 0.57446 0.0018856 0.42748 1.8032 1.8023 16.0073 144.991 0.00018372 -85.631 0.62196
0.726 0.98802 5.5211e-005 3.8182 0.01204 9.5624e-006 0.0011541 0.11797 0.0006575 0.11862 0.10744 0 0.039177 0.0389 0 0.87078 0.23823 0.062838 0.0088436 4.1512 0.05533 6.6205e-005 0.83474 0.0051596 0.0058968 0.0013911 0.98688 0.99166 3.0001e-006 1.2e-005 0.13091 0.92332 0.90445 0.0013996 0.98648 0.57461 0.0018855 0.42749 1.8037 1.8028 16.0073 144.991 0.00018357 -85.6313 0.62296
0.727 0.98802 5.5211e-005 3.8182 0.01204 9.5756e-006 0.0011541 0.11806 0.0006575 0.11871 0.10753 0 0.03917 0.0389 0 0.87084 0.23825 0.062847 0.0088448 4.1513 0.055337 6.6214e-005 0.83473 0.0051598 0.005897 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.13091 0.92351 0.90454 0.0013996 0.98654 0.57476 0.0018855 0.4275 1.8043 1.8034 16.0072 144.991 0.00018343 -85.6315 0.62396
0.728 0.98802 5.5211e-005 3.8182 0.01204 9.5888e-006 0.0011541 0.11816 0.0006575 0.11881 0.10762 0 0.039163 0.0389 0 0.8709 0.23828 0.062857 0.008846 4.1515 0.055344 6.6223e-005 0.83472 0.00516 0.0058972 0.0013909 0.98688 0.99166 2.9998e-006 1.1999e-005 0.13091 0.9237 0.90464 0.0013995 0.98661 0.57491 0.0018854 0.42751 1.8049 1.804 16.0072 144.9911 0.00018328 -85.6318 0.62496
0.729 0.98802 5.5211e-005 3.8182 0.01204 9.6019e-006 0.0011541 0.11825 0.00065751 0.1189 0.10771 0 0.039157 0.0389 0 0.87096 0.23831 0.062867 0.0088472 4.1517 0.055351 6.6232e-005 0.83472 0.0051602 0.0058974 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.13091 0.92389 0.90473 0.0013995 0.98668 0.57506 0.0018854 0.42753 1.8054 1.8045 16.0072 144.9911 0.00018313 -85.6321 0.62596
0.73 0.98802 5.5211e-005 3.8182 0.01204 9.6151e-006 0.0011541 0.11834 0.00065751 0.119 0.10779 0 0.03915 0.0389 0 0.87102 0.23833 0.062876 0.0088484 4.1519 0.055358 6.6241e-005 0.83471 0.0051604 0.0058976 0.0013908 0.98688 0.99167 2.9995e-006 1.1998e-005 0.13092 0.92407 0.90482 0.0013995 0.98675 0.5752 0.0018854 0.42754 1.806 1.8051 16.0072 144.9911 0.00018299 -85.6323 0.62696
0.731 0.98802 5.5211e-005 3.8182 0.01204 9.6282e-006 0.0011541 0.11844 0.00065751 0.11909 0.10788 0 0.039143 0.0389 0 0.87108 0.23836 0.062886 0.0088496 4.152 0.055365 6.625e-005 0.8347 0.0051606 0.0058978 0.0013908 0.98689 0.99167 2.9994e-006 1.1998e-005 0.13092 0.92426 0.90491 0.0013994 0.98682 0.57535 0.0018853 0.42755 1.8066 1.8057 16.0071 144.9911 0.00018284 -85.6326 0.62796
0.732 0.98802 5.5211e-005 3.8182 0.01204 9.6414e-006 0.0011541 0.11853 0.00065751 0.11918 0.10797 0 0.039136 0.0389 0 0.87114 0.23839 0.062896 0.0088508 4.1522 0.055372 6.6259e-005 0.83469 0.0051608 0.005898 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.13092 0.92444 0.90501 0.0013994 0.98689 0.5755 0.0018853 0.42757 1.8071 1.8062 16.0071 144.9911 0.00018269 -85.6329 0.62896
0.733 0.98802 5.5211e-005 3.8182 0.01204 9.6545e-006 0.0011541 0.11863 0.00065752 0.11928 0.10805 0 0.03913 0.0389 0 0.8712 0.23842 0.062905 0.008852 4.1524 0.05538 6.6268e-005 0.83469 0.005161 0.0058982 0.0013907 0.98689 0.99167 2.9991e-006 1.1996e-005 0.13092 0.92463 0.9051 0.0013994 0.98695 0.57565 0.0018852 0.42758 1.8077 1.8068 16.0071 144.9912 0.00018255 -85.6331 0.62996
0.734 0.98802 5.5211e-005 3.8182 0.01204 9.6677e-006 0.0011541 0.11872 0.00065752 0.11937 0.10814 0 0.039123 0.0389 0 0.87127 0.23844 0.062915 0.0088532 4.1526 0.055387 6.6278e-005 0.83468 0.0051612 0.0058984 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.13092 0.92481 0.90519 0.0013994 0.98702 0.57579 0.0018852 0.42759 1.8082 1.8074 16.0071 144.9912 0.00018241 -85.6334 0.63096
0.735 0.98802 5.5211e-005 3.8182 0.01204 9.6808e-006 0.0011541 0.11881 0.00065752 0.11947 0.10823 0 0.039116 0.0389 0 0.87133 0.23847 0.062925 0.0088544 4.1527 0.055394 6.6287e-005 0.83467 0.0051614 0.0058986 0.0013905 0.98689 0.99167 2.9989e-006 1.1995e-005 0.13092 0.925 0.90528 0.0013993 0.98708 0.57594 0.0018851 0.42761 1.8088 1.8079 16.0071 144.9912 0.00018226 -85.6336 0.63196
0.736 0.98802 5.5211e-005 3.8182 0.01204 9.694e-006 0.0011541 0.11891 0.00065753 0.11956 0.10832 0 0.03911 0.0389 0 0.87139 0.2385 0.062934 0.0088556 4.1529 0.055401 6.6296e-005 0.83467 0.0051616 0.0058988 0.0013905 0.98689 0.99167 2.9987e-006 1.1995e-005 0.13093 0.92518 0.90537 0.0013993 0.98715 0.57609 0.0018851 0.42762 1.8094 1.8085 16.007 144.9912 0.00018212 -85.6339 0.63296
0.737 0.98802 5.5211e-005 3.8182 0.01204 9.7072e-006 0.0011541 0.119 0.00065753 0.11965 0.1084 0 0.039103 0.0389 0 0.87145 0.23852 0.062944 0.0088569 4.1531 0.055408 6.6305e-005 0.83466 0.0051618 0.005899 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.13093 0.92536 0.90546 0.0013993 0.98722 0.57624 0.0018851 0.42763 1.8099 1.809 16.007 144.9912 0.00018198 -85.6341 0.63396
0.738 0.98802 5.5211e-005 3.8182 0.01204 9.7203e-006 0.0011541 0.11909 0.00065753 0.11975 0.10849 0 0.039096 0.0389 0 0.87151 0.23855 0.062954 0.0088581 4.1533 0.055416 6.6314e-005 0.83465 0.005162 0.0058992 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.13093 0.92554 0.90555 0.0013992 0.98728 0.57638 0.001885 0.42764 1.8105 1.8096 16.007 144.9913 0.00018183 -85.6344 0.63496
0.739 0.98802 5.5211e-005 3.8182 0.01204 9.7335e-006 0.0011541 0.11919 0.00065754 0.11984 0.10858 0 0.03909 0.0389 0 0.87157 0.23858 0.062964 0.0088593 4.1534 0.055423 6.6324e-005 0.83464 0.0051622 0.0058994 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.13093 0.92572 0.90564 0.0013992 0.98734 0.57653 0.001885 0.42766 1.811 1.8101 16.007 144.9913 0.00018169 -85.6346 0.63596
0.74 0.98802 5.521e-005 3.8182 0.01204 9.7466e-006 0.0011541 0.11928 0.00065754 0.11993 0.10866 0 0.039083 0.0389 0 0.87163 0.2386 0.062973 0.0088605 4.1536 0.05543 6.6333e-005 0.83464 0.0051624 0.0058996 0.0013902 0.98689 0.99167 2.9982e-006 1.1993e-005 0.13093 0.9259 0.90573 0.0013992 0.98741 0.57668 0.0018849 0.42767 1.8116 1.8107 16.0069 144.9913 0.00018155 -85.6349 0.63696
0.741 0.98802 5.521e-005 3.8182 0.01204 9.7598e-006 0.0011541 0.11937 0.00065754 0.12003 0.10875 0 0.039076 0.0389 0 0.87169 0.23863 0.062983 0.0088617 4.1538 0.055437 6.6342e-005 0.83463 0.0051627 0.0058998 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.13094 0.92608 0.90582 0.0013991 0.98747 0.57683 0.0018849 0.42768 1.8121 1.8112 16.0069 144.9913 0.00018141 -85.6351 0.63796
0.742 0.98802 5.521e-005 3.8182 0.01204 9.7729e-006 0.0011541 0.11947 0.00065754 0.12012 0.10884 0 0.03907 0.0389 0 0.87175 0.23866 0.062993 0.0088629 4.154 0.055445 6.6351e-005 0.83462 0.0051629 0.0059 0.0013901 0.98689 0.99167 2.9979e-006 1.1992e-005 0.13094 0.92626 0.90591 0.0013991 0.98753 0.57697 0.0018849 0.4277 1.8127 1.8118 16.0069 144.9913 0.00018127 -85.6354 0.63896
0.743 0.98802 5.521e-005 3.8182 0.01204 9.7861e-006 0.0011541 0.11956 0.00065755 0.12021 0.10892 0 0.039063 0.0389 0 0.87182 0.23869 0.063003 0.0088641 4.1541 0.055452 6.636e-005 0.83461 0.0051631 0.0059002 0.0013901 0.98689 0.99167 2.9978e-006 1.1991e-005 0.13094 0.92644 0.906 0.0013991 0.9876 0.57712 0.0018848 0.42771 1.8132 1.8123 16.0069 144.9914 0.00018113 -85.6356 0.63996
0.744 0.98802 5.521e-005 3.8182 0.01204 9.7992e-006 0.0011541 0.11965 0.00065755 0.12031 0.10901 0 0.039056 0.0389 0 0.87188 0.23871 0.063012 0.0088654 4.1543 0.055459 6.637e-005 0.83461 0.0051633 0.0059004 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.13094 0.92662 0.90609 0.001399 0.98766 0.57727 0.0018848 0.42772 1.8138 1.8129 16.0068 144.9914 0.00018099 -85.6359 0.64096
0.745 0.98802 5.521e-005 3.8182 0.01204 9.8124e-006 0.0011541 0.11975 0.00065755 0.1204 0.10909 0 0.03905 0.0389 0 0.87194 0.23874 0.063022 0.0088666 4.1545 0.055466 6.6379e-005 0.8346 0.0051635 0.0059006 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.13094 0.9268 0.90618 0.001399 0.98772 0.57741 0.0018848 0.42773 1.8143 1.8134 16.0068 144.9914 0.00018085 -85.6361 0.64196
0.746 0.98802 5.521e-005 3.8182 0.01204 9.8255e-006 0.0011541 0.11984 0.00065755 0.12049 0.10918 0 0.039043 0.0389 0 0.872 0.23877 0.063032 0.0088678 4.1547 0.055474 6.6388e-005 0.83459 0.0051637 0.0059009 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.13094 0.92698 0.90627 0.001399 0.98778 0.57756 0.0018847 0.42775 1.8148 1.814 16.0068 144.9914 0.00018072 -85.6364 0.64296
0.747 0.98802 5.521e-005 3.8182 0.01204 9.8387e-006 0.0011541 0.11993 0.00065756 0.12058 0.10927 0 0.039036 0.0389 0 0.87206 0.23879 0.063042 0.008869 4.1549 0.055481 6.6398e-005 0.83459 0.0051639 0.0059011 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.13095 0.92715 0.90635 0.001399 0.98784 0.57771 0.0018847 0.42776 1.8154 1.8145 16.0068 144.9914 0.00018058 -85.6366 0.64396
0.748 0.98802 5.521e-005 3.8182 0.01204 9.8519e-006 0.0011541 0.12002 0.00065756 0.12068 0.10935 0 0.03903 0.0389 0 0.87212 0.23882 0.063052 0.0088702 4.155 0.055488 6.6407e-005 0.83458 0.0051641 0.0059013 0.0013898 0.9869 0.99167 2.9972e-006 1.1989e-005 0.13095 0.92733 0.90644 0.0013989 0.9879 0.57785 0.0018846 0.42777 1.8159 1.8151 16.0068 144.9915 0.00018044 -85.6368 0.64496
0.749 0.98802 5.521e-005 3.8182 0.01204 9.865e-006 0.0011541 0.12012 0.00065756 0.12077 0.10944 0 0.039023 0.0389 0 0.87218 0.23885 0.063061 0.0088715 4.1552 0.055495 6.6416e-005 0.83457 0.0051643 0.0059015 0.0013897 0.9869 0.99167 2.997e-006 1.1988e-005 0.13095 0.9275 0.90653 0.0013989 0.98797 0.578 0.0018846 0.42779 1.8165 1.8156 16.0067 144.9915 0.00018031 -85.6371 0.64596
0.75 0.98802 5.521e-005 3.8182 0.01204 9.8782e-006 0.0011541 0.12021 0.00065757 0.12086 0.10953 0 0.039017 0.0389 0 0.87225 0.23888 0.063071 0.0088727 4.1554 0.055503 6.6425e-005 0.83456 0.0051645 0.0059017 0.0013897 0.9869 0.99168 2.9969e-006 1.1988e-005 0.13095 0.92768 0.90661 0.0013989 0.98802 0.57815 0.0018846 0.4278 1.817 1.8162 16.0067 144.9915 0.00018017 -85.6373 0.64696
0.751 0.98802 5.521e-005 3.8182 0.01204 9.8913e-006 0.0011541 0.1203 0.00065757 0.12095 0.10961 0 0.03901 0.0389 0 0.87231 0.2389 0.063081 0.0088739 4.1556 0.05551 6.6435e-005 0.83456 0.0051647 0.0059019 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.13095 0.92785 0.9067 0.0013988 0.98808 0.5783 0.0018845 0.42781 1.8175 1.8167 16.0067 144.9915 0.00018003 -85.6375 0.64796
0.752 0.98802 5.521e-005 3.8182 0.01204 9.9045e-006 0.0011541 0.12039 0.00065757 0.12105 0.1097 0 0.039004 0.0389 0 0.87237 0.23893 0.063091 0.0088751 4.1558 0.055517 6.6444e-005 0.83455 0.0051649 0.0059021 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.13095 0.92803 0.90679 0.0013988 0.98814 0.57844 0.0018845 0.42783 1.8181 1.8172 16.0067 144.9915 0.0001799 -85.6378 0.64896
0.753 0.98802 5.521e-005 3.8182 0.01204 9.9176e-006 0.0011541 0.12049 0.00065757 0.12114 0.10978 0 0.038997 0.0389 0 0.87243 0.23896 0.063101 0.0088764 4.156 0.055525 6.6453e-005 0.83454 0.0051652 0.0059023 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.13096 0.9282 0.90687 0.0013988 0.9882 0.57859 0.0018845 0.42784 1.8186 1.8178 16.0066 144.9916 0.00017976 -85.638 0.64996
0.754 0.98802 5.521e-005 3.8182 0.01204 9.9308e-006 0.0011541 0.12058 0.00065758 0.12123 0.10987 0 0.03899 0.0389 0 0.87249 0.23899 0.063111 0.0088776 4.1561 0.055532 6.6463e-005 0.83453 0.0051654 0.0059025 0.0013895 0.9869 0.99168 2.9964e-006 1.1986e-005 0.13096 0.92837 0.90696 0.0013988 0.98826 0.57874 0.0018844 0.42785 1.8191 1.8183 16.0066 144.9916 0.00017963 -85.6382 0.65096
0.755 0.98802 5.521e-005 3.8182 0.01204 9.9439e-006 0.0011541 0.12067 0.00065758 0.12132 0.10995 0 0.038984 0.0389 0 0.87256 0.23901 0.063121 0.0088788 4.1563 0.055539 6.6472e-005 0.83453 0.0051656 0.0059027 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.13096 0.92855 0.90704 0.0013987 0.98832 0.57888 0.0018844 0.42786 1.8197 1.8188 16.0066 144.9916 0.0001795 -85.6384 0.65196
0.756 0.98802 5.5209e-005 3.8182 0.01204 9.9571e-006 0.0011541 0.12076 0.00065758 0.12142 0.11004 0 0.038977 0.0389 0 0.87262 0.23904 0.06313 0.0088801 4.1565 0.055547 6.6481e-005 0.83452 0.0051658 0.0059029 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.13096 0.92872 0.90713 0.0013987 0.98838 0.57903 0.0018843 0.42788 1.8202 1.8194 16.0066 144.9916 0.00017936 -85.6387 0.65296
0.757 0.98802 5.5209e-005 3.8182 0.01204 9.9702e-006 0.0011541 0.12085 0.00065759 0.12151 0.11013 0 0.038971 0.0389 0 0.87268 0.23907 0.06314 0.0088813 4.1567 0.055554 6.6491e-005 0.83451 0.005166 0.0059032 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.13096 0.92889 0.90721 0.0013987 0.98843 0.57917 0.0018843 0.42789 1.8207 1.8199 16.0065 144.9916 0.00017923 -85.6389 0.65396
0.758 0.98802 5.5209e-005 3.8182 0.01204 9.9834e-006 0.0011541 0.12095 0.00065759 0.1216 0.11021 0 0.038964 0.0389 0 0.87274 0.23909 0.06315 0.0088825 4.1569 0.055561 6.65e-005 0.83451 0.0051662 0.0059034 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.13096 0.92906 0.9073 0.0013987 0.98849 0.57932 0.0018843 0.4279 1.8213 1.8204 16.0065 144.9917 0.0001791 -85.6391 0.65496
0.759 0.98802 5.5209e-005 3.8182 0.01204 9.9966e-006 0.0011541 0.12104 0.00065759 0.12169 0.1103 0 0.038958 0.0389 0 0.8728 0.23912 0.06316 0.0088837 4.1571 0.055569 6.651e-005 0.8345 0.0051664 0.0059036 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.13097 0.92923 0.90738 0.0013986 0.98855 0.57947 0.0018842 0.42792 1.8218 1.821 16.0065 144.9917 0.00017897 -85.6393 0.65596
0.76 0.98802 5.5209e-005 3.8182 0.01204 1.001e-005 0.0011541 0.12113 0.00065759 0.12178 0.11038 0 0.038951 0.0389 0 0.87287 0.23915 0.06317 0.008885 4.1572 0.055576 6.6519e-005 0.83449 0.0051666 0.0059038 0.0013892 0.98691 0.99168 2.9957e-006 1.1983e-005 0.13097 0.9294 0.90746 0.0013986 0.9886 0.57961 0.0018842 0.42793 1.8223 1.8215 16.0065 144.9917 0.00017883 -85.6395 0.65696
0.761 0.98802 5.5209e-005 3.8182 0.01204 1.0023e-005 0.0011541 0.12122 0.0006576 0.12188 0.11047 0 0.038945 0.0389 0 0.87293 0.23918 0.06318 0.0088862 4.1574 0.055583 6.6528e-005 0.83448 0.0051669 0.005904 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.13097 0.92957 0.90755 0.0013986 0.98866 0.57976 0.0018842 0.42794 1.8228 1.822 16.0064 144.9917 0.0001787 -85.6397 0.65796
0.762 0.98802 5.5209e-005 3.8182 0.01204 1.0036e-005 0.0011541 0.12131 0.0006576 0.12197 0.11055 0 0.038938 0.0389 0 0.87299 0.2392 0.06319 0.0088874 4.1576 0.055591 6.6538e-005 0.83448 0.0051671 0.0059042 0.0013891 0.98691 0.99168 2.9955e-006 1.1982e-005 0.13097 0.92974 0.90763 0.0013985 0.98871 0.57991 0.0018841 0.42795 1.8234 1.8225 16.0064 144.9917 0.00017857 -85.64 0.65896
0.763 0.98802 5.5209e-005 3.8182 0.01204 1.0049e-005 0.0011541 0.12141 0.0006576 0.12206 0.11064 0 0.038932 0.0389 0 0.87305 0.23923 0.0632 0.0088887 4.1578 0.055598 6.6547e-005 0.83447 0.0051673 0.0059044 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.13097 0.92991 0.90771 0.0013985 0.98877 0.58005 0.0018841 0.42797 1.8239 1.8231 16.0064 144.9918 0.00017844 -85.6402 0.65996
0.764 0.98802 5.5209e-005 3.8182 0.01204 1.0062e-005 0.0011541 0.1215 0.0006576 0.12215 0.11072 0 0.038925 0.0389 0 0.87311 0.23926 0.06321 0.0088899 4.158 0.055605 6.6557e-005 0.83446 0.0051675 0.0059046 0.001389 0.98691 0.99168 2.9953e-006 1.1981e-005 0.13098 0.93007 0.9078 0.0013985 0.98882 0.5802 0.0018841 0.42798 1.8244 1.8236 16.0064 144.9918 0.00017831 -85.6404 0.66096
0.765 0.98802 5.5209e-005 3.8182 0.01204 1.0075e-005 0.0011541 0.12159 0.00065761 0.12224 0.11081 0 0.038919 0.0389 0 0.87318 0.23929 0.06322 0.0088912 4.1582 0.055613 6.6566e-005 0.83445 0.0051677 0.0059049 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.13098 0.93024 0.90788 0.0013985 0.98888 0.58034 0.001884 0.42799 1.8249 1.8241 16.0063 144.9918 0.00017818 -85.6406 0.66196
0.766 0.98802 5.5209e-005 3.8182 0.01204 1.0089e-005 0.0011541 0.12168 0.00065761 0.12233 0.11089 0 0.038912 0.0389 0 0.87324 0.23931 0.06323 0.0088924 4.1584 0.05562 6.6575e-005 0.83445 0.0051679 0.0059051 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.13098 0.93041 0.90796 0.0013984 0.98893 0.58049 0.001884 0.42801 1.8254 1.8246 16.0063 144.9918 0.00017806 -85.6408 0.66296
0.767 0.98802 5.5209e-005 3.8182 0.01204 1.0102e-005 0.0011541 0.12177 0.00065761 0.12242 0.11098 0 0.038906 0.0389 0 0.8733 0.23934 0.06324 0.0088936 4.1585 0.055628 6.6585e-005 0.83444 0.0051682 0.0059053 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.13098 0.93057 0.90804 0.0013984 0.98899 0.58064 0.001884 0.42802 1.826 1.8252 16.0063 144.9918 0.00017793 -85.641 0.66396
0.768 0.98802 5.5209e-005 3.8182 0.01204 1.0115e-005 0.0011541 0.12186 0.00065762 0.12252 0.11106 0 0.038899 0.0389 0 0.87336 0.23937 0.06325 0.0088949 4.1587 0.055635 6.6594e-005 0.83443 0.0051684 0.0059055 0.0013888 0.98691 0.99168 2.9948e-006 1.1979e-005 0.13098 0.93074 0.90812 0.0013984 0.98904 0.58078 0.0018839 0.42803 1.8265 1.8257 16.0063 144.9919 0.0001778 -85.6412 0.66496
0.769 0.98802 5.5209e-005 3.8182 0.01204 1.0128e-005 0.0011541 0.12195 0.00065762 0.12261 0.11115 0 0.038893 0.0389 0 0.87343 0.2394 0.06326 0.0088961 4.1589 0.055642 6.6604e-005 0.83442 0.0051686 0.0059057 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.13098 0.9309 0.9082 0.0013984 0.98909 0.58093 0.0018839 0.42804 1.827 1.8262 16.0062 144.9919 0.00017767 -85.6414 0.66596
0.77 0.98802 5.5209e-005 3.8182 0.01204 1.0141e-005 0.0011541 0.12204 0.00065762 0.1227 0.11123 0 0.038887 0.0389 0 0.87349 0.23943 0.06327 0.0088974 4.1591 0.05565 6.6613e-005 0.83442 0.0051688 0.0059059 0.0013887 0.98691 0.99168 2.9946e-006 1.1978e-005 0.13099 0.93107 0.90828 0.0013983 0.98914 0.58107 0.0018839 0.42806 1.8275 1.8267 16.0062 144.9919 0.00017755 -85.6416 0.66696
0.771 0.98802 5.5209e-005 3.8182 0.01204 1.0154e-005 0.0011541 0.12214 0.00065762 0.12279 0.11132 0 0.03888 0.0389 0 0.87355 0.23945 0.06328 0.0088986 4.1593 0.055657 6.6623e-005 0.83441 0.005169 0.0059062 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.13099 0.93123 0.90836 0.0013983 0.9892 0.58122 0.0018838 0.42807 1.828 1.8272 16.0062 144.9919 0.00017742 -85.6418 0.66796
0.772 0.98802 5.5208e-005 3.8182 0.01204 1.0168e-005 0.0011541 0.12223 0.00065763 0.12288 0.1114 0 0.038874 0.0389 0 0.87362 0.23948 0.06329 0.0088998 4.1595 0.055665 6.6632e-005 0.8344 0.0051692 0.0059064 0.0013886 0.98691 0.99168 2.9944e-006 1.1978e-005 0.13099 0.93139 0.90844 0.0013983 0.98925 0.58137 0.0018838 0.42808 1.8285 1.8277 16.0062 144.9919 0.00017729 -85.642 0.66896
0.773 0.98802 5.5208e-005 3.8182 0.01204 1.0181e-005 0.0011541 0.12232 0.00065763 0.12297 0.11148 0 0.038867 0.0389 0 0.87368 0.23951 0.0633 0.0089011 4.1597 0.055672 6.6642e-005 0.83439 0.0051695 0.0059066 0.0013885 0.98691 0.99168 2.9943e-006 1.1977e-005 0.13099 0.93156 0.90852 0.0013983 0.9893 0.58151 0.0018838 0.4281 1.829 1.8282 16.0061 144.992 0.00017717 -85.6422 0.66996
0.774 0.98802 5.5208e-005 3.8182 0.01204 1.0194e-005 0.0011541 0.12241 0.00065763 0.12306 0.11157 0 0.038861 0.0389 0 0.87374 0.23954 0.06331 0.0089023 4.1599 0.05568 6.6651e-005 0.83439 0.0051697 0.0059068 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.13099 0.93172 0.9086 0.0013982 0.98935 0.58166 0.0018837 0.42811 1.8296 1.8288 16.0061 144.992 0.00017704 -85.6424 0.67096
0.775 0.98802 5.5208e-005 3.8182 0.01204 1.0207e-005 0.0011541 0.1225 0.00065763 0.12315 0.11165 0 0.038854 0.0389 0 0.8738 0.23956 0.06332 0.0089036 4.1601 0.055687 6.6661e-005 0.83438 0.0051699 0.005907 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.131 0.93188 0.90868 0.0013982 0.9894 0.5818 0.0018837 0.42812 1.8301 1.8293 16.0061 144.992 0.00017692 -85.6426 0.67196
0.776 0.98802 5.5208e-005 3.8182 0.01204 1.022e-005 0.0011541 0.12259 0.00065764 0.12324 0.11174 0 0.038848 0.0389 0 0.87387 0.23959 0.06333 0.0089048 4.1602 0.055694 6.667e-005 0.83437 0.0051701 0.0059073 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.131 0.93204 0.90876 0.0013982 0.98945 0.58195 0.0018837 0.42813 1.8306 1.8298 16.0061 144.992 0.00017679 -85.6428 0.67296
0.777 0.98802 5.5208e-005 3.8182 0.01204 1.0233e-005 0.0011541 0.12268 0.00065764 0.12333 0.11182 0 0.038842 0.0389 0 0.87393 0.23962 0.06334 0.0089061 4.1604 0.055702 6.668e-005 0.83436 0.0051703 0.0059075 0.0013883 0.98692 0.99169 2.9939e-006 1.1975e-005 0.131 0.9322 0.90884 0.0013982 0.9895 0.58209 0.0018836 0.42815 1.8311 1.8303 16.0061 144.992 0.00017667 -85.643 0.67396
0.778 0.98802 5.5208e-005 3.8182 0.01204 1.0246e-005 0.0011541 0.12277 0.00065764 0.12342 0.11191 0 0.038835 0.0389 0 0.87399 0.23965 0.06335 0.0089073 4.1606 0.055709 6.6689e-005 0.83436 0.0051706 0.0059077 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.131 0.93236 0.90892 0.0013981 0.98955 0.58224 0.0018836 0.42816 1.8316 1.8308 16.006 144.9921 0.00017655 -85.6432 0.67496
0.779 0.98802 5.5208e-005 3.8182 0.01204 1.026e-005 0.0011541 0.12286 0.00065764 0.12351 0.11199 0 0.038829 0.0389 0 0.87406 0.23968 0.06336 0.0089086 4.1608 0.055717 6.6699e-005 0.83435 0.0051708 0.0059079 0.0013882 0.98692 0.99169 2.9937e-006 1.1975e-005 0.131 0.93252 0.909 0.0013981 0.9896 0.58238 0.0018836 0.42817 1.8321 1.8313 16.006 144.9921 0.00017642 -85.6434 0.67596
0.78 0.98802 5.5208e-005 3.8182 0.01204 1.0273e-005 0.0011541 0.12295 0.00065765 0.1236 0.11207 0 0.038823 0.0389 0 0.87412 0.2397 0.06337 0.0089098 4.161 0.055724 6.6708e-005 0.83434 0.005171 0.0059081 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.131 0.93268 0.90908 0.0013981 0.98965 0.58253 0.0018836 0.42819 1.8326 1.8318 16.006 144.9921 0.0001763 -85.6436 0.67696
0.781 0.98802 5.5208e-005 3.8182 0.01204 1.0286e-005 0.0011541 0.12304 0.00065765 0.12369 0.11216 0 0.038816 0.0389 0 0.87418 0.23973 0.06338 0.0089111 4.1612 0.055732 6.6718e-005 0.83433 0.0051712 0.0059084 0.0013881 0.98692 0.99169 2.9935e-006 1.1974e-005 0.13101 0.93284 0.90915 0.0013981 0.9897 0.58267 0.0018835 0.4282 1.8331 1.8323 16.006 144.9921 0.00017618 -85.6438 0.67796
0.782 0.98802 5.5208e-005 3.8182 0.01204 1.0299e-005 0.0011541 0.12313 0.00065765 0.12379 0.11224 0 0.03881 0.0389 0 0.87425 0.23976 0.06339 0.0089123 4.1614 0.055739 6.6727e-005 0.83433 0.0051714 0.0059086 0.0013881 0.98692 0.99169 2.9934e-006 1.1973e-005 0.13101 0.933 0.90923 0.0013981 0.98975 0.58282 0.0018835 0.42821 1.8336 1.8328 16.0059 144.9921 0.00017606 -85.644 0.67896
0.783 0.98802 5.5208e-005 3.8182 0.01204 1.0312e-005 0.0011541 0.12322 0.00065765 0.12388 0.11233 0 0.038803 0.0389 0 0.87431 0.23979 0.0634 0.0089136 4.1616 0.055747 6.6737e-005 0.83432 0.0051717 0.0059088 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.13101 0.93316 0.90931 0.001398 0.9898 0.58296 0.0018835 0.42822 1.8341 1.8333 16.0059 144.9922 0.00017594 -85.6441 0.67996
0.784 0.98802 5.5208e-005 3.8182 0.01204 1.0325e-005 0.0011541 0.12331 0.00065766 0.12397 0.11241 0 0.038797 0.0389 0 0.87437 0.23982 0.06341 0.0089148 4.1618 0.055754 6.6747e-005 0.83431 0.0051719 0.005909 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.13101 0.93332 0.90938 0.001398 0.98984 0.58311 0.0018834 0.42824 1.8346 1.8338 16.0059 144.9922 0.00017582 -85.6443 0.68096
0.785 0.98802 5.5208e-005 3.8182 0.01204 1.0339e-005 0.0011541 0.1234 0.00065766 0.12406 0.11249 0 0.038791 0.0389 0 0.87444 0.23984 0.06342 0.0089161 4.162 0.055762 6.6756e-005 0.8343 0.0051721 0.0059092 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.13101 0.93347 0.90946 0.001398 0.98989 0.58325 0.0018834 0.42825 1.8351 1.8343 16.0059 144.9922 0.0001757 -85.6445 0.68196
0.786 0.98802 5.5208e-005 3.8182 0.01204 1.0352e-005 0.0011541 0.12349 0.00065766 0.12415 0.11258 0 0.038784 0.0389 0 0.8745 0.23987 0.06343 0.0089174 4.1622 0.055769 6.6766e-005 0.8343 0.0051723 0.0059095 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.13102 0.93363 0.90954 0.001398 0.98994 0.5834 0.0018834 0.42826 1.8356 1.8348 16.0058 144.9922 0.00017558 -85.6447 0.68296
0.787 0.98802 5.5208e-005 3.8182 0.01204 1.0365e-005 0.0011541 0.12358 0.00065766 0.12424 0.11266 0 0.038778 0.0389 0 0.87456 0.2399 0.06344 0.0089186 4.1624 0.055777 6.6775e-005 0.83429 0.0051726 0.0059097 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.13102 0.93379 0.90961 0.0013979 0.98999 0.58354 0.0018833 0.42827 1.8361 1.8353 16.0058 144.9923 0.00017546 -85.6449 0.68396
0.788 0.98802 5.5207e-005 3.8182 0.01204 1.0378e-005 0.0011541 0.12367 0.00065767 0.12432 0.11274 0 0.038772 0.0389 0 0.87463 0.23993 0.063451 0.0089199 4.1626 0.055784 6.6785e-005 0.83428 0.0051728 0.0059099 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.13102 0.93394 0.90969 0.0013979 0.99003 0.58369 0.0018833 0.42829 1.8366 1.8358 16.0058 144.9923 0.00017534 -85.6451 0.68496
0.789 0.98802 5.5207e-005 3.8182 0.01204 1.0391e-005 0.0011541 0.12376 0.00065767 0.12441 0.11283 0 0.038766 0.0389 0 0.87469 0.23996 0.063461 0.0089211 4.1628 0.055792 6.6795e-005 0.83427 0.005173 0.0059101 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.13102 0.9341 0.90977 0.0013979 0.99008 0.58383 0.0018833 0.4283 1.8371 1.8363 16.0057 144.9923 0.00017522 -85.6452 0.68596
0.79 0.98802 5.5207e-005 3.8182 0.01204 1.0404e-005 0.0011541 0.12385 0.00065767 0.1245 0.11291 0 0.038759 0.0389 0 0.87475 0.23998 0.063471 0.0089224 4.163 0.055799 6.6804e-005 0.83427 0.0051732 0.0059104 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.13102 0.93425 0.90984 0.0013979 0.99013 0.58398 0.0018833 0.42831 1.8376 1.8368 16.0057 144.9923 0.0001751 -85.6454 0.68696
0.791 0.98802 5.5207e-005 3.8182 0.01204 1.0417e-005 0.0011541 0.12394 0.00065767 0.12459 0.11299 0 0.038753 0.0389 0 0.87482 0.24001 0.063481 0.0089236 4.1632 0.055807 6.6814e-005 0.83426 0.0051735 0.0059106 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.13103 0.9344 0.90992 0.0013979 0.99017 0.58412 0.0018832 0.42833 1.8381 1.8373 16.0057 144.9923 0.00017498 -85.6456 0.68796
0.792 0.98802 5.5207e-005 3.8182 0.01204 1.0431e-005 0.0011541 0.12403 0.00065768 0.12468 0.11308 0 0.038747 0.0389 0 0.87488 0.24004 0.063491 0.0089249 4.1634 0.055815 6.6824e-005 0.83425 0.0051737 0.0059108 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.13103 0.93456 0.90999 0.0013978 0.99022 0.58427 0.0018832 0.42834 1.8386 1.8378 16.0057 144.9924 0.00017487 -85.6458 0.68896
0.793 0.98802 5.5207e-005 3.8182 0.012039 1.0444e-005 0.0011541 0.12412 0.00065768 0.12477 0.11316 0 0.03874 0.0389 0 0.87494 0.24007 0.063501 0.0089262 4.1636 0.055822 6.6833e-005 0.83424 0.0051739 0.005911 0.0013877 0.98693 0.99169 2.9923e-006 1.1969e-005 0.13103 0.93471 0.91006 0.0013978 0.99026 0.58441 0.0018832 0.42835 1.839 1.8383 16.0056 144.9924 0.00017475 -85.6459 0.68996
0.794 0.98802 5.5207e-005 3.8182 0.012039 1.0457e-005 0.0011541 0.12421 0.00065768 0.12486 0.11324 0 0.038734 0.0389 0 0.87501 0.2401 0.063511 0.0089274 4.1638 0.05583 6.6843e-005 0.83424 0.0051742 0.0059113 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.13103 0.93486 0.91014 0.0013978 0.99031 0.58456 0.0018832 0.42836 1.8395 1.8388 16.0056 144.9924 0.00017463 -85.6461 0.69096
0.795 0.98802 5.5207e-005 3.8182 0.012039 1.047e-005 0.0011541 0.1243 0.00065768 0.12495 0.11333 0 0.038728 0.0389 0 0.87507 0.24012 0.063522 0.0089287 4.164 0.055837 6.6853e-005 0.83423 0.0051744 0.0059115 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.13103 0.93502 0.91021 0.0013978 0.99035 0.5847 0.0018831 0.42838 1.84 1.8393 16.0056 144.9924 0.00017452 -85.6463 0.69196
0.796 0.98802 5.5207e-005 3.8182 0.012039 1.0483e-005 0.0011541 0.12439 0.00065769 0.12504 0.11341 0 0.038722 0.0389 0 0.87514 0.24015 0.063532 0.00893 4.1642 0.055845 6.6862e-005 0.83422 0.0051746 0.0059117 0.0013875 0.98693 0.99169 2.9921e-006 1.1968e-005 0.13103 0.93517 0.91029 0.0013978 0.9904 0.58485 0.0018831 0.42839 1.8405 1.8398 16.0056 144.9924 0.0001744 -85.6465 0.69296
0.797 0.98802 5.5207e-005 3.8182 0.012039 1.0496e-005 0.0011541 0.12448 0.00065769 0.12513 0.11349 0 0.038715 0.0389 0 0.8752 0.24018 0.063542 0.0089312 4.1644 0.055852 6.6872e-005 0.83421 0.0051748 0.0059119 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.13104 0.93532 0.91036 0.0013977 0.99044 0.58499 0.0018831 0.4284 1.841 1.8402 16.0055 144.9925 0.00017429 -85.6466 0.69396
0.798 0.98802 5.5207e-005 3.8182 0.012039 1.051e-005 0.0011541 0.12457 0.00065769 0.12522 0.11357 0 0.038709 0.0389 0 0.87526 0.24021 0.063552 0.0089325 4.1646 0.05586 6.6882e-005 0.83421 0.0051751 0.0059122 0.0013874 0.98693 0.99169 2.9919e-006 1.1967e-005 0.13104 0.93547 0.91043 0.0013977 0.99048 0.58514 0.001883 0.42841 1.8415 1.8407 16.0055 144.9925 0.00017417 -85.6468 0.69496
0.799 0.98802 5.5207e-005 3.8182 0.012039 1.0523e-005 0.0011541 0.12465 0.00065769 0.12531 0.11366 0 0.038703 0.0389 0 0.87533 0.24024 0.063562 0.0089338 4.1648 0.055868 6.6891e-005 0.8342 0.0051753 0.0059124 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.13104 0.93562 0.91051 0.0013977 0.99053 0.58528 0.001883 0.42843 1.842 1.8412 16.0055 144.9925 0.00017406 -85.647 0.69596
0.8 0.98802 5.5207e-005 3.8182 0.012039 1.0536e-005 0.0011541 0.12474 0.0006577 0.1254 0.11374 0 0.038697 0.0389 0 0.87539 0.24027 0.063573 0.008935 4.165 0.055875 6.6901e-005 0.83419 0.0051755 0.0059126 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.13104 0.93577 0.91058 0.0013977 0.99057 0.58542 0.001883 0.42844 1.8424 1.8417 16.0055 144.9925 0.00017394 -85.6471 0.69696
0.801 0.98802 5.5207e-005 3.8182 0.012039 1.0549e-005 0.0011541 0.12483 0.0006577 0.12549 0.11382 0 0.03869 0.0389 0 0.87546 0.24029 0.063583 0.0089363 4.1652 0.055883 6.6911e-005 0.83418 0.0051758 0.0059129 0.0013873 0.98693 0.99169 2.9916e-006 1.1966e-005 0.13104 0.93592 0.91065 0.0013976 0.99061 0.58557 0.001883 0.42845 1.8429 1.8422 16.0054 144.9925 0.00017383 -85.6473 0.69796
0.802 0.98802 5.5207e-005 3.8182 0.012039 1.0562e-005 0.0011541 0.12492 0.0006577 0.12557 0.11391 0 0.038684 0.0389 0 0.87552 0.24032 0.063593 0.0089376 4.1654 0.05589 6.692e-005 0.83418 0.005176 0.0059131 0.0013873 0.98693 0.99169 2.9915e-006 1.1966e-005 0.13105 0.93607 0.91072 0.0013976 0.99066 0.58571 0.0018829 0.42847 1.8434 1.8427 16.0054 144.9926 0.00017371 -85.6475 0.69896
0.803 0.98802 5.5207e-005 3.8182 0.012039 1.0575e-005 0.0011541 0.12501 0.0006577 0.12566 0.11399 0 0.038678 0.0389 0 0.87558 0.24035 0.063603 0.0089388 4.1656 0.055898 6.693e-005 0.83417 0.0051762 0.0059133 0.0013873 0.98693 0.9917 2.9914e-006 1.1966e-005 0.13105 0.93622 0.9108 0.0013976 0.9907 0.58586 0.0018829 0.42848 1.8439 1.8431 16.0054 144.9926 0.0001736 -85.6476 0.69996
0.804 0.98802 5.5206e-005 3.8182 0.012039 1.0588e-005 0.0011541 0.1251 0.00065771 0.12575 0.11407 0 0.038672 0.0389 0 0.87565 0.24038 0.063614 0.0089401 4.1658 0.055906 6.694e-005 0.83416 0.0051764 0.0059136 0.0013872 0.98693 0.9917 2.9914e-006 1.1965e-005 0.13105 0.93636 0.91087 0.0013976 0.99074 0.586 0.0018829 0.42849 1.8444 1.8436 16.0054 144.9926 0.00017349 -85.6478 0.70096
0.805 0.98802 5.5206e-005 3.8182 0.012039 1.0602e-005 0.0011541 0.12519 0.00065771 0.12584 0.11415 0 0.038666 0.0389 0 0.87571 0.24041 0.063624 0.0089414 4.166 0.055913 6.695e-005 0.83415 0.0051767 0.0059138 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.13105 0.93651 0.91094 0.0013976 0.99078 0.58615 0.0018829 0.4285 1.8448 1.8441 16.0053 144.9926 0.00017338 -85.6479 0.70196
0.806 0.98802 5.5206e-005 3.8182 0.012039 1.0615e-005 0.0011541 0.12528 0.00065771 0.12593 0.11424 0 0.038659 0.0389 0 0.87578 0.24044 0.063634 0.0089427 4.1662 0.055921 6.6959e-005 0.83415 0.0051769 0.005914 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.13105 0.93666 0.91101 0.0013975 0.99083 0.58629 0.0018828 0.42852 1.8453 1.8446 16.0053 144.9926 0.00017326 -85.6481 0.70296
0.807 0.98802 5.5206e-005 3.8182 0.012039 1.0628e-005 0.0011541 0.12536 0.00065771 0.12602 0.11432 0 0.038653 0.0389 0 0.87584 0.24046 0.063644 0.0089439 4.1664 0.055929 6.6969e-005 0.83414 0.0051771 0.0059142 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.13106 0.9368 0.91108 0.0013975 0.99087 0.58643 0.0018828 0.42853 1.8458 1.8451 16.0053 144.9927 0.00017315 -85.6483 0.70396
0.808 0.98802 5.5206e-005 3.8182 0.012039 1.0641e-005 0.0011541 0.12545 0.00065772 0.12611 0.1144 0 0.038647 0.0389 0 0.87591 0.24049 0.063655 0.0089452 4.1666 0.055936 6.6979e-005 0.83413 0.0051774 0.0059145 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.13106 0.93695 0.91115 0.0013975 0.99091 0.58658 0.0018828 0.42854 1.8463 1.8455 16.0053 144.9927 0.00017304 -85.6484 0.70496
0.809 0.98802 5.5206e-005 3.8182 0.012039 1.0654e-005 0.0011541 0.12554 0.00065772 0.12619 0.11448 0 0.038641 0.0389 0 0.87597 0.24052 0.063665 0.0089465 4.1668 0.055944 6.6989e-005 0.83412 0.0051776 0.0059147 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.13106 0.9371 0.91122 0.0013975 0.99095 0.58672 0.0018828 0.42855 1.8467 1.846 16.0052 144.9927 0.00017293 -85.6486 0.70596
0.81 0.98802 5.5206e-005 3.8182 0.012039 1.0667e-005 0.0011541 0.12563 0.00065772 0.12628 0.11456 0 0.038635 0.0389 0 0.87603 0.24055 0.063675 0.0089478 4.167 0.055952 6.6999e-005 0.83412 0.0051778 0.0059149 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.13106 0.93724 0.91129 0.0013975 0.99099 0.58686 0.0018827 0.42857 1.8472 1.8465 16.0052 144.9927 0.00017282 -85.6487 0.70696
0.811 0.98802 5.5206e-005 3.8182 0.012039 1.0681e-005 0.0011541 0.12572 0.00065772 0.12637 0.11465 0 0.038629 0.0389 0 0.8761 0.24058 0.063685 0.0089491 4.1672 0.055959 6.7008e-005 0.83411 0.0051781 0.0059152 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.13106 0.93739 0.91136 0.0013975 0.99103 0.58701 0.0018827 0.42858 1.8477 1.847 16.0052 144.9927 0.00017271 -85.6489 0.70796
0.812 0.98802 5.5206e-005 3.8182 0.012039 1.0694e-005 0.0011541 0.12581 0.00065773 0.12646 0.11473 0 0.038622 0.0389 0 0.87616 0.24061 0.063696 0.0089503 4.1674 0.055967 6.7018e-005 0.8341 0.0051783 0.0059154 0.0013869 0.98693 0.9917 2.9907e-006 1.1963e-005 0.13107 0.93753 0.91143 0.0013974 0.99107 0.58715 0.0018827 0.42859 1.8482 1.8474 16.0052 144.9928 0.0001726 -85.649 0.70896
0.813 0.98802 5.5206e-005 3.8182 0.012039 1.0707e-005 0.0011541 0.12589 0.00065773 0.12655 0.11481 0 0.038616 0.0389 0 0.87623 0.24064 0.063706 0.0089516 4.1676 0.055975 6.7028e-005 0.83409 0.0051785 0.0059156 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.13107 0.93767 0.9115 0.0013974 0.99111 0.5873 0.0018827 0.42861 1.8486 1.8479 16.0051 144.9928 0.00017249 -85.6492 0.70996
0.814 0.98802 5.5206e-005 3.8182 0.012039 1.072e-005 0.0011541 0.12598 0.00065773 0.12663 0.11489 0 0.03861 0.0389 0 0.87629 0.24066 0.063716 0.0089529 4.1678 0.055982 6.7038e-005 0.83408 0.0051788 0.0059159 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.13107 0.93782 0.91157 0.0013974 0.99115 0.58744 0.0018826 0.42862 1.8491 1.8484 16.0051 144.9928 0.00017238 -85.6493 0.71096
0.815 0.98802 5.5206e-005 3.8182 0.012039 1.0733e-005 0.0011541 0.12607 0.00065773 0.12672 0.11497 0 0.038604 0.0389 0 0.87636 0.24069 0.063727 0.0089542 4.168 0.05599 6.7048e-005 0.83408 0.005179 0.0059161 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.13107 0.93796 0.91164 0.0013974 0.99119 0.58758 0.0018826 0.42863 1.8496 1.8488 16.0051 144.9928 0.00017228 -85.6495 0.71196
0.816 0.98802 5.5206e-005 3.8182 0.012039 1.0746e-005 0.0011541 0.12616 0.00065774 0.12681 0.11505 0 0.038598 0.0389 0 0.87642 0.24072 0.063737 0.0089555 4.1682 0.055998 6.7057e-005 0.83407 0.0051793 0.0059164 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.13107 0.9381 0.91171 0.0013974 0.99123 0.58773 0.0018826 0.42864 1.85 1.8493 16.005 144.9928 0.00017217 -85.6496 0.71296
0.817 0.98802 5.5206e-005 3.8182 0.012039 1.0759e-005 0.0011541 0.12624 0.00065774 0.1269 0.11514 0 0.038592 0.0389 0 0.87649 0.24075 0.063747 0.0089567 4.1684 0.056005 6.7067e-005 0.83406 0.0051795 0.0059166 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.13108 0.93824 0.91178 0.0013973 0.99127 0.58787 0.0018826 0.42866 1.8505 1.8498 16.005 144.9929 0.00017206 -85.6498 0.71396
0.818 0.98802 5.5206e-005 3.8182 0.012039 1.0773e-005 0.0011541 0.12633 0.00065774 0.12699 0.11522 0 0.038586 0.0389 0 0.87655 0.24078 0.063758 0.008958 4.1686 0.056013 6.7077e-005 0.83405 0.0051797 0.0059168 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.13108 0.93839 0.91184 0.0013973 0.9913 0.58801 0.0018825 0.42867 1.851 1.8502 16.005 144.9929 0.00017195 -85.6499 0.71496
0.819 0.98802 5.5206e-005 3.8182 0.012039 1.0786e-005 0.0011541 0.12642 0.00065774 0.12707 0.1153 0 0.03858 0.0389 0 0.87662 0.24081 0.063768 0.0089593 4.1688 0.056021 6.7087e-005 0.83405 0.00518 0.0059171 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.13108 0.93853 0.91191 0.0013973 0.99134 0.58816 0.0018825 0.42868 1.8514 1.8507 16.005 144.9929 0.00017185 -85.6501 0.71596
0.82 0.98802 5.5205e-005 3.8182 0.012039 1.0799e-005 0.0011541 0.12651 0.00065775 0.12716 0.11538 0 0.038573 0.0389 0 0.87668 0.24084 0.063778 0.0089606 4.1691 0.056028 6.7097e-005 0.83404 0.0051802 0.0059173 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.13108 0.93867 0.91198 0.0013973 0.99138 0.5883 0.0018825 0.42869 1.8519 1.8512 16.0049 144.9929 0.00017174 -85.6502 0.71696
0.821 0.98802 5.5205e-005 3.8182 0.012039 1.0812e-005 0.0011541 0.12659 0.00065775 0.12725 0.11546 0 0.038567 0.0389 0 0.87675 0.24087 0.063789 0.0089619 4.1693 0.056036 6.7107e-005 0.83403 0.0051804 0.0059175 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.13108 0.93881 0.91205 0.0013973 0.99142 0.58844 0.0018825 0.42871 1.8523 1.8516 16.0049 144.9929 0.00017163 -85.6504 0.71796
0.822 0.98802 5.5205e-005 3.8182 0.012039 1.0825e-005 0.0011541 0.12668 0.00065775 0.12734 0.11554 0 0.038561 0.0389 0 0.87681 0.24089 0.063799 0.0089632 4.1695 0.056044 6.7117e-005 0.83402 0.0051807 0.0059178 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.13109 0.93895 0.91212 0.0013973 0.99145 0.58859 0.0018824 0.42872 1.8528 1.8521 16.0049 144.993 0.00017153 -85.6505 0.71896
0.823 0.98802 5.5205e-005 3.8182 0.012039 1.0838e-005 0.0011541 0.12677 0.00065775 0.12742 0.11562 0 0.038555 0.0389 0 0.87688 0.24092 0.06381 0.0089645 4.1697 0.056052 6.7126e-005 0.83402 0.0051809 0.005918 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.13109 0.93909 0.91218 0.0013972 0.99149 0.58873 0.0018824 0.42873 1.8533 1.8526 16.0049 144.993 0.00017142 -85.6507 0.71996
0.824 0.98802 5.5205e-005 3.8182 0.012039 1.0851e-005 0.0011541 0.12686 0.00065776 0.12751 0.11571 0 0.038549 0.0389 0 0.87694 0.24095 0.06382 0.0089657 4.1699 0.056059 6.7136e-005 0.83401 0.0051812 0.0059183 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.13109 0.93923 0.91225 0.0013972 0.99153 0.58887 0.0018824 0.42874 1.8537 1.853 16.0048 144.993 0.00017132 -85.6508 0.72096
0.825 0.98802 5.5205e-005 3.8182 0.012039 1.0865e-005 0.0011541 0.12694 0.00065776 0.1276 0.11579 0 0.038543 0.0389 0 0.87701 0.24098 0.06383 0.008967 4.1701 0.056067 6.7146e-005 0.834 0.0051814 0.0059185 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.13109 0.93936 0.91232 0.0013972 0.99157 0.58902 0.0018824 0.42876 1.8542 1.8535 16.0048 144.993 0.00017121 -85.6509 0.72196
0.826 0.98802 5.5205e-005 3.8182 0.012039 1.0878e-005 0.0011541 0.12703 0.00065776 0.12768 0.11587 0 0.038537 0.0389 0 0.87707 0.24101 0.063841 0.0089683 4.1703 0.056075 6.7156e-005 0.83399 0.0051816 0.0059187 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.13109 0.9395 0.91238 0.0013972 0.9916 0.58916 0.0018824 0.42877 1.8546 1.8539 16.0048 144.993 0.00017111 -85.6511 0.72296
0.827 0.98802 5.5205e-005 3.8182 0.012039 1.0891e-005 0.0011541 0.12712 0.00065776 0.12777 0.11595 0 0.038531 0.0389 0 0.87714 0.24104 0.063851 0.0089696 4.1705 0.056083 6.7166e-005 0.83398 0.0051819 0.005919 0.0013865 0.98694 0.9917 2.9895e-006 1.1958e-005 0.1311 0.93964 0.91245 0.0013972 0.99164 0.5893 0.0018823 0.42878 1.8551 1.8544 16.0048 144.9931 0.000171 -85.6512 0.72396
0.828 0.98802 5.5205e-005 3.8182 0.012039 1.0904e-005 0.0011541 0.1272 0.00065776 0.12786 0.11603 0 0.038525 0.0389 0 0.8772 0.24107 0.063862 0.0089709 4.1707 0.05609 6.7176e-005 0.83398 0.0051821 0.0059192 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.1311 0.93978 0.91251 0.0013972 0.99167 0.58945 0.0018823 0.42879 1.8556 1.8549 16.0047 144.9931 0.0001709 -85.6514 0.72496
0.829 0.98802 5.5205e-005 3.8182 0.012039 1.0917e-005 0.0011541 0.12729 0.00065777 0.12794 0.11611 0 0.038519 0.0389 0 0.87727 0.2411 0.063872 0.0089722 4.171 0.056098 6.7186e-005 0.83397 0.0051824 0.0059195 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.1311 0.93991 0.91258 0.0013971 0.99171 0.58959 0.0018823 0.42881 1.856 1.8553 16.0047 144.9931 0.0001708 -85.6515 0.72596
0.83 0.98802 5.5205e-005 3.8182 0.012039 1.093e-005 0.0011541 0.12738 0.00065777 0.12803 0.11619 0 0.038513 0.0389 0 0.87733 0.24112 0.063882 0.0089735 4.1712 0.056106 6.7196e-005 0.83396 0.0051826 0.0059197 0.0013864 0.98694 0.9917 2.9893e-006 1.1957e-005 0.1311 0.94005 0.91265 0.0013971 0.99175 0.58973 0.0018823 0.42882 1.8565 1.8558 16.0047 144.9931 0.00017069 -85.6516 0.72696
0.831 0.98802 5.5205e-005 3.8182 0.012039 1.0944e-005 0.0011541 0.12747 0.00065777 0.12812 0.11627 0 0.038507 0.0389 0 0.8774 0.24115 0.063893 0.0089748 4.1714 0.056114 6.7206e-005 0.83395 0.0051828 0.0059199 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.1311 0.94019 0.91271 0.0013971 0.99178 0.58987 0.0018822 0.42883 1.8569 1.8562 16.0046 144.9931 0.00017059 -85.6518 0.72796
0.832 0.98802 5.5205e-005 3.8182 0.012039 1.0957e-005 0.0011541 0.12755 0.00065777 0.12821 0.11635 0 0.038501 0.0389 0 0.87746 0.24118 0.063903 0.0089761 4.1716 0.056122 6.7216e-005 0.83395 0.0051831 0.0059202 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.13111 0.94032 0.91278 0.0013971 0.99182 0.59002 0.0018822 0.42885 1.8574 1.8567 16.0046 144.9932 0.00017049 -85.6519 0.72896
0.833 0.98802 5.5205e-005 3.8182 0.012039 1.097e-005 0.0011541 0.12764 0.00065778 0.12829 0.11643 0 0.038495 0.0389 0 0.87753 0.24121 0.063914 0.0089774 4.1718 0.056129 6.7226e-005 0.83394 0.0051833 0.0059204 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.13111 0.94046 0.91284 0.0013971 0.99185 0.59016 0.0018822 0.42886 1.8578 1.8571 16.0046 144.9932 0.00017039 -85.652 0.72996
0.834 0.98802 5.5205e-005 3.8182 0.012039 1.0983e-005 0.0011541 0.12773 0.00065778 0.12838 0.11651 0 0.038489 0.0389 0 0.8776 0.24124 0.063924 0.0089787 4.172 0.056137 6.7236e-005 0.83393 0.0051836 0.0059207 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.13111 0.94059 0.91291 0.0013971 0.99189 0.5903 0.0018822 0.42887 1.8583 1.8576 16.0046 144.9932 0.00017028 -85.6522 0.73096
0.835 0.98802 5.5205e-005 3.8182 0.012039 1.0996e-005 0.0011541 0.12781 0.00065778 0.12846 0.11659 0 0.038483 0.0389 0 0.87766 0.24127 0.063935 0.00898 4.1722 0.056145 6.7246e-005 0.83392 0.0051838 0.0059209 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.13111 0.94073 0.91297 0.001397 0.99192 0.59044 0.0018822 0.42888 1.8587 1.858 16.0045 144.9932 0.00017018 -85.6523 0.73196
0.836 0.98802 5.5204e-005 3.8182 0.012039 1.1009e-005 0.0011541 0.1279 0.00065778 0.12855 0.11667 0 0.038477 0.0389 0 0.87773 0.2413 0.063945 0.0089813 4.1725 0.056153 6.7256e-005 0.83391 0.0051841 0.0059211 0.0013862 0.98694 0.9917 2.9889e-006 1.1956e-005 0.13111 0.94086 0.91303 0.001397 0.99195 0.59059 0.0018821 0.4289 1.8592 1.8585 16.0045 144.9933 0.00017008 -85.6524 0.73296
0.837 0.98802 5.5204e-005 3.8182 0.012039 1.1022e-005 0.0011541 0.12798 0.00065779 0.12864 0.11676 0 0.038471 0.0389 0 0.87779 0.24133 0.063956 0.0089826 4.1727 0.056161 6.7266e-005 0.83391 0.0051843 0.0059214 0.0013861 0.98695 0.9917 2.9888e-006 1.1955e-005 0.13112 0.94099 0.9131 0.001397 0.99199 0.59073 0.0018821 0.42891 1.8596 1.8589 16.0045 144.9933 0.00016998 -85.6525 0.73396
0.838 0.98802 5.5204e-005 3.8182 0.012039 1.1036e-005 0.0011541 0.12807 0.00065779 0.12872 0.11684 0 0.038465 0.0389 0 0.87786 0.24136 0.063966 0.0089839 4.1729 0.056168 6.7276e-005 0.8339 0.0051846 0.0059216 0.0013861 0.98695 0.9917 2.9888e-006 1.1955e-005 0.13112 0.94113 0.91316 0.001397 0.99202 0.59087 0.0018821 0.42892 1.8601 1.8594 16.0045 144.9933 0.00016988 -85.6527 0.73496
0.839 0.98802 5.5204e-005 3.8182 0.012039 1.1049e-005 0.0011541 0.12816 0.00065779 0.12881 0.11692 0 0.038459 0.0389 0 0.87792 0.24139 0.063977 0.0089852 4.1731 0.056176 6.7286e-005 0.83389 0.0051848 0.0059219 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.13112 0.94126 0.91323 0.001397 0.99206 0.59101 0.0018821 0.42893 1.8605 1.8598 16.0044 144.9933 0.00016978 -85.6528 0.73596
0.84 0.98802 5.5204e-005 3.8182 0.012039 1.1062e-005 0.0011541 0.12824 0.00065779 0.1289 0.117 0 0.038453 0.0389 0 0.87799 0.24142 0.063987 0.0089865 4.1733 0.056184 6.7296e-005 0.83388 0.005185 0.0059221 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.13112 0.94139 0.91329 0.001397 0.99209 0.59116 0.0018821 0.42895 1.8609 1.8603 16.0044 144.9933 0.00016968 -85.6529 0.73696
0.841 0.98802 5.5204e-005 3.8182 0.012039 1.1075e-005 0.0011541 0.12833 0.00065779 0.12898 0.11708 0 0.038447 0.0389 0 0.87806 0.24144 0.063998 0.0089878 4.1735 0.056192 6.7306e-005 0.83388 0.0051853 0.0059224 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.13112 0.94152 0.91335 0.0013969 0.99212 0.5913 0.001882 0.42896 1.8614 1.8607 16.0044 144.9934 0.00016958 -85.6531 0.73796
0.842 0.98802 5.5204e-005 3.8182 0.012039 1.1088e-005 0.0011541 0.12841 0.0006578 0.12907 0.11716 0 0.038441 0.0389 0 0.87812 0.24147 0.064008 0.0089891 4.1738 0.0562 6.7316e-005 0.83387 0.0051855 0.0059226 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.13113 0.94165 0.91341 0.0013969 0.99216 0.59144 0.001882 0.42897 1.8618 1.8612 16.0043 144.9934 0.00016948 -85.6532 0.73896
0.843 0.98802 5.5204e-005 3.8182 0.012039 1.1101e-005 0.0011541 0.1285 0.0006578 0.12915 0.11724 0 0.038435 0.0389 0 0.87819 0.2415 0.064019 0.0089904 4.174 0.056208 6.7326e-005 0.83386 0.0051858 0.0059229 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.13113 0.94178 0.91348 0.0013969 0.99219 0.59158 0.001882 0.42898 1.8623 1.8616 16.0043 144.9934 0.00016939 -85.6533 0.73996
0.844 0.98802 5.5204e-005 3.8182 0.012039 1.1115e-005 0.0011541 0.12859 0.0006578 0.12924 0.11732 0 0.038429 0.0389 0 0.87825 0.24153 0.064029 0.0089917 4.1742 0.056216 6.7336e-005 0.83385 0.005186 0.0059231 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.13113 0.94191 0.91354 0.0013969 0.99222 0.59172 0.001882 0.429 1.8627 1.862 16.0043 144.9934 0.00016929 -85.6534 0.74096
0.845 0.98802 5.5204e-005 3.8182 0.012039 1.1128e-005 0.0011541 0.12867 0.0006578 0.12933 0.1174 0 0.038423 0.0389 0 0.87832 0.24156 0.06404 0.008993 4.1744 0.056223 6.7346e-005 0.83384 0.0051863 0.0059234 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.13113 0.94204 0.9136 0.0013969 0.99225 0.59187 0.001882 0.42901 1.8632 1.8625 16.0043 144.9934 0.00016919 -85.6535 0.74196
0.846 0.98802 5.5204e-005 3.8182 0.012039 1.1141e-005 0.0011541 0.12876 0.00065781 0.12941 0.11748 0 0.038417 0.0389 0 0.87839 0.24159 0.06405 0.0089943 4.1746 0.056231 6.7356e-005 0.83384 0.0051865 0.0059236 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.13113 0.94217 0.91366 0.0013969 0.99228 0.59201 0.0018819 0.42902 1.8636 1.8629 16.0042 144.9935 0.00016909 -85.6537 0.74296
0.847 0.98802 5.5204e-005 3.8182 0.012039 1.1154e-005 0.0011541 0.12884 0.00065781 0.1295 0.11756 0 0.038411 0.0389 0 0.87845 0.24162 0.064061 0.0089956 4.1748 0.056239 6.7366e-005 0.83383 0.0051868 0.0059239 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.13114 0.9423 0.91373 0.0013969 0.99232 0.59215 0.0018819 0.42903 1.864 1.8634 16.0042 144.9935 0.000169 -85.6538 0.74396
0.848 0.98802 5.5204e-005 3.8182 0.012039 1.1167e-005 0.0011541 0.12893 0.00065781 0.12958 0.11763 0 0.038405 0.0389 0 0.87852 0.24165 0.064071 0.0089969 4.1751 0.056247 6.7376e-005 0.83382 0.005187 0.0059241 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.13114 0.94243 0.91379 0.0013968 0.99235 0.59229 0.0018819 0.42905 1.8645 1.8638 16.0042 144.9935 0.0001689 -85.6539 0.74496
0.849 0.98802 5.5204e-005 3.8182 0.012039 1.118e-005 0.0011541 0.12901 0.00065781 0.12967 0.11771 0 0.0384 0.0389 0 0.87858 0.24168 0.064082 0.0089983 4.1753 0.056255 6.7386e-005 0.83381 0.0051873 0.0059244 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.13114 0.94256 0.91385 0.0013968 0.99238 0.59243 0.0018819 0.42906 1.8649 1.8642 16.0041 144.9935 0.0001688 -85.654 0.74596
0.85 0.98802 5.5204e-005 3.8182 0.012039 1.1193e-005 0.0011541 0.1291 0.00065781 0.12975 0.11779 0 0.038394 0.0389 0 0.87865 0.24171 0.064093 0.0089996 4.1755 0.056263 6.7396e-005 0.8338 0.0051875 0.0059246 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.13114 0.94269 0.91391 0.0013968 0.99241 0.59258 0.0018819 0.42907 1.8653 1.8647 16.0041 144.9935 0.00016871 -85.6541 0.74696
0.851 0.98802 5.5204e-005 3.8182 0.012039 1.1207e-005 0.0011541 0.12919 0.00065782 0.12984 0.11787 0 0.038388 0.0389 0 0.87872 0.24174 0.064103 0.0090009 4.1757 0.056271 6.7406e-005 0.8338 0.0051878 0.0059249 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.13114 0.94282 0.91397 0.0013968 0.99244 0.59272 0.0018818 0.42908 1.8658 1.8651 16.0041 144.9936 0.00016861 -85.6543 0.74796
0.852 0.98802 5.5203e-005 3.8182 0.012039 1.122e-005 0.0011541 0.12927 0.00065782 0.12992 0.11795 0 0.038382 0.0389 0 0.87878 0.24177 0.064114 0.0090022 4.176 0.056279 6.7417e-005 0.83379 0.005188 0.0059251 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.13115 0.94294 0.91403 0.0013968 0.99247 0.59286 0.0018818 0.4291 1.8662 1.8655 16.0041 144.9936 0.00016852 -85.6544 0.74896
0.853 0.98802 5.5203e-005 3.8182 0.012039 1.1233e-005 0.0011541 0.12936 0.00065782 0.13001 0.11803 0 0.038376 0.0389 0 0.87885 0.2418 0.064124 0.0090035 4.1762 0.056287 6.7427e-005 0.83378 0.0051883 0.0059254 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.13115 0.94307 0.91409 0.0013968 0.9925 0.593 0.0018818 0.42911 1.8666 1.866 16.004 144.9936 0.00016842 -85.6545 0.74996
0.854 0.98802 5.5203e-005 3.8182 0.012039 1.1246e-005 0.0011541 0.12944 0.00065782 0.13009 0.11811 0 0.03837 0.0389 0 0.87892 0.24183 0.064135 0.0090048 4.1764 0.056294 6.7437e-005 0.83377 0.0051885 0.0059256 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.13115 0.9432 0.91415 0.0013968 0.99253 0.59314 0.0018818 0.42912 1.8671 1.8664 16.004 144.9936 0.00016833 -85.6546 0.75096
0.855 0.98802 5.5203e-005 3.8182 0.012039 1.1259e-005 0.0011541 0.12953 0.00065783 0.13018 0.11819 0 0.038364 0.0389 0 0.87898 0.24185 0.064146 0.0090061 4.1766 0.056302 6.7447e-005 0.83377 0.0051888 0.0059259 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.13115 0.94332 0.91421 0.0013967 0.99256 0.59329 0.0018818 0.42913 1.8675 1.8668 16.004 144.9936 0.00016823 -85.6547 0.75196
0.856 0.98802 5.5203e-005 3.8182 0.012039 1.1272e-005 0.0011541 0.12961 0.00065783 0.13026 0.11827 0 0.038358 0.0389 0 0.87905 0.24188 0.064156 0.0090075 4.1768 0.05631 6.7457e-005 0.83376 0.005189 0.0059261 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.13115 0.94345 0.91427 0.0013967 0.99259 0.59343 0.0018818 0.42915 1.8679 1.8673 16.004 144.9937 0.00016814 -85.6548 0.75296
0.857 0.98802 5.5203e-005 3.8182 0.012039 1.1285e-005 0.0011541 0.1297 0.00065783 0.13035 0.11835 0 0.038353 0.0389 0 0.87912 0.24191 0.064167 0.0090088 4.1771 0.056318 6.7467e-005 0.83375 0.0051893 0.0059264 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.13116 0.94357 0.91433 0.0013967 0.99262 0.59357 0.0018817 0.42916 1.8684 1.8677 16.0039 144.9937 0.00016804 -85.655 0.75396
0.858 0.98802 5.5203e-005 3.8182 0.012039 1.1299e-005 0.0011541 0.12978 0.00065783 0.13043 0.11843 0 0.038347 0.0389 0 0.87918 0.24194 0.064177 0.0090101 4.1773 0.056326 6.7477e-005 0.83374 0.0051895 0.0059266 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.13116 0.9437 0.91439 0.0013967 0.99265 0.59371 0.0018817 0.42917 1.8688 1.8681 16.0039 144.9937 0.00016795 -85.6551 0.75496
0.859 0.98802 5.5203e-005 3.8182 0.012039 1.1312e-005 0.0011541 0.12987 0.00065783 0.13052 0.11851 0 0.038341 0.0389 0 0.87925 0.24197 0.064188 0.0090114 4.1775 0.056334 6.7488e-005 0.83373 0.0051898 0.0059269 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.13116 0.94382 0.91445 0.0013967 0.99268 0.59385 0.0018817 0.42918 1.8692 1.8686 16.0039 144.9937 0.00016786 -85.6552 0.75596
0.86 0.98802 5.5203e-005 3.8182 0.012039 1.1325e-005 0.0011541 0.12995 0.00065784 0.1306 0.11859 0 0.038335 0.0389 0 0.87932 0.242 0.064199 0.0090127 4.1777 0.056342 6.7498e-005 0.83373 0.0051901 0.0059271 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.13116 0.94395 0.91451 0.0013967 0.99271 0.59399 0.0018817 0.4292 1.8696 1.869 16.0038 144.9937 0.00016776 -85.6553 0.75696
0.861 0.98802 5.5203e-005 3.8182 0.012039 1.1338e-005 0.0011541 0.13004 0.00065784 0.13069 0.11866 0 0.038329 0.0389 0 0.87938 0.24203 0.064209 0.009014 4.178 0.05635 6.7508e-005 0.83372 0.0051903 0.0059274 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.13117 0.94407 0.91457 0.0013967 0.99274 0.59413 0.0018817 0.42921 1.8701 1.8694 16.0038 144.9938 0.00016767 -85.6554 0.75796
0.862 0.98802 5.5203e-005 3.8182 0.012039 1.1351e-005 0.0011541 0.13012 0.00065784 0.13077 0.11874 0 0.038323 0.0389 0 0.87945 0.24206 0.06422 0.0090154 4.1782 0.056358 6.7518e-005 0.83371 0.0051906 0.0059276 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.13117 0.94419 0.91463 0.0013966 0.99277 0.59427 0.0018816 0.42922 1.8705 1.8698 16.0038 144.9938 0.00016758 -85.6555 0.75896
0.863 0.98802 5.5203e-005 3.8182 0.012039 1.1364e-005 0.0011541 0.1302 0.00065784 0.13086 0.11882 0 0.038318 0.0389 0 0.87952 0.24209 0.064231 0.0090167 4.1784 0.056366 6.7528e-005 0.8337 0.0051908 0.0059279 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.13117 0.94432 0.91469 0.0013966 0.9928 0.59442 0.0018816 0.42923 1.8709 1.8703 16.0038 144.9938 0.00016749 -85.6556 0.75996
0.864 0.98802 5.5203e-005 3.8182 0.012039 1.1378e-005 0.0011541 0.13029 0.00065785 0.13094 0.1189 0 0.038312 0.0389 0 0.87958 0.24212 0.064241 0.009018 4.1786 0.056374 6.7538e-005 0.83369 0.0051911 0.0059281 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.13117 0.94444 0.91474 0.0013966 0.99283 0.59456 0.0018816 0.42925 1.8713 1.8707 16.0037 144.9938 0.00016739 -85.6557 0.76096
0.865 0.98802 5.5203e-005 3.8182 0.012039 1.1391e-005 0.0011541 0.13037 0.00065785 0.13103 0.11898 0 0.038306 0.0389 0 0.87965 0.24215 0.064252 0.0090193 4.1789 0.056382 6.7549e-005 0.83369 0.0051913 0.0059284 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.13117 0.94456 0.9148 0.0013966 0.99286 0.5947 0.0018816 0.42926 1.8718 1.8711 16.0037 144.9938 0.0001673 -85.6558 0.76196
0.866 0.98802 5.5203e-005 3.8182 0.012039 1.1404e-005 0.0011541 0.13046 0.00065785 0.13111 0.11906 0 0.0383 0.0389 0 0.87972 0.24218 0.064263 0.0090207 4.1791 0.05639 6.7559e-005 0.83368 0.0051916 0.0059287 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.13118 0.94468 0.91486 0.0013966 0.99288 0.59484 0.0018816 0.42927 1.8722 1.8715 16.0037 144.9939 0.00016721 -85.6559 0.76296
0.867 0.98802 5.5203e-005 3.8182 0.012038 1.1417e-005 0.0011541 0.13054 0.00065785 0.1312 0.11914 0 0.038294 0.0389 0 0.87978 0.24221 0.064273 0.009022 4.1793 0.056398 6.7569e-005 0.83367 0.0051918 0.0059289 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.13118 0.94481 0.91492 0.0013966 0.99291 0.59498 0.0018816 0.42928 1.8726 1.872 16.0036 144.9939 0.00016712 -85.656 0.76396
0.868 0.98802 5.5202e-005 3.8182 0.012038 1.143e-005 0.0011541 0.13063 0.00065785 0.13128 0.11921 0 0.038289 0.0389 0 0.87985 0.24224 0.064284 0.0090233 4.1796 0.056406 6.7579e-005 0.83366 0.0051921 0.0059292 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.13118 0.94493 0.91498 0.0013966 0.99294 0.59512 0.0018815 0.42929 1.873 1.8724 16.0036 144.9939 0.00016703 -85.6561 0.76496
0.869 0.98802 5.5202e-005 3.8182 0.012038 1.1443e-005 0.0011541 0.13071 0.00065786 0.13136 0.11929 0 0.038283 0.0389 0 0.87992 0.24227 0.064295 0.0090246 4.1798 0.056414 6.759e-005 0.83365 0.0051924 0.0059294 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.13118 0.94505 0.91503 0.0013966 0.99297 0.59526 0.0018815 0.42931 1.8735 1.8728 16.0036 144.9939 0.00016694 -85.6562 0.76596
0.87 0.98802 5.5202e-005 3.8182 0.012038 1.1456e-005 0.0011541 0.13079 0.00065786 0.13145 0.11937 0 0.038277 0.0389 0 0.87998 0.2423 0.064306 0.009026 4.18 0.056422 6.76e-005 0.83365 0.0051926 0.0059297 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.13118 0.94517 0.91509 0.0013965 0.99299 0.5954 0.0018815 0.42932 1.8739 1.8732 16.0036 144.9939 0.00016685 -85.6563 0.76696
0.871 0.98802 5.5202e-005 3.8182 0.012038 1.147e-005 0.0011541 0.13088 0.00065786 0.13153 0.11945 0 0.038271 0.0389 0 0.88005 0.24233 0.064316 0.0090273 4.1802 0.05643 6.761e-005 0.83364 0.0051929 0.0059299 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.13119 0.94529 0.91515 0.0013965 0.99302 0.59554 0.0018815 0.42933 1.8743 1.8737 16.0035 144.994 0.00016676 -85.6565 0.76796
0.872 0.98802 5.5202e-005 3.8182 0.012038 1.1483e-005 0.0011541 0.13096 0.00065786 0.13162 0.11953 0 0.038266 0.0389 0 0.88012 0.24236 0.064327 0.0090286 4.1805 0.056438 6.762e-005 0.83363 0.0051931 0.0059302 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.13119 0.94541 0.9152 0.0013965 0.99305 0.59568 0.0018815 0.42934 1.8747 1.8741 16.0035 144.994 0.00016667 -85.6566 0.76896
0.873 0.98802 5.5202e-005 3.8182 0.012038 1.1496e-005 0.0011541 0.13105 0.00065786 0.1317 0.11961 0 0.03826 0.0389 0 0.88019 0.24239 0.064338 0.0090299 4.1807 0.056446 6.7631e-005 0.83362 0.0051934 0.0059305 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.13119 0.94553 0.91526 0.0013965 0.99307 0.59583 0.0018815 0.42936 1.8751 1.8745 16.0035 144.994 0.00016658 -85.6567 0.76996
0.874 0.98802 5.5202e-005 3.8182 0.012038 1.1509e-005 0.0011541 0.13113 0.00065787 0.13178 0.11968 0 0.038254 0.0389 0 0.88025 0.24242 0.064348 0.0090313 4.1809 0.056454 6.7641e-005 0.83361 0.0051936 0.0059307 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.13119 0.94564 0.91532 0.0013965 0.9931 0.59597 0.0018814 0.42937 1.8755 1.8749 16.0034 144.994 0.00016649 -85.6568 0.77096
0.875 0.98802 5.5202e-005 3.8182 0.012038 1.1522e-005 0.0011541 0.13121 0.00065787 0.13187 0.11976 0 0.038248 0.0389 0 0.88032 0.24245 0.064359 0.0090326 4.1812 0.056462 6.7651e-005 0.83361 0.0051939 0.005931 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.1312 0.94576 0.91537 0.0013965 0.99313 0.59611 0.0018814 0.42938 1.876 1.8753 16.0034 144.994 0.00016641 -85.6569 0.77196
0.876 0.98802 5.5202e-005 3.8182 0.012038 1.1535e-005 0.0011541 0.1313 0.00065787 0.13195 0.11984 0 0.038243 0.0389 0 0.88039 0.24248 0.06437 0.0090339 4.1814 0.05647 6.7661e-005 0.8336 0.0051942 0.0059312 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.1312 0.94588 0.91543 0.0013965 0.99315 0.59625 0.0018814 0.42939 1.8764 1.8757 16.0034 144.9941 0.00016632 -85.657 0.77296
0.877 0.98802 5.5202e-005 3.8182 0.012038 1.1548e-005 0.0011541 0.13138 0.00065787 0.13203 0.11992 0 0.038237 0.0389 0 0.88046 0.24251 0.064381 0.0090353 4.1816 0.056478 6.7672e-005 0.83359 0.0051944 0.0059315 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.1312 0.946 0.91548 0.0013965 0.99318 0.59639 0.0018814 0.42941 1.8768 1.8761 16.0034 144.9941 0.00016623 -85.6571 0.77396
0.878 0.98802 5.5202e-005 3.8182 0.012038 1.1562e-005 0.0011541 0.13146 0.00065787 0.13212 0.12 0 0.038231 0.0389 0 0.88052 0.24254 0.064391 0.0090366 4.1819 0.056486 6.7682e-005 0.83358 0.0051947 0.0059318 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.1312 0.94612 0.91554 0.0013964 0.99321 0.59653 0.0018814 0.42942 1.8772 1.8766 16.0033 144.9941 0.00016614 -85.6571 0.77496
0.879 0.98802 5.5202e-005 3.8182 0.012038 1.1575e-005 0.0011541 0.13155 0.00065788 0.1322 0.12007 0 0.038225 0.0389 0 0.88059 0.24257 0.064402 0.0090379 4.1821 0.056494 6.7692e-005 0.83357 0.005195 0.005932 0.001385 0.98696 0.99171 2.9864e-006 1.1945e-005 0.1312 0.94623 0.9156 0.0013964 0.99323 0.59667 0.0018814 0.42943 1.8776 1.877 16.0033 144.9941 0.00016606 -85.6572 0.77596
0.88 0.98802 5.5202e-005 3.8182 0.012038 1.1588e-005 0.0011541 0.13163 0.00065788 0.13228 0.12015 0 0.03822 0.0389 0 0.88066 0.2426 0.064413 0.0090393 4.1823 0.056502 6.7703e-005 0.83357 0.0051952 0.0059323 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.13121 0.94635 0.91565 0.0013964 0.99326 0.59681 0.0018814 0.42944 1.878 1.8774 16.0033 144.9942 0.00016597 -85.6573 0.77696
0.881 0.98802 5.5202e-005 3.8182 0.012038 1.1601e-005 0.0011541 0.13171 0.00065788 0.13237 0.12023 0 0.038214 0.0389 0 0.88073 0.24263 0.064424 0.0090406 4.1826 0.05651 6.7713e-005 0.83356 0.0051955 0.0059325 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.13121 0.94647 0.91571 0.0013964 0.99328 0.59695 0.0018813 0.42946 1.8784 1.8778 16.0032 144.9942 0.00016588 -85.6574 0.77796
0.882 0.98802 5.5202e-005 3.8182 0.012038 1.1614e-005 0.0011541 0.1318 0.00065788 0.13245 0.12031 0 0.038208 0.0389 0 0.88079 0.24266 0.064435 0.0090419 4.1828 0.056518 6.7723e-005 0.83355 0.0051957 0.0059328 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.13121 0.94658 0.91576 0.0013964 0.99331 0.59709 0.0018813 0.42947 1.8788 1.8782 16.0032 144.9942 0.0001658 -85.6575 0.77896
0.883 0.98802 5.5202e-005 3.8182 0.012038 1.1627e-005 0.0011541 0.13188 0.00065789 0.13253 0.12038 0 0.038203 0.0389 0 0.88086 0.24269 0.064445 0.0090433 4.183 0.056526 6.7734e-005 0.83354 0.005196 0.0059331 0.001385 0.98696 0.99171 2.9861e-006 1.1944e-005 0.13121 0.9467 0.91582 0.0013964 0.99333 0.59723 0.0018813 0.42948 1.8792 1.8786 16.0032 144.9942 0.00016571 -85.6576 0.77996
0.884 0.98802 5.5201e-005 3.8182 0.012038 1.164e-005 0.0011541 0.13196 0.00065789 0.13262 0.12046 0 0.038197 0.0389 0 0.88093 0.24272 0.064456 0.0090446 4.1833 0.056535 6.7744e-005 0.83353 0.0051963 0.0059333 0.0013849 0.98696 0.99171 2.9861e-006 1.1944e-005 0.13121 0.94681 0.91587 0.0013964 0.99336 0.59737 0.0018813 0.42949 1.8797 1.879 16.0032 144.9942 0.00016562 -85.6577 0.78096
0.885 0.98802 5.5201e-005 3.8182 0.012038 1.1654e-005 0.0011541 0.13205 0.00065789 0.1327 0.12054 0 0.038191 0.0389 0 0.881 0.24275 0.064467 0.009046 4.1835 0.056543 6.7754e-005 0.83353 0.0051965 0.0059336 0.0013849 0.98696 0.99171 2.9861e-006 1.1944e-005 0.13122 0.94693 0.91592 0.0013964 0.99338 0.59751 0.0018813 0.42951 1.8801 1.8794 16.0031 144.9943 0.00016554 -85.6578 0.78196
0.886 0.98802 5.5201e-005 3.8182 0.012038 1.1667e-005 0.0011541 0.13213 0.00065789 0.13278 0.12062 0 0.038186 0.0389 0 0.88106 0.24278 0.064478 0.0090473 4.1837 0.056551 6.7765e-005 0.83352 0.0051968 0.0059339 0.0013849 0.98696 0.99171 2.986e-006 1.1944e-005 0.13122 0.94704 0.91598 0.0013964 0.99341 0.59765 0.0018813 0.42952 1.8805 1.8798 16.0031 144.9943 0.00016545 -85.6579 0.78296
0.887 0.98802 5.5201e-005 3.8182 0.012038 1.168e-005 0.0011541 0.13221 0.00065789 0.13287 0.12069 0 0.03818 0.0389 0 0.88113 0.24281 0.064489 0.0090486 4.184 0.056559 6.7775e-005 0.83351 0.0051971 0.0059341 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.13122 0.94716 0.91603 0.0013963 0.99343 0.59779 0.0018813 0.42953 1.8809 1.8802 16.0031 144.9943 0.00016537 -85.658 0.78396
0.888 0.98802 5.5201e-005 3.8182 0.012038 1.1693e-005 0.0011541 0.1323 0.0006579 0.13295 0.12077 0 0.038174 0.0389 0 0.8812 0.24284 0.0645 0.00905 4.1842 0.056567 6.7785e-005 0.8335 0.0051973 0.0059344 0.0013848 0.98696 0.99172 2.9859e-006 1.1944e-005 0.13122 0.94727 0.91609 0.0013963 0.99346 0.59793 0.0018812 0.42954 1.8813 1.8807 16.003 144.9943 0.00016528 -85.6581 0.78496
0.889 0.98802 5.5201e-005 3.8182 0.012038 1.1706e-005 0.0011541 0.13238 0.0006579 0.13303 0.12085 0 0.038169 0.0389 0 0.88127 0.24287 0.06451 0.0090513 4.1845 0.056575 6.7796e-005 0.83349 0.0051976 0.0059347 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.13123 0.94738 0.91614 0.0013963 0.99348 0.59807 0.0018812 0.42955 1.8817 1.8811 16.003 144.9943 0.0001652 -85.6582 0.78596
0.89 0.98802 5.5201e-005 3.8182 0.012038 1.1719e-005 0.0011541 0.13246 0.0006579 0.13312 0.12092 0 0.038163 0.0389 0 0.88134 0.2429 0.064521 0.0090527 4.1847 0.056583 6.7806e-005 0.83348 0.0051979 0.0059349 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.13123 0.9475 0.91619 0.0013963 0.99351 0.59821 0.0018812 0.42957 1.8821 1.8815 16.003 144.9944 0.00016512 -85.6583 0.78696
0.891 0.98802 5.5201e-005 3.8182 0.012038 1.1733e-005 0.0011541 0.13254 0.0006579 0.1332 0.121 0 0.038157 0.0389 0 0.8814 0.24293 0.064532 0.009054 4.1849 0.056591 6.7816e-005 0.83348 0.0051981 0.0059352 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.13123 0.94761 0.91625 0.0013963 0.99353 0.59835 0.0018812 0.42958 1.8825 1.8819 16.003 144.9944 0.00016503 -85.6584 0.78796
0.892 0.98802 5.5201e-005 3.8182 0.012038 1.1746e-005 0.0011541 0.13263 0.0006579 0.13328 0.12108 0 0.038152 0.0389 0 0.88147 0.24296 0.064543 0.0090554 4.1852 0.056599 6.7827e-005 0.83347 0.0051984 0.0059355 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.13123 0.94772 0.9163 0.0013963 0.99355 0.59849 0.0018812 0.42959 1.8829 1.8823 16.0029 144.9944 0.00016495 -85.6584 0.78896
0.893 0.98802 5.5201e-005 3.8182 0.012038 1.1759e-005 0.0011541 0.13271 0.00065791 0.13336 0.12116 0 0.038146 0.0389 0 0.88154 0.24299 0.064554 0.0090567 4.1854 0.056607 6.7837e-005 0.83346 0.0051987 0.0059357 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.13123 0.94783 0.91635 0.0013963 0.99358 0.59863 0.0018812 0.4296 1.8833 1.8827 16.0029 144.9944 0.00016487 -85.6585 0.78996
0.894 0.98802 5.5201e-005 3.8182 0.012038 1.1772e-005 0.0011541 0.13279 0.00065791 0.13345 0.12123 0 0.03814 0.0389 0 0.88161 0.24302 0.064565 0.009058 4.1856 0.056616 6.7848e-005 0.83345 0.0051989 0.005936 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.13124 0.94794 0.9164 0.0013963 0.9936 0.59877 0.0018812 0.42962 1.8837 1.8831 16.0029 144.9944 0.00016478 -85.6586 0.79096
0.895 0.98802 5.5201e-005 3.8182 0.012038 1.1785e-005 0.0011541 0.13287 0.00065791 0.13353 0.12131 0 0.038135 0.0389 0 0.88168 0.24305 0.064576 0.0090594 4.1859 0.056624 6.7858e-005 0.83344 0.0051992 0.0059363 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.13124 0.94806 0.91646 0.0013963 0.99362 0.59891 0.0018811 0.42963 1.8841 1.8835 16.0028 144.9945 0.0001647 -85.6587 0.79196
0.896 0.98802 5.5201e-005 3.8182 0.012038 1.1798e-005 0.0011541 0.13296 0.00065791 0.13361 0.12139 0 0.038129 0.0389 0 0.88174 0.24308 0.064586 0.0090607 4.1861 0.056632 6.7869e-005 0.83344 0.0051995 0.0059365 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.13124 0.94817 0.91651 0.0013962 0.99365 0.59905 0.0018811 0.42964 1.8845 1.8839 16.0028 144.9945 0.00016462 -85.6588 0.79296
0.897 0.98802 5.5201e-005 3.8182 0.012038 1.1811e-005 0.0011541 0.13304 0.00065791 0.13369 0.12146 0 0.038124 0.0389 0 0.88181 0.24311 0.064597 0.0090621 4.1864 0.05664 6.7879e-005 0.83343 0.0051997 0.0059368 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.13124 0.94828 0.91656 0.0013962 0.99367 0.59919 0.0018811 0.42965 1.8849 1.8843 16.0028 144.9945 0.00016454 -85.6589 0.79396
0.898 0.98802 5.5201e-005 3.8182 0.012038 1.1825e-005 0.0011541 0.13312 0.00065792 0.13377 0.12154 0 0.038118 0.0389 0 0.88188 0.24314 0.064608 0.0090634 4.1866 0.056648 6.7889e-005 0.83342 0.0052 0.0059371 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.13125 0.94839 0.91661 0.0013962 0.99369 0.59933 0.0018811 0.42967 1.8853 1.8847 16.0027 144.9945 0.00016446 -85.659 0.79496
0.899 0.98802 5.5201e-005 3.8182 0.012038 1.1838e-005 0.0011541 0.1332 0.00065792 0.13386 0.12162 0 0.038112 0.0389 0 0.88195 0.24317 0.064619 0.0090648 4.1868 0.056656 6.79e-005 0.83341 0.0052003 0.0059373 0.0013846 0.98696 0.99172 2.9854e-006 1.1941e-005 0.13125 0.9485 0.91667 0.0013962 0.99372 0.59947 0.0018811 0.42968 1.8857 1.8851 16.0027 144.9945 0.00016437 -85.659 0.79596
0.9 0.98802 5.5201e-005 3.8182 0.012038 1.1851e-005 0.0011541 0.13329 0.00065792 0.13394 0.12169 0 0.038107 0.0389 0 0.88202 0.2432 0.06463 0.0090661 4.1871 0.056665 6.791e-005 0.8334 0.0052005 0.0059376 0.0013846 0.98696 0.99172 2.9854e-006 1.1941e-005 0.13125 0.94861 0.91672 0.0013962 0.99374 0.59961 0.0018811 0.42969 1.8861 1.8855 16.0027 144.9946 0.00016429 -85.6591 0.79696
0.901 0.98802 5.52e-005 3.8182 0.012038 1.1864e-005 0.0011541 0.13337 0.00065792 0.13402 0.12177 0 0.038101 0.0389 0 0.88209 0.24323 0.064641 0.0090675 4.1873 0.056673 6.7921e-005 0.8334 0.0052008 0.0059379 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.13125 0.94872 0.91677 0.0013962 0.99376 0.59975 0.0018811 0.4297 1.8865 1.8859 16.0027 144.9946 0.00016421 -85.6592 0.79796
0.902 0.98802 5.52e-005 3.8182 0.012038 1.1877e-005 0.0011541 0.13345 0.00065792 0.1341 0.12184 0 0.038096 0.0389 0 0.88215 0.24326 0.064652 0.0090688 4.1876 0.056681 6.7931e-005 0.83339 0.0052011 0.0059381 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.13125 0.94882 0.91682 0.0013962 0.99378 0.59988 0.001881 0.42971 1.8869 1.8863 16.0026 144.9946 0.00016413 -85.6593 0.79896
0.903 0.98802 5.52e-005 3.8182 0.012038 1.189e-005 0.0011541 0.13353 0.00065793 0.13418 0.12192 0 0.03809 0.0389 0 0.88222 0.24329 0.064663 0.0090702 4.1878 0.056689 6.7942e-005 0.83338 0.0052014 0.0059384 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.13126 0.94893 0.91687 0.0013962 0.9938 0.60002 0.001881 0.42973 1.8872 1.8866 16.0026 144.9946 0.00016405 -85.6594 0.79996
0.904 0.98802 5.52e-005 3.8182 0.012038 1.1903e-005 0.0011541 0.13361 0.00065793 0.13427 0.122 0 0.038084 0.0389 0 0.88229 0.24332 0.064674 0.0090715 4.1881 0.056697 6.7952e-005 0.83337 0.0052016 0.0059387 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.13126 0.94904 0.91692 0.0013962 0.99383 0.60016 0.001881 0.42974 1.8876 1.887 16.0026 144.9946 0.00016397 -85.6595 0.80096
0.905 0.98802 5.52e-005 3.8182 0.012038 1.1917e-005 0.0011541 0.13369 0.00065793 0.13435 0.12207 0 0.038079 0.0389 0 0.88236 0.24335 0.064685 0.0090729 4.1883 0.056705 6.7963e-005 0.83336 0.0052019 0.005939 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.13126 0.94915 0.91697 0.0013962 0.99385 0.6003 0.001881 0.42975 1.888 1.8874 16.0025 144.9947 0.00016389 -85.6595 0.80196
0.906 0.98802 5.52e-005 3.8182 0.012038 1.193e-005 0.0011541 0.13378 0.00065793 0.13443 0.12215 0 0.038073 0.0389 0 0.88243 0.24338 0.064696 0.0090743 4.1885 0.056714 6.7973e-005 0.83335 0.0052022 0.0059392 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.13126 0.94926 0.91702 0.0013961 0.99387 0.60044 0.001881 0.42976 1.8884 1.8878 16.0025 144.9947 0.00016381 -85.6596 0.80296
0.907 0.98802 5.52e-005 3.8182 0.012038 1.1943e-005 0.0011541 0.13386 0.00065793 0.13451 0.12223 0 0.038068 0.0389 0 0.8825 0.24341 0.064707 0.0090756 4.1888 0.056722 6.7984e-005 0.83335 0.0052024 0.0059395 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.13127 0.94936 0.91707 0.0013961 0.99389 0.60058 0.001881 0.42978 1.8888 1.8882 16.0025 144.9947 0.00016373 -85.6597 0.80396
0.908 0.98802 5.52e-005 3.8182 0.012038 1.1956e-005 0.0011541 0.13394 0.00065794 0.13459 0.1223 0 0.038062 0.0389 0 0.88257 0.24344 0.064718 0.009077 4.189 0.05673 6.7994e-005 0.83334 0.0052027 0.0059398 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.13127 0.94947 0.91712 0.0013961 0.99391 0.60072 0.001881 0.42979 1.8892 1.8886 16.0024 144.9947 0.00016365 -85.6598 0.80496
0.909 0.98802 5.52e-005 3.8182 0.012038 1.1969e-005 0.0011541 0.13402 0.00065794 0.13467 0.12238 0 0.038057 0.0389 0 0.88263 0.24347 0.064729 0.0090783 4.1893 0.056738 6.8005e-005 0.83333 0.005203 0.00594 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.13127 0.94958 0.91717 0.0013961 0.99393 0.60086 0.001881 0.4298 1.8896 1.889 16.0024 144.9947 0.00016357 -85.6599 0.80596
0.91 0.98802 5.52e-005 3.8182 0.012038 1.1982e-005 0.0011541 0.1341 0.00065794 0.13476 0.12245 0 0.038051 0.0389 0 0.8827 0.2435 0.06474 0.0090797 4.1895 0.056747 6.8015e-005 0.83332 0.0052033 0.0059403 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.13127 0.94968 0.91722 0.0013961 0.99395 0.601 0.0018809 0.42981 1.89 1.8894 16.0024 144.9948 0.0001635 -85.6599 0.80696
0.911 0.98802 5.52e-005 3.8182 0.012038 1.1995e-005 0.0011541 0.13418 0.00065794 0.13484 0.12253 0 0.038046 0.0389 0 0.88277 0.24353 0.064751 0.009081 4.1898 0.056755 6.8026e-005 0.83331 0.0052035 0.0059406 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.13128 0.94979 0.91727 0.0013961 0.99398 0.60114 0.0018809 0.42982 1.8904 1.8898 16.0024 144.9948 0.00016342 -85.66 0.80796
0.912 0.98802 5.52e-005 3.8182 0.012038 1.2009e-005 0.0011541 0.13427 0.00065794 0.13492 0.12261 0 0.03804 0.0389 0 0.88284 0.24356 0.064762 0.0090824 4.19 0.056763 6.8036e-005 0.83331 0.0052038 0.0059409 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.13128 0.94989 0.91732 0.0013961 0.994 0.60127 0.0018809 0.42984 1.8908 1.8902 16.0023 144.9948 0.00016334 -85.6601 0.80896
0.913 0.98802 5.52e-005 3.8182 0.012038 1.2022e-005 0.0011541 0.13435 0.00065795 0.135 0.12268 0 0.038035 0.0389 0 0.88291 0.24359 0.064773 0.0090838 4.1903 0.056771 6.8047e-005 0.8333 0.0052041 0.0059411 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.13128 0.95 0.91737 0.0013961 0.99402 0.60141 0.0018809 0.42985 1.8911 1.8906 16.0023 144.9948 0.00016326 -85.6602 0.80996
0.914 0.98802 5.52e-005 3.8182 0.012038 1.2035e-005 0.0011541 0.13443 0.00065795 0.13508 0.12276 0 0.038029 0.0389 0 0.88298 0.24362 0.064784 0.0090851 4.1905 0.056779 6.8057e-005 0.83329 0.0052044 0.0059414 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.13128 0.9501 0.91742 0.0013961 0.99404 0.60155 0.0018809 0.42986 1.8915 1.8909 16.0023 144.9948 0.00016318 -85.6602 0.81096
0.915 0.98802 5.52e-005 3.8182 0.012038 1.2048e-005 0.0011541 0.13451 0.00065795 0.13516 0.12283 0 0.038024 0.0389 0 0.88305 0.24365 0.064795 0.0090865 4.1908 0.056788 6.8068e-005 0.83328 0.0052046 0.0059417 0.0013844 0.98697 0.99172 2.9847e-006 1.1939e-005 0.13128 0.95021 0.91747 0.0013961 0.99406 0.60169 0.0018809 0.42987 1.8919 1.8913 16.0022 144.9949 0.00016311 -85.6603 0.81196
0.916 0.98802 5.52e-005 3.8182 0.012038 1.2061e-005 0.0011541 0.13459 0.00065795 0.13524 0.12291 0 0.038018 0.0389 0 0.88312 0.24368 0.064806 0.0090879 4.191 0.056796 6.8078e-005 0.83327 0.0052049 0.005942 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.13129 0.95031 0.91752 0.001396 0.99408 0.60183 0.0018809 0.42989 1.8923 1.8917 16.0022 144.9949 0.00016303 -85.6604 0.81296
0.917 0.98802 5.5199e-005 3.8182 0.012038 1.2074e-005 0.0011541 0.13467 0.00065795 0.13532 0.12298 0 0.038013 0.0389 0 0.88319 0.24371 0.064817 0.0090892 4.1913 0.056804 6.8089e-005 0.83326 0.0052052 0.0059423 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.13129 0.95042 0.91757 0.001396 0.9941 0.60197 0.0018809 0.4299 1.8927 1.8921 16.0022 144.9949 0.00016295 -85.6605 0.81396
0.918 0.98802 5.5199e-005 3.8182 0.012038 1.2088e-005 0.0011541 0.13475 0.00065796 0.1354 0.12306 0 0.038007 0.0389 0 0.88325 0.24375 0.064828 0.0090906 4.1915 0.056812 6.81e-005 0.83326 0.0052055 0.0059425 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.13129 0.95052 0.91762 0.001396 0.99412 0.60211 0.0018808 0.42991 1.8931 1.8925 16.0021 144.9949 0.00016288 -85.6605 0.81496
0.919 0.98802 5.5199e-005 3.8182 0.012038 1.2101e-005 0.0011541 0.13483 0.00065796 0.13549 0.12313 0 0.038002 0.0389 0 0.88332 0.24378 0.064839 0.0090919 4.1918 0.056821 6.811e-005 0.83325 0.0052057 0.0059428 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.13129 0.95062 0.91766 0.001396 0.99414 0.60225 0.0018808 0.42992 1.8934 1.8929 16.0021 144.995 0.0001628 -85.6606 0.81596
0.92 0.98802 5.5199e-005 3.8182 0.012038 1.2114e-005 0.0011541 0.13491 0.00065796 0.13557 0.12321 0 0.037996 0.0389 0 0.88339 0.24381 0.06485 0.0090933 4.192 0.056829 6.8121e-005 0.83324 0.005206 0.0059431 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.1313 0.95073 0.91771 0.001396 0.99416 0.60238 0.0018808 0.42993 1.8938 1.8932 16.0021 144.995 0.00016273 -85.6607 0.81696
0.921 0.98802 5.5199e-005 3.8182 0.012038 1.2127e-005 0.0011541 0.13499 0.00065796 0.13565 0.12328 0 0.037991 0.0389 0 0.88346 0.24384 0.064861 0.0090947 4.1923 0.056837 6.8131e-005 0.83323 0.0052063 0.0059434 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.1313 0.95083 0.91776 0.001396 0.99418 0.60252 0.0018808 0.42995 1.8942 1.8936 16.0021 144.995 0.00016265 -85.6608 0.81796
0.922 0.98802 5.5199e-005 3.8182 0.012038 1.214e-005 0.0011541 0.13507 0.00065796 0.13573 0.12336 0 0.037985 0.0389 0 0.88353 0.24387 0.064872 0.009096 4.1925 0.056846 6.8142e-005 0.83322 0.0052066 0.0059436 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.1313 0.95093 0.91781 0.001396 0.9942 0.60266 0.0018808 0.42996 1.8946 1.894 16.002 144.995 0.00016257 -85.6608 0.81896
0.923 0.98802 5.5199e-005 3.8182 0.012038 1.2153e-005 0.0011541 0.13515 0.00065796 0.13581 0.12343 0 0.03798 0.0389 0 0.8836 0.2439 0.064883 0.0090974 4.1928 0.056854 6.8153e-005 0.83321 0.0052069 0.0059439 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.1313 0.95103 0.91786 0.001396 0.99422 0.6028 0.0018808 0.42997 1.895 1.8944 16.002 144.995 0.0001625 -85.6609 0.81996
0.924 0.98802 5.5199e-005 3.8182 0.012038 1.2166e-005 0.0011541 0.13524 0.00065797 0.13589 0.12351 0 0.037974 0.0389 0 0.88367 0.24393 0.064894 0.0090988 4.193 0.056862 6.8163e-005 0.83321 0.0052071 0.0059442 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.13131 0.95113 0.9179 0.001396 0.99424 0.60294 0.0018808 0.42998 1.8953 1.8948 16.002 144.9951 0.00016242 -85.661 0.82096
0.925 0.98802 5.5199e-005 3.8182 0.012038 1.218e-005 0.0011541 0.13532 0.00065797 0.13597 0.12358 0 0.037969 0.0389 0 0.88374 0.24396 0.064905 0.0091001 4.1933 0.05687 6.8174e-005 0.8332 0.0052074 0.0059445 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.13131 0.95124 0.91795 0.001396 0.99426 0.60308 0.0018808 0.42999 1.8957 1.8951 16.0019 144.9951 0.00016235 -85.661 0.82196
0.926 0.98802 5.5199e-005 3.8182 0.012038 1.2193e-005 0.0011541 0.1354 0.00065797 0.13605 0.12366 0 0.037964 0.0389 0 0.88381 0.24399 0.064916 0.0091015 4.1935 0.056879 6.8184e-005 0.83319 0.0052077 0.0059448 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.13131 0.95134 0.918 0.001396 0.99427 0.60321 0.0018808 0.43001 1.8961 1.8955 16.0019 144.9951 0.00016227 -85.6611 0.82296
0.927 0.98802 5.5199e-005 3.8182 0.012038 1.2206e-005 0.0011541 0.13548 0.00065797 0.13613 0.12373 0 0.037958 0.0389 0 0.88388 0.24402 0.064927 0.0091029 4.1938 0.056887 6.8195e-005 0.83318 0.005208 0.005945 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.13131 0.95144 0.91805 0.001396 0.99429 0.60335 0.0018807 0.43002 1.8965 1.8959 16.0019 144.9951 0.0001622 -85.6612 0.82396
0.928 0.98802 5.5199e-005 3.8182 0.012038 1.2219e-005 0.0011541 0.13556 0.00065797 0.13621 0.12381 0 0.037953 0.0389 0 0.88395 0.24405 0.064938 0.0091043 4.194 0.056895 6.8206e-005 0.83317 0.0052083 0.0059453 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.13131 0.95154 0.91809 0.0013959 0.99431 0.60349 0.0018807 0.43003 1.8968 1.8963 16.0018 144.9951 0.00016213 -85.6612 0.82496
0.929 0.98802 5.5199e-005 3.8182 0.012038 1.2232e-005 0.0011541 0.13564 0.00065798 0.13629 0.12388 0 0.037947 0.0389 0 0.88402 0.24408 0.064949 0.0091056 4.1943 0.056904 6.8216e-005 0.83316 0.0052085 0.0059456 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.13132 0.95164 0.91814 0.0013959 0.99433 0.60363 0.0018807 0.43004 1.8972 1.8967 16.0018 144.9952 0.00016205 -85.6613 0.82596
0.93 0.98802 5.5199e-005 3.8182 0.012038 1.2245e-005 0.0011541 0.13572 0.00065798 0.13637 0.12396 0 0.037942 0.0389 0 0.88409 0.24411 0.064961 0.009107 4.1945 0.056912 6.8227e-005 0.83316 0.0052088 0.0059459 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.13132 0.95174 0.91819 0.0013959 0.99435 0.60377 0.0018807 0.43006 1.8976 1.897 16.0018 144.9952 0.00016198 -85.6614 0.82696
0.931 0.98802 5.5199e-005 3.8182 0.012038 1.2258e-005 0.0011541 0.1358 0.00065798 0.13645 0.12403 0 0.037936 0.0389 0 0.88416 0.24414 0.064972 0.0091084 4.1948 0.05692 6.8238e-005 0.83315 0.0052091 0.0059462 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.13132 0.95184 0.91823 0.0013959 0.99437 0.6039 0.0018807 0.43007 1.898 1.8974 16.0018 144.9952 0.00016191 -85.6614 0.82796
0.932 0.98802 5.5199e-005 3.8182 0.012038 1.2272e-005 0.0011541 0.13588 0.00065798 0.13653 0.12411 0 0.037931 0.0389 0 0.88423 0.24418 0.064983 0.0091098 4.195 0.056929 6.8248e-005 0.83314 0.0052094 0.0059465 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.13132 0.95194 0.91828 0.0013959 0.99439 0.60404 0.0018807 0.43008 1.8983 1.8978 16.0017 144.9952 0.00016183 -85.6615 0.82896
0.933 0.98802 5.5198e-005 3.8182 0.012038 1.2285e-005 0.0011541 0.13596 0.00065798 0.13661 0.12418 0 0.037926 0.0389 0 0.8843 0.24421 0.064994 0.0091111 4.1953 0.056937 6.8259e-005 0.83313 0.0052097 0.0059467 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.13133 0.95204 0.91833 0.0013959 0.9944 0.60418 0.0018807 0.43009 1.8987 1.8981 16.0017 144.9952 0.00016176 -85.6616 0.82996
0.934 0.98802 5.5198e-005 3.8182 0.012038 1.2298e-005 0.0011541 0.13604 0.00065799 0.13669 0.12426 0 0.03792 0.0389 0 0.88436 0.24424 0.065005 0.0091125 4.1956 0.056945 6.827e-005 0.83312 0.00521 0.005947 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.13133 0.95213 0.91837 0.0013959 0.99442 0.60432 0.0018807 0.4301 1.8991 1.8985 16.0017 144.9953 0.00016169 -85.6616 0.83096
0.935 0.98802 5.5198e-005 3.8182 0.012038 1.2311e-005 0.0011541 0.13612 0.00065799 0.13677 0.12433 0 0.037915 0.0389 0 0.88443 0.24427 0.065016 0.0091139 4.1958 0.056954 6.828e-005 0.83311 0.0052102 0.0059473 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.13133 0.95223 0.91842 0.0013959 0.99444 0.60445 0.0018807 0.43012 1.8995 1.8989 16.0016 144.9953 0.00016162 -85.6617 0.83196
0.936 0.98802 5.5198e-005 3.8182 0.012038 1.2324e-005 0.0011541 0.1362 0.00065799 0.13685 0.12441 0 0.03791 0.0389 0 0.8845 0.2443 0.065027 0.0091153 4.1961 0.056962 6.8291e-005 0.83311 0.0052105 0.0059476 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.13133 0.95233 0.91846 0.0013959 0.99446 0.60459 0.0018806 0.43013 1.8998 1.8993 16.0016 144.9953 0.00016154 -85.6618 0.83296
0.937 0.98802 5.5198e-005 3.8182 0.012038 1.2337e-005 0.0011541 0.13628 0.00065799 0.13693 0.12448 0 0.037904 0.0389 0 0.88457 0.24433 0.065039 0.0091166 4.1963 0.05697 6.8302e-005 0.8331 0.0052108 0.0059479 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.13134 0.95243 0.91851 0.0013959 0.99448 0.60473 0.0018806 0.43014 1.9002 1.8996 16.0016 144.9953 0.00016147 -85.6618 0.83396
0.938 0.98802 5.5198e-005 3.8182 0.012038 1.235e-005 0.0011541 0.13636 0.00065799 0.13701 0.12455 0 0.037899 0.0389 0 0.88464 0.24436 0.06505 0.009118 4.1966 0.056979 6.8313e-005 0.83309 0.0052111 0.0059482 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.13134 0.95252 0.91855 0.0013959 0.99449 0.60487 0.0018806 0.43015 1.9006 1.9 16.0015 144.9953 0.0001614 -85.6619 0.83496
0.939 0.98802 5.5198e-005 3.8182 0.012038 1.2364e-005 0.0011541 0.13644 0.00065799 0.13709 0.12463 0 0.037893 0.0389 0 0.88471 0.24439 0.065061 0.0091194 4.1968 0.056987 6.8323e-005 0.83308 0.0052114 0.0059484 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.13134 0.95262 0.9186 0.0013959 0.99451 0.605 0.0018806 0.43016 1.9009 1.9004 16.0015 144.9954 0.00016133 -85.662 0.83596
0.94 0.98802 5.5198e-005 3.8182 0.012038 1.2377e-005 0.0011541 0.13651 0.000658 0.13717 0.1247 0 0.037888 0.0389 0 0.88478 0.24442 0.065072 0.0091208 4.1971 0.056996 6.8334e-005 0.83307 0.0052117 0.0059487 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.13134 0.95272 0.91864 0.0013958 0.99453 0.60514 0.0018806 0.43018 1.9013 1.9007 16.0015 144.9954 0.00016126 -85.662 0.83696
0.941 0.98802 5.5198e-005 3.8182 0.012038 1.239e-005 0.0011541 0.13659 0.000658 0.13725 0.12478 0 0.037883 0.0389 0 0.88485 0.24445 0.065083 0.0091222 4.1974 0.057004 6.8345e-005 0.83306 0.005212 0.005949 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.13135 0.95281 0.91869 0.0013958 0.99455 0.60528 0.0018806 0.43019 1.9017 1.9011 16.0015 144.9954 0.00016119 -85.6621 0.83796
0.942 0.98802 5.5198e-005 3.8182 0.012037 1.2403e-005 0.0011541 0.13667 0.000658 0.13733 0.12485 0 0.037877 0.0389 0 0.88492 0.24448 0.065094 0.0091235 4.1976 0.057012 6.8355e-005 0.83306 0.0052122 0.0059493 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.13135 0.95291 0.91873 0.0013958 0.99456 0.60542 0.0018806 0.4302 1.902 1.9015 16.0014 144.9954 0.00016112 -85.6622 0.83896
0.943 0.98802 5.5198e-005 3.8182 0.012037 1.2416e-005 0.0011541 0.13675 0.000658 0.13741 0.12492 0 0.037872 0.0389 0 0.88499 0.24452 0.065106 0.0091249 4.1979 0.057021 6.8366e-005 0.83305 0.0052125 0.0059496 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13135 0.95301 0.91878 0.0013958 0.99458 0.60555 0.0018806 0.43021 1.9024 1.9018 16.0014 144.9954 0.00016105 -85.6622 0.83996
0.944 0.98802 5.5198e-005 3.8182 0.012037 1.2429e-005 0.0011541 0.13683 0.000658 0.13749 0.125 0 0.037867 0.0389 0 0.88506 0.24455 0.065117 0.0091263 4.1981 0.057029 6.8377e-005 0.83304 0.0052128 0.0059499 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13135 0.9531 0.91882 0.0013958 0.9946 0.60569 0.0018806 0.43022 1.9028 1.9022 16.0014 144.9955 0.00016098 -85.6623 0.84096
0.945 0.98802 5.5198e-005 3.8182 0.012037 1.2442e-005 0.0011541 0.13691 0.00065801 0.13756 0.12507 0 0.037861 0.0389 0 0.88513 0.24458 0.065128 0.0091277 4.1984 0.057037 6.8388e-005 0.83303 0.0052131 0.0059502 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13135 0.9532 0.91887 0.0013958 0.99461 0.60583 0.0018806 0.43024 1.9031 1.9026 16.0013 144.9955 0.00016091 -85.6623 0.84196
0.946 0.98802 5.5198e-005 3.8182 0.012037 1.2456e-005 0.0011541 0.13699 0.00065801 0.13764 0.12515 0 0.037856 0.0389 0 0.8852 0.24461 0.065139 0.0091291 4.1987 0.057046 6.8398e-005 0.83302 0.0052134 0.0059505 0.0013839 0.98697 0.99172 2.9836e-006 1.1934e-005 0.13136 0.95329 0.91891 0.0013958 0.99463 0.60597 0.0018805 0.43025 1.9035 1.9029 16.0013 144.9955 0.00016084 -85.6624 0.84296
0.947 0.98802 5.5198e-005 3.8182 0.012037 1.2469e-005 0.0011541 0.13707 0.00065801 0.13772 0.12522 0 0.037851 0.0389 0 0.88527 0.24464 0.06515 0.0091305 4.1989 0.057054 6.8409e-005 0.83301 0.0052137 0.0059507 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.13136 0.95339 0.91896 0.0013958 0.99465 0.6061 0.0018805 0.43026 1.9039 1.9033 16.0013 144.9955 0.00016077 -85.6625 0.84396
0.948 0.98802 5.5198e-005 3.8182 0.012037 1.2482e-005 0.0011541 0.13715 0.00065801 0.1378 0.12529 0 0.037845 0.0389 0 0.88534 0.24467 0.065162 0.0091318 4.1992 0.057063 6.842e-005 0.83301 0.005214 0.005951 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.13136 0.95348 0.919 0.0013958 0.99466 0.60624 0.0018805 0.43027 1.9042 1.9037 16.0012 144.9955 0.0001607 -85.6625 0.84496
0.949 0.98802 5.5197e-005 3.8182 0.012037 1.2495e-005 0.0011541 0.13723 0.00065801 0.13788 0.12537 0 0.03784 0.0389 0 0.88541 0.2447 0.065173 0.0091332 4.1994 0.057071 6.8431e-005 0.833 0.0052143 0.0059513 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13136 0.95357 0.91904 0.0013958 0.99468 0.60638 0.0018805 0.43028 1.9046 1.904 16.0012 144.9956 0.00016063 -85.6626 0.84596
0.95 0.98802 5.5197e-005 3.8182 0.012037 1.2508e-005 0.0011541 0.13731 0.00065801 0.13796 0.12544 0 0.037835 0.0389 0 0.88549 0.24473 0.065184 0.0091346 4.1997 0.05708 6.8442e-005 0.83299 0.0052145 0.0059516 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13137 0.95367 0.91909 0.0013958 0.9947 0.60651 0.0018805 0.4303 1.9049 1.9044 16.0012 144.9956 0.00016056 -85.6626 0.84696
0.951 0.98802 5.5197e-005 3.8182 0.012037 1.2521e-005 0.0011541 0.13738 0.00065802 0.13804 0.12551 0 0.03783 0.0389 0 0.88556 0.24476 0.065195 0.009136 4.2 0.057088 6.8452e-005 0.83298 0.0052148 0.0059519 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13137 0.95376 0.91913 0.0013958 0.99471 0.60665 0.0018805 0.43031 1.9053 1.9048 16.0011 144.9956 0.00016049 -85.6627 0.84796
0.952 0.98802 5.5197e-005 3.8182 0.012037 1.2535e-005 0.0011541 0.13746 0.00065802 0.13812 0.12559 0 0.037824 0.0389 0 0.88563 0.2448 0.065207 0.0091374 4.2002 0.057096 6.8463e-005 0.83297 0.0052151 0.0059522 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.13137 0.95385 0.91917 0.0013958 0.99473 0.60679 0.0018805 0.43032 1.9057 1.9051 16.0011 144.9956 0.00016042 -85.6628 0.84896
0.953 0.98802 5.5197e-005 3.8182 0.012037 1.2548e-005 0.0011541 0.13754 0.00065802 0.1382 0.12566 0 0.037819 0.0389 0 0.8857 0.24483 0.065218 0.0091388 4.2005 0.057105 6.8474e-005 0.83296 0.0052154 0.0059525 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.13137 0.95395 0.91922 0.0013958 0.99474 0.60692 0.0018805 0.43033 1.906 1.9055 16.0011 144.9956 0.00016036 -85.6628 0.84996
0.954 0.98802 5.5197e-005 3.8182 0.012037 1.2561e-005 0.0011541 0.13762 0.00065802 0.13827 0.12573 0 0.037814 0.0389 0 0.88577 0.24486 0.065229 0.0091402 4.2008 0.057113 6.8485e-005 0.83296 0.0052157 0.0059528 0.0013838 0.98698 0.99172 2.9834e-006 1.1933e-005 0.13138 0.95404 0.91926 0.0013957 0.99476 0.60706 0.0018805 0.43034 1.9064 1.9058 16.0011 144.9957 0.00016029 -85.6629 0.85096
0.955 0.98802 5.5197e-005 3.8182 0.012037 1.2574e-005 0.0011541 0.1377 0.00065802 0.13835 0.12581 0 0.037808 0.0389 0 0.88584 0.24489 0.06524 0.0091416 4.201 0.057122 6.8496e-005 0.83295 0.005216 0.0059531 0.0013837 0.98698 0.99172 2.9834e-006 1.1933e-005 0.13138 0.95413 0.9193 0.0013957 0.99477 0.6072 0.0018805 0.43036 1.9067 1.9062 16.001 144.9957 0.00016022 -85.6629 0.85196
0.956 0.98802 5.5197e-005 3.8182 0.012037 1.2587e-005 0.0011541 0.13778 0.00065803 0.13843 0.12588 0 0.037803 0.0389 0 0.88591 0.24492 0.065252 0.009143 4.2013 0.05713 6.8506e-005 0.83294 0.0052163 0.0059534 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.13138 0.95422 0.91935 0.0013957 0.99479 0.60733 0.0018805 0.43037 1.9071 1.9066 16.001 144.9957 0.00016015 -85.663 0.85296
0.957 0.98802 5.5197e-005 3.8182 0.012037 1.26e-005 0.0011541 0.13786 0.00065803 0.13851 0.12595 0 0.037798 0.0389 0 0.88598 0.24495 0.065263 0.0091444 4.2016 0.057139 6.8517e-005 0.83293 0.0052166 0.0059537 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.13138 0.95432 0.91939 0.0013957 0.99481 0.60747 0.0018804 0.43038 1.9074 1.9069 16.001 144.9957 0.00016009 -85.663 0.85396
0.958 0.98802 5.5197e-005 3.8182 0.012037 1.2613e-005 0.0011541 0.13793 0.00065803 0.13859 0.12603 0 0.037793 0.0389 0 0.88605 0.24498 0.065274 0.0091457 4.2018 0.057147 6.8528e-005 0.83292 0.0052169 0.005954 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.13139 0.95441 0.91943 0.0013957 0.99482 0.60761 0.0018804 0.43039 1.9078 1.9073 16.0009 144.9958 0.00016002 -85.6631 0.85496
0.959 0.98802 5.5197e-005 3.8182 0.012037 1.2627e-005 0.0011541 0.13801 0.00065803 0.13867 0.1261 0 0.037787 0.0389 0 0.88612 0.24501 0.065286 0.0091471 4.2021 0.057156 6.8539e-005 0.83291 0.0052172 0.0059542 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13139 0.9545 0.91947 0.0013957 0.99484 0.60774 0.0018804 0.4304 1.9082 1.9076 16.0009 144.9958 0.00015995 -85.6631 0.85596
0.96 0.98802 5.5197e-005 3.8182 0.012037 1.264e-005 0.0011541 0.13809 0.00065803 0.13874 0.12617 0 0.037782 0.0389 0 0.88619 0.24505 0.065297 0.0091485 4.2024 0.057164 6.855e-005 0.8329 0.0052175 0.0059545 0.0013836 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13139 0.95459 0.91952 0.0013957 0.99485 0.60788 0.0018804 0.43042 1.9085 1.908 16.0009 144.9958 0.00015989 -85.6632 0.85696
0.961 0.98802 5.5197e-005 3.8182 0.012037 1.2653e-005 0.0011541 0.13817 0.00065803 0.13882 0.12625 0 0.037777 0.0389 0 0.88626 0.24508 0.065308 0.0091499 4.2026 0.057172 6.8561e-005 0.8329 0.0052178 0.0059548 0.0013836 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13139 0.95468 0.91956 0.0013957 0.99487 0.60802 0.0018804 0.43043 1.9089 1.9083 16.0008 144.9958 0.00015982 -85.6633 0.85796
0.962 0.98802 5.5197e-005 3.8182 0.012037 1.2666e-005 0.0011541 0.13825 0.00065804 0.1389 0.12632 0 0.037772 0.0389 0 0.88633 0.24511 0.065319 0.0091513 4.2029 0.057181 6.8572e-005 0.83289 0.0052181 0.0059551 0.0013836 0.98698 0.99173 2.9832e-006 1.1933e-005 0.1314 0.95477 0.9196 0.0013957 0.99488 0.60815 0.0018804 0.43044 1.9092 1.9087 16.0008 144.9958 0.00015975 -85.6633 0.85896
0.963 0.98802 5.5197e-005 3.8182 0.012037 1.2679e-005 0.0011541 0.13833 0.00065804 0.13898 0.12639 0 0.037767 0.0389 0 0.8864 0.24514 0.065331 0.0091527 4.2032 0.057189 6.8582e-005 0.83288 0.0052184 0.0059554 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.1314 0.95486 0.91964 0.0013957 0.9949 0.60829 0.0018804 0.43045 1.9096 1.909 16.0008 144.9959 0.00015969 -85.6634 0.85996
0.964 0.98802 5.5197e-005 3.8182 0.012037 1.2692e-005 0.0011541 0.1384 0.00065804 0.13906 0.12646 0 0.037761 0.0389 0 0.88647 0.24517 0.065342 0.0091541 4.2034 0.057198 6.8593e-005 0.83287 0.0052186 0.0059557 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.1314 0.95495 0.91968 0.0013957 0.99491 0.60843 0.0018804 0.43046 1.9099 1.9094 16.0007 144.9959 0.00015962 -85.6634 0.86096
0.965 0.98802 5.5196e-005 3.8182 0.012037 1.2705e-005 0.0011541 0.13848 0.00065804 0.13913 0.12654 0 0.037756 0.0389 0 0.88654 0.2452 0.065353 0.0091555 4.2037 0.057206 6.8604e-005 0.83286 0.0052189 0.005956 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.1314 0.95504 0.91973 0.0013957 0.99493 0.60856 0.0018804 0.43048 1.9103 1.9097 16.0007 144.9959 0.00015956 -85.6635 0.86196
0.966 0.98802 5.5196e-005 3.8182 0.012037 1.2719e-005 0.0011541 0.13856 0.00065804 0.13921 0.12661 0 0.037751 0.0389 0 0.88662 0.24523 0.065365 0.0091569 4.204 0.057215 6.8615e-005 0.83285 0.0052192 0.0059563 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13141 0.95513 0.91977 0.0013957 0.99494 0.6087 0.0018804 0.43049 1.9106 1.9101 16.0007 144.9959 0.00015949 -85.6635 0.86296
0.967 0.98802 5.5196e-005 3.8182 0.012037 1.2732e-005 0.0011541 0.13864 0.00065804 0.13929 0.12668 0 0.037746 0.0389 0 0.88669 0.24527 0.065376 0.0091583 4.2042 0.057223 6.8626e-005 0.83285 0.0052195 0.0059566 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13141 0.95522 0.91981 0.0013957 0.99496 0.60884 0.0018804 0.4305 1.911 1.9105 16.0006 144.9959 0.00015943 -85.6636 0.86396
0.968 0.98802 5.5196e-005 3.8182 0.012037 1.2745e-005 0.0011541 0.13871 0.00065805 0.13937 0.12675 0 0.037741 0.0389 0 0.88676 0.2453 0.065387 0.0091597 4.2045 0.057232 6.8637e-005 0.83284 0.0052198 0.0059569 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13141 0.9553 0.91985 0.0013957 0.99497 0.60897 0.0018804 0.43051 1.9113 1.9108 16.0006 144.996 0.00015936 -85.6636 0.86496
0.969 0.98802 5.5196e-005 3.8182 0.012037 1.2758e-005 0.0011541 0.13879 0.00065805 0.13945 0.12683 0 0.037735 0.0389 0 0.88683 0.24533 0.065399 0.0091611 4.2048 0.05724 6.8648e-005 0.83283 0.0052201 0.0059572 0.0013835 0.98698 0.99173 2.983e-006 1.1932e-005 0.13141 0.95539 0.91989 0.0013956 0.99498 0.60911 0.0018803 0.43052 1.9117 1.9112 16.0006 144.996 0.0001593 -85.6637 0.86596
0.97 0.98802 5.5196e-005 3.8182 0.012037 1.2771e-005 0.0011541 0.13887 0.00065805 0.13952 0.1269 0 0.03773 0.0389 0 0.8869 0.24536 0.06541 0.0091625 4.2051 0.057249 6.8659e-005 0.83282 0.0052204 0.0059575 0.0013835 0.98698 0.99173 2.9829e-006 1.1932e-005 0.13142 0.95548 0.91993 0.0013956 0.995 0.60924 0.0018803 0.43054 1.912 1.9115 16.0006 144.996 0.00015923 -85.6637 0.86696
0.971 0.98802 5.5196e-005 3.8182 0.012037 1.2784e-005 0.0011541 0.13895 0.00065805 0.1396 0.12697 0 0.037725 0.0389 0 0.88697 0.24539 0.065422 0.0091639 4.2053 0.057258 6.867e-005 0.83281 0.0052207 0.0059578 0.0013835 0.98698 0.99173 2.9829e-006 1.1932e-005 0.13142 0.95557 0.91997 0.0013956 0.99501 0.60938 0.0018803 0.43055 1.9124 1.9119 16.0005 144.996 0.00015917 -85.6638 0.86796
0.972 0.98802 5.5196e-005 3.8182 0.012037 1.2797e-005 0.0011541 0.13902 0.00065805 0.13968 0.12704 0 0.03772 0.0389 0 0.88704 0.24542 0.065433 0.0091653 4.2056 0.057266 6.8681e-005 0.8328 0.005221 0.0059581 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.13142 0.95566 0.92001 0.0013956 0.99503 0.60952 0.0018803 0.43056 1.9127 1.9122 16.0005 144.996 0.00015911 -85.6638 0.86896
0.973 0.98802 5.5196e-005 3.8182 0.012037 1.2811e-005 0.0011541 0.1391 0.00065806 0.13976 0.12712 0 0.037715 0.0389 0 0.88711 0.24545 0.065444 0.0091667 4.2059 0.057275 6.8691e-005 0.83279 0.0052213 0.0059584 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.13142 0.95574 0.92005 0.0013956 0.99504 0.60965 0.0018803 0.43057 1.9131 1.9125 16.0005 144.9961 0.00015904 -85.6639 0.86996
0.974 0.98802 5.5196e-005 3.8182 0.012037 1.2824e-005 0.0011541 0.13918 0.00065806 0.13983 0.12719 0 0.037709 0.0389 0 0.88718 0.24549 0.065456 0.0091681 4.2061 0.057283 6.8702e-005 0.83279 0.0052216 0.0059587 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13143 0.95583 0.92009 0.0013956 0.99505 0.60979 0.0018803 0.43058 1.9134 1.9129 16.0004 144.9961 0.00015898 -85.6639 0.87096
0.975 0.98802 5.5196e-005 3.8182 0.012037 1.2837e-005 0.0011541 0.13926 0.00065806 0.13991 0.12726 0 0.037704 0.0389 0 0.88726 0.24552 0.065467 0.0091695 4.2064 0.057292 6.8713e-005 0.83278 0.0052219 0.005959 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13143 0.95592 0.92013 0.0013956 0.99507 0.60992 0.0018803 0.4306 1.9138 1.9132 16.0004 144.9961 0.00015892 -85.664 0.87196
0.976 0.98802 5.5196e-005 3.8182 0.012037 1.285e-005 0.0011541 0.13933 0.00065806 0.13999 0.12733 0 0.037699 0.0389 0 0.88733 0.24555 0.065478 0.0091709 4.2067 0.0573 6.8724e-005 0.83277 0.0052222 0.0059593 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13143 0.956 0.92017 0.0013956 0.99508 0.61006 0.0018803 0.43061 1.9141 1.9136 16.0004 144.9961 0.00015885 -85.664 0.87296
0.977 0.98802 5.5196e-005 3.8182 0.012037 1.2863e-005 0.0011541 0.13941 0.00065806 0.14006 0.1274 0 0.037694 0.0389 0 0.8874 0.24558 0.06549 0.0091723 4.207 0.057309 6.8735e-005 0.83276 0.0052225 0.0059596 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13143 0.95609 0.92021 0.0013956 0.9951 0.61019 0.0018803 0.43062 1.9145 1.9139 16.0003 144.9961 0.00015879 -85.6641 0.87396
0.978 0.98802 5.5196e-005 3.8182 0.012037 1.2876e-005 0.0011541 0.13949 0.00065806 0.14014 0.12748 0 0.037689 0.0389 0 0.88747 0.24561 0.065501 0.0091738 4.2072 0.057317 6.8746e-005 0.83275 0.0052228 0.0059599 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13144 0.95617 0.92025 0.0013956 0.99511 0.61033 0.0018803 0.43063 1.9148 1.9143 16.0003 144.9962 0.00015873 -85.6641 0.87496
0.979 0.98802 5.5196e-005 3.8182 0.012037 1.2889e-005 0.0011541 0.13957 0.00065807 0.14022 0.12755 0 0.037684 0.0389 0 0.88754 0.24564 0.065513 0.0091752 4.2075 0.057326 6.8757e-005 0.83274 0.0052231 0.0059602 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13144 0.95626 0.92029 0.0013956 0.99512 0.61047 0.0018803 0.43064 1.9151 1.9146 16.0003 144.9962 0.00015867 -85.6642 0.87596
0.98 0.98802 5.5196e-005 3.8182 0.012037 1.2903e-005 0.0011541 0.13964 0.00065807 0.1403 0.12762 0 0.037679 0.0389 0 0.88761 0.24568 0.065524 0.0091766 4.2078 0.057334 6.8768e-005 0.83273 0.0052234 0.0059605 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13144 0.95635 0.92033 0.0013956 0.99514 0.6106 0.0018803 0.43065 1.9155 1.915 16.0002 144.9962 0.0001586 -85.6642 0.87696
0.981 0.98802 5.5195e-005 3.8182 0.012037 1.2916e-005 0.0011541 0.13972 0.00065807 0.14037 0.12769 0 0.037673 0.0389 0 0.88768 0.24571 0.065536 0.009178 4.2081 0.057343 6.8779e-005 0.83273 0.0052237 0.0059608 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13144 0.95643 0.92037 0.0013956 0.99515 0.61074 0.0018803 0.43067 1.9158 1.9153 16.0002 144.9962 0.00015854 -85.6642 0.87796
0.982 0.98802 5.5195e-005 3.8182 0.012037 1.2929e-005 0.0011541 0.1398 0.00065807 0.14045 0.12776 0 0.037668 0.0389 0 0.88776 0.24574 0.065547 0.0091794 4.2083 0.057352 6.879e-005 0.83272 0.005224 0.0059611 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13145 0.95652 0.92041 0.0013956 0.99516 0.61087 0.0018802 0.43068 1.9162 1.9157 16.0002 144.9962 0.00015848 -85.6643 0.87896
0.983 0.98802 5.5195e-005 3.8182 0.012037 1.2942e-005 0.0011541 0.13987 0.00065807 0.14053 0.12784 0 0.037663 0.0389 0 0.88783 0.24577 0.065558 0.0091808 4.2086 0.05736 6.8801e-005 0.83271 0.0052243 0.0059614 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13145 0.9566 0.92045 0.0013956 0.99518 0.61101 0.0018802 0.43069 1.9165 1.916 16.0001 144.9963 0.00015842 -85.6643 0.87996
0.984 0.98802 5.5195e-005 3.8182 0.012037 1.2955e-005 0.0011541 0.13995 0.00065807 0.1406 0.12791 0 0.037658 0.0389 0 0.8879 0.2458 0.06557 0.0091822 4.2089 0.057369 6.8812e-005 0.8327 0.0052246 0.0059617 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13145 0.95668 0.92049 0.0013956 0.99519 0.61114 0.0018802 0.4307 1.9168 1.9163 16.0001 144.9963 0.00015836 -85.6644 0.88096
0.985 0.98802 5.5195e-005 3.8182 0.012037 1.2968e-005 0.0011541 0.14003 0.00065808 0.14068 0.12798 0 0.037653 0.0389 0 0.88797 0.24583 0.065581 0.0091836 4.2092 0.057377 6.8823e-005 0.83269 0.0052249 0.005962 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13145 0.95677 0.92053 0.0013956 0.9952 0.61128 0.0018802 0.43071 1.9172 1.9167 16.0001 144.9963 0.0001583 -85.6644 0.88196
0.986 0.98802 5.5195e-005 3.8182 0.012037 1.2981e-005 0.0011541 0.1401 0.00065808 0.14076 0.12805 0 0.037648 0.0389 0 0.88804 0.24587 0.065593 0.009185 4.2094 0.057386 6.8834e-005 0.83268 0.0052252 0.0059623 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.13146 0.95685 0.92057 0.0013955 0.99521 0.61141 0.0018802 0.43073 1.9175 1.917 16 144.9963 0.00015823 -85.6645 0.88296
0.987 0.98802 5.5195e-005 3.8182 0.012037 1.2995e-005 0.0011541 0.14018 0.00065808 0.14083 0.12812 0 0.037643 0.0389 0 0.88811 0.2459 0.065604 0.0091864 4.2097 0.057395 6.8845e-005 0.83267 0.0052256 0.0059626 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.13146 0.95693 0.92061 0.0013955 0.99523 0.61155 0.0018802 0.43074 1.9179 1.9174 16 144.9963 0.00015817 -85.6645 0.88396
0.988 0.98802 5.5195e-005 3.8182 0.012037 1.3008e-005 0.0011541 0.14026 0.00065808 0.14091 0.12819 0 0.037638 0.0389 0 0.88819 0.24593 0.065616 0.0091879 4.21 0.057403 6.8856e-005 0.83267 0.0052259 0.005963 0.0013833 0.98698 0.99173 2.9825e-006 1.193e-005 0.13146 0.95702 0.92064 0.0013955 0.99524 0.61168 0.0018802 0.43075 1.9182 1.9177 16 144.9964 0.00015811 -85.6646 0.88496
0.989 0.98802 5.5195e-005 3.8182 0.012037 1.3021e-005 0.0011541 0.14033 0.00065808 0.14099 0.12826 0 0.037633 0.0389 0 0.88826 0.24596 0.065627 0.0091893 4.2103 0.057412 6.8867e-005 0.83266 0.0052262 0.0059633 0.0013833 0.98698 0.99173 2.9825e-006 1.193e-005 0.13146 0.9571 0.92068 0.0013955 0.99525 0.61182 0.0018802 0.43076 1.9185 1.918 15.9999 144.9964 0.00015805 -85.6646 0.88596
0.99 0.98802 5.5195e-005 3.8182 0.012037 1.3034e-005 0.0011541 0.14041 0.00065808 0.14106 0.12834 0 0.037628 0.0389 0 0.88833 0.24599 0.065639 0.0091907 4.2106 0.05742 6.8878e-005 0.83265 0.0052265 0.0059636 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.13147 0.95718 0.92072 0.0013955 0.99526 0.61195 0.0018802 0.43077 1.9189 1.9184 15.9999 144.9964 0.00015799 -85.6647 0.88696
0.991 0.98802 5.5195e-005 3.8182 0.012037 1.3047e-005 0.0011541 0.14048 0.00065809 0.14114 0.12841 0 0.037623 0.0389 0 0.8884 0.24603 0.06565 0.0091921 4.2108 0.057429 6.8889e-005 0.83264 0.0052268 0.0059639 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.13147 0.95727 0.92076 0.0013955 0.99528 0.61209 0.0018802 0.43078 1.9192 1.9187 15.9999 144.9964 0.00015793 -85.6647 0.88796
0.992 0.98802 5.5195e-005 3.8182 0.012037 1.306e-005 0.0011541 0.14056 0.00065809 0.14121 0.12848 0 0.037617 0.0389 0 0.88847 0.24606 0.065662 0.0091935 4.2111 0.057438 6.89e-005 0.83263 0.0052271 0.0059642 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.13147 0.95735 0.9208 0.0013955 0.99529 0.61222 0.0018802 0.4308 1.9196 1.919 15.9999 144.9964 0.00015787 -85.6647 0.88896
0.993 0.98802 5.5195e-005 3.8182 0.012037 1.3073e-005 0.0011541 0.14064 0.00065809 0.14129 0.12855 0 0.037612 0.0389 0 0.88854 0.24609 0.065673 0.0091949 4.2114 0.057446 6.8912e-005 0.83262 0.0052274 0.0059645 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.13147 0.95743 0.92083 0.0013955 0.9953 0.61236 0.0018802 0.43081 1.9199 1.9194 15.9998 144.9965 0.00015781 -85.6648 0.88996
0.994 0.98802 5.5195e-005 3.8182 0.012037 1.3087e-005 0.0011541 0.14071 0.00065809 0.14137 0.12862 0 0.037607 0.0389 0 0.88862 0.24612 0.065685 0.0091964 4.2117 0.057455 6.8923e-005 0.83261 0.0052277 0.0059648 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.13148 0.95751 0.92087 0.0013955 0.99531 0.61249 0.0018802 0.43082 1.9202 1.9197 15.9998 144.9965 0.00015775 -85.6648 0.89096
0.995 0.98802 5.5195e-005 3.8182 0.012037 1.31e-005 0.0011541 0.14079 0.00065809 0.14144 0.12869 0 0.037602 0.0389 0 0.88869 0.24615 0.065696 0.0091978 4.212 0.057464 6.8934e-005 0.83261 0.005228 0.0059651 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13148 0.95759 0.92091 0.0013955 0.99533 0.61263 0.0018802 0.43083 1.9206 1.9201 15.9998 144.9965 0.00015769 -85.6649 0.89196
0.996 0.98802 5.5194e-005 3.8182 0.012037 1.3113e-005 0.0011541 0.14087 0.00065809 0.14152 0.12876 0 0.037597 0.0389 0 0.88876 0.24618 0.065708 0.0091992 4.2123 0.057472 6.8945e-005 0.8326 0.0052283 0.0059654 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13148 0.95767 0.92095 0.0013955 0.99534 0.61276 0.0018801 0.43084 1.9209 1.9204 15.9997 144.9965 0.00015764 -85.6649 0.89296
0.997 0.98802 5.5194e-005 3.8182 0.012037 1.3126e-005 0.0011541 0.14094 0.0006581 0.14159 0.12883 0 0.037592 0.0389 0 0.88883 0.24622 0.065719 0.0092006 4.2125 0.057481 6.8956e-005 0.83259 0.0052286 0.0059657 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13148 0.95775 0.92098 0.0013955 0.99535 0.6129 0.0018801 0.43086 1.9212 1.9207 15.9997 144.9966 0.00015758 -85.6649 0.89396
0.998 0.98802 5.5194e-005 3.8182 0.012037 1.3139e-005 0.0011541 0.14102 0.0006581 0.14167 0.1289 0 0.037587 0.0389 0 0.8889 0.24625 0.065731 0.009202 4.2128 0.057489 6.8967e-005 0.83258 0.0052289 0.005966 0.0013832 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13149 0.95784 0.92102 0.0013955 0.99536 0.61303 0.0018801 0.43087 1.9216 1.9211 15.9997 144.9966 0.00015752 -85.665 0.89496
0.999 0.98802 5.5194e-005 3.8182 0.012037 1.3152e-005 0.0011541 0.14109 0.0006581 0.14175 0.12897 0 0.037582 0.0389 0 0.88898 0.24628 0.065742 0.0092035 4.2131 0.057498 6.8978e-005 0.83257 0.0052292 0.0059663 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13149 0.95792 0.92106 0.0013955 0.99537 0.61317 0.0018801 0.43088 1.9219 1.9214 15.9996 144.9966 0.00015746 -85.665 0.89596
1 0.98802 5.5194e-005 3.8182 0.012037 1.3165e-005 0.0011541 0.14117 0.0006581 0.14182 0.12905 0 0.037577 0.0389 0 0.88905 0.24631 0.065754 0.0092049 4.2134 0.057507 6.8989e-005 0.83256 0.0052295 0.0059667 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13149 0.958 0.9211 0.0013955 0.99539 0.6133 0.0018801 0.43089 1.9222 1.9217 15.9996 144.9966 0.0001574 -85.6651 0.89696
1.001 0.98802 5.5194e-005 3.8182 0.012037 1.3179e-005 0.0011541 0.14124 0.0006581 0.1419 0.12912 0 0.037572 0.0389 0 0.88912 0.24634 0.065765 0.0092063 4.2137 0.057515 6.9e-005 0.83255 0.0052299 0.005967 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13149 0.95808 0.92113 0.0013955 0.9954 0.61344 0.0018801 0.4309 1.9226 1.9221 15.9996 144.9966 0.00015734 -85.6651 0.89796
1.002 0.98802 5.5194e-005 3.8182 0.012037 1.3192e-005 0.0011541 0.14132 0.0006581 0.14197 0.12919 0 0.037567 0.0389 0 0.88919 0.24638 0.065777 0.0092077 4.214 0.057524 6.9011e-005 0.83254 0.0052302 0.0059673 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.1315 0.95816 0.92117 0.0013955 0.99541 0.61357 0.0018801 0.43091 1.9229 1.9224 15.9995 144.9967 0.00015729 -85.6651 0.89896
1.003 0.98802 5.5194e-005 3.8182 0.012037 1.3205e-005 0.0011541 0.1414 0.00065811 0.14205 0.12926 0 0.037562 0.0389 0 0.88927 0.24641 0.065788 0.0092091 4.2142 0.057533 6.9023e-005 0.83254 0.0052305 0.0059676 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.1315 0.95823 0.92121 0.0013955 0.99542 0.61371 0.0018801 0.43093 1.9232 1.9227 15.9995 144.9967 0.00015723 -85.6652 0.89996
1.004 0.98802 5.5194e-005 3.8182 0.012037 1.3218e-005 0.0011541 0.14147 0.00065811 0.14212 0.12933 0 0.037557 0.0389 0 0.88934 0.24644 0.0658 0.0092106 4.2145 0.057541 6.9034e-005 0.83253 0.0052308 0.0059679 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.1315 0.95831 0.92124 0.0013955 0.99543 0.61384 0.0018801 0.43094 1.9235 1.9231 15.9995 144.9967 0.00015717 -85.6652 0.90096
1.005 0.98802 5.5194e-005 3.8182 0.012037 1.3231e-005 0.0011541 0.14155 0.00065811 0.1422 0.1294 0 0.037552 0.0389 0 0.88941 0.24647 0.065812 0.009212 4.2148 0.05755 6.9045e-005 0.83252 0.0052311 0.0059682 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.1315 0.95839 0.92128 0.0013955 0.99544 0.61398 0.0018801 0.43095 1.9239 1.9234 15.9994 144.9967 0.00015711 -85.6653 0.90196
1.006 0.98802 5.5194e-005 3.8182 0.012037 1.3244e-005 0.0011541 0.14162 0.00065811 0.14228 0.12947 0 0.037547 0.0389 0 0.88948 0.2465 0.065823 0.0092134 4.2151 0.057559 6.9056e-005 0.83251 0.0052314 0.0059685 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13151 0.95847 0.92131 0.0013954 0.99545 0.61411 0.0018801 0.43096 1.9242 1.9237 15.9994 144.9967 0.00015706 -85.6653 0.90296
1.007 0.98802 5.5194e-005 3.8182 0.012037 1.3257e-005 0.0011541 0.1417 0.00065811 0.14235 0.12954 0 0.037542 0.0389 0 0.88955 0.24654 0.065835 0.0092149 4.2154 0.057568 6.9067e-005 0.8325 0.0052317 0.0059688 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13151 0.95855 0.92135 0.0013954 0.99547 0.61424 0.0018801 0.43097 1.9245 1.924 15.9994 144.9968 0.000157 -85.6653 0.90396
1.008 0.98802 5.5194e-005 3.8182 0.012037 1.3271e-005 0.0011541 0.14177 0.00065811 0.14243 0.12961 0 0.037537 0.0389 0 0.88963 0.24657 0.065846 0.0092163 4.2157 0.057576 6.9078e-005 0.83249 0.005232 0.0059692 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13151 0.95863 0.92139 0.0013954 0.99548 0.61438 0.0018801 0.43098 1.9249 1.9244 15.9993 144.9968 0.00015694 -85.6654 0.90496
1.009 0.98802 5.5194e-005 3.8182 0.012037 1.3284e-005 0.0011541 0.14185 0.00065812 0.1425 0.12968 0 0.037532 0.0389 0 0.8897 0.2466 0.065858 0.0092177 4.216 0.057585 6.9089e-005 0.83248 0.0052324 0.0059695 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.13151 0.95871 0.92142 0.0013954 0.99549 0.61451 0.0018801 0.431 1.9252 1.9247 15.9993 144.9968 0.00015689 -85.6654 0.90596
1.01 0.98803 5.5194e-005 3.8182 0.012037 1.3297e-005 0.0011541 0.14192 0.00065812 0.14258 0.12975 0 0.037527 0.0389 0 0.88977 0.24663 0.06587 0.0092191 4.2163 0.057594 6.9101e-005 0.83248 0.0052327 0.0059698 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.13152 0.95878 0.92146 0.0013954 0.9955 0.61465 0.0018801 0.43101 1.9255 1.925 15.9993 144.9968 0.00015683 -85.6655 0.90696
1.011 0.98803 5.5194e-005 3.8182 0.012037 1.331e-005 0.0011541 0.142 0.00065812 0.14265 0.12982 0 0.037522 0.0389 0 0.88985 0.24667 0.065881 0.0092206 4.2165 0.057602 6.9112e-005 0.83247 0.005233 0.0059701 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.13152 0.95886 0.92149 0.0013954 0.99551 0.61478 0.0018801 0.43102 1.9258 1.9253 15.9992 144.9968 0.00015677 -85.6655 0.90796
1.012 0.98803 5.5193e-005 3.8182 0.012037 1.3323e-005 0.0011541 0.14207 0.00065812 0.14273 0.12989 0 0.037517 0.0389 0 0.88992 0.2467 0.065893 0.009222 4.2168 0.057611 6.9123e-005 0.83246 0.0052333 0.0059704 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.13152 0.95894 0.92153 0.0013954 0.99552 0.61491 0.00188 0.43103 1.9262 1.9257 15.9992 144.9969 0.00015672 -85.6655 0.90896
1.013 0.98803 5.5193e-005 3.8182 0.012037 1.3336e-005 0.0011541 0.14215 0.00065812 0.1428 0.12996 0 0.037512 0.0389 0 0.88999 0.24673 0.065904 0.0092234 4.2171 0.05762 6.9134e-005 0.83245 0.0052336 0.0059707 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.13153 0.95901 0.92157 0.0013954 0.99553 0.61505 0.00188 0.43104 1.9265 1.926 15.9992 144.9969 0.00015666 -85.6656 0.90996
1.014 0.98803 5.5193e-005 3.8182 0.012037 1.3349e-005 0.0011541 0.14222 0.00065812 0.14288 0.13003 0 0.037507 0.0389 0 0.89006 0.24676 0.065916 0.0092249 4.2174 0.057628 6.9145e-005 0.83244 0.0052339 0.0059711 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.13153 0.95909 0.9216 0.0013954 0.99554 0.61518 0.00188 0.43105 1.9268 1.9263 15.9991 144.9969 0.00015661 -85.6656 0.91096
1.015 0.98803 5.5193e-005 3.8182 0.012037 1.3363e-005 0.0011541 0.1423 0.00065813 0.14295 0.1301 0 0.037502 0.0389 0 0.89014 0.24679 0.065928 0.0092263 4.2177 0.057637 6.9156e-005 0.83243 0.0052342 0.0059714 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.13153 0.95917 0.92164 0.0013954 0.99555 0.61532 0.00188 0.43107 1.9271 1.9267 15.9991 144.9969 0.00015655 -85.6656 0.91196
1.016 0.98803 5.5193e-005 3.8182 0.012036 1.3376e-005 0.0011541 0.14237 0.00065813 0.14303 0.13017 0 0.037497 0.0389 0 0.89021 0.24683 0.065939 0.0092277 4.218 0.057646 6.9168e-005 0.83242 0.0052346 0.0059717 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.13153 0.95924 0.92167 0.0013954 0.99556 0.61545 0.00188 0.43108 1.9275 1.927 15.9991 144.9969 0.0001565 -85.6657 0.91296
1.017 0.98803 5.5193e-005 3.8182 0.012036 1.3389e-005 0.0011541 0.14245 0.00065813 0.1431 0.13024 0 0.037493 0.0389 0 0.89028 0.24686 0.065951 0.0092292 4.2183 0.057655 6.9179e-005 0.83241 0.0052349 0.005972 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.13154 0.95932 0.92171 0.0013954 0.99557 0.61558 0.00188 0.43109 1.9278 1.9273 15.999 144.997 0.00015644 -85.6657 0.91396
1.018 0.98803 5.5193e-005 3.8182 0.012036 1.3402e-005 0.0011541 0.14252 0.00065813 0.14317 0.13031 0 0.037488 0.0389 0 0.89035 0.24689 0.065963 0.0092306 4.2186 0.057663 6.919e-005 0.83241 0.0052352 0.0059723 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.13154 0.9594 0.92174 0.0013954 0.99558 0.61572 0.00188 0.4311 1.9281 1.9276 15.999 144.997 0.00015639 -85.6657 0.91496
1.019 0.98803 5.5193e-005 3.8182 0.012036 1.3415e-005 0.0011541 0.1426 0.00065813 0.14325 0.13038 0 0.037483 0.0389 0 0.89043 0.24692 0.065974 0.009232 4.2189 0.057672 6.9201e-005 0.8324 0.0052355 0.0059726 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13154 0.95947 0.92178 0.0013954 0.99559 0.61585 0.00188 0.43111 1.9284 1.9279 15.999 144.997 0.00015633 -85.6658 0.91596
1.02 0.98803 5.5193e-005 3.8182 0.012036 1.3428e-005 0.0011541 0.14267 0.00065813 0.14332 0.13045 0 0.037478 0.0389 0 0.8905 0.24696 0.065986 0.0092335 4.2192 0.057681 6.9213e-005 0.83239 0.0052358 0.005973 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13154 0.95955 0.92181 0.0013954 0.9956 0.61599 0.00188 0.43113 1.9287 1.9283 15.999 144.997 0.00015628 -85.6658 0.91696
1.021 0.98803 5.5193e-005 3.8182 0.012036 1.3441e-005 0.0011541 0.14274 0.00065813 0.1434 0.13052 0 0.037473 0.0389 0 0.89057 0.24699 0.065997 0.0092349 4.2195 0.05769 6.9224e-005 0.83238 0.0052361 0.0059733 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13155 0.95962 0.92184 0.0013954 0.99561 0.61612 0.00188 0.43114 1.9291 1.9286 15.9989 144.997 0.00015622 -85.6658 0.91796
1.022 0.98803 5.5193e-005 3.8182 0.012036 1.3455e-005 0.0011541 0.14282 0.00065814 0.14347 0.13059 0 0.037468 0.0389 0 0.89065 0.24702 0.066009 0.0092363 4.2197 0.057698 6.9235e-005 0.83237 0.0052365 0.0059736 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13155 0.9597 0.92188 0.0013954 0.99562 0.61625 0.00188 0.43115 1.9294 1.9289 15.9989 144.9971 0.00015617 -85.6659 0.91896
1.023 0.98803 5.5193e-005 3.8182 0.012036 1.3468e-005 0.0011541 0.14289 0.00065814 0.14355 0.13066 0 0.037463 0.0389 0 0.89072 0.24705 0.066021 0.0092378 4.22 0.057707 6.9246e-005 0.83236 0.0052368 0.0059739 0.0013831 0.98699 0.99173 2.9818e-006 1.1927e-005 0.13155 0.95977 0.92191 0.0013954 0.99563 0.61639 0.00188 0.43116 1.9297 1.9292 15.9989 144.9971 0.00015611 -85.6659 0.91996
1.024 0.98803 5.5193e-005 3.8182 0.012036 1.3481e-005 0.0011541 0.14297 0.00065814 0.14362 0.13073 0 0.037458 0.0389 0 0.89079 0.24708 0.066033 0.0092392 4.2203 0.057716 6.9258e-005 0.83235 0.0052371 0.0059742 0.0013831 0.98699 0.99173 2.9818e-006 1.1927e-005 0.13155 0.95984 0.92195 0.0013954 0.99564 0.61652 0.00188 0.43117 1.93 1.9295 15.9988 144.9971 0.00015606 -85.6659 0.92096
1.025 0.98803 5.5193e-005 3.8182 0.012036 1.3494e-005 0.0011541 0.14304 0.00065814 0.1437 0.1308 0 0.037453 0.0389 0 0.89086 0.24712 0.066044 0.0092406 4.2206 0.057725 6.9269e-005 0.83234 0.0052374 0.0059746 0.0013831 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13156 0.95992 0.92198 0.0013954 0.99565 0.61665 0.00188 0.43118 1.9303 1.9299 15.9988 144.9971 0.00015601 -85.666 0.92196
1.026 0.98803 5.5193e-005 3.8182 0.012036 1.3507e-005 0.0011541 0.14312 0.00065814 0.14377 0.13086 0 0.037448 0.0389 0 0.89094 0.24715 0.066056 0.0092421 4.2209 0.057734 6.928e-005 0.83234 0.0052377 0.0059749 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13156 0.95999 0.92202 0.0013954 0.99566 0.61679 0.00188 0.43119 1.9307 1.9302 15.9988 144.9971 0.00015595 -85.666 0.92296
1.027 0.98803 5.5193e-005 3.8182 0.012036 1.352e-005 0.0011541 0.14319 0.00065814 0.14384 0.13093 0 0.037443 0.0389 0 0.89101 0.24718 0.066068 0.0092435 4.2212 0.057742 6.9291e-005 0.83233 0.0052381 0.0059752 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13156 0.96007 0.92205 0.0013954 0.99567 0.61692 0.00188 0.43121 1.931 1.9305 15.9987 144.9972 0.0001559 -85.666 0.92396
1.028 0.98803 5.5192e-005 3.8182 0.012036 1.3533e-005 0.0011541 0.14326 0.00065815 0.14392 0.131 0 0.037439 0.0389 0 0.89108 0.24721 0.066079 0.009245 4.2215 0.057751 6.9303e-005 0.83232 0.0052384 0.0059755 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13156 0.96014 0.92208 0.0013954 0.99568 0.61705 0.00188 0.43122 1.9313 1.9308 15.9987 144.9972 0.00015585 -85.6661 0.92496
1.029 0.98803 5.5192e-005 3.8182 0.012036 1.3547e-005 0.0011541 0.14334 0.00065815 0.14399 0.13107 0 0.037434 0.0389 0 0.89116 0.24725 0.066091 0.0092464 4.2218 0.05776 6.9314e-005 0.83231 0.0052387 0.0059758 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13157 0.96021 0.92212 0.0013954 0.99569 0.61719 0.00188 0.43123 1.9316 1.9311 15.9987 144.9972 0.00015579 -85.6661 0.92596
1.03 0.98803 5.5192e-005 3.8182 0.012036 1.356e-005 0.0011541 0.14341 0.00065815 0.14407 0.13114 0 0.037429 0.0389 0 0.89123 0.24728 0.066103 0.0092478 4.2221 0.057769 6.9325e-005 0.8323 0.005239 0.0059762 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13157 0.96029 0.92215 0.0013953 0.9957 0.61732 0.00188 0.43124 1.9319 1.9315 15.9986 144.9972 0.00015574 -85.6661 0.92696
1.031 0.98803 5.5192e-005 3.8182 0.012036 1.3573e-005 0.0011541 0.14349 0.00065815 0.14414 0.13121 0 0.037424 0.0389 0 0.8913 0.24731 0.066114 0.0092493 4.2224 0.057777 6.9336e-005 0.83229 0.0052393 0.0059765 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13157 0.96036 0.92218 0.0013953 0.99571 0.61745 0.0018799 0.43125 1.9322 1.9318 15.9986 144.9972 0.00015569 -85.6662 0.92796
1.032 0.98803 5.5192e-005 3.8182 0.012036 1.3586e-005 0.0011541 0.14356 0.00065815 0.14421 0.13128 0 0.037419 0.0389 0 0.89138 0.24734 0.066126 0.0092507 4.2227 0.057786 6.9348e-005 0.83228 0.0052397 0.0059768 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13158 0.96043 0.92222 0.0013953 0.99572 0.61759 0.0018799 0.43126 1.9326 1.9321 15.9986 144.9973 0.00015564 -85.6662 0.92896
1.033 0.98803 5.5192e-005 3.8182 0.012036 1.3599e-005 0.0011541 0.14363 0.00065815 0.14429 0.13135 0 0.037414 0.0389 0 0.89145 0.24738 0.066138 0.0092522 4.223 0.057795 6.9359e-005 0.83227 0.00524 0.0059771 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13158 0.9605 0.92225 0.0013953 0.99573 0.61772 0.0018799 0.43128 1.9329 1.9324 15.9985 144.9973 0.00015558 -85.6662 0.92996
1.034 0.98803 5.5192e-005 3.8182 0.012036 1.3612e-005 0.0011541 0.14371 0.00065815 0.14436 0.13142 0 0.037409 0.0389 0 0.89152 0.24741 0.06615 0.0092536 4.2233 0.057804 6.937e-005 0.83227 0.0052403 0.0059775 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13158 0.96057 0.92228 0.0013953 0.99574 0.61785 0.0018799 0.43129 1.9332 1.9327 15.9985 144.9973 0.00015553 -85.6663 0.93096
1.035 0.98803 5.5192e-005 3.8182 0.012036 1.3625e-005 0.0011541 0.14378 0.00065816 0.14443 0.13149 0 0.037405 0.0389 0 0.8916 0.24744 0.066161 0.0092551 4.2236 0.057813 6.9382e-005 0.83226 0.0052406 0.0059778 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13158 0.96065 0.92232 0.0013953 0.99575 0.61798 0.0018799 0.4313 1.9335 1.933 15.9985 144.9973 0.00015548 -85.6663 0.93196
1.036 0.98803 5.5192e-005 3.8182 0.012036 1.3639e-005 0.0011541 0.14385 0.00065816 0.14451 0.13155 0 0.0374 0.0389 0 0.89167 0.24747 0.066173 0.0092565 4.2239 0.057822 6.9393e-005 0.83225 0.005241 0.0059781 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13159 0.96072 0.92235 0.0013953 0.99576 0.61812 0.0018799 0.43131 1.9338 1.9333 15.9984 144.9974 0.00015543 -85.6663 0.93296
1.037 0.98803 5.5192e-005 3.8182 0.012036 1.3652e-005 0.0011541 0.14393 0.00065816 0.14458 0.13162 0 0.037395 0.0389 0 0.89174 0.24751 0.066185 0.0092579 4.2242 0.05783 6.9404e-005 0.83224 0.0052413 0.0059784 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13159 0.96079 0.92238 0.0013953 0.99577 0.61825 0.0018799 0.43132 1.9341 1.9337 15.9984 144.9974 0.00015538 -85.6663 0.93396
1.038 0.98803 5.5192e-005 3.8182 0.012036 1.3665e-005 0.0011541 0.144 0.00065816 0.14466 0.13169 0 0.03739 0.0389 0 0.89182 0.24754 0.066197 0.0092594 4.2245 0.057839 6.9416e-005 0.83223 0.0052416 0.0059788 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13159 0.96086 0.92241 0.0013953 0.99578 0.61838 0.0018799 0.43133 1.9344 1.934 15.9984 144.9974 0.00015532 -85.6664 0.93496
1.039 0.98803 5.5192e-005 3.8182 0.012036 1.3678e-005 0.0011541 0.14408 0.00065816 0.14473 0.13176 0 0.037385 0.0389 0 0.89189 0.24757 0.066208 0.0092608 4.2248 0.057848 6.9427e-005 0.83222 0.0052419 0.0059791 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13159 0.96093 0.92245 0.0013953 0.99579 0.61852 0.0018799 0.43135 1.9348 1.9343 15.9983 144.9974 0.00015527 -85.6664 0.93596
1.04 0.98803 5.5192e-005 3.8182 0.012036 1.3691e-005 0.0011541 0.14415 0.00065816 0.1448 0.13183 0 0.03738 0.0389 0 0.89196 0.24761 0.06622 0.0092623 4.2251 0.057857 6.9438e-005 0.83221 0.0052423 0.0059794 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.1316 0.961 0.92248 0.0013953 0.9958 0.61865 0.0018799 0.43136 1.9351 1.9346 15.9983 144.9974 0.00015522 -85.6664 0.93696
1.041 0.98803 5.5192e-005 3.8182 0.012036 1.3704e-005 0.0011541 0.14422 0.00065817 0.14488 0.1319 0 0.037376 0.0389 0 0.89204 0.24764 0.066232 0.0092637 4.2254 0.057866 6.945e-005 0.8322 0.0052426 0.0059797 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.1316 0.96107 0.92251 0.0013953 0.99581 0.61878 0.0018799 0.43137 1.9354 1.9349 15.9983 144.9975 0.00015517 -85.6665 0.93796
1.042 0.98803 5.5192e-005 3.8182 0.012036 1.3717e-005 0.0011541 0.1443 0.00065817 0.14495 0.13197 0 0.037371 0.0389 0 0.89211 0.24767 0.066244 0.0092652 4.2257 0.057875 6.9461e-005 0.83219 0.0052429 0.0059801 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.1316 0.96114 0.92254 0.0013953 0.99581 0.61891 0.0018799 0.43138 1.9357 1.9352 15.9982 144.9975 0.00015512 -85.6665 0.93896
1.043 0.98803 5.5192e-005 3.8182 0.012036 1.3731e-005 0.0011541 0.14437 0.00065817 0.14502 0.13203 0 0.037366 0.0389 0 0.89219 0.2477 0.066256 0.0092666 4.226 0.057883 6.9472e-005 0.83219 0.0052432 0.0059804 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13161 0.96121 0.92258 0.0013953 0.99582 0.61905 0.0018799 0.43139 1.936 1.9355 15.9982 144.9975 0.00015507 -85.6665 0.93996
1.044 0.98803 5.5191e-005 3.8182 0.012036 1.3744e-005 0.0011541 0.14444 0.00065817 0.14509 0.1321 0 0.037361 0.0389 0 0.89226 0.24774 0.066267 0.0092681 4.2263 0.057892 6.9484e-005 0.83218 0.0052436 0.0059807 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13161 0.96128 0.92261 0.0013953 0.99583 0.61918 0.0018799 0.4314 1.9363 1.9358 15.9982 144.9975 0.00015502 -85.6665 0.94096
1.045 0.98803 5.5191e-005 3.8182 0.012036 1.3757e-005 0.0011541 0.14451 0.00065817 0.14517 0.13217 0 0.037356 0.0389 0 0.89233 0.24777 0.066279 0.0092695 4.2266 0.057901 6.9495e-005 0.83217 0.0052439 0.0059811 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13161 0.96135 0.92264 0.0013953 0.99584 0.61931 0.0018799 0.43141 1.9366 1.9362 15.9981 144.9975 0.00015497 -85.6666 0.94196
1.046 0.98803 5.5191e-005 3.8182 0.012036 1.377e-005 0.0011541 0.14459 0.00065817 0.14524 0.13224 0 0.037352 0.0389 0 0.89241 0.2478 0.066291 0.009271 4.2269 0.05791 6.9506e-005 0.83216 0.0052442 0.0059814 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13161 0.96142 0.92267 0.0013953 0.99585 0.61944 0.0018799 0.43143 1.9369 1.9365 15.9981 144.9976 0.00015492 -85.6666 0.94296
1.047 0.98803 5.5191e-005 3.8182 0.012036 1.3783e-005 0.0011541 0.14466 0.00065817 0.14531 0.13231 0 0.037347 0.0389 0 0.89248 0.24783 0.066303 0.0092724 4.2272 0.057919 6.9518e-005 0.83215 0.0052445 0.0059817 0.0013829 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13162 0.96149 0.9227 0.0013953 0.99586 0.61958 0.0018799 0.43144 1.9372 1.9368 15.9981 144.9976 0.00015487 -85.6666 0.94396
1.048 0.98803 5.5191e-005 3.8182 0.012036 1.3796e-005 0.0011541 0.14473 0.00065818 0.14539 0.13238 0 0.037342 0.0389 0 0.89255 0.24787 0.066315 0.0092739 4.2275 0.057928 6.9529e-005 0.83214 0.0052449 0.005982 0.0013828 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13162 0.96156 0.92274 0.0013953 0.99587 0.61971 0.0018799 0.43145 1.9375 1.9371 15.998 144.9976 0.00015482 -85.6667 0.94496
1.049 0.98803 5.5191e-005 3.8182 0.012036 1.3809e-005 0.0011541 0.14481 0.00065818 0.14546 0.13244 0 0.037337 0.0389 0 0.89263 0.2479 0.066326 0.0092753 4.2278 0.057937 6.9541e-005 0.83213 0.0052452 0.0059824 0.0013828 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13162 0.96163 0.92277 0.0013953 0.99588 0.61984 0.0018799 0.43146 1.9378 1.9374 15.998 144.9976 0.00015477 -85.6667 0.94596
1.05 0.98803 5.5191e-005 3.8182 0.012036 1.3823e-005 0.0011541 0.14488 0.00065818 0.14553 0.13251 0 0.037333 0.0389 0 0.8927 0.24793 0.066338 0.0092768 4.2281 0.057946 6.9552e-005 0.83212 0.0052455 0.0059827 0.0013828 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13162 0.9617 0.9228 0.0013953 0.99588 0.61997 0.0018799 0.43147 1.9381 1.9377 15.998 144.9976 0.00015472 -85.6667 0.94696
1.051 0.98803 5.5191e-005 3.8182 0.012036 1.3836e-005 0.0011541 0.14495 0.00065818 0.14561 0.13258 0 0.037328 0.0389 0 0.89278 0.24796 0.06635 0.0092783 4.2285 0.057954 6.9563e-005 0.83212 0.0052459 0.005983 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13163 0.96177 0.92283 0.0013953 0.99589 0.62011 0.0018799 0.43148 1.9385 1.938 15.9979 144.9977 0.00015467 -85.6667 0.94796
1.052 0.98803 5.5191e-005 3.8182 0.012036 1.3849e-005 0.0011541 0.14502 0.00065818 0.14568 0.13265 0 0.037323 0.0389 0 0.89285 0.248 0.066362 0.0092797 4.2288 0.057963 6.9575e-005 0.83211 0.0052462 0.0059834 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13163 0.96183 0.92286 0.0013953 0.9959 0.62024 0.0018798 0.4315 1.9388 1.9383 15.9979 144.9977 0.00015462 -85.6668 0.94896
1.053 0.98803 5.5191e-005 3.8182 0.012036 1.3862e-005 0.0011541 0.1451 0.00065818 0.14575 0.13272 0 0.037318 0.0389 0 0.89292 0.24803 0.066374 0.0092812 4.2291 0.057972 6.9586e-005 0.8321 0.0052465 0.0059837 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13163 0.9619 0.92289 0.0013953 0.99591 0.62037 0.0018798 0.43151 1.9391 1.9386 15.9979 144.9977 0.00015457 -85.6668 0.94996
1.054 0.98803 5.5191e-005 3.8182 0.012036 1.3875e-005 0.0011541 0.14517 0.00065819 0.14582 0.13278 0 0.037314 0.0389 0 0.893 0.24806 0.066386 0.0092826 4.2294 0.057981 6.9598e-005 0.83209 0.0052468 0.005984 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13164 0.96197 0.92292 0.0013953 0.99592 0.6205 0.0018798 0.43152 1.9394 1.9389 15.9978 144.9977 0.00015452 -85.6668 0.95096
1.055 0.98803 5.5191e-005 3.8182 0.012036 1.3888e-005 0.0011541 0.14524 0.00065819 0.1459 0.13285 0 0.037309 0.0389 0 0.89307 0.2481 0.066397 0.0092841 4.2297 0.05799 6.9609e-005 0.83208 0.0052472 0.0059844 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13164 0.96204 0.92295 0.0013953 0.99592 0.62063 0.0018798 0.43153 1.9397 1.9392 15.9978 144.9977 0.00015448 -85.6668 0.95196
1.056 0.98803 5.5191e-005 3.8182 0.012036 1.3901e-005 0.0011541 0.14531 0.00065819 0.14597 0.13292 0 0.037304 0.0389 0 0.89315 0.24813 0.066409 0.0092855 4.23 0.057999 6.9621e-005 0.83207 0.0052475 0.0059847 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13164 0.9621 0.92298 0.0013953 0.99593 0.62077 0.0018798 0.43154 1.94 1.9395 15.9978 144.9978 0.00015443 -85.6669 0.95296
1.057 0.98803 5.5191e-005 3.8182 0.012036 1.3915e-005 0.0011541 0.14539 0.00065819 0.14604 0.13299 0 0.037299 0.0389 0 0.89322 0.24816 0.066421 0.009287 4.2303 0.058008 6.9632e-005 0.83206 0.0052478 0.005985 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13164 0.96217 0.92302 0.0013953 0.99594 0.6209 0.0018798 0.43155 1.9403 1.9398 15.9977 144.9978 0.00015438 -85.6669 0.95396
1.058 0.98803 5.5191e-005 3.8182 0.012036 1.3928e-005 0.0011541 0.14546 0.00065819 0.14611 0.13305 0 0.037295 0.0389 0 0.89329 0.2482 0.066433 0.0092885 4.2306 0.058017 6.9643e-005 0.83205 0.0052482 0.0059854 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13165 0.96224 0.92305 0.0013953 0.99595 0.62103 0.0018798 0.43156 1.9406 1.9401 15.9977 144.9978 0.00015433 -85.6669 0.95496
1.059 0.98803 5.5191e-005 3.8182 0.012036 1.3941e-005 0.0011541 0.14553 0.00065819 0.14618 0.13312 0 0.03729 0.0389 0 0.89337 0.24823 0.066445 0.0092899 4.2309 0.058026 6.9655e-005 0.83204 0.0052485 0.0059857 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13165 0.9623 0.92308 0.0013952 0.99596 0.62116 0.0018798 0.43158 1.9409 1.9404 15.9977 144.9978 0.00015428 -85.6669 0.95596
1.06 0.98803 5.519e-005 3.8182 0.012036 1.3954e-005 0.0011541 0.1456 0.00065819 0.14626 0.13319 0 0.037285 0.0389 0 0.89344 0.24826 0.066457 0.0092914 4.2312 0.058035 6.9666e-005 0.83204 0.0052488 0.005986 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13165 0.96237 0.92311 0.0013952 0.99596 0.62129 0.0018798 0.43159 1.9412 1.9407 15.9976 144.9978 0.00015424 -85.667 0.95696
1.061 0.98803 5.519e-005 3.8182 0.012036 1.3967e-005 0.0011541 0.14568 0.0006582 0.14633 0.13326 0 0.03728 0.0389 0 0.89352 0.24829 0.066469 0.0092928 4.2315 0.058043 6.9678e-005 0.83203 0.0052492 0.0059864 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13165 0.96244 0.92314 0.0013952 0.99597 0.62143 0.0018798 0.4316 1.9415 1.941 15.9976 144.9979 0.00015419 -85.667 0.95796
1.062 0.98803 5.519e-005 3.8182 0.012036 1.398e-005 0.0011541 0.14575 0.0006582 0.1464 0.13332 0 0.037276 0.0389 0 0.89359 0.24833 0.066481 0.0092943 4.2319 0.058052 6.9689e-005 0.83202 0.0052495 0.0059867 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13166 0.9625 0.92317 0.0013952 0.99598 0.62156 0.0018798 0.43161 1.9418 1.9413 15.9976 144.9979 0.00015414 -85.667 0.95896
1.063 0.98803 5.519e-005 3.8182 0.012036 1.3993e-005 0.0011541 0.14582 0.0006582 0.14647 0.13339 0 0.037271 0.0389 0 0.89367 0.24836 0.066492 0.0092958 4.2322 0.058061 6.9701e-005 0.83201 0.0052498 0.005987 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13166 0.96257 0.9232 0.0013952 0.99599 0.62169 0.0018798 0.43162 1.9421 1.9416 15.9975 144.9979 0.00015409 -85.667 0.95996
1.064 0.98803 5.519e-005 3.8182 0.012036 1.4007e-005 0.0011541 0.14589 0.0006582 0.14654 0.13346 0 0.037266 0.0389 0 0.89374 0.24839 0.066504 0.0092972 4.2325 0.05807 6.9712e-005 0.832 0.0052502 0.0059874 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13166 0.96263 0.92323 0.0013952 0.996 0.62182 0.0018798 0.43163 1.9424 1.9419 15.9975 144.9979 0.00015405 -85.6671 0.96096
1.065 0.98803 5.519e-005 3.8182 0.012036 1.402e-005 0.0011541 0.14596 0.0006582 0.14662 0.13352 0 0.037262 0.0389 0 0.89381 0.24843 0.066516 0.0092987 4.2328 0.058079 6.9724e-005 0.83199 0.0052505 0.0059877 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13167 0.9627 0.92326 0.0013952 0.996 0.62195 0.0018798 0.43164 1.9427 1.9422 15.9975 144.9979 0.000154 -85.6671 0.96196
1.066 0.98803 5.519e-005 3.8182 0.012036 1.4033e-005 0.0011541 0.14604 0.0006582 0.14669 0.13359 0 0.037257 0.0389 0 0.89389 0.24846 0.066528 0.0093001 4.2331 0.058088 6.9735e-005 0.83198 0.0052508 0.0059881 0.0013828 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13167 0.96276 0.92329 0.0013952 0.99601 0.62208 0.0018798 0.43166 1.943 1.9425 15.9974 144.998 0.00015395 -85.6671 0.96296
1.067 0.98803 5.519e-005 3.8182 0.012036 1.4046e-005 0.0011541 0.14611 0.0006582 0.14676 0.13366 0 0.037252 0.0389 0 0.89396 0.24849 0.06654 0.0093016 4.2334 0.058097 6.9747e-005 0.83197 0.0052512 0.0059884 0.0013828 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13167 0.96283 0.92332 0.0013952 0.99602 0.62222 0.0018798 0.43167 1.9433 1.9428 15.9974 144.998 0.00015391 -85.6671 0.96396
1.068 0.98803 5.519e-005 3.8182 0.012036 1.4059e-005 0.0011541 0.14618 0.00065821 0.14683 0.13373 0 0.037248 0.0389 0 0.89404 0.24852 0.066552 0.0093031 4.2337 0.058106 6.9758e-005 0.83196 0.0052515 0.0059887 0.0013827 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13167 0.96289 0.92335 0.0013952 0.99603 0.62235 0.0018798 0.43168 1.9436 1.9431 15.9974 144.998 0.00015386 -85.6672 0.96496
1.069 0.98803 5.519e-005 3.8182 0.012036 1.4072e-005 0.0011541 0.14625 0.00065821 0.1469 0.13379 0 0.037243 0.0389 0 0.89411 0.24856 0.066564 0.0093045 4.234 0.058115 6.977e-005 0.83195 0.0052519 0.0059891 0.0013827 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13168 0.96296 0.92338 0.0013952 0.99603 0.62248 0.0018798 0.43169 1.9439 1.9434 15.9973 144.998 0.00015381 -85.6672 0.96596
1.07 0.98803 5.519e-005 3.8182 0.012036 1.4085e-005 0.0011541 0.14632 0.00065821 0.14698 0.13386 0 0.037238 0.0389 0 0.89419 0.24859 0.066576 0.009306 4.2344 0.058124 6.9781e-005 0.83195 0.0052522 0.0059894 0.0013827 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13168 0.96302 0.9234 0.0013952 0.99604 0.62261 0.0018798 0.4317 1.9442 1.9437 15.9973 144.9981 0.00015377 -85.6672 0.96696
1.071 0.98803 5.519e-005 3.8182 0.012036 1.4099e-005 0.0011541 0.14639 0.00065821 0.14705 0.13393 0 0.037234 0.0389 0 0.89426 0.24862 0.066588 0.0093075 4.2347 0.058133 6.9793e-005 0.83194 0.0052525 0.0059898 0.0013827 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13168 0.96309 0.92343 0.0013952 0.99605 0.62274 0.0018798 0.43171 1.9445 1.944 15.9973 144.9981 0.00015372 -85.6672 0.96796
1.072 0.98803 5.519e-005 3.8182 0.012036 1.4112e-005 0.0011541 0.14646 0.00065821 0.14712 0.13399 0 0.037229 0.0389 0 0.89434 0.24866 0.0666 0.0093089 4.235 0.058142 6.9804e-005 0.83193 0.0052529 0.0059901 0.0013827 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13169 0.96315 0.92346 0.0013952 0.99606 0.62287 0.0018798 0.43172 1.9448 1.9443 15.9972 144.9981 0.00015367 -85.6672 0.96896
1.073 0.98803 5.519e-005 3.8182 0.012036 1.4125e-005 0.0011541 0.14654 0.00065821 0.14719 0.13406 0 0.037224 0.0389 0 0.89441 0.24869 0.066612 0.0093104 4.2353 0.058151 6.9816e-005 0.83192 0.0052532 0.0059904 0.0013827 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13169 0.96321 0.92349 0.0013952 0.99606 0.623 0.0018798 0.43174 1.9451 1.9446 15.9972 144.9981 0.00015363 -85.6673 0.96996
1.074 0.98803 5.519e-005 3.8182 0.012036 1.4138e-005 0.0011541 0.14661 0.00065821 0.14726 0.13413 0 0.03722 0.0389 0 0.89449 0.24872 0.066624 0.0093119 4.2356 0.05816 6.9827e-005 0.83191 0.0052535 0.0059908 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.13169 0.96328 0.92352 0.0013952 0.99607 0.62314 0.0018798 0.43175 1.9454 1.9449 15.9972 144.9981 0.00015358 -85.6673 0.97096
1.075 0.98803 5.519e-005 3.8182 0.012036 1.4151e-005 0.0011541 0.14668 0.00065822 0.14733 0.13419 0 0.037215 0.0389 0 0.89456 0.24876 0.066636 0.0093133 4.2359 0.058169 6.9839e-005 0.8319 0.0052539 0.0059911 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.13169 0.96334 0.92355 0.0013952 0.99608 0.62327 0.0018798 0.43176 1.9457 1.9452 15.9971 144.9982 0.00015354 -85.6673 0.97196
1.076 0.98803 5.5189e-005 3.8182 0.012036 1.4164e-005 0.0011541 0.14675 0.00065822 0.1474 0.13426 0 0.03721 0.0389 0 0.89464 0.24879 0.066648 0.0093148 4.2363 0.058178 6.9851e-005 0.83189 0.0052542 0.0059915 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.1317 0.9634 0.92358 0.0013952 0.99608 0.6234 0.0018798 0.43177 1.946 1.9455 15.9971 144.9982 0.00015349 -85.6673 0.97296
1.077 0.98803 5.5189e-005 3.8182 0.012036 1.4177e-005 0.0011541 0.14682 0.00065822 0.14748 0.13433 0 0.037206 0.0389 0 0.89471 0.24882 0.06666 0.0093163 4.2366 0.058187 6.9862e-005 0.83188 0.0052546 0.0059918 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.1317 0.96347 0.92361 0.0013952 0.99609 0.62353 0.0018798 0.43178 1.9463 1.9458 15.9971 144.9982 0.00015345 -85.6674 0.97396
1.078 0.98803 5.5189e-005 3.8182 0.012036 1.4191e-005 0.0011541 0.14689 0.00065822 0.14755 0.13439 0 0.037201 0.0389 0 0.89479 0.24886 0.066672 0.0093178 4.2369 0.058196 6.9874e-005 0.83187 0.0052549 0.0059921 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.1317 0.96353 0.92364 0.0013952 0.9961 0.62366 0.0018798 0.43179 1.9465 1.9461 15.997 144.9982 0.0001534 -85.6674 0.97496
1.079 0.98803 5.5189e-005 3.8182 0.012036 1.4204e-005 0.0011541 0.14696 0.00065822 0.14762 0.13446 0 0.037196 0.0389 0 0.89486 0.24889 0.066684 0.0093192 4.2372 0.058205 6.9885e-005 0.83186 0.0052552 0.0059925 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.1317 0.96359 0.92367 0.0013952 0.99611 0.62379 0.0018797 0.4318 1.9468 1.9464 15.997 144.9982 0.00015336 -85.6674 0.97596
1.08 0.98803 5.5189e-005 3.8182 0.012036 1.4217e-005 0.0011541 0.14703 0.00065822 0.14769 0.13453 0 0.037192 0.0389 0 0.89494 0.24892 0.066696 0.0093207 4.2375 0.058214 6.9897e-005 0.83186 0.0052556 0.0059928 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.13171 0.96365 0.92369 0.0013952 0.99611 0.62392 0.0018797 0.43181 1.9471 1.9467 15.997 144.9983 0.00015331 -85.6674 0.97696
1.081 0.98803 5.5189e-005 3.8182 0.012036 1.423e-005 0.0011541 0.14711 0.00065822 0.14776 0.13459 0 0.037187 0.0389 0 0.89501 0.24896 0.066708 0.0093222 4.2378 0.058223 6.9908e-005 0.83185 0.0052559 0.0059932 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.13171 0.96372 0.92372 0.0013952 0.99612 0.62405 0.0018797 0.43183 1.9474 1.947 15.9969 144.9983 0.00015327 -85.6674 0.97796
1.082 0.98803 5.5189e-005 3.8182 0.012036 1.4243e-005 0.0011541 0.14718 0.00065823 0.14783 0.13466 0 0.037183 0.0389 0 0.89509 0.24899 0.06672 0.0093236 4.2382 0.058232 6.992e-005 0.83184 0.0052563 0.0059935 0.0013827 0.98699 0.99173 2.981e-006 1.1924e-005 0.13171 0.96378 0.92375 0.0013952 0.99613 0.62418 0.0018797 0.43184 1.9477 1.9473 15.9969 144.9983 0.00015322 -85.6675 0.97896
1.083 0.98803 5.5189e-005 3.8182 0.012036 1.4256e-005 0.0011541 0.14725 0.00065823 0.1479 0.13473 0 0.037178 0.0389 0 0.89516 0.24902 0.066732 0.0093251 4.2385 0.058241 6.9932e-005 0.83183 0.0052566 0.0059939 0.0013827 0.98699 0.99173 2.9809e-006 1.1924e-005 0.13172 0.96384 0.92378 0.0013952 0.99613 0.62431 0.0018797 0.43185 1.948 1.9476 15.9969 144.9983 0.00015318 -85.6675 0.97996
1.084 0.98803 5.5189e-005 3.8182 0.012036 1.4269e-005 0.0011541 0.14732 0.00065823 0.14797 0.13479 0 0.037173 0.0389 0 0.89524 0.24906 0.066744 0.0093266 4.2388 0.05825 6.9943e-005 0.83182 0.0052569 0.0059942 0.0013827 0.98699 0.99173 2.9809e-006 1.1924e-005 0.13172 0.9639 0.92381 0.0013952 0.99614 0.62444 0.0018797 0.43186 1.9483 1.9479 15.9968 144.9983 0.00015313 -85.6675 0.98096
1.085 0.98803 5.5189e-005 3.8182 0.012036 1.4283e-005 0.0011541 0.14739 0.00065823 0.14804 0.13486 0 0.037169 0.0389 0 0.89531 0.24909 0.066756 0.0093281 4.2391 0.058259 6.9955e-005 0.83181 0.0052573 0.0059945 0.0013827 0.98699 0.99173 2.9809e-006 1.1924e-005 0.13172 0.96396 0.92383 0.0013952 0.99615 0.62458 0.0018797 0.43187 1.9486 1.9482 15.9968 144.9984 0.00015309 -85.6675 0.98196
1.086 0.98803 5.5189e-005 3.8182 0.012036 1.4296e-005 0.0011541 0.14746 0.00065823 0.14811 0.13492 0 0.037164 0.0389 0 0.89539 0.24912 0.066768 0.0093295 4.2394 0.058268 6.9966e-005 0.8318 0.0052576 0.0059949 0.0013827 0.98699 0.99173 2.9809e-006 1.1924e-005 0.13172 0.96402 0.92386 0.0013952 0.99615 0.62471 0.0018797 0.43188 1.9489 1.9485 15.9968 144.9984 0.00015305 -85.6675 0.98296
1.087 0.98803 5.5189e-005 3.8182 0.012036 1.4309e-005 0.0011541 0.14753 0.00065823 0.14818 0.13499 0 0.03716 0.0389 0 0.89546 0.24916 0.06678 0.009331 4.2398 0.058277 6.9978e-005 0.83179 0.005258 0.0059952 0.0013827 0.98699 0.99173 2.9809e-006 1.1924e-005 0.13173 0.96409 0.92389 0.0013952 0.99616 0.62484 0.0018797 0.43189 1.9492 1.9487 15.9967 144.9984 0.000153 -85.6676 0.98396
1.088 0.98803 5.5189e-005 3.8182 0.012036 1.4322e-005 0.0011541 0.1476 0.00065823 0.14825 0.13506 0 0.037155 0.0389 0 0.89554 0.24919 0.066792 0.0093325 4.2401 0.058286 6.999e-005 0.83178 0.0052583 0.0059956 0.0013826 0.98699 0.99173 2.9809e-006 1.1923e-005 0.13173 0.96415 0.92392 0.0013952 0.99617 0.62497 0.0018797 0.43191 1.9495 1.949 15.9967 144.9984 0.00015296 -85.6676 0.98496
1.089 0.98803 5.5189e-005 3.8182 0.012036 1.4335e-005 0.0011542 0.14767 0.00065824 0.14832 0.13512 0 0.03715 0.0389 0 0.89561 0.24922 0.066804 0.009334 4.2404 0.058295 7.0001e-005 0.83177 0.0052587 0.0059959 0.0013826 0.98699 0.99173 2.9809e-006 1.1923e-005 0.13173 0.96421 0.92395 0.0013952 0.99617 0.6251 0.0018797 0.43192 1.9498 1.9493 15.9967 144.9984 0.00015291 -85.6676 0.98596
1.09 0.98803 5.5189e-005 3.8182 0.012036 1.4348e-005 0.0011542 0.14774 0.00065824 0.1484 0.13519 0 0.037146 0.0389 0 0.89569 0.24926 0.066816 0.0093355 4.2407 0.058304 7.0013e-005 0.83177 0.005259 0.0059963 0.0013826 0.98699 0.99173 2.9809e-006 1.1923e-005 0.13174 0.96427 0.92397 0.0013952 0.99618 0.62523 0.0018797 0.43193 1.95 1.9496 15.9966 144.9985 0.00015287 -85.6676 0.98696
1.091 0.98803 5.5189e-005 3.8182 0.012035 1.4361e-005 0.0011542 0.14781 0.00065824 0.14847 0.13525 0 0.037141 0.0389 0 0.89576 0.24929 0.066828 0.0093369 4.2411 0.058313 7.0024e-005 0.83176 0.0052594 0.0059966 0.0013826 0.98699 0.99173 2.9809e-006 1.1923e-005 0.13174 0.96433 0.924 0.0013952 0.99619 0.62536 0.0018797 0.43194 1.9503 1.9499 15.9966 144.9985 0.00015283 -85.6676 0.98796
1.092 0.98803 5.5188e-005 3.8182 0.012035 1.4374e-005 0.0011542 0.14788 0.00065824 0.14854 0.13532 0 0.037137 0.0389 0 0.89584 0.24932 0.06684 0.0093384 4.2414 0.058322 7.0036e-005 0.83175 0.0052597 0.005997 0.0013827 0.98699 0.99173 2.9809e-006 1.1923e-005 0.13174 0.96439 0.92403 0.0013952 0.99619 0.62549 0.0018797 0.43195 1.9506 1.9502 15.9966 144.9985 0.00015279 -85.6676 0.98896
1.093 0.98803 5.5188e-005 3.8182 0.012035 1.4388e-005 0.0011542 0.14795 0.00065824 0.14861 0.13538 0 0.037132 0.0389 0 0.89591 0.24936 0.066852 0.0093399 4.2417 0.058331 7.0048e-005 0.83174 0.00526 0.0059973 0.0013827 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13174 0.96445 0.92406 0.0013952 0.9962 0.62562 0.0018797 0.43196 1.9509 1.9505 15.9965 144.9985 0.00015274 -85.6677 0.98996
1.094 0.98803 5.5188e-005 3.8182 0.012035 1.4401e-005 0.0011542 0.14802 0.00065824 0.14868 0.13545 0 0.037128 0.0389 0 0.89599 0.24939 0.066864 0.0093414 4.242 0.05834 7.0059e-005 0.83173 0.0052604 0.0059977 0.0013827 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13175 0.96451 0.92408 0.0013952 0.99621 0.62575 0.0018797 0.43197 1.9512 1.9508 15.9965 144.9985 0.0001527 -85.6677 0.99096
1.095 0.98803 5.5188e-005 3.8182 0.012035 1.4414e-005 0.0011542 0.14809 0.00065824 0.14875 0.13552 0 0.037123 0.0389 0 0.89606 0.24942 0.066876 0.0093429 4.2424 0.05835 7.0071e-005 0.83172 0.0052607 0.005998 0.0013827 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13175 0.96457 0.92411 0.0013952 0.99621 0.62588 0.0018797 0.43198 1.9515 1.9511 15.9965 144.9986 0.00015266 -85.6677 0.99196
1.096 0.98803 5.5188e-005 3.8182 0.012035 1.4427e-005 0.0011542 0.14816 0.00065825 0.14882 0.13558 0 0.037119 0.0389 0 0.89614 0.24946 0.066888 0.0093443 4.2427 0.058359 7.0083e-005 0.83171 0.0052611 0.0059984 0.0013827 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13175 0.96463 0.92414 0.0013952 0.99622 0.62601 0.0018797 0.432 1.9518 1.9513 15.9964 144.9986 0.00015261 -85.6677 0.99296
1.097 0.98803 5.5188e-005 3.8182 0.012035 1.444e-005 0.0011542 0.14823 0.00065825 0.14889 0.13565 0 0.037114 0.0389 0 0.89621 0.24949 0.0669 0.0093458 4.243 0.058368 7.0094e-005 0.8317 0.0052614 0.0059987 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13176 0.96469 0.92416 0.0013952 0.99622 0.62614 0.0018797 0.43201 1.9521 1.9516 15.9964 144.9986 0.00015257 -85.6677 0.99396
1.098 0.98803 5.5188e-005 3.8182 0.012035 1.4453e-005 0.0011542 0.1483 0.00065825 0.14896 0.13571 0 0.037109 0.0389 0 0.89629 0.24952 0.066912 0.0093473 4.2433 0.058377 7.0106e-005 0.83169 0.0052618 0.0059991 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13176 0.96474 0.92419 0.0013951 0.99623 0.62627 0.0018797 0.43202 1.9523 1.9519 15.9964 144.9986 0.00015253 -85.6678 0.99496
1.099 0.98803 5.5188e-005 3.8182 0.012035 1.4466e-005 0.0011542 0.14837 0.00065825 0.14903 0.13578 0 0.037105 0.0389 0 0.89636 0.24956 0.066924 0.0093488 4.2437 0.058386 7.0118e-005 0.83168 0.0052621 0.0059994 0.0013826 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13176 0.9648 0.92422 0.0013951 0.99624 0.6264 0.0018797 0.43203 1.9526 1.9522 15.9963 144.9986 0.00015249 -85.6678 0.99596
1.1 0.98803 5.5188e-005 3.8182 0.012035 1.448e-005 0.0011542 0.14844 0.00065825 0.1491 0.13584 0 0.0371 0.0389 0 0.89644 0.24959 0.066937 0.0093503 4.244 0.058395 7.0129e-005 0.83168 0.0052625 0.0059998 0.0013827 0.98699 0.99173 2.9808e-006 1.1923e-005 0.13176 0.96486 0.92424 0.0013951 0.99624 0.62653 0.0018797 0.43204 1.9529 1.9525 15.9963 144.9987 0.00015245 -85.6646 0.99696
1.101 0.98803 5.5188e-005 3.8182 0.012035 1.4493e-005 0.0011542 0.14851 0.00065825 0.14917 0.13591 0 0.037096 0.0389 0 0.89652 0.24962 0.066949 0.0093518 4.2443 0.058404 7.0141e-005 0.83167 0.0052628 0.0060001 0.0064718 0.98324 0.991 1.4514e-005 5.332e-005 0.13177 0.96487 0.92427 0.0027729 0.99623 0.62664 0.002395 0.432 1.9532 1.9528 15.9962 144.9987 0.00015241 -76.162 0.99796
1.102 0.98803 5.5188e-005 3.8182 0.012035 1.4506e-005 0.0011542 0.14858 0.00065825 0.14924 0.13597 0 0.037091 0.0389 0 0.89659 0.24966 0.066961 0.0093532 4.2447 0.058413 7.0153e-005 0.83166 0.0052632 0.0060005 0.026215 0.97172 0.98767 6.596e-005 0.00022944 0.13177 0.96466 0.9243 0.0053002 0.99618 0.62674 0.0033358 0.43188 1.9535 1.9531 15.9962 144.9986 0.0001524 -67.1482 0.99896
1.103 0.98803 5.5188e-005 3.8182 0.012035 1.4519e-005 0.0011542 0.14865 0.00065825 0.14931 0.13604 0 0.037087 0.0389 0 0.89667 0.24969 0.066973 0.0093547 4.245 0.058422 7.0164e-005 0.83165 0.0052635 0.0060008 0.094853 0.94723 0.97734 0.00028432 0.00091291 0.13177 0.9639 0.92432 0.0092468 0.99592 0.62682 0.0044246 0.43171 1.9538 1.9533 15.9961 144.9986 0.00015241 -58.017 0.99996
1.104 0.98803 5.5188e-005 3.8182 0.012035 1.4532e-005 0.0011542 0.14872 0.00065826 0.14938 0.1361 0 0.037082 0.0389 0 0.89674 0.24972 0.066985 0.0093562 4.2453 0.058431 7.0176e-005 0.83164 0.0052639 0.0060012 0.48775 0.85644 0.93876 0.0021772 0.0054714 0.13178 0.96187 0.92434 0.01575 0.99181 0.62683 0.0056234 0.43152 1.954 1.9536 15.9968 144.9986 0.00015245 -37.2335 0.1564
1.105 0.98803 5.5188e-005 3.8182 0.012035 1.4545e-005 0.0011542 0.14879 0.00065826 0.14945 0.13617 0 0.037078 0.0389 0 0.89682 0.24976 0.066997 0.0093577 4.2456 0.05844 7.0188e-005 0.83163 0.0052642 0.0060015 0.99959 0.0021826 0.71218 0.93591 0.9957 0.13178 0.92831 0.9214 0.33179 0.96439 0.61307 0.043959 0.43132 1.9134 0.96878 16.0007 144.9983 0.0002317 23.8159 0.0019501
1.106 0.98803 5.5188e-005 3.8182 0.012035 1.4558e-005 0.0011542 0.14886 0.00065826 0.14952 0.13623 0 0.037073 0.0389 0 0.89689 0.24979 0.067009 0.0093592 4.246 0.05845 7.02e-005 0.83162 0.0052646 0.0060019 0.99924 1.4699e-006 0.52841 0.99594 0.99917 0.13178 0.88826 0.90352 0.59542 0.93723 0.596 0.093559 0.43111 1.7309 0.58831 16.0004 144.997 0.00034055 17.4443 0.0029501
1.107 0.98803 5.5188e-005 3.8182 0.012035 1.4572e-005 0.0011542 0.14893 0.00065826 0.14958 0.1363 0 0.037069 0.0389 0 0.89697 0.24983 0.067021 0.0093607 4.2463 0.058459 7.0211e-005 0.83161 0.0052649 0.0060022 0.99852 1.247e-008 0.39262 0.99224 0.99769 0.13179 0.85132 0.8804 0.70434 0.91083 0.57989 0.12897 0.43091 1.5556 0.56005 16 144.9954 0.00040818 11.2953 0.0039501
1.108 0.98803 5.5187e-005 3.8182 0.012035 1.4585e-005 0.0011542 0.149 0.00065826 0.14965 0.13636 0 0.037064 0.0389 0 0.89705 0.24986 0.067034 0.0093622 4.2466 0.058468 7.0223e-005 0.8316 0.0052653 0.0060026 0.99768 -2.1896e-009 0.29228 0.98466 0.99528 0.13179 0.81821 0.85497 0.74913 0.88519 0.56506 0.15556 0.4307 1.4089 0.5958 15.9997 144.9937 0.0004581 7.2143 0.0049501
1.109 0.98803 5.5187e-005 3.8182 0.012035 1.4598e-005 0.0011542 0.14907 0.00065826 0.14972 0.13643 0 0.03706 0.0389 0 0.89712 0.24989 0.067046 0.0093637 4.247 0.058477 7.0235e-005 0.83159 0.0052656 0.0060029 0.99685 -4.5295e-010 0.21799 0.97495 0.99226 0.13179 0.78853 0.82864 0.76537 0.86027 0.55156 0.17707 0.4305 1.2921 0.65187 15.9994 144.9922 0.00049602 4.471 0.0059501
1.11 0.98803 5.5187e-005 3.8182 0.012035 1.4611e-005 0.0011542 0.14914 0.00065826 0.14979 0.13649 0 0.037055 0.0389 0 0.8972 0.24993 0.067058 0.0093651 4.2473 0.058486 7.0246e-005 0.83158 0.005266 0.0060033 0.99603 -1.257e-010 0.16287 0.96373 0.98877 0.13179 0.7617 0.80235 0.76716 0.83606 0.53928 0.19524 0.43029 1.2023 0.71284 15.9991 144.9906 0.0005247 2.373 0.0069501
1.111 0.98803 5.5187e-005 3.8182 0.012035 1.4624e-005 0.0011542 0.14921 0.00065827 0.14986 0.13656 0 0.037051 0.0389 0 0.89727 0.24996 0.06707 0.0093666 4.2476 0.058495 7.0258e-005 0.83158 0.0052663 0.0060037 0.99515 -5.8357e-011 0.1219 0.95095 0.98471 0.1318 0.73732 0.77677 0.76069 0.81255 0.52813 0.21089 0.43009 1.1353 0.77089 15.9988 144.9892 0.00054623 0.56388 0.0079501
1.112 0.98803 5.5187e-005 3.8182 0.012035 1.4637e-005 0.0011542 0.14928 0.00065827 0.14993 0.13662 0 0.037046 0.0389 0 0.89735 0.24999 0.067082 0.0093681 4.248 0.058504 7.027e-005 0.83157 0.0052667 0.006004 0.99414 1.4055e-011 0.091401 0.93618 0.97986 0.1318 0.71515 0.75238 0.74892 0.7897 0.51804 0.22446 0.42988 1.087 0.82185 15.9985 144.9879 0.00056235 -1.1365 0.0089501
1.113 0.98803 5.5187e-005 3.8182 0.012035 1.465e-005 0.0011542 0.14935 0.00065827 0.15 0.13669 0 0.037042 0.0389 0 0.89743 0.25003 0.067094 0.0093696 4.2483 0.058513 7.0282e-005 0.83156 0.005267 0.0060044 0.99293 2.9946e-011 0.068681 0.91873 0.97386 0.1318 0.69505 0.72951 0.73335 0.76751 0.50902 0.23617 0.42968 1.0531 0.86398 15.9983 144.9866 0.00057446 -2.8369 0.0099501
1.114 0.98803 5.5187e-005 3.8182 0.012035 1.4664e-005 0.0011542 0.14942 0.00065827 0.15007 0.13675 0 0.037037 0.0389 0 0.8975 0.25006 0.067107 0.0093711 4.2486 0.058523 7.0293e-005 0.83155 0.0052674 0.0060047 0.99138 -1.9804e-011 0.05174 0.8976 0.96619 0.13181 0.67695 0.70845 0.71465 0.74596 0.50105 0.24619 0.42947 1.0302 0.89724 15.998 144.9854 0.00058366 -4.6236 0.01095
1.115 0.98803 5.5187e-005 3.8182 0.012035 1.4677e-005 0.0011542 0.14948 0.00065827 0.15014 0.13682 0 0.037033 0.0389 0 0.89758 0.2501 0.067119 0.0093726 4.249 0.058532 7.0305e-005 0.83154 0.0052677 0.0060051 0.98928 3.1276e-012 0.039104 0.87134 0.95603 0.13181 0.66083 0.68944 0.69304 0.72503 0.49416 0.25456 0.42927 1.0151 0.92264 15.9978 144.9843 0.00059069 -6.5864 0.01195
1.116 0.98803 5.5187e-005 3.8182 0.012035 1.469e-005 0.0011542 0.14955 0.00065827 0.15021 0.13688 0 0.037029 0.0389 0 0.89765 0.25013 0.067131 0.0093741 4.2493 0.058541 7.0317e-005 0.83153 0.0052681 0.0060054 0.98623 6.0401e-012 0.02968 0.8378 0.94209 0.13181 0.64671 0.67273 0.66839 0.70473 0.48839 0.26133 0.42907 1.0058 0.94161 15.9975 144.9834 0.00059608 -8.8372 0.01295
1.117 0.98803 5.5187e-005 3.8182 0.012035 1.4703e-005 0.0011542 0.14962 0.00065827 0.15028 0.13695 0 0.037024 0.0389 0 0.89773 0.25016 0.067143 0.0093756 4.2496 0.05855 7.0329e-005 0.83152 0.0052685 0.0060058 0.98143 -9.5273e-012 0.022665 0.79375 0.92218 0.13181 0.63468 0.65857 0.64037 0.68505 0.48377 0.26648 0.42886 1.0003 0.95563 15.9973 144.9825 0.00060011 -11.5283 0.01395
1.118 0.98803 5.5187e-005 3.8182 0.012035 1.4716e-005 0.0011542 0.14969 0.00065828 0.15035 0.13701 0 0.03702 0.0389 0 0.89781 0.2502 0.067155 0.0093771 4.25 0.058559 7.034e-005 0.83151 0.0052688 0.0060061 0.97307 7.2519e-012 0.017469 0.73425 0.89257 0.13182 0.6248 0.64721 0.60855 0.66602 0.4803 0.26998 0.42866 0.99756 0.96602 15.9971 144.9817 0.0006029 -14.8664 0.01495
1.119 0.98803 5.5187e-005 3.8182 0.012035 1.4729e-005 0.0011542 0.14976 0.00065828 0.15041 0.13708 0 0.037015 0.0389 0 0.89788 0.25023 0.067167 0.0093786 4.2503 0.058568 7.0352e-005 0.8315 0.0052692 0.0060065 0.95689 -6.4107e-012 0.013666 0.65215 0.84691 0.13182 0.61713 0.63885 0.57266 0.64772 0.47792 0.27187 0.42845 0.99659 0.97395 15.9969 144.981 0.00060446 -19.0978 0.01595
1.12 0.98803 5.5187e-005 3.8182 0.012035 1.4742e-005 0.0011542 0.14983 0.00065828 0.15048 0.13714 0 0.037011 0.0389 0 0.89796 0.25026 0.06718 0.0093801 4.2506 0.058578 7.0364e-005 0.83149 0.0052695 0.0060069 0.92256 1.4451e-012 0.010956 0.53887 0.77505 0.13182 0.61152 0.63346 0.53278 0.63038 0.47647 0.27225 0.42825 0.99686 0.98048 15.9967 144.9804 0.00060469 -24.3882 0.01695
1.121 0.98803 5.5187e-005 3.8182 0.012035 1.4756e-005 0.0011542 0.1499 0.00065828 0.15055 0.1372 0 0.037006 0.0389 0 0.89803 0.2503 0.067192 0.0093816 4.251 0.058587 7.0376e-005 0.83148 0.0052699 0.0060072 0.84954 6.0192e-013 0.0091182 0.39118 0.66433 0.13183 0.60759 0.63052 0.4887 0.61469 0.47569 0.27138 0.42805 0.99798 0.98566 15.9966 144.9799 0.00060383 -30.5075 0.01795
1.122 0.98803 5.5187e-005 3.8182 0.012035 1.4769e-005 0.0011542 0.14997 0.00065828 0.15062 0.13727 0 0.037002 0.0389 0 0.89811 0.25033 0.067204 0.0093831 4.2513 0.058596 7.0388e-005 0.83147 0.0052702 0.0060076 0.71964 1.6942e-012 0.0079421 0.22897 0.51047 0.13183 0.60479 0.629 0.43823 0.60219 0.47532 0.26938 0.42785 0.99962 0.98972 15.9964 144.9795 0.00060236 -36.6101 0.01895
1.123 0.98803 5.5187e-005 3.8182 0.012035 1.4782e-005 0.0011542 0.15004 0.00065828 0.15069 0.13733 0 0.036998 0.0389 0 0.89819 0.25037 0.067216 0.0093846 4.2517 0.058605 7.0399e-005 0.83147 0.0052706 0.0060079 0.55489 0.0001495 0.0072449 0.099188 0.336 0.13183 0.60271 0.62809 0.37811 0.59474 0.47518 0.26611 0.42765 1.0016 0.99309 15.9963 144.9792 0.00060067 -41.8686 0.01995
1.124 0.98803 5.5186e-005 3.8182 0.012035 1.4795e-005 0.0011542 0.1501 0.00065828 0.15076 0.1374 0 0.036993 0.0389 0 0.89826 0.2504 0.067229 0.0093861 4.252 0.058614 7.0411e-005 0.83146 0.0052709 0.0060083 0.40406 0.00077534 0.0070435 0.030608 0.18376 0.13184 0.60115 0.62773 0.30845 0.59205 0.47517 0.26123 0.42745 1.0037 0.99606 15.9963 144.979 0.00059891 -46.111 0.02095
1.125 0.98803 5.5186e-005 3.8182 0.012035 1.4808e-005 0.0011542 0.15017 0.00065828 0.15083 0.13746 0 0.036989 0.0389 0 0.89834 0.25043 0.067241 0.0093876 4.2523 0.058623 7.0423e-005 0.83145 0.0052713 0.0060087 0.29267 0.0018586 0.0072939 0.0073437 0.082925 0.13184 0.6 0.62817 0.23497 0.592 0.47522 0.2545 0.42726 1.0059 0.9988 15.9962 144.9789 0.00059712 -49.4637 0.02195
1.126 0.98803 5.5186e-005 3.8182 0.012035 1.4821e-005 0.0011542 0.15024 0.00065829 0.15089 0.13753 0 0.036984 0.0389 0 0.89842 0.25047 0.067253 0.0093891 4.2527 0.058633 7.0435e-005 0.83144 0.0052717 0.006009 0.21846 0.0035327 0.0079726 0.0020156 0.031801 0.13184 0.59919 0.62931 0.16664 0.59293 0.4753 0.24584 0.42707 1.0082 1.0014 15.9962 144.9787 0.0005953 -52.091 0.02295
1.127 0.98803 5.5186e-005 3.8182 0.012035 1.4834e-005 0.0011542 0.15031 0.00065829 0.15096 0.13759 0 0.03698 0.0389 0 0.89849 0.2505 0.067265 0.0093906 4.253 0.058642 7.0447e-005 0.83143 0.005272 0.0060094 0.16988 0.0058819 0.0090525 0.00095971 0.011387 0.13184 0.59865 0.63082 0.11094 0.59415 0.47541 0.23541 0.42688 1.0105 1.0039 15.9961 144.9787 0.00059345 -54.1667 0.02395
1.128 0.98803 5.5186e-005 3.8182 0.012035 1.4847e-005 0.0011542 0.15038 0.00065829 0.15103 0.13765 0 0.036976 0.0389 0 0.89857 0.25054 0.067277 0.0093921 4.2534 0.058651 7.0459e-005 0.83142 0.0052724 0.0060098 0.13695 0.0089538 0.010507 0.00064731 0.0045865 0.13185 0.59833 0.63247 0.070766 0.59542 0.47552 0.22349 0.4267 1.0129 1.0064 15.9961 144.9786 0.0005916 -55.8554 0.02495
1.129 0.98803 5.5186e-005 3.8182 0.012035 1.4861e-005 0.0011542 0.15045 0.00065829 0.1511 0.13772 0 0.036971 0.0389 0 0.89865 0.25057 0.06729 0.0093936 4.2537 0.05866 7.047e-005 0.83141 0.0052727 0.0060101 0.11326 0.012785 0.012318 0.00048703 0.0024652 0.13185 0.59818 0.63416 0.044674 0.59668 0.47564 0.21038 0.42652 1.0152 1.0088 15.9961 144.9786 0.00058973 -57.2926 0.02595
1.13 0.98803 5.5186e-005 3.8182 0.012035 1.4874e-005 0.0011542 0.15051 0.00065829 0.15117 0.13778 0 0.036967 0.0389 0 0.89872 0.2506 0.067302 0.0093951 4.254 0.058669 7.0482e-005 0.8314 0.0052731 0.0060105 0.095165 0.017425 0.014479 0.0003822 0.0016975 0.13185 0.59817 0.63584 0.029111 0.59789 0.47576 0.19637 0.42634 1.0176 1.0112 15.9961 144.9785 0.00058786 -58.5756 0.02695
1.131 0.98803 5.5186e-005 3.8182 0.012035 1.4887e-005 0.0011542 0.15058 0.00065829 0.15124 0.13784 0 0.036962 0.0389 0 0.8988 0.25064 0.067314 0.0093966 4.2544 0.058679 7.0494e-005 0.83139 0.0052735 0.0060108 0.080686 0.022949 0.016997 0.00030665 0.0013081 0.13186 0.5983 0.63752 0.020371 0.59906 0.47588 0.1817 0.42617 1.0199 1.0136 15.9961 144.9785 0.00058598 -59.7667 0.02795
1.132 0.98803 5.5186e-005 3.8182 0.012035 1.49e-005 0.0011542 0.15065 0.00065829 0.1513 0.13791 0 0.036958 0.0389 0 0.89887 0.25067 0.067327 0.0093981 4.2547 0.058688 7.0506e-005 0.83138 0.0052738 0.0060112 0.068742 0.029457 0.019891 0.00024922 0.0010484 0.13186 0.59853 0.63919 0.015573 0.60018 0.47601 0.16659 0.42599 1.0223 1.016 15.9961 144.9785 0.0005841 -60.9016 0.02895
1.133 0.98803 5.5186e-005 3.8182 0.012035 1.4913e-005 0.0011542 0.15072 0.00065829 0.15137 0.13797 0 0.036954 0.0389 0 0.89895 0.25071 0.067339 0.0093996 4.2551 0.058697 7.0518e-005 0.83137 0.0052742 0.0060116 0.058726 0.037076 0.023186 0.0002042 0.00085276 0.13186 0.59887 0.64084 0.012848 0.60127 0.47614 0.15125 0.42583 1.0247 1.0184 15.9961 144.9785 0.00058222 -61.9992 0.02995
1.134 0.98803 5.5186e-005 3.8182 0.012035 1.4926e-005 0.0011542 0.15079 0.0006583 0.15144 0.13804 0 0.036949 0.0389 0 0.89903 0.25074 0.067351 0.0094011 4.2554 0.058706 7.053e-005 0.83136 0.0052745 0.0060119 0.05026 0.04595 0.026914 0.00016829 0.00069928 0.13187 0.5993 0.64248 0.01114 0.60231 0.47626 0.13588 0.42566 1.027 1.0207 15.9961 144.9784 0.00058033 -63.0687 0.03095
1.135 0.98803 5.5186e-005 3.8182 0.012035 1.4939e-005 0.0011542 0.15085 0.0006583 0.15151 0.1381 0 0.036945 0.0389 0 0.8991 0.25077 0.067363 0.0094026 4.2557 0.058716 7.0541e-005 0.83135 0.0052749 0.0060123 0.04308 0.05624 0.031112 0.00013939 0.00057669 0.13187 0.59981 0.64411 0.0099193 0.60333 0.47639 0.12071 0.4255 1.0294 1.0231 15.9961 144.9784 0.00057844 -64.1142 0.03195
1.136 0.98803 5.5186e-005 3.8182 0.012035 1.4953e-005 0.0011542 0.15092 0.0006583 0.15158 0.13816 0 0.03694 0.0389 0 0.89918 0.25081 0.067376 0.0094041 4.2561 0.058725 7.0553e-005 0.83135 0.0052753 0.0060127 0.036984 0.068114 0.035819 0.00011593 0.00047805 0.13187 0.60039 0.64572 0.0089473 0.60432 0.47652 0.10595 0.42535 1.0317 1.0255 15.9962 144.9784 0.00057655 -65.1372 0.03295
1.137 0.98803 5.5186e-005 3.8182 0.012035 1.4966e-005 0.0011542 0.15099 0.0006583 0.15164 0.13823 0 0.036936 0.0389 0 0.89926 0.25084 0.067388 0.0094056 4.2564 0.058734 7.0565e-005 0.83134 0.0052756 0.006013 0.031805 0.08175 0.04108 9.6862e-005 0.00039809 0.13187 0.60104 0.64732 0.0081238 0.60529 0.47665 0.09182 0.4252 1.0341 1.0279 15.9962 144.9784 0.00057465 -66.1386 0.03395
1.138 0.98803 5.5186e-005 3.8182 0.012035 1.4979e-005 0.0011542 0.15106 0.0006583 0.15171 0.13829 0 0.036932 0.0389 0 0.89933 0.25088 0.0674 0.0094071 4.2568 0.058743 7.0577e-005 0.83133 0.005276 0.0060134 0.027404 0.097324 0.046945 8.1239e-005 0.00033304 0.13188 0.60176 0.6489 0.0074056 0.60624 0.47678 0.078522 0.42505 1.0364 1.0302 15.9962 144.9783 0.00057276 -67.118 0.03495
1.139 0.98803 5.5186e-005 3.8182 0.012035 1.4992e-005 0.0011542 0.15113 0.0006583 0.15178 0.13835 0 0.036927 0.0389 0 0.89941 0.25091 0.067413 0.0094086 4.2571 0.058752 7.0589e-005 0.83132 0.0052764 0.0060138 0.023664 0.11501 0.053468 6.8438e-005 0.00027985 0.13188 0.60252 0.65048 0.0067722 0.60719 0.47691 0.066231 0.42491 1.0388 1.0326 15.9962 144.9783 0.00057086 -68.0752 0.03595
1.14 0.98803 5.5185e-005 3.8182 0.012035 1.5005e-005 0.0011542 0.15119 0.0006583 0.15185 0.13842 0 0.036923 0.0389 0 0.89949 0.25094 0.067425 0.0094101 4.2575 0.058762 7.0601e-005 0.83131 0.0052767 0.0060141 0.020485 0.13496 0.060709 5.7888e-005 0.00023625 0.13188 0.60333 0.65203 0.0062105 0.60813 0.47704 0.055088 0.42477 1.0411 1.035 15.9963 144.9783 0.00056897 -69.0093 0.03695
1.141 0.98803 5.5185e-005 3.8182 0.012035 1.5018e-005 0.0011542 0.15126 0.00065831 0.15191 0.13848 0 0.036919 0.0389 0 0.89957 0.25098 0.067437 0.0094116 4.2578 0.058771 7.0613e-005 0.8313 0.0052771 0.0060145 0.017783 0.15732 0.068736 4.9196e-005 0.00020037 0.13189 0.60419 0.65358 0.0057112 0.60907 0.47717 0.04519 0.42464 1.0434 1.0373 15.9963 144.9782 0.00056707 -69.9194 0.03795
1.142 0.98803 5.5185e-005 3.8182 0.012035 1.5031e-005 0.0011542 0.15133 0.00065831 0.15198 0.13854 0 0.036914 0.0389 0 0.89964 0.25101 0.067449 0.0094131 4.2582 0.05878 7.0625e-005 0.83129 0.0052774 0.0060149 0.015485 0.18218 0.077623 4.2e-005 0.00017075 0.13189 0.60508 0.65511 0.0052664 0.61002 0.47731 0.036586 0.42451 1.0458 1.0397 15.9964 144.9782 0.00056517 -70.804 0.03895
1.143 0.98803 5.5185e-005 3.8182 0.012035 1.5045e-005 0.0011542 0.1514 0.00065831 0.15205 0.13861 0 0.03691 0.0389 0 0.89972 0.25105 0.067462 0.0094146 4.2585 0.058789 7.0637e-005 0.83128 0.0052778 0.0060152 0.01353 0.20961 0.087449 3.6032e-005 0.00014626 0.13189 0.606 0.65663 0.0048699 0.61098 0.47744 0.029273 0.42439 1.0481 1.042 15.9964 144.9782 0.00056328 -71.6618 0.03995
1.144 0.98803 5.5185e-005 3.8182 0.012035 1.5058e-005 0.0011542 0.15146 0.00065831 0.15212 0.13867 0 0.036906 0.0389 0 0.8998 0.25108 0.067474 0.0094161 4.2589 0.058799 7.0648e-005 0.83127 0.0052782 0.0060156 0.011868 0.23959 0.098298 3.1073e-005 0.00012595 0.1319 0.60695 0.65814 0.0045162 0.61195 0.47758 0.0232 0.42428 1.0504 1.0444 15.9965 144.9782 0.00056138 -72.4912 0.04095
1.145 0.98803 5.5185e-005 3.8182 0.012035 1.5071e-005 0.0011542 0.15153 0.00065831 0.15218 0.13873 0 0.036901 0.0389 0 0.89987 0.25111 0.067486 0.0094176 4.2592 0.058808 7.066e-005 0.83126 0.0052785 0.006016 0.010453 0.27207 0.11025 2.694e-005 0.00010906 0.1319 0.60792 0.65963 0.0042006 0.61295 0.47771 0.018277 0.42417 1.0528 1.0467 15.9965 144.9781 0.00055949 -73.2905 0.04195
1.146 0.98803 5.5185e-005 3.8182 0.012035 1.5084e-005 0.0011542 0.1516 0.00065831 0.15225 0.1388 0 0.036897 0.0389 0 0.89995 0.25115 0.067499 0.0094191 4.2596 0.058817 7.0672e-005 0.83125 0.0052789 0.0060163 0.0092481 0.30688 0.12339 2.3494e-005 9.4994e-005 0.1319 0.60892 0.66112 0.0039191 0.61396 0.47785 0.01438 0.42406 1.0551 1.0491 15.9966 144.9781 0.00055759 -74.0581 0.04295
1.147 0.98803 5.5185e-005 3.8182 0.012035 1.5097e-005 0.0011542 0.15167 0.00065831 0.15232 0.13886 0 0.036893 0.0389 0 0.90003 0.25118 0.067511 0.0094207 4.2599 0.058827 7.0684e-005 0.83124 0.0052793 0.0060167 0.0082227 0.34379 0.13778 2.0611e-005 8.3242e-005 0.1319 0.60993 0.66259 0.003668 0.61501 0.47799 0.011366 0.42397 1.0574 1.0514 15.9967 144.9781 0.0005557 -74.7925 0.04395
1.148 0.98803 5.5185e-005 3.8182 0.012035 1.511e-005 0.0011542 0.15173 0.00065831 0.15239 0.13892 0 0.036888 0.0389 0 0.9001 0.25122 0.067523 0.0094222 4.2602 0.058836 7.0696e-005 0.83123 0.0052796 0.0060171 0.007348 0.38249 0.15347 1.8192e-005 7.3407e-005 0.13191 0.61095 0.66404 0.0034441 0.61608 0.47813 0.0090856 0.42387 1.0597 1.0537 15.9967 144.978 0.00055382 -75.4923 0.04495
1.149 0.98803 5.5185e-005 3.8182 0.012035 1.5123e-005 0.0011542 0.1518 0.00065832 0.15245 0.13898 0 0.036884 0.0389 0 0.90018 0.25125 0.067536 0.0094237 4.2606 0.058845 7.0708e-005 0.83123 0.00528 0.0060174 0.0066022 0.42257 0.17047 1.6162e-005 6.5155e-005 0.13191 0.61199 0.66549 0.0032446 0.61719 0.47827 0.007394 0.42379 1.062 1.0561 15.9968 144.978 0.00055193 -76.1565 0.04595
1.15 0.98803 5.5185e-005 3.8182 0.012035 1.5137e-005 0.0011542 0.15187 0.00065832 0.15252 0.13905 0 0.03688 0.0389 0 0.90026 0.25129 0.067548 0.0094252 4.2609 0.058854 7.072e-005 0.83122 0.0052804 0.0060178 0.0059651 0.46358 0.18878 1.4451e-005 5.8213e-005 0.13191 0.61304 0.66692 0.003067 0.61833 0.47842 0.0061587 0.42371 1.0643 1.0584 15.9969 144.978 0.00055005 -76.7842 0.04695
1.151 0.98803 5.5185e-005 3.8182 0.012035 1.515e-005 0.0011542 0.15193 0.00065832 0.15259 0.13911 0 0.036876 0.0389 0 0.90034 0.25132 0.067561 0.0094267 4.2613 0.058864 7.0732e-005 0.83121 0.0052807 0.0060182 0.0054207 0.50499 0.20833 1.3008e-005 5.2359e-005 0.13192 0.6141 0.66834 0.0029089 0.61951 0.47856 0.005266 0.42363 1.0666 1.0607 15.9969 144.978 0.00054817 -77.375 0.04795
1.152 0.98803 5.5185e-005 3.8182 0.012035 1.5163e-005 0.0011542 0.152 0.00065832 0.15266 0.13917 0 0.036871 0.0389 0 0.90041 0.25135 0.067573 0.0094282 4.2616 0.058873 7.0744e-005 0.8312 0.0052811 0.0060186 0.004954 0.54629 0.22905 1.1786e-005 4.7411e-005 0.13192 0.61517 0.66975 0.0027683 0.62073 0.47871 0.0046229 0.42356 1.069 1.0631 15.997 144.9779 0.0005463 -77.9289 0.04895
1.153 0.98803 5.5185e-005 3.8182 0.012035 1.5176e-005 0.0011542 0.15207 0.00065832 0.15272 0.13924 0 0.036867 0.0389 0 0.90049 0.25139 0.067585 0.0094297 4.262 0.058882 7.0756e-005 0.83119 0.0052815 0.0060189 0.0045537 0.58691 0.25082 1.0749e-005 4.3215e-005 0.13192 0.61624 0.67115 0.0026433 0.62198 0.47885 0.0041571 0.4235 1.0713 1.0654 15.9971 144.9779 0.00054444 -78.446 0.04995
1.154 0.98803 5.5185e-005 3.8182 0.012035 1.5189e-005 0.0011542 0.15214 0.00065832 0.15279 0.1393 0 0.036863 0.0389 0 0.90057 0.25142 0.067598 0.0094312 4.2624 0.058892 7.0768e-005 0.83118 0.0052818 0.0060193 0.0042103 0.62637 0.27349 9.8672e-006 3.9646e-005 0.13193 0.61731 0.67254 0.0025323 0.62328 0.479 0.003815 0.42344 1.0736 1.0677 15.9972 144.9779 0.00054257 -78.9271 0.05095
1.155 0.98803 5.5185e-005 3.8182 0.012035 1.5202e-005 0.0011542 0.1522 0.00065832 0.15286 0.13936 0 0.036858 0.0389 0 0.90064 0.25146 0.06761 0.0094328 4.2627 0.058901 7.078e-005 0.83117 0.0052822 0.0060197 0.0039142 0.66419 0.2969 9.1144e-006 3.6604e-005 0.13193 0.61839 0.67391 0.0024336 0.62461 0.47915 0.0035579 0.42338 1.0758 1.07 15.9973 144.9779 0.00054072 -79.373 0.05195
1.156 0.98803 5.5184e-005 3.8182 0.012035 1.5215e-005 0.0011542 0.15227 0.00065832 0.15292 0.13942 0 0.036854 0.0389 0 0.90072 0.25149 0.067622 0.0094343 4.2631 0.05891 7.0792e-005 0.83116 0.0052826 0.00602 0.003659 0.69999 0.32087 8.4702e-006 3.4002e-005 0.13193 0.61948 0.67528 0.0023459 0.62599 0.47931 0.0033595 0.42333 1.0781 1.0723 15.9974 144.9779 0.00053887 -79.7849 0.05295
1.157 0.98803 5.5184e-005 3.8182 0.012035 1.5228e-005 0.0011542 0.15234 0.00065833 0.15299 0.13949 0 0.03685 0.0389 0 0.9008 0.25153 0.067635 0.0094358 4.2634 0.058919 7.0804e-005 0.83115 0.005283 0.0060204 0.0034385 0.73346 0.34523 7.9174e-006 3.1771e-005 0.13194 0.62056 0.67663 0.002268 0.6274 0.47946 0.0032017 0.42329 1.0804 1.0746 15.9974 144.9779 0.00053702 -80.1642 0.05395
1.158 0.98803 5.5184e-005 3.8182 0.012035 1.5242e-005 0.0011542 0.1524 0.00065833 0.15306 0.13955 0 0.036846 0.0389 0 0.90088 0.25156 0.067647 0.0094373 4.2638 0.058929 7.0816e-005 0.83114 0.0052833 0.0060208 0.0032473 0.76438 0.36982 7.4415e-006 2.9851e-005 0.13194 0.62165 0.67797 0.0021987 0.62885 0.47962 0.0030728 0.42324 1.0827 1.0769 15.9975 144.9778 0.00053519 -80.5126 0.05495
1.159 0.98803 5.5184e-005 3.8182 0.012035 1.5255e-005 0.0011542 0.15247 0.00065833 0.15312 0.13961 0 0.036841 0.0389 0 0.90095 0.25159 0.06766 0.0094388 4.2641 0.058938 7.0828e-005 0.83113 0.0052837 0.0060212 0.0030814 0.79262 0.39446 7.0308e-006 2.8195e-005 0.13194 0.62273 0.67931 0.0021372 0.63033 0.47977 0.002965 0.4232 1.085 1.0792 15.9976 144.9778 0.00053336 -80.8318 0.05595
1.16 0.98803 5.5184e-005 3.8182 0.012035 1.5268e-005 0.0011542 0.15254 0.00065833 0.15319 0.13967 0 0.036837 0.0389 0 0.90103 0.25163 0.067672 0.0094403 4.2645 0.058947 7.084e-005 0.83112 0.0052841 0.0060215 0.0029369 0.81814 0.419 6.6753e-006 2.6762e-005 0.13194 0.62382 0.68063 0.0020825 0.63184 0.47993 0.0028731 0.42317 1.0873 1.0815 15.9977 144.9778 0.00053153 -81.1235 0.05695
1.161 0.98803 5.5184e-005 3.8182 0.012035 1.5281e-005 0.0011542 0.1526 0.00065833 0.15326 0.13974 0 0.036833 0.0389 0 0.90111 0.25166 0.067684 0.0094419 4.2648 0.058957 7.0852e-005 0.83111 0.0052844 0.0060219 0.0028111 0.84097 0.44332 6.3669e-006 2.5519e-005 0.13195 0.62491 0.68194 0.0020339 0.63339 0.48009 0.002794 0.42313 1.0895 1.0838 15.9978 144.9778 0.00052972 -81.3895 0.05795
1.162 0.98803 5.5184e-005 3.8182 0.012035 1.5294e-005 0.0011542 0.15267 0.00065833 0.15332 0.1398 0 0.036829 0.0389 0 0.90119 0.2517 0.067697 0.0094434 4.2652 0.058966 7.0864e-005 0.8311 0.0052848 0.0060223 0.0027011 0.86119 0.4673 6.0985e-006 2.4438e-005 0.13195 0.62599 0.68324 0.0019906 0.63496 0.48025 0.0027252 0.4231 1.0918 1.0861 15.9979 144.9778 0.00052791 -81.6318 0.05895
1.163 0.98803 5.5184e-005 3.8182 0.012035 1.5307e-005 0.0011542 0.15274 0.00065833 0.15339 0.13986 0 0.036824 0.0389 0 0.90126 0.25173 0.067709 0.0094449 4.2655 0.058975 7.0876e-005 0.8311 0.0052852 0.0060227 0.0026046 0.87895 0.49083 5.8642e-006 2.3495e-005 0.13195 0.62708 0.68453 0.0019521 0.63656 0.48041 0.002665 0.42308 1.0941 1.0884 15.998 144.9778 0.00052611 -81.8521 0.05995
1.164 0.98803 5.5184e-005 3.8182 0.012035 1.532e-005 0.0011542 0.1528 0.00065833 0.15346 0.13992 0 0.03682 0.0389 0 0.90134 0.25177 0.067722 0.0094464 4.2659 0.058985 7.0888e-005 0.83109 0.0052856 0.006023 0.0025201 0.89443 0.51382 5.6594e-006 2.267e-005 0.13196 0.62816 0.68581 0.0019178 0.63819 0.48057 0.002612 0.42305 1.0964 1.0907 15.9981 144.9778 0.00052432 -82.0521 0.06095
1.165 0.98803 5.5184e-005 3.8182 0.012034 1.5334e-005 0.0011542 0.15287 0.00065834 0.15352 0.13998 0 0.036816 0.0389 0 0.90142 0.2518 0.067734 0.0094479 4.2662 0.058994 7.09e-005 0.83108 0.0052859 0.0060234 0.0024457 0.90781 0.53622 5.4797e-006 2.1947e-005 0.13196 0.62925 0.68709 0.0018872 0.63983 0.48073 0.0025651 0.42303 1.0986 1.093 15.9982 144.9778 0.00052254 -82.2336 0.06195
1.166 0.98803 5.5184e-005 3.8182 0.012034 1.5347e-005 0.0011542 0.15293 0.00065834 0.15359 0.14005 0 0.036812 0.0389 0 0.9015 0.25184 0.067747 0.0094494 4.2666 0.059003 7.0912e-005 0.83107 0.0052863 0.0060238 0.00238 0.91931 0.55796 5.3218e-006 2.1311e-005 0.13196 0.63033 0.68835 0.0018598 0.64149 0.48089 0.0025236 0.423 1.1009 1.0952 15.9982 144.9778 0.00052077 -82.3982 0.06295
1.167 0.98803 5.5184e-005 3.8182 0.012034 1.536e-005 0.0011542 0.153 0.00065834 0.15365 0.14011 0 0.036807 0.0389 0 0.90157 0.25187 0.067759 0.009451 4.267 0.059013 7.0924e-005 0.83106 0.0052867 0.0060242 0.002322 0.92913 0.579 5.1826e-006 2.0752e-005 0.13197 0.63141 0.6896 0.0018354 0.64317 0.48106 0.0024869 0.42298 1.1031 1.0975 15.9983 144.9778 0.000519 -82.5473 0.06395
1.168 0.98803 5.5184e-005 3.8182 0.012034 1.5373e-005 0.0011542 0.15307 0.00065834 0.15372 0.14017 0 0.036803 0.0389 0 0.90165 0.2519 0.067771 0.0094525 4.2673 0.059022 7.0936e-005 0.83105 0.005287 0.0060245 0.0022707 0.93747 0.59931 5.0596e-006 2.0257e-005 0.13197 0.63249 0.69084 0.0018136 0.64487 0.48122 0.0024542 0.42296 1.1054 1.0998 15.9984 144.9778 0.00051724 -82.6824 0.06495
1.169 0.98803 5.5184e-005 3.8182 0.012034 1.5386e-005 0.0011542 0.15313 0.00065834 0.15379 0.14023 0 0.036799 0.0389 0 0.90173 0.25194 0.067784 0.009454 4.2677 0.059031 7.0948e-005 0.83104 0.0052874 0.0060249 0.0022253 0.94452 0.61888 4.9508e-006 1.9819e-005 0.13197 0.63356 0.69207 0.0017941 0.64657 0.48139 0.0024251 0.42295 1.1076 1.1021 15.9985 144.9778 0.0005155 -82.8048 0.06595
1.17 0.98803 5.5184e-005 3.8182 0.012034 1.5399e-005 0.0011542 0.1532 0.00065834 0.15385 0.14029 0 0.036795 0.0389 0 0.90181 0.25197 0.067796 0.0094555 4.268 0.059041 7.096e-005 0.83103 0.0052878 0.0060253 0.0021847 0.95046 0.63768 4.8542e-006 1.9431e-005 0.13198 0.63463 0.6933 0.0017765 0.64829 0.48155 0.0023991 0.42293 1.1099 1.1043 15.9986 144.9778 0.00051376 -82.9157 0.06695
1.171 0.98803 5.5184e-005 3.8182 0.012034 1.5412e-005 0.0011542 0.15327 0.00065834 0.15392 0.14036 0 0.036791 0.0389 0 0.90188 0.25201 0.067809 0.0094571 4.2684 0.05905 7.0972e-005 0.83102 0.0052882 0.0060257 0.0021485 0.95544 0.65572 4.7682e-006 1.9086e-005 0.13198 0.6357 0.69451 0.0017608 0.65002 0.48172 0.0023759 0.42292 1.1121 1.1066 15.9987 144.9778 0.00051203 -83.0162 0.06795
1.172 0.98803 5.5183e-005 3.8182 0.012034 1.5426e-005 0.0011542 0.15333 0.00065834 0.15398 0.14042 0 0.036786 0.0389 0 0.90196 0.25204 0.067821 0.0094586 4.2688 0.05906 7.0984e-005 0.83101 0.0052885 0.0060261 0.0021163 0.9596 0.673 4.6915e-006 1.8777e-005 0.13198 0.63677 0.69572 0.0017466 0.65175 0.48188 0.0023551 0.4229 1.1143 1.1088 15.9988 144.9778 0.00051031 -83.1075 0.06895
1.173 0.98803 5.5183e-005 3.8182 0.012034 1.5439e-005 0.0011542 0.1534 0.00065834 0.15405 0.14048 0 0.036782 0.0389 0 0.90204 0.25208 0.067834 0.0094601 4.2691 0.059069 7.0996e-005 0.831 0.0052889 0.0060264 0.0020877 0.96308 0.68953 4.6231e-006 1.8502e-005 0.13198 0.63784 0.69691 0.0017339 0.65349 0.48205 0.0023364 0.42289 1.1166 1.1111 15.9989 144.9778 0.00050859 -83.1903 0.06995
1.174 0.98803 5.5183e-005 3.8182 0.012034 1.5452e-005 0.0011542 0.15346 0.00065835 0.15412 0.14054 0 0.036778 0.0389 0 0.90212 0.25211 0.067846 0.0094616 4.2695 0.059078 7.1008e-005 0.83099 0.0052893 0.0060268 0.0020615 0.96598 0.70531 4.5616e-006 1.8255e-005 0.13199 0.6389 0.6981 0.0017224 0.65524 0.48222 0.0023197 0.42288 1.1188 1.1133 15.999 144.9778 0.00050689 -83.2656 0.07095
1.175 0.98803 5.5183e-005 3.8182 0.012034 1.5465e-005 0.0011542 0.15353 0.00065835 0.15418 0.1406 0 0.036774 0.0389 0 0.9022 0.25215 0.067859 0.0094632 4.2698 0.059088 7.102e-005 0.83098 0.0052897 0.0060272 0.0020385 0.96839 0.72037 4.5065e-006 1.8034e-005 0.13199 0.63996 0.69928 0.001712 0.65698 0.48238 0.0023046 0.42287 1.121 1.1156 15.9991 144.9778 0.0005052 -83.3341 0.07195
1.176 0.98803 5.5183e-005 3.8182 0.012034 1.5478e-005 0.0011542 0.15359 0.00065835 0.15425 0.14066 0 0.03677 0.0389 0 0.90227 0.25218 0.067871 0.0094647 4.2702 0.059097 7.1032e-005 0.83097 0.0052901 0.0060276 0.0020175 0.9704 0.73472 4.4568e-006 1.7834e-005 0.13199 0.64102 0.70045 0.0017026 0.65873 0.48255 0.002291 0.42286 1.1233 1.1178 15.9992 144.9778 0.00050351 -83.3966 0.07295
1.177 0.98803 5.5183e-005 3.8182 0.012034 1.5491e-005 0.0011542 0.15366 0.00065835 0.15431 0.14073 0 0.036765 0.0389 0 0.90235 0.25222 0.067884 0.0094662 4.2706 0.059106 7.1044e-005 0.83096 0.0052904 0.006028 0.001998 0.97207 0.74838 4.4118e-006 1.7654e-005 0.132 0.64207 0.70161 0.001694 0.66049 0.48272 0.0022786 0.42285 1.1255 1.1201 15.9992 144.9778 0.00050183 -83.4536 0.07395
1.178 0.98803 5.5183e-005 3.8182 0.012034 1.5504e-005 0.0011542 0.15373 0.00065835 0.15438 0.14079 0 0.036761 0.0389 0 0.90243 0.25225 0.067896 0.0094677 4.2709 0.059116 7.1056e-005 0.83096 0.0052908 0.0060283 0.0019811 0.97347 0.76137 4.3712e-006 1.749e-005 0.132 0.64313 0.70277 0.0016862 0.66224 0.48289 0.0022674 0.42284 1.1277 1.1223 15.9993 144.9778 0.00050017 -83.5058 0.07495
1.179 0.98803 5.5183e-005 3.8182 0.012034 1.5517e-005 0.0011542 0.15379 0.00065835 0.15445 0.14085 0 0.036757 0.0389 0 0.90251 0.25228 0.067909 0.0094693 4.2713 0.059125 7.1069e-005 0.83095 0.0052912 0.0060287 0.0019656 0.97463 0.77372 4.3342e-006 1.7342e-005 0.132 0.64417 0.70391 0.0016791 0.66399 0.48305 0.0022573 0.42283 1.1299 1.1245 15.9994 144.9778 0.00049851 -83.5536 0.07595
1.18 0.98803 5.5183e-005 3.8182 0.012034 1.5531e-005 0.0011542 0.15386 0.00065835 0.15451 0.14091 0 0.036753 0.0389 0 0.90259 0.25232 0.067921 0.0094708 4.2717 0.059135 7.1081e-005 0.83094 0.0052916 0.0060291 0.0019511 0.9756 0.78545 4.3005e-006 1.7207e-005 0.13201 0.64522 0.70505 0.0016726 0.66574 0.48322 0.002248 0.42282 1.1321 1.1267 15.9995 144.9778 0.00049686 -83.5976 0.07695
1.181 0.98803 5.5183e-005 3.8182 0.012034 1.5544e-005 0.0011542 0.15392 0.00065835 0.15458 0.14097 0 0.036749 0.0389 0 0.90266 0.25235 0.067934 0.0094723 4.272 0.059144 7.1093e-005 0.83093 0.0052919 0.0060295 0.0019379 0.97641 0.79658 4.2697e-006 1.7083e-005 0.13201 0.64626 0.70617 0.0016667 0.66749 0.48339 0.0022396 0.42281 1.1343 1.129 15.9996 144.9778 0.00049522 -83.6381 0.07795
1.182 0.98803 5.5183e-005 3.8182 0.012034 1.5557e-005 0.0011542 0.15399 0.00065836 0.15464 0.14103 0 0.036745 0.0389 0 0.90274 0.25239 0.067946 0.0094738 4.2724 0.059153 7.1105e-005 0.83092 0.0052923 0.0060299 0.0019265 0.9771 0.80715 4.2415e-006 1.697e-005 0.13201 0.6473 0.70729 0.0016612 0.66923 0.48356 0.0022318 0.42281 1.1365 1.1312 15.9997 144.9778 0.00049359 -83.6755 0.07895
1.183 0.98803 5.5183e-005 3.8182 0.012034 1.557e-005 0.0011542 0.15405 0.00065836 0.15471 0.14109 0 0.03674 0.0389 0 0.90282 0.25242 0.067959 0.0094754 4.2727 0.059163 7.1117e-005 0.83091 0.0052927 0.0060303 0.0019153 0.97767 0.81717 4.2155e-006 1.6865e-005 0.13202 0.64834 0.70841 0.0016561 0.67098 0.48373 0.0022247 0.4228 1.1387 1.1334 15.9998 144.9778 0.00049196 -83.7101 0.07995
1.184 0.98803 5.5183e-005 3.8182 0.012034 1.5583e-005 0.0011542 0.15412 0.00065836 0.15477 0.14115 0 0.036736 0.0389 0 0.9029 0.25246 0.067971 0.0094769 4.2731 0.059172 7.1129e-005 0.8309 0.0052931 0.0060306 0.0019051 0.97816 0.82666 4.1915e-006 1.6769e-005 0.13202 0.64938 0.70951 0.0016514 0.67272 0.4839 0.0022181 0.42279 1.1409 1.1356 15.9999 144.9779 0.00049035 -83.7423 0.08095
1.185 0.98803 5.5183e-005 3.8182 0.012034 1.5596e-005 0.0011542 0.15418 0.00065836 0.15484 0.14122 0 0.036732 0.0389 0 0.90298 0.25249 0.067984 0.0094784 4.2735 0.059182 7.1141e-005 0.83089 0.0052935 0.006031 0.0018956 0.97857 0.83566 4.1693e-006 1.668e-005 0.13202 0.65041 0.71061 0.0016471 0.67445 0.48406 0.002212 0.42279 1.1431 1.1378 15.9999 144.9779 0.00048874 -83.7722 0.08195
1.186 0.98803 5.5183e-005 3.8182 0.012034 1.5609e-005 0.0011542 0.15425 0.00065836 0.1549 0.14128 0 0.036728 0.0389 0 0.90305 0.25253 0.067996 0.00948 4.2738 0.059191 7.1153e-005 0.83088 0.0052938 0.0060314 0.0018867 0.97893 0.84417 4.1486e-006 1.6597e-005 0.13203 0.65143 0.71169 0.001643 0.67618 0.48423 0.0022064 0.42278 1.1453 1.14 16 144.9779 0.00048715 -83.8002 0.08295
1.187 0.98803 5.5183e-005 3.8182 0.012034 1.5623e-005 0.0011542 0.15431 0.00065836 0.15497 0.14134 0 0.036724 0.0389 0 0.90313 0.25256 0.068009 0.0094815 4.2742 0.0592 7.1165e-005 0.83087 0.0052942 0.0060318 0.0018784 0.97923 0.85224 4.1294e-006 1.652e-005 0.13203 0.65246 0.71277 0.0016392 0.67791 0.4844 0.0022011 0.42278 1.1475 1.1422 16.0001 144.9779 0.00048556 -83.8264 0.08395
1.188 0.98803 5.5182e-005 3.8182 0.012034 1.5636e-005 0.0011542 0.15438 0.00065836 0.15503 0.1414 0 0.03672 0.0389 0 0.90321 0.2526 0.068021 0.009483 4.2746 0.05921 7.1177e-005 0.83086 0.0052946 0.0060322 0.0018708 0.9795 0.85987 4.1114e-006 1.6448e-005 0.13203 0.65348 0.71385 0.0016357 0.67963 0.48457 0.0021962 0.42277 1.1496 1.1444 16.0002 144.9779 0.00048398 -83.851 0.08495
1.189 0.98803 5.5182e-005 3.8182 0.012034 1.5649e-005 0.0011542 0.15444 0.00065836 0.1551 0.14146 0 0.036716 0.0389 0 0.90329 0.25263 0.068034 0.0094846 4.2749 0.059219 7.119e-005 0.83085 0.005295 0.0060326 0.0018636 0.97973 0.8671 4.0945e-006 1.638e-005 0.13203 0.6545 0.71491 0.0016323 0.68135 0.48474 0.0021916 0.42277 1.1518 1.1466 16.0003 144.9779 0.00048241 -83.8742 0.08595
1.19 0.98803 5.5182e-005 3.8182 0.012034 1.5662e-005 0.0011542 0.15451 0.00065837 0.15516 0.14152 0 0.036711 0.0389 0 0.90337 0.25267 0.068046 0.0094861 4.2753 0.059229 7.1202e-005 0.83084 0.0052954 0.006033 0.0018569 0.97993 0.87393 4.0786e-006 1.6316e-005 0.13204 0.65552 0.71597 0.0016292 0.68306 0.48491 0.0021873 0.42276 1.154 1.1488 16.0004 144.9779 0.00048085 -83.8962 0.08695
1.191 0.98803 5.5182e-005 3.8182 0.012034 1.5675e-005 0.0011542 0.15457 0.00065837 0.15523 0.14158 0 0.036707 0.0389 0 0.90344 0.2527 0.068059 0.0094876 4.2757 0.059238 7.1214e-005 0.83083 0.0052957 0.0060333 0.0018505 0.98011 0.88039 4.0636e-006 1.6256e-005 0.13204 0.65653 0.71702 0.0016262 0.68477 0.48508 0.0021832 0.42276 1.1561 1.151 16.0005 144.9779 0.0004793 -83.917 0.08795
1.192 0.98803 5.5182e-005 3.8182 0.012034 1.5688e-005 0.0011542 0.15464 0.00065837 0.15529 0.14164 0 0.036703 0.0389 0 0.90352 0.25274 0.068072 0.0094892 4.276 0.059248 7.1226e-005 0.83082 0.0052961 0.0060337 0.0018444 0.98026 0.8865 4.0493e-006 1.6199e-005 0.13204 0.65754 0.71806 0.0016234 0.68647 0.48525 0.0021793 0.42275 1.1583 1.1532 16.0005 144.9779 0.00047775 -83.9368 0.08895
1.193 0.98803 5.5182e-005 3.8182 0.012034 1.5701e-005 0.0011542 0.1547 0.00065837 0.15536 0.1417 0 0.036699 0.0389 0 0.9036 0.25277 0.068084 0.0094907 4.2764 0.059257 7.1238e-005 0.83081 0.0052965 0.0060341 0.0018385 0.98041 0.89227 4.0357e-006 1.6144e-005 0.13205 0.65855 0.7191 0.0016207 0.68816 0.48542 0.0021757 0.42275 1.1605 1.1553 16.0006 144.9779 0.00047621 -83.9557 0.08995
1.194 0.98803 5.5182e-005 3.8182 0.012034 1.5715e-005 0.0011542 0.15477 0.00065837 0.15542 0.14176 0 0.036695 0.0389 0 0.90368 0.25281 0.068097 0.0094922 4.2768 0.059266 7.125e-005 0.8308 0.0052969 0.0060345 0.0018329 0.98054 0.89773 4.0227e-006 1.6093e-005 0.13205 0.65955 0.72013 0.0016181 0.68985 0.48559 0.0021722 0.42275 1.1626 1.1575 16.0007 144.9779 0.00047469 -83.9738 0.09095
1.195 0.98803 5.5182e-005 3.8182 0.012034 1.5728e-005 0.0011542 0.15483 0.00065837 0.15549 0.14182 0 0.036691 0.0389 0 0.90376 0.25284 0.068109 0.0094938 4.2772 0.059276 7.1263e-005 0.8308 0.0052973 0.0060349 0.0018275 0.98065 0.90289 4.0103e-006 1.6043e-005 0.13205 0.66055 0.72115 0.0016156 0.69153 0.48576 0.0021688 0.42274 1.1648 1.1597 16.0008 144.9779 0.00047317 -83.9912 0.09195
1.196 0.98803 5.5182e-005 3.8182 0.012034 1.5741e-005 0.0011542 0.1549 0.00065837 0.15555 0.14189 0 0.036687 0.0389 0 0.90384 0.25288 0.068122 0.0094953 4.2775 0.059285 7.1275e-005 0.83079 0.0052977 0.0060353 0.0018225 0.98076 0.90776 3.9984e-006 1.5995e-005 0.13206 0.66155 0.72217 0.0016133 0.6932 0.48593 0.0021656 0.42274 1.1669 1.1618 16.0009 144.9779 0.00047166 -84.0079 0.09295
1.197 0.98803 5.5182e-005 3.8182 0.012034 1.5754e-005 0.0011542 0.15496 0.00065837 0.15562 0.14195 0 0.036683 0.0389 0 0.90392 0.25291 0.068134 0.0094968 4.2779 0.059295 7.1287e-005 0.83078 0.0052981 0.0060357 0.0018176 0.98086 0.91236 3.9871e-006 1.595e-005 0.13206 0.66255 0.72317 0.001611 0.69487 0.4861 0.0021626 0.42274 1.1691 1.164 16.0009 144.9779 0.00047015 -84.024 0.09395
1.198 0.98803 5.5182e-005 3.8182 0.012034 1.5767e-005 0.0011542 0.15503 0.00065837 0.15568 0.14201 0 0.036679 0.0389 0 0.90399 0.25295 0.068147 0.0094984 4.2783 0.059304 7.1299e-005 0.83077 0.0052984 0.0060361 0.001813 0.98095 0.91671 3.9761e-006 1.5906e-005 0.13206 0.66354 0.72418 0.0016088 0.69654 0.48627 0.0021596 0.42273 1.1712 1.1662 16.001 144.978 0.00046866 -84.0396 0.09495
1.199 0.98803 5.5182e-005 3.8182 0.012034 1.578e-005 0.0011542 0.15509 0.00065838 0.15575 0.14207 0 0.036674 0.0389 0 0.90407 0.25298 0.06816 0.0094999 4.2786 0.059314 7.1311e-005 0.83076 0.0052988 0.0060364 0.0018086 0.98104 0.92082 3.9656e-006 1.5864e-005 0.13207 0.66453 0.72517 0.0016067 0.69819 0.48644 0.0021568 0.42273 1.1733 1.1683 16.0011 144.978 0.00046717 -84.0547 0.09595
1.2 0.98803 5.5182e-005 3.8182 0.012034 1.5793e-005 0.0011542 0.15516 0.00065838 0.15581 0.14213 0 0.03667 0.0389 0 0.90415 0.25302 0.068172 0.0095014 4.279 0.059323 7.1323e-005 0.83075 0.0052992 0.0060368 0.0018043 0.98112 0.9247 3.9553e-006 1.5823e-005 0.13207 0.66552 0.72616 0.0016046 0.69984 0.48661 0.002154 0.42273 1.1755 1.1705 16.0012 144.978 0.00046569 -84.0694 0.09695
1.201 0.98803 5.5182e-005 3.8182 0.012034 1.5806e-005 0.0011542 0.15522 0.00065838 0.15588 0.14219 0 0.036666 0.0389 0 0.90423 0.25305 0.068185 0.009503 4.2794 0.059333 7.1336e-005 0.83074 0.0052996 0.0060372 0.0018001 0.9812 0.92837 3.9454e-006 1.5783e-005 0.13207 0.6665 0.72714 0.0016026 0.70148 0.48678 0.0021513 0.42272 1.1776 1.1726 16.0013 144.978 0.00046422 -84.0836 0.09795
1.202 0.98803 5.5182e-005 3.8182 0.012034 1.582e-005 0.0011542 0.15529 0.00065838 0.15594 0.14225 0 0.036662 0.0389 0 0.90431 0.25309 0.068197 0.0095045 4.2798 0.059342 7.1348e-005 0.83073 0.0053 0.0060376 0.0017958 0.98127 0.93183 3.9356e-006 1.5744e-005 0.13208 0.66748 0.72811 0.0016007 0.70312 0.48695 0.0021487 0.42272 1.1797 1.1747 16.0013 144.978 0.00046276 -84.0975 0.09895
1.203 0.98803 5.5181e-005 3.8182 0.012034 1.5833e-005 0.0011542 0.15535 0.00065838 0.156 0.14231 0 0.036658 0.0389 0 0.90439 0.25312 0.06821 0.0095061 4.2801 0.059352 7.136e-005 0.83072 0.0053004 0.006038 0.0017918 0.98134 0.93509 3.9262e-006 1.5706e-005 0.13208 0.66846 0.72908 0.0015988 0.70475 0.48711 0.0021462 0.42272 1.1818 1.1769 16.0014 144.978 0.0004613 -84.1111 0.09995
1.204 0.98803 5.5181e-005 3.8182 0.012034 1.5846e-005 0.0011542 0.15541 0.00065838 0.15607 0.14237 0 0.036654 0.0389 0 0.90447 0.25316 0.068223 0.0095076 4.2805 0.059361 7.1372e-005 0.83071 0.0053008 0.0060384 0.0017879 0.9814 0.93818 3.917e-006 1.5669e-005 0.13208 0.66943 0.73004 0.0015969 0.70637 0.48728 0.0021438 0.42272 1.1839 1.179 16.0015 144.978 0.00045986 -84.1243 0.10095
1.205 0.98803 5.5181e-005 3.8182 0.012034 1.5859e-005 0.0011542 0.15548 0.00065838 0.15613 0.14243 0 0.03665 0.0389 0 0.90454 0.25319 0.068235 0.0095091 4.2809 0.05937 7.1384e-005 0.8307 0.0053011 0.0060388 0.0017841 0.98147 0.94109 3.9081e-006 1.5634e-005 0.13209 0.6704 0.731 0.0015951 0.70799 0.48745 0.0021414 0.42272 1.1861 1.1811 16.0016 144.978 0.00045842 -84.1373 0.10195
1.206 0.98803 5.5181e-005 3.8182 0.012034 1.5872e-005 0.0011542 0.15554 0.00065838 0.1562 0.14249 0 0.036646 0.0389 0 0.90462 0.25323 0.068248 0.0095107 4.2813 0.05938 7.1397e-005 0.83069 0.0053015 0.0060392 0.0017804 0.98153 0.94383 3.8994e-006 1.5598e-005 0.13209 0.67137 0.73194 0.0015933 0.70959 0.48762 0.002139 0.42272 1.1882 1.1833 16.0016 144.978 0.00045698 -84.15 0.10295
1.207 0.98803 5.5181e-005 3.8182 0.012034 1.5885e-005 0.0011542 0.15561 0.00065838 0.15626 0.14255 0 0.036642 0.0389 0 0.9047 0.25326 0.06826 0.0095122 4.2816 0.059389 7.1409e-005 0.83068 0.0053019 0.0060396 0.0017767 0.98159 0.94643 3.8908e-006 1.5564e-005 0.13209 0.67234 0.73289 0.0015916 0.7112 0.48779 0.0021367 0.42271 1.1903 1.1854 16.0017 144.978 0.00045556 -84.1625 0.10395
1.208 0.98803 5.5181e-005 3.8182 0.012034 1.5898e-005 0.0011542 0.15567 0.00065839 0.15632 0.14261 0 0.036638 0.0389 0 0.90478 0.2533 0.068273 0.0095138 4.282 0.059399 7.1421e-005 0.83067 0.0053023 0.00604 0.001773 0.98164 0.94888 3.8823e-006 1.553e-005 0.1321 0.6733 0.73382 0.0015899 0.71279 0.48796 0.0021345 0.42271 1.1924 1.1875 16.0018 144.978 0.00045414 -84.1747 0.10495
1.209 0.98803 5.5181e-005 3.8182 0.012034 1.5912e-005 0.0011542 0.15573 0.00065839 0.15639 0.14267 0 0.036634 0.0389 0 0.90486 0.25333 0.068286 0.0095153 4.2824 0.059408 7.1433e-005 0.83066 0.0053027 0.0060404 0.0017694 0.9817 0.95119 3.874e-006 1.5497e-005 0.1321 0.67426 0.73475 0.0015882 0.71438 0.48813 0.0021322 0.42271 1.1945 1.1896 16.0019 144.9781 0.00045274 -84.1868 0.10595
1.21 0.98803 5.5181e-005 3.8182 0.012034 1.5925e-005 0.0011542 0.1558 0.00065839 0.15645 0.14273 0 0.03663 0.0389 0 0.90494 0.25337 0.068298 0.0095169 4.2828 0.059418 7.1446e-005 0.83065 0.0053031 0.0060408 0.0017659 0.98175 0.95337 3.8659e-006 1.5465e-005 0.1321 0.67522 0.73568 0.0015865 0.71596 0.4883 0.0021301 0.42271 1.1966 1.1917 16.0019 144.9781 0.00045134 -84.1986 0.10695
1.211 0.98803 5.5181e-005 3.8182 0.012034 1.5938e-005 0.0011542 0.15586 0.00065839 0.15652 0.14279 0 0.036626 0.0389 0 0.90502 0.2534 0.068311 0.0095184 4.2831 0.059427 7.1458e-005 0.83064 0.0053035 0.0060411 0.0017626 0.9818 0.95542 3.8579e-006 1.5433e-005 0.13211 0.67617 0.73659 0.0015849 0.71753 0.48847 0.0021279 0.42271 1.1986 1.1938 16.002 144.9781 0.00044994 -84.2103 0.10795
1.212 0.98803 5.5181e-005 3.8182 0.012034 1.5951e-005 0.0011542 0.15593 0.00065839 0.15658 0.14285 0 0.036622 0.0389 0 0.9051 0.25344 0.068324 0.0095199 4.2835 0.059437 7.147e-005 0.83063 0.0053039 0.0060415 0.0017592 0.98185 0.95736 3.8501e-006 1.5401e-005 0.13211 0.67712 0.7375 0.0015833 0.7191 0.48864 0.0021258 0.42271 1.2007 1.1959 16.0021 144.9781 0.00044856 -84.2218 0.10895
1.213 0.98803 5.5181e-005 3.8182 0.012034 1.5964e-005 0.0011542 0.15599 0.00065839 0.15664 0.14291 0 0.036618 0.0389 0 0.90517 0.25347 0.068336 0.0095215 4.2839 0.059446 7.1482e-005 0.83063 0.0053043 0.0060419 0.0017557 0.9819 0.95919 3.8423e-006 1.537e-005 0.13211 0.67807 0.73841 0.0015817 0.72066 0.48881 0.0021238 0.42271 1.2028 1.198 16.0022 144.9781 0.00044718 -84.2331 0.10995
1.214 0.98803 5.5181e-005 3.8182 0.012034 1.5977e-005 0.0011542 0.15605 0.00065839 0.15671 0.14297 0 0.036614 0.0389 0 0.90525 0.25351 0.068349 0.009523 4.2843 0.059456 7.1494e-005 0.83062 0.0053046 0.0060423 0.0017523 0.98195 0.96092 3.8347e-006 1.534e-005 0.13212 0.67902 0.73931 0.0015802 0.72221 0.48898 0.0021217 0.42271 1.2049 1.2001 16.0022 144.9781 0.00044581 -84.2443 0.11095
1.215 0.98803 5.5181e-005 3.8182 0.012034 1.599e-005 0.0011542 0.15612 0.00065839 0.15677 0.14303 0 0.03661 0.0389 0 0.90533 0.25354 0.068362 0.0095246 4.2846 0.059465 7.1507e-005 0.83061 0.005305 0.0060427 0.0017491 0.982 0.96255 3.8272e-006 1.531e-005 0.13212 0.67996 0.7402 0.0015787 0.72376 0.48915 0.0021197 0.42271 1.2069 1.2022 16.0023 144.9781 0.00044444 -84.2554 0.11195
1.216 0.98803 5.5181e-005 3.8182 0.012034 1.6003e-005 0.0011542 0.15618 0.00065839 0.15684 0.14309 0 0.036606 0.0389 0 0.90541 0.25358 0.068374 0.0095261 4.285 0.059475 7.1519e-005 0.8306 0.0053054 0.0060431 0.0017459 0.98205 0.96409 3.8198e-006 1.528e-005 0.13212 0.6809 0.74109 0.0015772 0.7253 0.48932 0.0021177 0.42271 1.209 1.2043 16.0024 144.9781 0.00044309 -84.2663 0.11295
1.217 0.98803 5.5181e-005 3.8182 0.012034 1.6017e-005 0.0011542 0.15625 0.0006584 0.1569 0.14315 0 0.036602 0.0389 0 0.90549 0.25361 0.068387 0.0095277 4.2854 0.059484 7.1531e-005 0.83059 0.0053058 0.0060435 0.0017429 0.98209 0.96554 3.8125e-006 1.5251e-005 0.13212 0.68184 0.74198 0.0015757 0.72683 0.48949 0.0021158 0.42271 1.2111 1.2064 16.0024 144.9781 0.00044174 -84.2771 0.11395
1.218 0.98803 5.5181e-005 3.8182 0.012034 1.603e-005 0.0011542 0.15631 0.0006584 0.15696 0.14321 0 0.036598 0.0389 0 0.90557 0.25365 0.0684 0.0095292 4.2858 0.059494 7.1544e-005 0.83058 0.0053062 0.0060439 0.0017399 0.98214 0.96691 3.8053e-006 1.5222e-005 0.13213 0.68277 0.74285 0.0015742 0.72835 0.48966 0.0021139 0.42271 1.2131 1.2084 16.0025 144.9781 0.00044039 -84.2878 0.11495
1.219 0.98803 5.518e-005 3.8182 0.012034 1.6043e-005 0.0011542 0.15637 0.0006584 0.15703 0.14327 0 0.036593 0.0389 0 0.90565 0.25368 0.068412 0.0095308 4.2862 0.059504 7.1556e-005 0.83057 0.0053066 0.0060443 0.0017369 0.98218 0.9682 3.7982e-006 1.5194e-005 0.13213 0.6837 0.74372 0.0015728 0.72987 0.48983 0.002112 0.42271 1.2152 1.2105 16.0026 144.9781 0.00043906 -84.2984 0.11595
1.22 0.98803 5.518e-005 3.8182 0.012034 1.6056e-005 0.0011542 0.15644 0.0006584 0.15709 0.14333 0 0.036589 0.0389 0 0.90573 0.25372 0.068425 0.0095323 4.2865 0.059513 7.1568e-005 0.83056 0.005307 0.0060447 0.001734 0.98223 0.96942 3.7912e-006 1.5166e-005 0.13213 0.68463 0.74459 0.0015713 0.73138 0.49 0.0021101 0.42271 1.2172 1.2126 16.0027 144.9782 0.00043773 -84.3088 0.11695
1.221 0.98803 5.518e-005 3.8182 0.012034 1.6069e-005 0.0011542 0.1565 0.0006584 0.15715 0.14338 0 0.036585 0.0389 0 0.90581 0.25375 0.068438 0.0095339 4.2869 0.059523 7.158e-005 0.83055 0.0053074 0.0060451 0.001731 0.98227 0.97057 3.7843e-006 1.5138e-005 0.13214 0.68555 0.74545 0.0015699 0.73289 0.49017 0.0021082 0.42271 1.2193 1.2146 16.0027 144.9782 0.00043641 -84.3192 0.11795
1.222 0.98803 5.518e-005 3.8182 0.012034 1.6082e-005 0.0011542 0.15656 0.0006584 0.15722 0.14344 0 0.036581 0.0389 0 0.90589 0.25379 0.06845 0.0095354 4.2873 0.059532 7.1593e-005 0.83054 0.0053078 0.0060455 0.001728 0.98231 0.97165 3.7774e-006 1.511e-005 0.13214 0.68648 0.74631 0.0015685 0.73438 0.49034 0.0021064 0.42271 1.2213 1.2167 16.0028 144.9782 0.0004351 -84.3294 0.11895
1.223 0.98803 5.518e-005 3.8182 0.012034 1.6095e-005 0.0011542 0.15663 0.0006584 0.15728 0.1435 0 0.036577 0.0389 0 0.90597 0.25382 0.068463 0.009537 4.2877 0.059542 7.1605e-005 0.83053 0.0053082 0.0060459 0.0017249 0.98235 0.97268 3.7706e-006 1.5083e-005 0.13214 0.6874 0.74716 0.0015671 0.73587 0.49051 0.0021045 0.42271 1.2234 1.2188 16.0029 144.9782 0.00043379 -84.3395 0.11995
1.224 0.98803 5.518e-005 3.8182 0.012034 1.6109e-005 0.0011542 0.15669 0.0006584 0.15734 0.14356 0 0.036574 0.0389 0 0.90605 0.25386 0.068476 0.0095385 4.2881 0.059551 7.1617e-005 0.83052 0.0053086 0.0060463 0.001722 0.9824 0.97364 3.7639e-006 1.5056e-005 0.13215 0.68831 0.748 0.0015657 0.73736 0.49068 0.0021027 0.42271 1.2254 1.2208 16.0029 144.9782 0.00043249 -84.3496 0.12095
1.225 0.98803 5.518e-005 3.8182 0.012034 1.6122e-005 0.0011542 0.15675 0.00065841 0.15741 0.14362 0 0.03657 0.0389 0 0.90612 0.25389 0.068489 0.0095401 4.2885 0.059561 7.163e-005 0.83051 0.005309 0.0060467 0.0017191 0.98244 0.97455 3.7573e-006 1.503e-005 0.13215 0.68923 0.74884 0.0015643 0.73883 0.49085 0.002101 0.42271 1.2274 1.2229 16.003 144.9782 0.0004312 -84.3595 0.12195
1.226 0.98803 5.518e-005 3.8182 0.012034 1.6135e-005 0.0011542 0.15682 0.00065841 0.15747 0.14368 0 0.036566 0.0389 0 0.9062 0.25393 0.068501 0.0095416 4.2888 0.05957 7.1642e-005 0.8305 0.0053094 0.0060471 0.0017164 0.98248 0.97541 3.7508e-006 1.5004e-005 0.13215 0.69014 0.74967 0.001563 0.7403 0.49102 0.0020992 0.42271 1.2295 1.2249 16.0031 144.9782 0.00042991 -84.3694 0.12295
1.227 0.98803 5.518e-005 3.8182 0.012034 1.6148e-005 0.0011542 0.15688 0.00065841 0.15753 0.14374 0 0.036562 0.0389 0 0.90628 0.25396 0.068514 0.0095432 4.2892 0.05958 7.1654e-005 0.83049 0.0053098 0.0060475 0.0017137 0.98252 0.97622 3.7443e-006 1.4978e-005 0.13216 0.69105 0.7505 0.0015617 0.74177 0.49119 0.0020974 0.42271 1.2315 1.2269 16.0031 144.9782 0.00042863 -84.3791 0.12395
1.228 0.98803 5.518e-005 3.8182 0.012034 1.6161e-005 0.0011542 0.15694 0.00065841 0.1576 0.1438 0 0.036558 0.0389 0 0.90636 0.254 0.068527 0.0095447 4.2896 0.059589 7.1666e-005 0.83048 0.0053102 0.0060479 0.001711 0.98256 0.97698 3.7379e-006 1.4952e-005 0.13216 0.69195 0.75132 0.0015603 0.74322 0.49136 0.0020957 0.42271 1.2335 1.229 16.0032 144.9782 0.00042736 -84.3888 0.12495
1.229 0.98803 5.518e-005 3.8182 0.012034 1.6174e-005 0.0011542 0.157 0.00065841 0.15766 0.14386 0 0.036554 0.0389 0 0.90644 0.25403 0.06854 0.0095463 4.29 0.059599 7.1679e-005 0.83047 0.0053105 0.0060483 0.0017083 0.98259 0.9777 3.7316e-006 1.4927e-005 0.13216 0.69286 0.75214 0.001559 0.74467 0.49153 0.002094 0.42271 1.2355 1.231 16.0033 144.9783 0.00042609 -84.3984 0.12595
1.23 0.98803 5.518e-005 3.8182 0.012034 1.6187e-005 0.0011542 0.15707 0.00065841 0.15772 0.14392 0 0.03655 0.0389 0 0.90652 0.25407 0.068552 0.0095478 4.2904 0.059609 7.1691e-005 0.83046 0.0053109 0.0060487 0.0017055 0.98263 0.97838 3.7253e-006 1.4902e-005 0.13217 0.69376 0.75296 0.0015577 0.74611 0.4917 0.0020923 0.42271 1.2375 1.233 16.0033 144.9783 0.00042483 -84.4079 0.12695
1.231 0.98803 5.518e-005 3.8182 0.012034 1.62e-005 0.0011542 0.15713 0.00065841 0.15778 0.14398 0 0.036546 0.0389 0 0.9066 0.2541 0.068565 0.0095494 4.2908 0.059618 7.1703e-005 0.83045 0.0053113 0.0060491 0.0017028 0.98267 0.97903 3.7191e-006 1.4877e-005 0.13217 0.69466 0.75377 0.0015565 0.74755 0.49187 0.0020906 0.42272 1.2395 1.235 16.0034 144.9783 0.00042358 -84.4173 0.12795
1.232 0.98803 5.518e-005 3.8182 0.012034 1.6214e-005 0.0011542 0.15719 0.00065841 0.15785 0.14404 0 0.036542 0.0389 0 0.90668 0.25414 0.068578 0.0095509 4.2912 0.059628 7.1716e-005 0.83044 0.0053117 0.0060495 0.0017002 0.98271 0.97963 3.7129e-006 1.4852e-005 0.13217 0.69555 0.75457 0.0015552 0.74898 0.49204 0.002089 0.42272 1.2415 1.2371 16.0035 144.9783 0.00042234 -84.4267 0.12895
1.233 0.98803 5.518e-005 3.8182 0.012034 1.6227e-005 0.0011542 0.15726 0.00065841 0.15791 0.14409 0 0.036538 0.0389 0 0.90676 0.25417 0.068591 0.0095525 4.2915 0.059637 7.1728e-005 0.83043 0.0053121 0.0060499 0.0016976 0.98275 0.9802 3.7069e-006 1.4828e-005 0.13218 0.69644 0.75537 0.0015539 0.7504 0.49221 0.0020873 0.42272 1.2435 1.2391 16.0035 144.9783 0.0004211 -84.4359 0.12995
1.234 0.98803 5.518e-005 3.8182 0.012034 1.624e-005 0.0011542 0.15732 0.00065841 0.15797 0.14415 0 0.036534 0.0389 0 0.90684 0.25421 0.068603 0.009554 4.2919 0.059647 7.174e-005 0.83042 0.0053125 0.0060503 0.001695 0.98278 0.98074 3.7009e-006 1.4804e-005 0.13218 0.69733 0.75616 0.0015527 0.75181 0.49238 0.0020857 0.42272 1.2455 1.2411 16.0036 144.9783 0.00041986 -84.4451 0.13095
1.235 0.98803 5.5179e-005 3.8182 0.012034 1.6253e-005 0.0011542 0.15738 0.00065842 0.15804 0.14421 0 0.03653 0.0389 0 0.90692 0.25425 0.068616 0.0095556 4.2923 0.059656 7.1753e-005 0.83042 0.0053129 0.0060507 0.0016924 0.98282 0.98125 3.6949e-006 1.478e-005 0.13218 0.69822 0.75695 0.0015514 0.75322 0.49255 0.0020841 0.42272 1.2475 1.2431 16.0036 144.9783 0.00041864 -84.4542 0.13195
1.236 0.98803 5.5179e-005 3.8182 0.012034 1.6266e-005 0.0011542 0.15744 0.00065842 0.1581 0.14427 0 0.036526 0.0389 0 0.907 0.25428 0.068629 0.0095571 4.2927 0.059666 7.1765e-005 0.83041 0.0053133 0.0060511 0.0016899 0.98285 0.98173 3.689e-006 1.4757e-005 0.13219 0.6991 0.75773 0.0015502 0.75462 0.49272 0.0020825 0.42272 1.2495 1.2451 16.0037 144.9783 0.00041742 -84.4632 0.13295
1.237 0.98803 5.5179e-005 3.8182 0.012034 1.6279e-005 0.0011542 0.15751 0.00065842 0.15816 0.14433 0 0.036522 0.0389 0 0.90708 0.25432 0.068642 0.0095587 4.2931 0.059676 7.1778e-005 0.8304 0.0053137 0.0060515 0.0016873 0.98289 0.98218 3.6831e-006 1.4733e-005 0.13219 0.69998 0.75851 0.001549 0.75602 0.49289 0.0020809 0.42273 1.2515 1.2471 16.0038 144.9783 0.0004162 -84.4722 0.13395
1.238 0.98803 5.5179e-005 3.8182 0.012033 1.6292e-005 0.0011542 0.15757 0.00065842 0.15822 0.14439 0 0.036518 0.0389 0 0.90716 0.25435 0.068654 0.0095603 4.2935 0.059685 7.179e-005 0.83039 0.0053141 0.0060519 0.0016849 0.98292 0.98261 3.6774e-006 1.471e-005 0.13219 0.70086 0.75929 0.0015478 0.7574 0.49306 0.0020793 0.42273 1.2534 1.2491 16.0038 144.9784 0.000415 -84.4811 0.13495
1.239 0.98803 5.5179e-005 3.8182 0.012033 1.6306e-005 0.0011542 0.15763 0.00065842 0.15829 0.14445 0 0.036514 0.0389 0 0.90724 0.25439 0.068667 0.0095618 4.2939 0.059695 7.1802e-005 0.83038 0.0053145 0.0060523 0.0016824 0.98296 0.98302 3.6716e-006 1.4687e-005 0.1322 0.70174 0.76006 0.0015466 0.75878 0.49323 0.0020777 0.42273 1.2554 1.2511 16.0039 144.9784 0.00041379 -84.4899 0.13595
1.24 0.98803 5.5179e-005 3.8182 0.012033 1.6319e-005 0.0011542 0.15769 0.00065842 0.15835 0.14451 0 0.03651 0.0389 0 0.90732 0.25442 0.06868 0.0095634 4.2943 0.059704 7.1815e-005 0.83037 0.0053149 0.0060527 0.00168 0.98299 0.9834 3.666e-006 1.4664e-005 0.1322 0.70261 0.76082 0.0015454 0.76016 0.4934 0.0020762 0.42273 1.2574 1.253 16.004 144.9784 0.0004126 -84.4986 0.13695
1.241 0.98803 5.5179e-005 3.8182 0.012033 1.6332e-005 0.0011542 0.15776 0.00065842 0.15841 0.14456 0 0.036506 0.0389 0 0.9074 0.25446 0.068693 0.0095649 4.2947 0.059714 7.1827e-005 0.83036 0.0053153 0.0060531 0.0016775 0.98303 0.98376 3.6603e-006 1.4642e-005 0.1322 0.70348 0.76158 0.0015443 0.76153 0.49357 0.0020747 0.42273 1.2594 1.255 16.004 144.9784 0.00041141 -84.5073 0.13795
1.242 0.98803 5.5179e-005 3.8182 0.012033 1.6345e-005 0.0011542 0.15782 0.00065842 0.15847 0.14462 0 0.036502 0.0389 0 0.90748 0.25449 0.068705 0.0095665 4.295 0.059724 7.1839e-005 0.83035 0.0053157 0.0060536 0.0016751 0.98306 0.9841 3.6548e-006 1.462e-005 0.13221 0.70435 0.76234 0.0015431 0.76289 0.49374 0.0020731 0.42274 1.2613 1.257 16.0041 144.9784 0.00041023 -84.5159 0.13895
1.243 0.98803 5.5179e-005 3.8182 0.012033 1.6358e-005 0.0011542 0.15788 0.00065842 0.15854 0.14468 0 0.036498 0.0389 0 0.90756 0.25453 0.068718 0.009568 4.2954 0.059733 7.1852e-005 0.83034 0.0053161 0.006054 0.0016728 0.98309 0.98442 3.6493e-006 1.4598e-005 0.13221 0.70522 0.76309 0.0015419 0.76424 0.49391 0.0020716 0.42274 1.2633 1.259 16.0041 144.9784 0.00040905 -84.5244 0.13995
1.244 0.98803 5.5179e-005 3.8182 0.012033 1.6371e-005 0.0011542 0.15794 0.00065843 0.1586 0.14474 0 0.036495 0.0389 0 0.90764 0.25456 0.068731 0.0095696 4.2958 0.059743 7.1864e-005 0.83033 0.0053165 0.0060544 0.0016704 0.98313 0.98472 3.6438e-006 1.4576e-005 0.13221 0.70608 0.76384 0.0015408 0.76559 0.49408 0.0020701 0.42274 1.2652 1.2609 16.0042 144.9784 0.00040788 -84.5329 0.14095
1.245 0.98803 5.5179e-005 3.8182 0.012033 1.6384e-005 0.0011542 0.15801 0.00065843 0.15866 0.1448 0 0.036491 0.0389 0 0.90772 0.2546 0.068744 0.0095712 4.2962 0.059752 7.1877e-005 0.83032 0.0053169 0.0060548 0.0016681 0.98316 0.98501 3.6384e-006 1.4554e-005 0.13222 0.70694 0.76458 0.0015397 0.76693 0.49425 0.0020687 0.42275 1.2672 1.2629 16.0043 144.9784 0.00040672 -84.5413 0.14195
1.246 0.98803 5.5179e-005 3.8182 0.012033 1.6397e-005 0.0011542 0.15807 0.00065843 0.15872 0.14486 0 0.036487 0.0389 0 0.9078 0.25464 0.068757 0.0095727 4.2966 0.059762 7.1889e-005 0.83031 0.0053173 0.0060552 0.0016658 0.98319 0.98528 3.633e-006 1.4533e-005 0.13222 0.7078 0.76532 0.0015385 0.76826 0.49442 0.0020672 0.42275 1.2691 1.2649 16.0043 144.9784 0.00040556 -84.5496 0.14295
1.247 0.98803 5.5179e-005 3.8182 0.012033 1.6411e-005 0.0011542 0.15813 0.00065843 0.15878 0.14491 0 0.036483 0.0389 0 0.90788 0.25467 0.068769 0.0095743 4.297 0.059772 7.1901e-005 0.8303 0.0053177 0.0060556 0.0016635 0.98322 0.98553 3.6277e-006 1.4512e-005 0.13222 0.70865 0.76606 0.0015374 0.76959 0.49459 0.0020658 0.42275 1.271 1.2668 16.0044 144.9785 0.00040441 -84.5579 0.14395
1.248 0.98803 5.5179e-005 3.8182 0.012033 1.6424e-005 0.0011542 0.15819 0.00065843 0.15885 0.14497 0 0.036479 0.0389 0 0.90795 0.25471 0.068782 0.0095758 4.2974 0.059781 7.1914e-005 0.83029 0.0053181 0.006056 0.0016612 0.98326 0.98578 3.6225e-006 1.4491e-005 0.13223 0.7095 0.76679 0.0015363 0.77091 0.49476 0.0020643 0.42275 1.273 1.2688 16.0044 144.9785 0.00040326 -84.566 0.14495
1.249 0.98803 5.5179e-005 3.8182 0.012033 1.6437e-005 0.0011542 0.15825 0.00065843 0.15891 0.14503 0 0.036475 0.0389 0 0.90803 0.25474 0.068795 0.0095774 4.2978 0.059791 7.1926e-005 0.83028 0.0053185 0.0060564 0.001659 0.98329 0.986 3.6173e-006 1.447e-005 0.13223 0.71035 0.76751 0.0015352 0.77223 0.49493 0.0020629 0.42276 1.2749 1.2707 16.0045 144.9785 0.00040212 -84.5742 0.14595
1.25 0.98803 5.5179e-005 3.8182 0.012033 1.645e-005 0.0011542 0.15832 0.00065843 0.15897 0.14509 0 0.036471 0.0389 0 0.90811 0.25478 0.068808 0.009579 4.2982 0.0598 7.1939e-005 0.83027 0.005319 0.0060568 0.0016568 0.98332 0.98622 3.6121e-006 1.4449e-005 0.13223 0.7112 0.76823 0.0015342 0.77354 0.4951 0.0020615 0.42276 1.2768 1.2726 16.0045 144.9785 0.00040099 -84.5822 0.14695
1.251 0.98803 5.5178e-005 3.8182 0.012033 1.6463e-005 0.0011542 0.15838 0.00065843 0.15903 0.14515 0 0.036467 0.0389 0 0.90819 0.25481 0.068821 0.0095805 4.2986 0.05981 7.1951e-005 0.83026 0.0053194 0.0060572 0.0016546 0.98335 0.98642 3.607e-006 1.4429e-005 0.13224 0.71204 0.76895 0.0015331 0.77484 0.49527 0.0020601 0.42276 1.2788 1.2746 16.0046 144.9785 0.00039986 -84.5902 0.14795
1.252 0.98803 5.5178e-005 3.8182 0.012033 1.6476e-005 0.0011542 0.15844 0.00065843 0.15909 0.1452 0 0.036463 0.0389 0 0.90827 0.25485 0.068834 0.0095821 4.299 0.05982 7.1963e-005 0.83025 0.0053198 0.0060576 0.0016524 0.98338 0.98662 3.6019e-006 1.4408e-005 0.13224 0.71289 0.76967 0.001532 0.77613 0.49543 0.0020587 0.42277 1.2807 1.2765 16.0047 144.9785 0.00039874 -84.5982 0.14895
1.253 0.98803 5.5178e-005 3.8182 0.012033 1.6489e-005 0.0011542 0.1585 0.00065844 0.15916 0.14526 0 0.03646 0.0389 0 0.90835 0.25488 0.068846 0.0095837 4.2994 0.059829 7.1976e-005 0.83024 0.0053202 0.006058 0.0016502 0.98341 0.9868 3.5969e-006 1.4388e-005 0.13224 0.71372 0.77037 0.001531 0.77742 0.4956 0.0020573 0.42277 1.2826 1.2784 16.0047 144.9785 0.00039762 -84.606 0.14995
1.254 0.98803 5.5178e-005 3.8182 0.012033 1.6503e-005 0.0011542 0.15856 0.00065844 0.15922 0.14532 0 0.036456 0.0389 0 0.90843 0.25492 0.068859 0.0095852 4.2998 0.059839 7.1988e-005 0.83023 0.0053206 0.0060585 0.0016481 0.98344 0.98697 3.592e-006 1.4368e-005 0.13225 0.71456 0.77108 0.0015299 0.7787 0.49577 0.0020559 0.42277 1.2845 1.2804 16.0048 144.9785 0.00039651 -84.6139 0.15095
1.255 0.98803 5.5178e-005 3.8182 0.012033 1.6516e-005 0.0011542 0.15863 0.00065844 0.15928 0.14538 0 0.036452 0.0389 0 0.90851 0.25496 0.068872 0.0095868 4.3002 0.059849 7.2001e-005 0.83022 0.005321 0.0060589 0.0016459 0.98347 0.98714 3.587e-006 1.4349e-005 0.13225 0.7154 0.77178 0.0015289 0.77998 0.49594 0.0020546 0.42278 1.2864 1.2823 16.0048 144.9786 0.0003954 -84.6216 0.15195
1.256 0.98803 5.5178e-005 3.8182 0.012033 1.6529e-005 0.0011542 0.15869 0.00065844 0.15934 0.14544 0 0.036448 0.0389 0 0.9086 0.25499 0.068885 0.0095883 4.3006 0.059858 7.2013e-005 0.83021 0.0053214 0.0060593 0.0016438 0.9835 0.98729 3.5822e-006 1.4329e-005 0.13225 0.71623 0.77248 0.0015279 0.78125 0.49611 0.0020532 0.42278 1.2883 1.2842 16.0049 144.9786 0.0003943 -84.6293 0.15295
1.257 0.98803 5.5178e-005 3.8182 0.012033 1.6542e-005 0.0011542 0.15875 0.00065844 0.1594 0.14549 0 0.036444 0.0389 0 0.90868 0.25503 0.068898 0.0095899 4.301 0.059868 7.2026e-005 0.8302 0.0053218 0.0060597 0.0016418 0.98353 0.98744 3.5773e-006 1.431e-005 0.13226 0.71706 0.77317 0.0015268 0.78251 0.49628 0.0020519 0.42279 1.2902 1.2861 16.0049 144.9786 0.00039321 -84.6369 0.15395
1.258 0.98803 5.5178e-005 3.8182 0.012033 1.6555e-005 0.0011542 0.15881 0.00065844 0.15946 0.14555 0 0.03644 0.0389 0 0.90876 0.25506 0.068911 0.0095915 4.3014 0.059878 7.2038e-005 0.83019 0.0053222 0.0060601 0.0016397 0.98356 0.98758 3.5725e-006 1.4291e-005 0.13226 0.71788 0.77386 0.0015258 0.78377 0.49645 0.0020506 0.42279 1.2921 1.288 16.005 144.9786 0.00039212 -84.6445 0.15495
1.259 0.98803 5.5178e-005 3.8182 0.012033 1.6568e-005 0.0011542 0.15887 0.00065844 0.15953 0.14561 0 0.036436 0.0389 0 0.90884 0.2551 0.068924 0.009593 4.3018 0.059887 7.205e-005 0.83018 0.0053226 0.0060605 0.0016376 0.98358 0.98771 3.5678e-006 1.4272e-005 0.13226 0.71871 0.77454 0.0015248 0.78502 0.49662 0.0020493 0.42279 1.294 1.2899 16.005 144.9786 0.00039104 -84.652 0.15595
1.26 0.98803 5.5178e-005 3.8182 0.012033 1.6581e-005 0.0011542 0.15893 0.00065844 0.15959 0.14567 0 0.036433 0.0389 0 0.90892 0.25513 0.068936 0.0095946 4.3022 0.059897 7.2063e-005 0.83018 0.005323 0.0060609 0.0016356 0.98361 0.98783 3.5631e-006 1.4253e-005 0.13227 0.71953 0.77523 0.0015238 0.78626 0.49679 0.002048 0.4228 1.2959 1.2918 16.0051 144.9786 0.00038996 -84.6595 0.15695
1.261 0.98803 5.5178e-005 3.8182 0.012033 1.6594e-005 0.0011542 0.15899 0.00065844 0.15965 0.14572 0 0.036429 0.0389 0 0.909 0.25517 0.068949 0.0095962 4.3026 0.059907 7.2075e-005 0.83017 0.0053234 0.0060613 0.0016336 0.98364 0.98795 3.5584e-006 1.4234e-005 0.13227 0.72035 0.7759 0.0015228 0.7875 0.49696 0.0020467 0.4228 1.2977 1.2937 16.0051 144.9786 0.00038889 -84.6668 0.15795
1.262 0.98803 5.5178e-005 3.8182 0.012033 1.6608e-005 0.0011542 0.15906 0.00065844 0.15971 0.14578 0 0.036425 0.0389 0 0.90908 0.25521 0.068962 0.0095977 4.303 0.059916 7.2088e-005 0.83016 0.0053238 0.0060617 0.0016316 0.98367 0.98806 3.5538e-006 1.4216e-005 0.13227 0.72116 0.77658 0.0015219 0.78873 0.49713 0.0020454 0.42281 1.2996 1.2956 16.0052 144.9786 0.00038782 -84.6742 0.15895
1.263 0.98803 5.5178e-005 3.8182 0.012033 1.6621e-005 0.0011542 0.15912 0.00065845 0.15977 0.14584 0 0.036421 0.0389 0 0.90916 0.25524 0.068975 0.0095993 4.3034 0.059926 7.21e-005 0.83015 0.0053242 0.0060622 0.0016296 0.98369 0.98817 3.5492e-006 1.4197e-005 0.13228 0.72198 0.77725 0.0015209 0.78995 0.4973 0.0020441 0.42281 1.3015 1.2975 16.0052 144.9787 0.00038676 -84.6815 0.15995
1.264 0.98803 5.5178e-005 3.8182 0.012033 1.6634e-005 0.0011542 0.15918 0.00065845 0.15983 0.1459 0 0.036417 0.0389 0 0.90924 0.25528 0.068988 0.0096009 4.3038 0.059936 7.2113e-005 0.83014 0.0053246 0.0060626 0.0016277 0.98372 0.98827 3.5447e-006 1.4179e-005 0.13228 0.72279 0.77791 0.0015199 0.79117 0.49747 0.0020429 0.42281 1.3034 1.2994 16.0053 144.9787 0.0003857 -84.6887 0.16095
1.265 0.98803 5.5178e-005 3.8182 0.012033 1.6647e-005 0.0011542 0.15924 0.00065845 0.15989 0.14595 0 0.036413 0.0389 0 0.90932 0.25531 0.069001 0.0096024 4.3042 0.059945 7.2125e-005 0.83013 0.0053251 0.006063 0.0016257 0.98375 0.98836 3.5402e-006 1.4161e-005 0.13228 0.7236 0.77858 0.001519 0.79238 0.49764 0.0020416 0.42282 1.3052 1.3012 16.0053 144.9787 0.00038465 -84.6959 0.16195
1.266 0.98803 5.5178e-005 3.8182 0.012033 1.666e-005 0.0011542 0.1593 0.00065845 0.15996 0.14601 0 0.03641 0.0389 0 0.9094 0.25535 0.069014 0.009604 4.3046 0.059955 7.2138e-005 0.83012 0.0053255 0.0060634 0.0016238 0.98377 0.98845 3.5358e-006 1.4144e-005 0.13229 0.7244 0.77923 0.001518 0.79359 0.49781 0.0020404 0.42282 1.3071 1.3031 16.0054 144.9787 0.00038361 -84.703 0.16295
1.267 0.98803 5.5177e-005 3.8182 0.012033 1.6673e-005 0.0011542 0.15936 0.00065845 0.16002 0.14607 0 0.036406 0.0389 0 0.90948 0.25538 0.069027 0.0096056 4.305 0.059965 7.215e-005 0.83011 0.0053259 0.0060638 0.0016219 0.9838 0.98854 3.5314e-006 1.4126e-005 0.13229 0.72521 0.77989 0.0015171 0.79479 0.49798 0.0020392 0.42283 1.3089 1.305 16.0054 144.9787 0.00038257 -84.71 0.16395
1.268 0.98803 5.5177e-005 3.8182 0.012033 1.6686e-005 0.0011542 0.15942 0.00065845 0.16008 0.14613 0 0.036402 0.0389 0 0.90956 0.25542 0.06904 0.0096072 4.3054 0.059974 7.2163e-005 0.8301 0.0053263 0.0060642 0.00162 0.98383 0.98862 3.527e-006 1.4108e-005 0.13229 0.72601 0.78054 0.0015162 0.79598 0.49815 0.0020379 0.42283 1.3108 1.3068 16.0055 144.9787 0.00038153 -84.717 0.16495
1.269 0.98803 5.5177e-005 3.8182 0.012033 1.67e-005 0.0011542 0.15948 0.00065845 0.16014 0.14618 0 0.036398 0.0389 0 0.90964 0.25546 0.069053 0.0096087 4.3058 0.059984 7.2175e-005 0.83009 0.0053267 0.0060647 0.0016181 0.98385 0.9887 3.5226e-006 1.4091e-005 0.1323 0.72681 0.78119 0.0015153 0.79717 0.49832 0.0020367 0.42284 1.3126 1.3087 16.0055 144.9787 0.00038051 -84.724 0.16595
1.27 0.98803 5.5177e-005 3.8182 0.012033 1.6713e-005 0.0011542 0.15955 0.00065845 0.1602 0.14624 0 0.036394 0.0389 0 0.90972 0.25549 0.069065 0.0096103 4.3062 0.059994 7.2188e-005 0.83008 0.0053271 0.0060651 0.0016163 0.98388 0.98878 3.5184e-006 1.4074e-005 0.1323 0.7276 0.78183 0.0015143 0.79835 0.49849 0.0020356 0.42284 1.3145 1.3106 16.0056 144.9787 0.00037948 -84.7309 0.16695
1.271 0.98803 5.5177e-005 3.8182 0.012033 1.6726e-005 0.0011542 0.15961 0.00065845 0.16026 0.1463 0 0.03639 0.0389 0 0.9098 0.25553 0.069078 0.0096119 4.3066 0.060003 7.22e-005 0.83007 0.0053275 0.0060655 0.0016144 0.9839 0.98885 3.5141e-006 1.4057e-005 0.1323 0.7284 0.78247 0.0015134 0.79953 0.49866 0.0020344 0.42285 1.3163 1.3124 16.0056 144.9788 0.00037846 -84.7377 0.16795
1.272 0.98803 5.5177e-005 3.8182 0.012033 1.6739e-005 0.0011542 0.15967 0.00065846 0.16032 0.14635 0 0.036387 0.0389 0 0.90988 0.25556 0.069091 0.0096134 4.307 0.060013 7.2213e-005 0.83006 0.0053279 0.0060659 0.0016126 0.98393 0.98891 3.5099e-006 1.404e-005 0.13231 0.72919 0.78311 0.0015125 0.80069 0.49882 0.0020332 0.42285 1.3181 1.3143 16.0057 144.9788 0.00037745 -84.7445 0.16895
1.273 0.98803 5.5177e-005 3.8182 0.012033 1.6752e-005 0.0011542 0.15973 0.00065846 0.16038 0.14641 0 0.036383 0.0389 0 0.90996 0.2556 0.069104 0.009615 4.3074 0.060023 7.2225e-005 0.83005 0.0053283 0.0060663 0.0016108 0.98395 0.98898 3.5057e-006 1.4023e-005 0.13231 0.72998 0.78374 0.0015116 0.80186 0.49899 0.002032 0.42286 1.32 1.3161 16.0057 144.9788 0.00037644 -84.7512 0.16995
1.274 0.98803 5.5177e-005 3.8182 0.012033 1.6765e-005 0.0011542 0.15979 0.00065846 0.16044 0.14647 0 0.036379 0.0389 0 0.91004 0.25563 0.069117 0.0096166 4.3078 0.060032 7.2238e-005 0.83004 0.0053288 0.0060667 0.001609 0.98398 0.98904 3.5016e-006 1.4007e-005 0.13232 0.73077 0.78438 0.0015108 0.80301 0.49916 0.0020309 0.42286 1.3218 1.3179 16.0058 144.9788 0.00037544 -84.7579 0.17095
1.275 0.98803 5.5177e-005 3.8182 0.012033 1.6778e-005 0.0011542 0.15985 0.00065846 0.1605 0.14652 0 0.036375 0.0389 0 0.91012 0.25567 0.06913 0.0096182 4.3082 0.060042 7.225e-005 0.83003 0.0053292 0.0060672 0.0016073 0.984 0.9891 3.4974e-006 1.399e-005 0.13232 0.73155 0.785 0.0015099 0.80416 0.49933 0.0020297 0.42287 1.3236 1.3198 16.0058 144.9788 0.00037444 -84.7645 0.17195
1.276 0.98803 5.5177e-005 3.8182 0.012033 1.6791e-005 0.0011542 0.15991 0.00065846 0.16056 0.14658 0 0.036372 0.0389 0 0.9102 0.25571 0.069143 0.0096197 4.3086 0.060052 7.2263e-005 0.83002 0.0053296 0.0060676 0.0016055 0.98403 0.98915 3.4934e-006 1.3974e-005 0.13232 0.73233 0.78563 0.001509 0.80531 0.4995 0.0020286 0.42287 1.3254 1.3216 16.0059 144.9788 0.00037344 -84.7711 0.17295
1.277 0.98803 5.5177e-005 3.8182 0.012033 1.6805e-005 0.0011542 0.15997 0.00065846 0.16062 0.14664 0 0.036368 0.0389 0 0.91028 0.25574 0.069156 0.0096213 4.309 0.060062 7.2275e-005 0.83001 0.00533 0.006068 0.0016037 0.98405 0.98921 3.4893e-006 1.3958e-005 0.13233 0.73311 0.78625 0.0015082 0.80645 0.49967 0.0020275 0.42288 1.3272 1.3234 16.0059 144.9788 0.00037246 -84.7776 0.17395
1.278 0.98803 5.5177e-005 3.8182 0.012033 1.6818e-005 0.0011542 0.16003 0.00065846 0.16069 0.1467 0 0.036364 0.0389 0 0.91036 0.25578 0.069169 0.0096229 4.3094 0.060071 7.2288e-005 0.83 0.0053304 0.0060684 0.001602 0.98407 0.98926 3.4853e-006 1.3942e-005 0.13233 0.73389 0.78686 0.0015073 0.80758 0.49984 0.0020263 0.42288 1.329 1.3253 16.006 144.9789 0.00037147 -84.7841 0.17495
1.279 0.98803 5.5177e-005 3.8182 0.012033 1.6831e-005 0.0011542 0.16009 0.00065846 0.16075 0.14675 0 0.03636 0.0389 0 0.91044 0.25581 0.069182 0.0096245 4.3098 0.060081 7.23e-005 0.82999 0.0053308 0.0060688 0.0016003 0.9841 0.9893 3.4814e-006 1.3926e-005 0.13233 0.73466 0.78748 0.0015064 0.80871 0.50001 0.0020252 0.42289 1.3308 1.3271 16.006 144.9789 0.00037049 -84.7906 0.17595
1.28 0.98803 5.5177e-005 3.8182 0.012033 1.6844e-005 0.0011542 0.16015 0.00065846 0.16081 0.14681 0 0.036356 0.0389 0 0.91053 0.25585 0.069195 0.009626 4.3102 0.060091 7.2313e-005 0.82998 0.0053312 0.0060693 0.0015986 0.98412 0.98935 3.4775e-006 1.391e-005 0.13234 0.73544 0.78809 0.0015056 0.80983 0.50018 0.0020241 0.4229 1.3326 1.3289 16.0061 144.9789 0.00036952 -84.7969 0.17695
1.281 0.98803 5.5177e-005 3.8182 0.012033 1.6857e-005 0.0011542 0.16021 0.00065846 0.16087 0.14687 0 0.036353 0.0389 0 0.91061 0.25589 0.069208 0.0096276 4.3107 0.060101 7.2326e-005 0.82997 0.0053316 0.0060697 0.0015969 0.98414 0.9894 3.4736e-006 1.3895e-005 0.13234 0.73621 0.78869 0.0015048 0.81094 0.50035 0.002023 0.4229 1.3344 1.3307 16.0061 144.9789 0.00036855 -84.8033 0.17795
1.282 0.98803 5.5177e-005 3.8182 0.012033 1.687e-005 0.0011542 0.16027 0.00065847 0.16093 0.14692 0 0.036349 0.0389 0 0.91069 0.25592 0.069221 0.0096292 4.3111 0.06011 7.2338e-005 0.82996 0.0053321 0.0060701 0.0015953 0.98417 0.98944 3.4697e-006 1.3879e-005 0.13234 0.73697 0.7893 0.0015039 0.81205 0.50052 0.002022 0.42291 1.3362 1.3325 16.0062 144.9789 0.00036759 -84.8095 0.17895
1.283 0.98803 5.5176e-005 3.8182 0.012033 1.6883e-005 0.0011542 0.16033 0.00065847 0.16099 0.14698 0 0.036345 0.0389 0 0.91077 0.25596 0.069234 0.0096308 4.3115 0.06012 7.2351e-005 0.82995 0.0053325 0.0060705 0.0015936 0.98419 0.98948 3.4659e-006 1.3864e-005 0.13235 0.73774 0.7899 0.0015031 0.81315 0.50069 0.0020209 0.42291 1.338 1.3343 16.0062 144.9789 0.00036663 -84.8158 0.17995
1.284 0.98803 5.5176e-005 3.8182 0.012033 1.6896e-005 0.0011542 0.16039 0.00065847 0.16105 0.14704 0 0.036341 0.0389 0 0.91085 0.25599 0.069247 0.0096323 4.3119 0.06013 7.2363e-005 0.82994 0.0053329 0.0060709 0.001592 0.98421 0.98952 3.4621e-006 1.3849e-005 0.13235 0.7385 0.79049 0.0015023 0.81425 0.50085 0.0020198 0.42292 1.3398 1.3361 16.0062 144.9789 0.00036568 -84.822 0.18095
1.285 0.98803 5.5176e-005 3.8182 0.012033 1.691e-005 0.0011542 0.16045 0.00065847 0.16111 0.14709 0 0.036338 0.0389 0 0.91093 0.25603 0.06926 0.0096339 4.3123 0.060139 7.2376e-005 0.82993 0.0053333 0.0060714 0.0015903 0.98423 0.98955 3.4583e-006 1.3834e-005 0.13235 0.73926 0.79109 0.0015015 0.81534 0.50102 0.0020188 0.42293 1.3416 1.3379 16.0063 144.979 0.00036473 -84.8281 0.18195
1.286 0.98803 5.5176e-005 3.8182 0.012033 1.6923e-005 0.0011542 0.16051 0.00065847 0.16117 0.14715 0 0.036334 0.0389 0 0.91101 0.25607 0.069273 0.0096355 4.3127 0.060149 7.2388e-005 0.82992 0.0053337 0.0060718 0.0015887 0.98426 0.98959 3.4546e-006 1.3819e-005 0.13236 0.74002 0.79168 0.0015007 0.81643 0.50119 0.0020177 0.42293 1.3433 1.3397 16.0063 144.979 0.00036378 -84.8342 0.18295
1.287 0.98803 5.5176e-005 3.8182 0.012033 1.6936e-005 0.0011542 0.16057 0.00065847 0.16123 0.1472 0 0.03633 0.0389 0 0.91109 0.2561 0.069286 0.0096371 4.3131 0.060159 7.2401e-005 0.82991 0.0053341 0.0060722 0.0015871 0.98428 0.98963 3.4509e-006 1.3804e-005 0.13236 0.74078 0.79227 0.0014999 0.81751 0.50136 0.0020167 0.42294 1.3451 1.3414 16.0064 144.979 0.00036284 -84.8402 0.18395
1.288 0.98803 5.5176e-005 3.8182 0.012033 1.6949e-005 0.0011542 0.16063 0.00065847 0.16129 0.14726 0 0.036326 0.0389 0 0.91117 0.25614 0.069299 0.0096387 4.3135 0.060169 7.2414e-005 0.8299 0.0053346 0.0060726 0.0015855 0.9843 0.98966 3.4472e-006 1.3789e-005 0.13236 0.74153 0.79285 0.0014991 0.81858 0.50153 0.0020157 0.42294 1.3469 1.3432 16.0064 144.979 0.00036191 -84.8462 0.18495
1.289 0.98803 5.5176e-005 3.8182 0.012033 1.6962e-005 0.0011542 0.16069 0.00065847 0.16135 0.14732 0 0.036323 0.0389 0 0.91125 0.25617 0.069312 0.0096402 4.3139 0.060178 7.2426e-005 0.82989 0.005335 0.0060731 0.001584 0.98432 0.98969 3.4436e-006 1.3775e-005 0.13237 0.74228 0.79343 0.0014983 0.81965 0.5017 0.0020146 0.42295 1.3486 1.345 16.0065 144.979 0.00036097 -84.8522 0.18595
1.29 0.98803 5.5176e-005 3.8182 0.012033 1.6975e-005 0.0011542 0.16075 0.00065847 0.16141 0.14737 0 0.036319 0.0389 0 0.91133 0.25621 0.069325 0.0096418 4.3143 0.060188 7.2439e-005 0.82988 0.0053354 0.0060735 0.0015824 0.98434 0.98972 3.44e-006 1.376e-005 0.13237 0.74303 0.79401 0.0014976 0.82071 0.50187 0.0020136 0.42296 1.3504 1.3468 16.0065 144.979 0.00036005 -84.8581 0.18695
1.291 0.98803 5.5176e-005 3.8182 0.012033 1.6988e-005 0.0011542 0.16081 0.00065847 0.16147 0.14743 0 0.036315 0.0389 0 0.91142 0.25625 0.069338 0.0096434 4.3148 0.060198 7.2451e-005 0.82987 0.0053358 0.0060739 0.0015809 0.98436 0.98975 3.4364e-006 1.3746e-005 0.13237 0.74378 0.79458 0.0014968 0.82177 0.50204 0.0020126 0.42296 1.3522 1.3485 16.0065 144.979 0.00035913 -84.864 0.18795
1.292 0.98803 5.5176e-005 3.8182 0.012033 1.7002e-005 0.0011542 0.16087 0.00065848 0.16153 0.14749 0 0.036311 0.0389 0 0.9115 0.25628 0.069351 0.009645 4.3152 0.060208 7.2464e-005 0.82986 0.0053362 0.0060743 0.0015793 0.98438 0.98978 3.4329e-006 1.3732e-005 0.13238 0.74452 0.79516 0.001496 0.82282 0.50221 0.0020116 0.42297 1.3539 1.3503 16.0066 144.9791 0.00035821 -84.8698 0.18895
1.293 0.98803 5.5176e-005 3.8182 0.012033 1.7015e-005 0.0011542 0.16093 0.00065848 0.16159 0.14754 0 0.036308 0.0389 0 0.91158 0.25632 0.069364 0.0096466 4.3156 0.060217 7.2476e-005 0.82986 0.0053367 0.0060747 0.0015778 0.98441 0.98981 3.4294e-006 1.3718e-005 0.13238 0.74527 0.79573 0.0014953 0.82387 0.50238 0.0020106 0.42298 1.3556 1.3521 16.0066 144.9791 0.0003573 -84.8756 0.18995
1.294 0.98803 5.5176e-005 3.8182 0.012033 1.7028e-005 0.0011542 0.16099 0.00065848 0.16165 0.1476 0 0.036304 0.0389 0 0.91166 0.25635 0.069377 0.0096481 4.316 0.060227 7.2489e-005 0.82985 0.0053371 0.0060752 0.0015763 0.98443 0.98983 3.4259e-006 1.3704e-005 0.13238 0.74601 0.79629 0.0014945 0.8249 0.50254 0.0020097 0.42298 1.3574 1.3538 16.0067 144.9791 0.00035639 -84.8813 0.19095
1.295 0.98803 5.5176e-005 3.8182 0.012033 1.7041e-005 0.0011542 0.16105 0.00065848 0.16171 0.14765 0 0.0363 0.0389 0 0.91174 0.25639 0.06939 0.0096497 4.3164 0.060237 7.2502e-005 0.82984 0.0053375 0.0060756 0.0015748 0.98445 0.98986 3.4225e-006 1.369e-005 0.13239 0.74674 0.79686 0.0014938 0.82594 0.50271 0.0020087 0.42299 1.3591 1.3556 16.0067 144.9791 0.00035549 -84.887 0.19195
1.296 0.98803 5.5176e-005 3.8182 0.012033 1.7054e-005 0.0011542 0.16111 0.00065848 0.16177 0.14771 0 0.036297 0.0389 0 0.91182 0.25643 0.069403 0.0096513 4.3168 0.060247 7.2514e-005 0.82983 0.0053379 0.006076 0.0015733 0.98447 0.98988 3.4191e-006 1.3677e-005 0.13239 0.74748 0.79742 0.0014931 0.82697 0.50288 0.0020077 0.42299 1.3609 1.3573 16.0068 144.9791 0.00035459 -84.8926 0.19295
1.297 0.98803 5.5176e-005 3.8182 0.012033 1.7067e-005 0.0011542 0.16117 0.00065848 0.16183 0.14777 0 0.036293 0.0389 0 0.9119 0.25646 0.069416 0.0096529 4.3173 0.060257 7.2527e-005 0.82982 0.0053383 0.0060765 0.0015719 0.98449 0.98991 3.4157e-006 1.3663e-005 0.13239 0.74821 0.79797 0.0014923 0.82799 0.50305 0.0020068 0.423 1.3626 1.359 16.0068 144.9791 0.00035369 -84.8982 0.19395
1.298 0.98803 5.5175e-005 3.8182 0.012033 1.708e-005 0.0011542 0.16123 0.00065848 0.16189 0.14782 0 0.036289 0.0389 0 0.91198 0.2565 0.069429 0.0096545 4.3177 0.060266 7.254e-005 0.82981 0.0053388 0.0060769 0.0015704 0.98451 0.98993 3.4123e-006 1.365e-005 0.1324 0.74894 0.79853 0.0014916 0.82901 0.50322 0.0020058 0.42301 1.3643 1.3608 16.0068 144.9791 0.0003528 -84.9038 0.19495
1.299 0.98803 5.5175e-005 3.8182 0.012033 1.7093e-005 0.0011542 0.16129 0.00065848 0.16195 0.14788 0 0.036285 0.0389 0 0.91206 0.25653 0.069442 0.0096561 4.3181 0.060276 7.2552e-005 0.8298 0.0053392 0.0060773 0.001569 0.98453 0.98995 3.409e-006 1.3636e-005 0.1324 0.74967 0.79908 0.0014909 0.83002 0.50339 0.0020049 0.42302 1.366 1.3625 16.0069 144.9792 0.00035192 -84.9093 0.19595
1.3 0.98803 5.5175e-005 3.8182 0.012033 1.7107e-005 0.0011542 0.16135 0.00065848 0.16201 0.14793 0 0.036282 0.0389 0 0.91215 0.25657 0.069455 0.0096576 4.3185 0.060286 7.2565e-005 0.82979 0.0053396 0.0060777 0.0015675 0.98455 0.98998 3.4057e-006 1.3623e-005 0.13241 0.7504 0.79963 0.0014902 0.83103 0.50356 0.0020039 0.42302 1.3677 1.3642 16.0069 144.9792 0.00035104 -84.9148 0.19695
1.301 0.98803 5.5175e-005 3.8182 0.012033 1.712e-005 0.0011542 0.16141 0.00065848 0.16207 0.14799 0 0.036278 0.0389 0 0.91223 0.25661 0.069468 0.0096592 4.3189 0.060296 7.2577e-005 0.82978 0.00534 0.0060782 0.0015661 0.98456 0.99 3.4024e-006 1.361e-005 0.13241 0.75112 0.80018 0.0014895 0.83203 0.50373 0.002003 0.42303 1.3694 1.366 16.007 144.9792 0.00035016 -84.9202 0.19795
1.302 0.98803 5.5175e-005 3.8182 0.012033 1.7133e-005 0.0011542 0.16147 0.00065849 0.16212 0.14805 0 0.036274 0.0389 0 0.91231 0.25664 0.069481 0.0096608 4.3193 0.060305 7.259e-005 0.82977 0.0053404 0.0060786 0.0015647 0.98458 0.99002 3.3992e-006 1.3597e-005 0.13241 0.75184 0.80072 0.0014888 0.83302 0.50389 0.0020021 0.42304 1.3712 1.3677 16.007 144.9792 0.00034929 -84.9256 0.19895
1.303 0.98803 5.5175e-005 3.8182 0.012033 1.7146e-005 0.0011542 0.16153 0.00065849 0.16218 0.1481 0 0.036271 0.0389 0 0.91239 0.25668 0.069494 0.0096624 4.3198 0.060315 7.2603e-005 0.82976 0.0053409 0.006079 0.0015633 0.9846 0.99004 3.396e-006 1.3584e-005 0.13242 0.75256 0.80126 0.0014881 0.83401 0.50406 0.0020012 0.42304 1.3729 1.3694 16.007 144.9792 0.00034842 -84.9309 0.19995
1.304 0.98803 5.5175e-005 3.8182 0.012033 1.7159e-005 0.0011542 0.16159 0.00065849 0.16224 0.14816 0 0.036267 0.0389 0 0.91247 0.25672 0.069507 0.009664 4.3202 0.060325 7.2615e-005 0.82975 0.0053413 0.0060794 0.001562 0.98462 0.99006 3.3928e-006 1.3571e-005 0.13242 0.75328 0.8018 0.0014874 0.835 0.50423 0.0020003 0.42305 1.3746 1.3711 16.0071 144.9792 0.00034755 -84.9362 0.20095
1.305 0.98803 5.5175e-005 3.8182 0.012033 1.7172e-005 0.0011542 0.16165 0.00065849 0.1623 0.14821 0 0.036263 0.0389 0 0.91255 0.25675 0.06952 0.0096656 4.3206 0.060335 7.2628e-005 0.82974 0.0053417 0.0060799 0.0015606 0.98464 0.99008 3.3896e-006 1.3559e-005 0.13242 0.754 0.80233 0.0014867 0.83598 0.5044 0.0019994 0.42306 1.3762 1.3728 16.0071 144.9792 0.00034669 -84.9415 0.20195
1.306 0.98803 5.5175e-005 3.8182 0.012033 1.7185e-005 0.0011542 0.16171 0.00065849 0.16236 0.14827 0 0.03626 0.0389 0 0.91263 0.25679 0.069533 0.0096672 4.321 0.060345 7.2641e-005 0.82973 0.0053421 0.0060803 0.0015592 0.98466 0.9901 3.3865e-006 1.3546e-005 0.13243 0.75471 0.80286 0.001486 0.83695 0.50457 0.0019985 0.42306 1.3779 1.3745 16.0071 144.9793 0.00034584 -84.9467 0.20295
1.307 0.98803 5.5175e-005 3.8182 0.012033 1.7199e-005 0.0011542 0.16177 0.00065849 0.16242 0.14832 0 0.036256 0.0389 0 0.91271 0.25682 0.069546 0.0096687 4.3214 0.060354 7.2653e-005 0.82972 0.0053426 0.0060807 0.0015579 0.98468 0.99011 3.3834e-006 1.3534e-005 0.13243 0.75542 0.80339 0.0014853 0.83792 0.50474 0.0019976 0.42307 1.3796 1.3762 16.0072 144.9793 0.00034499 -84.9519 0.20395
1.308 0.98803 5.5175e-005 3.8182 0.012033 1.7212e-005 0.0011542 0.16183 0.00065849 0.16248 0.14838 0 0.036252 0.0389 0 0.9128 0.25686 0.069559 0.0096703 4.3219 0.060364 7.2666e-005 0.82971 0.005343 0.0060812 0.0015565 0.98469 0.99013 3.3803e-006 1.3521e-005 0.13243 0.75613 0.80392 0.0014847 0.83888 0.50491 0.0019967 0.42308 1.3813 1.3779 16.0072 144.9793 0.00034414 -84.9571 0.20495
1.309 0.98803 5.5175e-005 3.8182 0.012033 1.7225e-005 0.0011542 0.16189 0.00065849 0.16254 0.14843 0 0.036249 0.0389 0 0.91288 0.2569 0.069572 0.0096719 4.3223 0.060374 7.2679e-005 0.8297 0.0053434 0.0060816 0.0015552 0.98471 0.99015 3.3772e-006 1.3509e-005 0.13244 0.75684 0.80444 0.001484 0.83984 0.50507 0.0019959 0.42309 1.383 1.3796 16.0073 144.9793 0.0003433 -84.9622 0.20595
1.31 0.98803 5.5175e-005 3.8182 0.012033 1.7238e-005 0.0011542 0.16194 0.00065849 0.1626 0.14849 0 0.036245 0.0389 0 0.91296 0.25693 0.069586 0.0096735 4.3227 0.060384 7.2691e-005 0.82969 0.0053438 0.006082 0.0015539 0.98473 0.99016 3.3742e-006 1.3497e-005 0.13244 0.75754 0.80497 0.0014833 0.84079 0.50524 0.001995 0.42309 1.3847 1.3813 16.0073 144.9793 0.00034246 -84.9673 0.20695
1.311 0.98803 5.5175e-005 3.8182 0.012033 1.7251e-005 0.0011542 0.162 0.00065849 0.16266 0.14855 0 0.036241 0.0389 0 0.91304 0.25697 0.069599 0.0096751 4.3231 0.060394 7.2704e-005 0.82968 0.0053443 0.0060825 0.0015526 0.98475 0.99018 3.3712e-006 1.3485e-005 0.13244 0.75824 0.80549 0.0014827 0.84174 0.50541 0.0019942 0.4231 1.3863 1.383 16.0073 144.9793 0.00034162 -84.9723 0.20795
1.312 0.98803 5.5175e-005 3.8182 0.012032 1.7264e-005 0.0011542 0.16206 0.0006585 0.16272 0.1486 0 0.036238 0.0389 0 0.91312 0.25701 0.069612 0.0096767 4.3235 0.060403 7.2717e-005 0.82967 0.0053447 0.0060829 0.0015513 0.98477 0.9902 3.3682e-006 1.3473e-005 0.13245 0.75894 0.806 0.001482 0.84268 0.50558 0.0019933 0.42311 1.388 1.3846 16.0074 144.9793 0.00034079 -84.9773 0.20895
1.313 0.98803 5.5175e-005 3.8182 0.012032 1.7277e-005 0.0011542 0.16212 0.0006585 0.16278 0.14866 0 0.036234 0.0389 0 0.9132 0.25704 0.069625 0.0096783 4.324 0.060413 7.2729e-005 0.82966 0.0053451 0.0060833 0.00155 0.98478 0.99021 3.3652e-006 1.3461e-005 0.13245 0.75964 0.80652 0.0014814 0.84362 0.50575 0.0019925 0.42312 1.3896 1.3863 16.0074 144.9794 0.00033996 -84.9823 0.20995
1.314 0.98803 5.5174e-005 3.8182 0.012032 1.729e-005 0.0011542 0.16218 0.0006585 0.16283 0.14871 0 0.03623 0.0389 0 0.91329 0.25708 0.069638 0.0096799 4.3244 0.060423 7.2742e-005 0.82965 0.0053455 0.0060838 0.0015488 0.9848 0.99023 3.3623e-006 1.345e-005 0.13245 0.76034 0.80703 0.0014807 0.84455 0.50592 0.0019916 0.42312 1.3913 1.388 16.0074 144.9794 0.00033914 -84.9872 0.21095
1.315 0.98803 5.5174e-005 3.8182 0.012032 1.7304e-005 0.0011542 0.16224 0.0006585 0.16289 0.14877 0 0.036227 0.0389 0 0.91337 0.25711 0.069651 0.0096815 4.3248 0.060433 7.2755e-005 0.82964 0.005346 0.0060842 0.0015475 0.98482 0.99024 3.3594e-006 1.3438e-005 0.13246 0.76103 0.80753 0.0014801 0.84547 0.50608 0.0019908 0.42313 1.393 1.3896 16.0075 144.9794 0.00033832 -84.9921 0.21195
1.316 0.98803 5.5174e-005 3.8182 0.012032 1.7317e-005 0.0011542 0.1623 0.0006585 0.16295 0.14882 0 0.036223 0.0389 0 0.91345 0.25715 0.069664 0.009683 4.3252 0.060443 7.2767e-005 0.82963 0.0053464 0.0060846 0.0015462 0.98483 0.99026 3.3565e-006 1.3426e-005 0.13246 0.76172 0.80804 0.0014795 0.8464 0.50625 0.00199 0.42314 1.3946 1.3913 16.0075 144.9794 0.00033751 -84.9969 0.21295
1.317 0.98803 5.5174e-005 3.8182 0.012032 1.733e-005 0.0011542 0.16236 0.0006585 0.16301 0.14888 0 0.036219 0.0389 0 0.91353 0.25719 0.069677 0.0096846 4.3257 0.060453 7.278e-005 0.82962 0.0053468 0.0060851 0.001545 0.98485 0.99027 3.3537e-006 1.3415e-005 0.13247 0.76241 0.80854 0.0014789 0.84731 0.50642 0.0019892 0.42315 1.3962 1.393 16.0075 144.9794 0.0003367 -85.0017 0.21395
1.318 0.98803 5.5174e-005 3.8182 0.012032 1.7343e-005 0.0011542 0.16242 0.0006585 0.16307 0.14893 0 0.036216 0.0389 0 0.91361 0.25722 0.06969 0.0096862 4.3261 0.060462 7.2793e-005 0.82961 0.0053472 0.0060855 0.0015438 0.98487 0.99029 3.3508e-006 1.3404e-005 0.13247 0.7631 0.80905 0.0014782 0.84822 0.50659 0.0019884 0.42316 1.3979 1.3946 16.0076 144.9794 0.00033589 -85.0065 0.21495
1.319 0.98803 5.5174e-005 3.8182 0.012032 1.7356e-005 0.0011542 0.16247 0.0006585 0.16313 0.14899 0 0.036212 0.0389 0 0.91369 0.25726 0.069704 0.0096878 4.3265 0.060472 7.2806e-005 0.8296 0.0053477 0.0060859 0.0015426 0.98488 0.9903 3.348e-006 1.3392e-005 0.13247 0.76378 0.80954 0.0014776 0.84913 0.50676 0.0019876 0.42316 1.3995 1.3962 16.0076 144.9795 0.00033509 -85.0113 0.21595
1.32 0.98803 5.5174e-005 3.8182 0.012032 1.7369e-005 0.0011542 0.16253 0.0006585 0.16319 0.14904 0 0.036209 0.0389 0 0.91378 0.2573 0.069717 0.0096894 4.3269 0.060482 7.2818e-005 0.82959 0.0053481 0.0060864 0.0015414 0.9849 0.99031 3.3452e-006 1.3381e-005 0.13248 0.76447 0.81004 0.001477 0.85003 0.50692 0.0019868 0.42317 1.4012 1.3979 16.0076 144.9795 0.00033429 -85.016 0.21695
1.321 0.98803 5.5174e-005 3.8182 0.012032 1.7382e-005 0.0011542 0.16259 0.0006585 0.16324 0.1491 0 0.036205 0.0389 0 0.91386 0.25733 0.06973 0.009691 4.3274 0.060492 7.2831e-005 0.82958 0.0053485 0.0060868 0.0015402 0.98492 0.99033 3.3425e-006 1.337e-005 0.13248 0.76515 0.81053 0.0014764 0.85093 0.50709 0.001986 0.42318 1.4028 1.3995 16.0077 144.9795 0.00033349 -85.0206 0.21795
1.322 0.98803 5.5174e-005 3.8182 0.012032 1.7395e-005 0.0011542 0.16265 0.0006585 0.1633 0.14915 0 0.036201 0.0389 0 0.91394 0.25737 0.069743 0.0096926 4.3278 0.060502 7.2844e-005 0.82957 0.005349 0.0060872 0.001539 0.98493 0.99034 3.3397e-006 1.3359e-005 0.13248 0.76582 0.81102 0.0014758 0.85182 0.50726 0.0019852 0.42319 1.4044 1.4012 16.0077 144.9795 0.0003327 -85.0253 0.21895
1.323 0.98803 5.5174e-005 3.8182 0.012032 1.7409e-005 0.0011542 0.16271 0.00065851 0.16336 0.14921 0 0.036198 0.0389 0 0.91402 0.25741 0.069756 0.0096942 4.3282 0.060512 7.2856e-005 0.82956 0.0053494 0.0060877 0.0015378 0.98495 0.99035 3.337e-006 1.3348e-005 0.13249 0.7665 0.81151 0.0014752 0.8527 0.50743 0.0019844 0.4232 1.406 1.4028 16.0077 144.9795 0.00033191 -85.0299 0.21995
1.324 0.98803 5.5174e-005 3.8182 0.012032 1.7422e-005 0.0011542 0.16277 0.00065851 0.16342 0.14926 0 0.036194 0.0389 0 0.9141 0.25744 0.069769 0.0096958 4.3287 0.060522 7.2869e-005 0.82955 0.0053498 0.0060881 0.0015366 0.98496 0.99036 3.3343e-006 1.3338e-005 0.13249 0.76718 0.812 0.0014746 0.85358 0.5076 0.0019836 0.4232 1.4076 1.4044 16.0078 144.9795 0.00033113 -85.0344 0.22095
1.325 0.98803 5.5174e-005 3.8182 0.012032 1.7435e-005 0.0011542 0.16282 0.00065851 0.16348 0.14932 0 0.036191 0.0389 0 0.91418 0.25748 0.069782 0.0096974 4.3291 0.060531 7.2882e-005 0.82954 0.0053502 0.0060885 0.0015355 0.98498 0.99038 3.3317e-006 1.3327e-005 0.13249 0.76785 0.81248 0.0014741 0.85446 0.50776 0.0019829 0.42321 1.4092 1.406 16.0078 144.9795 0.00033035 -85.039 0.22195
1.326 0.98803 5.5174e-005 3.8182 0.012032 1.7448e-005 0.0011542 0.16288 0.00065851 0.16354 0.14937 0 0.036187 0.0389 0 0.91427 0.25752 0.069795 0.009699 4.3295 0.060541 7.2895e-005 0.82953 0.0053507 0.006089 0.0015343 0.98499 0.99039 3.329e-006 1.3316e-005 0.1325 0.76852 0.81297 0.0014735 0.85533 0.50793 0.0019821 0.42322 1.4109 1.4077 16.0078 144.9796 0.00032957 -85.0434 0.22295
1.327 0.98803 5.5174e-005 3.8182 0.012032 1.7461e-005 0.0011542 0.16294 0.00065851 0.1636 0.14942 0 0.036183 0.0389 0 0.91435 0.25755 0.069809 0.0097006 4.3299 0.060551 7.2907e-005 0.82952 0.0053511 0.0060894 0.0015332 0.98501 0.9904 3.3264e-006 1.3306e-005 0.1325 0.76919 0.81344 0.0014729 0.8562 0.5081 0.0019814 0.42323 1.4125 1.4093 16.0079 144.9796 0.0003288 -85.0479 0.22395
1.328 0.98803 5.5174e-005 3.8182 0.012032 1.7474e-005 0.0011543 0.163 0.00065851 0.16365 0.14948 0 0.03618 0.0389 0 0.91443 0.25759 0.069822 0.0097022 4.3304 0.060561 7.292e-005 0.82951 0.0053515 0.0060899 0.001532 0.98503 0.99041 3.3238e-006 1.3295e-005 0.1325 0.76985 0.81392 0.0014723 0.85706 0.50827 0.0019806 0.42324 1.4141 1.4109 16.0079 144.9796 0.00032803 -85.0523 0.22495
1.329 0.98803 5.5174e-005 3.8182 0.012032 1.7487e-005 0.0011543 0.16306 0.00065851 0.16371 0.14953 0 0.036176 0.0389 0 0.91451 0.25762 0.069835 0.0097038 4.3308 0.060571 7.2933e-005 0.8295 0.005352 0.0060903 0.0015309 0.98504 0.99042 3.3212e-006 1.3285e-005 0.13251 0.77052 0.8144 0.0014718 0.85791 0.50844 0.0019799 0.42325 1.4157 1.4125 16.0079 144.9796 0.00032726 -85.0567 0.22595
1.33 0.98803 5.5173e-005 3.8182 0.012032 1.75e-005 0.0011543 0.16312 0.00065851 0.16377 0.14959 0 0.036173 0.0389 0 0.91459 0.25766 0.069848 0.0097054 4.3312 0.060581 7.2946e-005 0.82949 0.0053524 0.0060907 0.0015298 0.98506 0.99044 3.3186e-006 1.3275e-005 0.13251 0.77118 0.81487 0.0014712 0.85876 0.5086 0.0019792 0.42325 1.4172 1.4141 16.0079 144.9796 0.0003265 -85.0611 0.22695
1.331 0.98803 5.5173e-005 3.8182 0.012032 1.7514e-005 0.0011543 0.16317 0.00065851 0.16383 0.14964 0 0.036169 0.0389 0 0.91468 0.2577 0.069861 0.009707 4.3317 0.060591 7.2958e-005 0.82948 0.0053528 0.0060912 0.0015287 0.98507 0.99045 3.3161e-006 1.3265e-005 0.13251 0.77184 0.81534 0.0014706 0.85961 0.50877 0.0019784 0.42326 1.4188 1.4157 16.008 144.9796 0.00032574 -85.0654 0.22795
1.332 0.98803 5.5173e-005 3.8182 0.012032 1.7527e-005 0.0011543 0.16323 0.00065851 0.16389 0.1497 0 0.036165 0.0389 0 0.91476 0.25773 0.069874 0.0097086 4.3321 0.0606 7.2971e-005 0.82947 0.0053533 0.0060916 0.0015276 0.98508 0.99046 3.3136e-006 1.3254e-005 0.13252 0.7725 0.81581 0.0014701 0.86045 0.50894 0.0019777 0.42327 1.4204 1.4173 16.008 144.9797 0.00032499 -85.0697 0.22895
1.333 0.98803 5.5173e-005 3.8182 0.012032 1.754e-005 0.0011543 0.16329 0.00065852 0.16394 0.14975 0 0.036162 0.0389 0 0.91484 0.25777 0.069888 0.0097102 4.3325 0.06061 7.2984e-005 0.82946 0.0053537 0.006092 0.0015265 0.9851 0.99047 3.3111e-006 1.3244e-005 0.13252 0.77315 0.81627 0.0014695 0.86129 0.50911 0.001977 0.42328 1.422 1.4189 16.008 144.9797 0.00032424 -85.074 0.22995
1.334 0.98803 5.5173e-005 3.8182 0.012032 1.7553e-005 0.0011543 0.16335 0.00065852 0.164 0.14981 0 0.036158 0.0389 0 0.91492 0.25781 0.069901 0.0097118 4.333 0.06062 7.2997e-005 0.82945 0.0053541 0.0060925 0.0015254 0.98511 0.99048 3.3086e-006 1.3234e-005 0.13253 0.77381 0.81673 0.001469 0.86212 0.50927 0.0019763 0.42329 1.4236 1.4205 16.0081 144.9797 0.00032349 -85.0782 0.23095
1.335 0.98803 5.5173e-005 3.8182 0.012032 1.7566e-005 0.0011543 0.16341 0.00065852 0.16406 0.14986 0 0.036155 0.0389 0 0.915 0.25784 0.069914 0.0097134 4.3334 0.06063 7.3009e-005 0.82944 0.0053546 0.0060929 0.0015244 0.98513 0.99049 3.3061e-006 1.3225e-005 0.13253 0.77446 0.8172 0.0014685 0.86295 0.50944 0.0019756 0.4233 1.4251 1.422 16.0081 144.9797 0.00032275 -85.0824 0.23195
1.336 0.98803 5.5173e-005 3.8182 0.012032 1.7579e-005 0.0011543 0.16346 0.00065852 0.16412 0.14991 0 0.036151 0.0389 0 0.91509 0.25788 0.069927 0.009715 4.3338 0.06064 7.3022e-005 0.82943 0.005355 0.0060934 0.0015233 0.98514 0.9905 3.3037e-006 1.3215e-005 0.13253 0.77511 0.81765 0.0014679 0.86377 0.50961 0.0019749 0.42331 1.4267 1.4236 16.0081 144.9797 0.00032201 -85.0866 0.23295
1.337 0.98803 5.5173e-005 3.8182 0.012032 1.7592e-005 0.0011543 0.16352 0.00065852 0.16418 0.14997 0 0.036148 0.0389 0 0.91517 0.25792 0.06994 0.0097166 4.3343 0.06065 7.3035e-005 0.82942 0.0053554 0.0060938 0.0015223 0.98516 0.99051 3.3013e-006 1.3205e-005 0.13254 0.77576 0.81811 0.0014674 0.86459 0.50978 0.0019742 0.42332 1.4283 1.4252 16.0082 144.9797 0.00032127 -85.0908 0.23395
1.338 0.98803 5.5173e-005 3.8182 0.012032 1.7606e-005 0.0011543 0.16358 0.00065852 0.16423 0.15002 0 0.036144 0.0389 0 0.91525 0.25795 0.069954 0.0097182 4.3347 0.06066 7.3048e-005 0.82941 0.0053559 0.0060942 0.0015212 0.98517 0.99052 3.2989e-006 1.3196e-005 0.13254 0.7764 0.81856 0.0014669 0.8654 0.50994 0.0019735 0.42332 1.4298 1.4268 16.0082 144.9798 0.00032054 -85.0949 0.23495
1.339 0.98803 5.5173e-005 3.8182 0.012032 1.7619e-005 0.0011543 0.16364 0.00065852 0.16429 0.15008 0 0.03614 0.0389 0 0.91533 0.25799 0.069967 0.0097198 4.3351 0.06067 7.306e-005 0.8294 0.0053563 0.0060947 0.0015202 0.98518 0.99053 3.2965e-006 1.3186e-005 0.13254 0.77705 0.81902 0.0014663 0.86621 0.51011 0.0019728 0.42333 1.4314 1.4283 16.0082 144.9798 0.00031981 -85.0989 0.23595
1.34 0.98803 5.5173e-005 3.8182 0.012032 1.7632e-005 0.0011543 0.16369 0.00065852 0.16435 0.15013 0 0.036137 0.0389 0 0.91542 0.25803 0.06998 0.0097214 4.3356 0.06068 7.3073e-005 0.82939 0.0053567 0.0060951 0.0015192 0.9852 0.99054 3.2941e-006 1.3177e-005 0.13255 0.77769 0.81947 0.0014658 0.86702 0.51028 0.0019721 0.42334 1.4329 1.4299 16.0082 144.9798 0.00031908 -85.103 0.23695
1.341 0.98803 5.5173e-005 3.8182 0.012032 1.7645e-005 0.0011543 0.16375 0.00065852 0.16441 0.15019 0 0.036133 0.0389 0 0.9155 0.25806 0.069993 0.009723 4.336 0.060689 7.3086e-005 0.82938 0.0053572 0.0060956 0.0015181 0.98521 0.99055 3.2918e-006 1.3167e-005 0.13255 0.77833 0.81991 0.0014653 0.86782 0.51045 0.0019714 0.42335 1.4345 1.4314 16.0083 144.9798 0.00031836 -85.107 0.23795
1.342 0.98803 5.5173e-005 3.8182 0.012032 1.7658e-005 0.0011543 0.16381 0.00065852 0.16446 0.15024 0 0.03613 0.0389 0 0.91558 0.2581 0.070006 0.0097246 4.3364 0.060699 7.3099e-005 0.82937 0.0053576 0.006096 0.0015171 0.98523 0.99056 3.2894e-006 1.3158e-005 0.13255 0.77897 0.82036 0.0014648 0.86861 0.51061 0.0019708 0.42336 1.436 1.433 16.0083 144.9798 0.00031764 -85.111 0.23895
1.343 0.98803 5.5173e-005 3.8182 0.012032 1.7671e-005 0.0011543 0.16387 0.00065852 0.16452 0.15029 0 0.036126 0.0389 0 0.91566 0.25814 0.07002 0.0097262 4.3369 0.060709 7.3112e-005 0.82936 0.005358 0.0060965 0.0015161 0.98524 0.99057 3.2871e-006 1.3149e-005 0.13256 0.77961 0.8208 0.0014643 0.8694 0.51078 0.0019701 0.42337 1.4376 1.4346 16.0083 144.9798 0.00031692 -85.115 0.23995
1.344 0.98803 5.5173e-005 3.8182 0.012032 1.7684e-005 0.0011543 0.16392 0.00065853 0.16458 0.15035 0 0.036123 0.0389 0 0.91574 0.25817 0.070033 0.0097278 4.3373 0.060719 7.3124e-005 0.82935 0.0053585 0.0060969 0.0015151 0.98525 0.99058 3.2849e-006 1.314e-005 0.13256 0.78024 0.82124 0.0014638 0.87019 0.51095 0.0019694 0.42338 1.4391 1.4361 16.0083 144.9799 0.00031621 -85.1189 0.24095
1.345 0.98803 5.5173e-005 3.8182 0.012032 1.7697e-005 0.0011543 0.16398 0.00065853 0.16464 0.1504 0 0.036119 0.0389 0 0.91583 0.25821 0.070046 0.0097294 4.3377 0.060729 7.3137e-005 0.82934 0.0053589 0.0060973 0.0015142 0.98527 0.99059 3.2826e-006 1.3131e-005 0.13257 0.78087 0.82168 0.0014633 0.87097 0.51112 0.0019688 0.42339 1.4406 1.4376 16.0084 144.9799 0.0003155 -85.1228 0.24195
1.346 0.98803 5.5172e-005 3.8182 0.012032 1.7711e-005 0.0011543 0.16404 0.00065853 0.16469 0.15045 0 0.036116 0.0389 0 0.91591 0.25825 0.070059 0.009731 4.3382 0.060739 7.315e-005 0.82933 0.0053594 0.0060978 0.0015132 0.98528 0.9906 3.2803e-006 1.3122e-005 0.13257 0.7815 0.82212 0.0014628 0.87175 0.51128 0.0019681 0.4234 1.4421 1.4392 16.0084 144.9799 0.0003148 -85.1267 0.24295
1.347 0.98803 5.5172e-005 3.8182 0.012032 1.7724e-005 0.0011543 0.1641 0.00065853 0.16475 0.15051 0 0.036112 0.0389 0 0.91599 0.25828 0.070073 0.0097326 4.3386 0.060749 7.3163e-005 0.82932 0.0053598 0.0060982 0.0015122 0.98529 0.99061 3.2781e-006 1.3113e-005 0.13257 0.78213 0.82256 0.0014623 0.87252 0.51145 0.0019675 0.42341 1.4437 1.4407 16.0084 144.9799 0.00031409 -85.1305 0.24395
1.348 0.98803 5.5172e-005 3.8182 0.012032 1.7737e-005 0.0011543 0.16415 0.00065853 0.16481 0.15056 0 0.036109 0.0389 0 0.91607 0.25832 0.070086 0.0097342 4.3391 0.060759 7.3176e-005 0.82931 0.0053602 0.0060987 0.0015113 0.9853 0.99062 3.2759e-006 1.3104e-005 0.13258 0.78276 0.82299 0.0014618 0.87329 0.51162 0.0019669 0.42341 1.4452 1.4422 16.0085 144.9799 0.0003134 -85.1343 0.24495
1.349 0.98803 5.5172e-005 3.8182 0.012032 1.775e-005 0.0011543 0.16421 0.00065853 0.16486 0.15062 0 0.036105 0.0389 0 0.91616 0.25836 0.070099 0.0097358 4.3395 0.060769 7.3189e-005 0.8293 0.0053607 0.0060991 0.0015103 0.98532 0.99063 3.2737e-006 1.3095e-005 0.13258 0.78338 0.82342 0.0014613 0.87405 0.51178 0.0019662 0.42342 1.4467 1.4438 16.0085 144.9799 0.0003127 -85.1381 0.24595
1.35 0.98803 5.5172e-005 3.8182 0.012032 1.7763e-005 0.0011543 0.16427 0.00065853 0.16492 0.15067 0 0.036102 0.0389 0 0.91624 0.25839 0.070112 0.0097374 4.3399 0.060779 7.3201e-005 0.82929 0.0053611 0.0060996 0.0015094 0.98533 0.99063 3.2715e-006 1.3086e-005 0.13258 0.784 0.82385 0.0014608 0.87481 0.51195 0.0019656 0.42343 1.4482 1.4453 16.0085 144.9799 0.00031201 -85.1419 0.24695
1.351 0.98803 5.5172e-005 3.8182 0.012032 1.7776e-005 0.0011543 0.16433 0.00065853 0.16498 0.15072 0 0.036098 0.0389 0 0.91632 0.25843 0.070126 0.009739 4.3404 0.060789 7.3214e-005 0.82928 0.0053615 0.0061 0.0015084 0.98534 0.99064 3.2694e-006 1.3078e-005 0.13259 0.78462 0.82428 0.0014604 0.87557 0.51212 0.001965 0.42344 1.4497 1.4468 16.0085 144.98 0.00031132 -85.1456 0.24795
1.352 0.98803 5.5172e-005 3.8182 0.012032 1.7789e-005 0.0011543 0.16438 0.00065853 0.16504 0.15078 0 0.036094 0.0389 0 0.9164 0.25847 0.070139 0.0097406 4.3408 0.060799 7.3227e-005 0.82927 0.005362 0.0061005 0.0015075 0.98535 0.99065 3.2672e-006 1.3069e-005 0.13259 0.78524 0.8247 0.0014599 0.87632 0.51229 0.0019644 0.42345 1.4512 1.4483 16.0086 144.98 0.00031063 -85.1493 0.24895
1.353 0.98803 5.5172e-005 3.8182 0.012032 1.7802e-005 0.0011543 0.16444 0.00065853 0.16509 0.15083 0 0.036091 0.0389 0 0.91649 0.2585 0.070152 0.0097422 4.3413 0.060809 7.324e-005 0.82926 0.0053624 0.0061009 0.0015066 0.98537 0.99066 3.2651e-006 1.3061e-005 0.13259 0.78586 0.82512 0.0014594 0.87706 0.51245 0.0019637 0.42346 1.4527 1.4498 16.0086 144.98 0.00030995 -85.153 0.24995
1.354 0.98803 5.5172e-005 3.8182 0.012032 1.7816e-005 0.0011543 0.1645 0.00065853 0.16515 0.15088 0 0.036087 0.0389 0 0.91657 0.25854 0.070165 0.0097438 4.3417 0.060818 7.3253e-005 0.82925 0.0053629 0.0061014 0.0015056 0.98538 0.99067 3.263e-006 1.3052e-005 0.1326 0.78647 0.82555 0.001459 0.8778 0.51262 0.0019631 0.42347 1.4542 1.4513 16.0086 144.98 0.00030927 -85.1566 0.25095
1.355 0.98803 5.5172e-005 3.8182 0.012032 1.7829e-005 0.0011543 0.16455 0.00065854 0.16521 0.15094 0 0.036084 0.0389 0 0.91665 0.25858 0.070179 0.0097454 4.3421 0.060828 7.3266e-005 0.82924 0.0053633 0.0061018 0.0015047 0.98539 0.99068 3.2609e-006 1.3044e-005 0.1326 0.78709 0.82596 0.0014585 0.87854 0.51279 0.0019625 0.42348 1.4557 1.4528 16.0086 144.98 0.00030859 -85.1603 0.25195
1.356 0.98803 5.5172e-005 3.8182 0.012032 1.7842e-005 0.0011543 0.16461 0.00065854 0.16526 0.15099 0 0.03608 0.0389 0 0.91673 0.25861 0.070192 0.009747 4.3426 0.060838 7.3278e-005 0.82923 0.0053637 0.0061023 0.0015038 0.9854 0.99069 3.2588e-006 1.3035e-005 0.13261 0.7877 0.82638 0.001458 0.87927 0.51295 0.0019619 0.42349 1.4572 1.4543 16.0086 144.98 0.00030792 -85.1639 0.25295
1.357 0.98803 5.5172e-005 3.8182 0.012032 1.7855e-005 0.0011543 0.16467 0.00065854 0.16532 0.15104 0 0.036077 0.0389 0 0.91682 0.25865 0.070205 0.0097486 4.343 0.060848 7.3291e-005 0.82923 0.0053642 0.0061027 0.0015029 0.98541 0.99069 3.2568e-006 1.3027e-005 0.13261 0.78831 0.8268 0.0014576 0.88 0.51312 0.0019613 0.4235 1.4587 1.4558 16.0087 144.9801 0.00030725 -85.1674 0.25395
1.358 0.98803 5.5172e-005 3.8182 0.012032 1.7868e-005 0.0011543 0.16472 0.00065854 0.16538 0.1511 0 0.036073 0.0389 0 0.9169 0.25869 0.070218 0.0097503 4.3435 0.060858 7.3304e-005 0.82922 0.0053646 0.0061032 0.0015021 0.98543 0.9907 3.2547e-006 1.3019e-005 0.13261 0.78892 0.82721 0.0014571 0.88073 0.51329 0.0019607 0.42351 1.4602 1.4573 16.0087 144.9801 0.00030658 -85.171 0.25495
1.359 0.98803 5.5172e-005 3.8182 0.012032 1.7881e-005 0.0011543 0.16478 0.00065854 0.16543 0.15115 0 0.03607 0.0389 0 0.91698 0.25873 0.070232 0.0097519 4.3439 0.060868 7.3317e-005 0.82921 0.0053651 0.0061036 0.0015012 0.98544 0.99071 3.2527e-006 1.3011e-005 0.13262 0.78952 0.82762 0.0014567 0.88145 0.51345 0.0019602 0.42352 1.4616 1.4588 16.0087 144.9801 0.00030592 -85.1745 0.25595
1.36 0.98803 5.5172e-005 3.8182 0.012032 1.7894e-005 0.0011543 0.16484 0.00065854 0.16549 0.1512 0 0.036067 0.0389 0 0.91706 0.25876 0.070245 0.0097535 4.3444 0.060878 7.333e-005 0.8292 0.0053655 0.006104 0.0015003 0.98545 0.99072 3.2507e-006 1.3003e-005 0.13262 0.79012 0.82803 0.0014562 0.88216 0.51362 0.0019596 0.42353 1.4631 1.4603 16.0087 144.9801 0.00030526 -85.178 0.25695
1.361 0.98803 5.5171e-005 3.8182 0.012032 1.7907e-005 0.0011543 0.16489 0.00065854 0.16555 0.15126 0 0.036063 0.0389 0 0.91715 0.2588 0.070258 0.0097551 4.3448 0.060888 7.3343e-005 0.82919 0.005366 0.0061045 0.0014994 0.98546 0.99073 3.2487e-006 1.2995e-005 0.13262 0.79073 0.82844 0.0014558 0.88288 0.51379 0.001959 0.42354 1.4646 1.4618 16.0088 144.9801 0.0003046 -85.1814 0.25795
1.362 0.98803 5.5171e-005 3.8182 0.012032 1.7921e-005 0.0011543 0.16495 0.00065854 0.1656 0.15131 0 0.03606 0.0389 0 0.91723 0.25884 0.070272 0.0097567 4.3453 0.060898 7.3356e-005 0.82918 0.0053664 0.0061049 0.0014986 0.98547 0.99073 3.2467e-006 1.2987e-005 0.13263 0.79133 0.82884 0.0014554 0.88359 0.51395 0.0019584 0.42355 1.466 1.4632 16.0088 144.9801 0.00030395 -85.1849 0.25895
1.363 0.98803 5.5171e-005 3.8182 0.012032 1.7934e-005 0.0011543 0.16501 0.00065854 0.16566 0.15136 0 0.036056 0.0389 0 0.91731 0.25887 0.070285 0.0097583 4.3457 0.060908 7.3369e-005 0.82917 0.0053668 0.0061054 0.0014977 0.98548 0.99074 3.2448e-006 1.2979e-005 0.13263 0.79192 0.82925 0.0014549 0.88429 0.51412 0.0019579 0.42356 1.4675 1.4647 16.0088 144.9802 0.00030329 -85.1883 0.25995
1.364 0.98803 5.5171e-005 3.8182 0.012032 1.7947e-005 0.0011543 0.16506 0.00065854 0.16572 0.15142 0 0.036053 0.0389 0 0.9174 0.25891 0.070298 0.0097599 4.3461 0.060918 7.3381e-005 0.82916 0.0053673 0.0061059 0.0014969 0.9855 0.99075 3.2428e-006 1.2971e-005 0.13263 0.79252 0.82965 0.0014545 0.88499 0.51429 0.0019573 0.42357 1.4689 1.4662 16.0088 144.9802 0.00030265 -85.1917 0.26095
1.365 0.98803 5.5171e-005 3.8182 0.012032 1.796e-005 0.0011543 0.16512 0.00065854 0.16577 0.15147 0 0.036049 0.0389 0 0.91748 0.25895 0.070312 0.0097615 4.3466 0.060928 7.3394e-005 0.82915 0.0053677 0.0061063 0.001496 0.98551 0.99076 3.2409e-006 1.2964e-005 0.13264 0.79311 0.83005 0.0014541 0.88568 0.51445 0.0019567 0.42358 1.4704 1.4676 16.0089 144.9802 0.000302 -85.1951 0.26195
1.366 0.98803 5.5171e-005 3.8182 0.012032 1.7973e-005 0.0011543 0.16518 0.00065855 0.16583 0.15152 0 0.036046 0.0389 0 0.91756 0.25898 0.070325 0.0097631 4.347 0.060938 7.3407e-005 0.82914 0.0053682 0.0061068 0.0014952 0.98552 0.99076 3.239e-006 1.2956e-005 0.13264 0.79371 0.83045 0.0014536 0.88638 0.51462 0.0019562 0.42359 1.4718 1.4691 16.0089 144.9802 0.00030136 -85.1984 0.26295
1.367 0.98803 5.5171e-005 3.8182 0.012032 1.7986e-005 0.0011543 0.16523 0.00065855 0.16589 0.15158 0 0.036042 0.0389 0 0.91764 0.25902 0.070338 0.0097647 4.3475 0.060948 7.342e-005 0.82913 0.0053686 0.0061072 0.0014944 0.98553 0.99077 3.2371e-006 1.2948e-005 0.13265 0.7943 0.83084 0.0014532 0.88706 0.51479 0.0019556 0.4236 1.4733 1.4705 16.0089 144.9802 0.00030072 -85.2017 0.26395
1.368 0.98803 5.5171e-005 3.8182 0.012032 1.7999e-005 0.0011543 0.16529 0.00065855 0.16594 0.15163 0 0.036039 0.0389 0 0.91773 0.25906 0.070351 0.0097664 4.3479 0.060958 7.3433e-005 0.82912 0.0053691 0.0061077 0.0014936 0.98554 0.99078 3.2352e-006 1.2941e-005 0.13265 0.79489 0.83124 0.0014528 0.88775 0.51495 0.0019551 0.42361 1.4747 1.472 16.0089 144.9802 0.00030008 -85.205 0.26495
1.369 0.98803 5.5171e-005 3.8182 0.012032 1.8012e-005 0.0011543 0.16535 0.00065855 0.166 0.15168 0 0.036035 0.0389 0 0.91781 0.25909 0.070365 0.009768 4.3484 0.060968 7.3446e-005 0.82911 0.0053695 0.0061081 0.0014927 0.98555 0.99079 3.2333e-006 1.2933e-005 0.13265 0.79547 0.83163 0.0014524 0.88843 0.51512 0.0019545 0.42362 1.4762 1.4734 16.0089 144.9803 0.00029945 -85.2083 0.26595
1.37 0.98803 5.5171e-005 3.8182 0.012032 1.8026e-005 0.0011543 0.1654 0.00065855 0.16606 0.15173 0 0.036032 0.0389 0 0.91789 0.25913 0.070378 0.0097696 4.3488 0.060978 7.3459e-005 0.8291 0.0053699 0.0061086 0.0014919 0.98556 0.99079 3.2315e-006 1.2926e-005 0.13266 0.79606 0.83202 0.001452 0.8891 0.51529 0.001954 0.42363 1.4776 1.4749 16.009 144.9803 0.00029882 -85.2115 0.26695
1.371 0.98803 5.5171e-005 3.8182 0.012032 1.8039e-005 0.0011543 0.16546 0.00065855 0.16611 0.15179 0 0.036028 0.0389 0 0.91798 0.25917 0.070391 0.0097712 4.3493 0.060988 7.3472e-005 0.82909 0.0053704 0.006109 0.0014911 0.98557 0.9908 3.2296e-006 1.2919e-005 0.13266 0.79664 0.83241 0.0014516 0.88977 0.51545 0.0019535 0.42364 1.479 1.4763 16.009 144.9803 0.00029819 -85.2147 0.26795
1.372 0.98803 5.5171e-005 3.8182 0.012032 1.8052e-005 0.0011543 0.16551 0.00065855 0.16617 0.15184 0 0.036025 0.0389 0 0.91806 0.2592 0.070405 0.0097728 4.3497 0.060998 7.3485e-005 0.82908 0.0053708 0.0061095 0.0014903 0.98558 0.99081 3.2278e-006 1.2911e-005 0.13266 0.79722 0.8328 0.0014512 0.89044 0.51562 0.0019529 0.42365 1.4805 1.4778 16.009 144.9803 0.00029756 -85.2179 0.26895
1.373 0.98803 5.5171e-005 3.8182 0.012032 1.8065e-005 0.0011543 0.16557 0.00065855 0.16622 0.15189 0 0.036022 0.0389 0 0.91814 0.25924 0.070418 0.0097744 4.3502 0.061008 7.3498e-005 0.82907 0.0053713 0.0061099 0.0014896 0.98559 0.99082 3.226e-006 1.2904e-005 0.13267 0.7978 0.83318 0.0014508 0.89111 0.51578 0.0019524 0.42366 1.4819 1.4792 16.009 144.9803 0.00029694 -85.2211 0.26995
1.374 0.98803 5.5171e-005 3.8182 0.012032 1.8078e-005 0.0011543 0.16563 0.00065855 0.16628 0.15194 0 0.036018 0.0389 0 0.91822 0.25928 0.070431 0.009776 4.3506 0.061018 7.351e-005 0.82906 0.0053717 0.0061104 0.0014888 0.9856 0.99082 3.2242e-006 1.2897e-005 0.13267 0.79838 0.83357 0.0014504 0.89176 0.51595 0.0019519 0.42367 1.4833 1.4806 16.009 144.9803 0.00029632 -85.2242 0.27095
1.375 0.98803 5.5171e-005 3.8182 0.012032 1.8091e-005 0.0011543 0.16568 0.00065855 0.16634 0.152 0 0.036015 0.0389 0 0.91831 0.25932 0.070445 0.0097777 4.3511 0.061028 7.3523e-005 0.82905 0.0053722 0.0061108 0.001488 0.98561 0.99083 3.2224e-006 1.289e-005 0.13268 0.79896 0.83395 0.00145 0.89242 0.51612 0.0019514 0.42368 1.4847 1.482 16.0091 144.9804 0.00029571 -85.2274 0.27195
1.376 0.98803 5.5171e-005 3.8182 0.012032 1.8104e-005 0.0011543 0.16574 0.00065855 0.16639 0.15205 0 0.036011 0.0389 0 0.91839 0.25935 0.070458 0.0097793 4.3515 0.061038 7.3536e-005 0.82904 0.0053726 0.0061113 0.0014872 0.98562 0.99084 3.2206e-006 1.2883e-005 0.13268 0.79953 0.83433 0.0014496 0.89307 0.51628 0.0019509 0.42369 1.4861 1.4835 16.0091 144.9804 0.00029509 -85.2305 0.27295
1.377 0.98803 5.517e-005 3.8182 0.012032 1.8118e-005 0.0011543 0.16579 0.00065856 0.16645 0.1521 0 0.036008 0.0389 0 0.91847 0.25939 0.070472 0.0097809 4.352 0.061048 7.3549e-005 0.82903 0.0053731 0.0061117 0.0014865 0.98563 0.99084 3.2189e-006 1.2876e-005 0.13268 0.8001 0.83471 0.0014492 0.89372 0.51645 0.0019503 0.4237 1.4875 1.4849 16.0091 144.9804 0.00029448 -85.2336 0.27395
1.378 0.98803 5.517e-005 3.8182 0.012032 1.8131e-005 0.0011543 0.16585 0.00065856 0.1665 0.15215 0 0.036004 0.0389 0 0.91856 0.25943 0.070485 0.0097825 4.3524 0.061058 7.3562e-005 0.82902 0.0053735 0.0061122 0.0014857 0.98564 0.99085 3.2171e-006 1.2869e-005 0.13269 0.80068 0.83509 0.0014488 0.89437 0.51662 0.0019498 0.42371 1.4889 1.4863 16.0091 144.9804 0.00029387 -85.2366 0.27495
1.379 0.98803 5.517e-005 3.8182 0.012032 1.8144e-005 0.0011543 0.16591 0.00065856 0.16656 0.15221 0 0.036001 0.0389 0 0.91864 0.25946 0.070498 0.0097841 4.3529 0.061068 7.3575e-005 0.82901 0.005374 0.0061127 0.001485 0.98565 0.99086 3.2154e-006 1.2862e-005 0.13269 0.80124 0.83546 0.0014484 0.89501 0.51678 0.0019493 0.42372 1.4903 1.4877 16.0091 144.9804 0.00029327 -85.2396 0.27595
1.38 0.98803 5.517e-005 3.8182 0.012032 1.8157e-005 0.0011543 0.16596 0.00065856 0.16662 0.15226 0 0.035998 0.0389 0 0.91872 0.2595 0.070512 0.0097857 4.3533 0.061078 7.3588e-005 0.829 0.0053744 0.0061131 0.0014842 0.98566 0.99086 3.2137e-006 1.2855e-005 0.13269 0.80181 0.83583 0.001448 0.89564 0.51695 0.0019488 0.42373 1.4917 1.4891 16.0091 144.9805 0.00029267 -85.2427 0.27695
1.381 0.98803 5.517e-005 3.8182 0.012032 1.817e-005 0.0011543 0.16602 0.00065856 0.16667 0.15231 0 0.035994 0.0389 0 0.91881 0.25954 0.070525 0.0097874 4.3538 0.061088 7.3601e-005 0.82899 0.0053749 0.0061136 0.0014835 0.98567 0.99087 3.212e-006 1.2848e-005 0.1327 0.80238 0.83621 0.0014476 0.89628 0.51711 0.0019483 0.42374 1.4931 1.4905 16.0092 144.9805 0.00029207 -85.2457 0.27795
1.382 0.98803 5.517e-005 3.8182 0.012032 1.8183e-005 0.0011543 0.16607 0.00065856 0.16673 0.15236 0 0.035991 0.0389 0 0.91889 0.25958 0.070538 0.009789 4.3543 0.061098 7.3614e-005 0.82898 0.0053753 0.006114 0.0014827 0.98568 0.99088 3.2103e-006 1.2841e-005 0.1327 0.80294 0.83658 0.0014473 0.89691 0.51728 0.0019478 0.42375 1.4945 1.4919 16.0092 144.9805 0.00029147 -85.2486 0.27895
1.383 0.98803 5.517e-005 3.8182 0.012032 1.8196e-005 0.0011543 0.16613 0.00065856 0.16678 0.15242 0 0.035987 0.0389 0 0.91897 0.25961 0.070552 0.0097906 4.3547 0.061108 7.3627e-005 0.82897 0.0053758 0.0061145 0.001482 0.98569 0.99088 3.2086e-006 1.2835e-005 0.13271 0.8035 0.83694 0.0014469 0.89753 0.51744 0.0019474 0.42376 1.4959 1.4933 16.0092 144.9805 0.00029088 -85.2516 0.27995
1.384 0.98803 5.517e-005 3.8182 0.012032 1.8209e-005 0.0011543 0.16618 0.00065856 0.16684 0.15247 0 0.035984 0.0389 0 0.91906 0.25965 0.070565 0.0097922 4.3552 0.061118 7.364e-005 0.82896 0.0053762 0.0061149 0.0014813 0.9857 0.99089 3.207e-006 1.2828e-005 0.13271 0.80406 0.83731 0.0014465 0.89815 0.51761 0.0019469 0.42377 1.4973 1.4947 16.0092 144.9805 0.00029029 -85.2545 0.28095
1.385 0.98803 5.517e-005 3.8182 0.012031 1.8223e-005 0.0011543 0.16624 0.00065856 0.16689 0.15252 0 0.035981 0.0389 0 0.91914 0.25969 0.070579 0.0097938 4.3556 0.061128 7.3653e-005 0.82895 0.0053767 0.0061154 0.0014806 0.98571 0.9909 3.2053e-006 1.2821e-005 0.13271 0.80462 0.83768 0.0014461 0.89877 0.51778 0.0019464 0.42378 1.4987 1.4961 16.0092 144.9805 0.0002897 -85.2574 0.28195
1.386 0.98803 5.517e-005 3.8182 0.012031 1.8236e-005 0.0011543 0.1663 0.00065856 0.16695 0.15257 0 0.035977 0.0389 0 0.91922 0.25972 0.070592 0.0097954 4.3561 0.061138 7.3666e-005 0.82894 0.0053771 0.0061159 0.0014799 0.98572 0.9909 3.2037e-006 1.2815e-005 0.13272 0.80518 0.83804 0.0014458 0.89939 0.51794 0.0019459 0.42379 1.5 1.4974 16.0093 144.9806 0.00028911 -85.2603 0.28295
1.387 0.98803 5.517e-005 3.8182 0.012031 1.8249e-005 0.0011543 0.16635 0.00065856 0.16701 0.15263 0 0.035974 0.0389 0 0.91931 0.25976 0.070605 0.0097971 4.3565 0.061148 7.3679e-005 0.82893 0.0053776 0.0061163 0.0014792 0.98573 0.99091 3.2021e-006 1.2808e-005 0.13272 0.80573 0.8384 0.0014454 0.9 0.51811 0.0019454 0.4238 1.5014 1.4988 16.0093 144.9806 0.00028853 -85.2632 0.28395
1.388 0.98803 5.517e-005 3.8182 0.012031 1.8262e-005 0.0011543 0.16641 0.00065856 0.16706 0.15268 0 0.03597 0.0389 0 0.91939 0.2598 0.070619 0.0097987 4.357 0.061158 7.3692e-005 0.82892 0.005378 0.0061168 0.0014785 0.98574 0.99091 3.2004e-006 1.2802e-005 0.13272 0.80629 0.83876 0.0014451 0.9006 0.51827 0.001945 0.42381 1.5028 1.5002 16.0093 144.9806 0.00028795 -85.266 0.28495
1.389 0.98803 5.517e-005 3.8182 0.012031 1.8275e-005 0.0011543 0.16646 0.00065857 0.16712 0.15273 0 0.035967 0.0389 0 0.91947 0.25984 0.070632 0.0098003 4.3575 0.061168 7.3705e-005 0.82891 0.0053785 0.0061172 0.0014778 0.98575 0.99092 3.1988e-006 1.2795e-005 0.13273 0.80684 0.83912 0.0014447 0.90121 0.51844 0.0019445 0.42382 1.5041 1.5016 16.0093 144.9806 0.00028737 -85.2688 0.28595
1.39 0.98803 5.517e-005 3.8182 0.012031 1.8288e-005 0.0011543 0.16652 0.00065857 0.16717 0.15278 0 0.035964 0.0389 0 0.91956 0.25987 0.070645 0.0098019 4.3579 0.061178 7.3718e-005 0.8289 0.0053789 0.0061177 0.0014771 0.98576 0.99093 3.1973e-006 1.2789e-005 0.13273 0.80739 0.83948 0.0014444 0.90181 0.5186 0.001944 0.42383 1.5055 1.5029 16.0093 144.9806 0.00028679 -85.2716 0.28695
1.391 0.98803 5.517e-005 3.8182 0.012031 1.8301e-005 0.0011543 0.16657 0.00065857 0.16723 0.15283 0 0.03596 0.0389 0 0.91964 0.25991 0.070659 0.0098035 4.3584 0.061188 7.3731e-005 0.82889 0.0053794 0.0061182 0.0014764 0.98577 0.99093 3.1957e-006 1.2783e-005 0.13274 0.80794 0.83983 0.001444 0.9024 0.51877 0.0019436 0.42384 1.5068 1.5043 16.0093 144.9806 0.00028622 -85.2744 0.28795
1.392 0.98803 5.517e-005 3.8182 0.012031 1.8314e-005 0.0011543 0.16663 0.00065857 0.16728 0.15289 0 0.035957 0.0389 0 0.91972 0.25995 0.070672 0.0098052 4.3588 0.061198 7.3744e-005 0.82888 0.0053798 0.0061186 0.0014757 0.98578 0.99094 3.1941e-006 1.2777e-005 0.13274 0.80848 0.84019 0.0014437 0.903 0.51894 0.0019431 0.42385 1.5082 1.5057 16.0093 144.9807 0.00028565 -85.2772 0.28895
1.393 0.98803 5.5169e-005 3.8182 0.012031 1.8328e-005 0.0011543 0.16668 0.00065857 0.16734 0.15294 0 0.035953 0.0389 0 0.91981 0.25998 0.070686 0.0098068 4.3593 0.061208 7.3757e-005 0.82887 0.0053803 0.0061191 0.001475 0.98579 0.99094 3.1926e-006 1.277e-005 0.13274 0.80903 0.84054 0.0014433 0.90359 0.5191 0.0019427 0.42387 1.5095 1.507 16.0094 144.9807 0.00028508 -85.2799 0.28995
1.394 0.98803 5.5169e-005 3.8182 0.012031 1.8341e-005 0.0011543 0.16674 0.00065857 0.16739 0.15299 0 0.03595 0.0389 0 0.91989 0.26002 0.070699 0.0098084 4.3597 0.061218 7.377e-005 0.82886 0.0053807 0.0061195 0.0014744 0.98579 0.99095 3.191e-006 1.2764e-005 0.13275 0.80957 0.84089 0.001443 0.90417 0.51927 0.0019422 0.42388 1.5109 1.5084 16.0094 144.9807 0.00028452 -85.2826 0.29095
1.395 0.98803 5.5169e-005 3.8182 0.012031 1.8354e-005 0.0011543 0.16679 0.00065857 0.16745 0.15304 0 0.035947 0.0389 0 0.91997 0.26006 0.070713 0.00981 4.3602 0.061228 7.3783e-005 0.82885 0.0053812 0.00612 0.0014737 0.9858 0.99096 3.1895e-006 1.2758e-005 0.13275 0.81011 0.84124 0.0014426 0.90475 0.51943 0.0019418 0.42389 1.5122 1.5097 16.0094 144.9807 0.00028396 -85.2853 0.29195
1.396 0.98803 5.5169e-005 3.8182 0.012031 1.8367e-005 0.0011543 0.16685 0.00065857 0.1675 0.15309 0 0.035943 0.0389 0 0.92006 0.2601 0.070726 0.0098117 4.3607 0.061238 7.3796e-005 0.82884 0.0053816 0.0061205 0.001473 0.98581 0.99096 3.188e-006 1.2752e-005 0.13275 0.81065 0.84159 0.0014423 0.90533 0.5196 0.0019413 0.4239 1.5136 1.5111 16.0094 144.9807 0.0002834 -85.288 0.29295
1.397 0.98803 5.5169e-005 3.8182 0.012031 1.838e-005 0.0011543 0.1669 0.00065857 0.16756 0.15314 0 0.03594 0.0389 0 0.92014 0.26013 0.070739 0.0098133 4.3611 0.061248 7.3809e-005 0.82883 0.0053821 0.0061209 0.0014724 0.98582 0.99097 3.1865e-006 1.2746e-005 0.13276 0.81119 0.84193 0.0014419 0.90591 0.51976 0.0019409 0.42391 1.5149 1.5124 16.0094 144.9807 0.00028284 -85.2907 0.29395
1.398 0.98803 5.5169e-005 3.8182 0.012031 1.8393e-005 0.0011543 0.16696 0.00065857 0.16761 0.1532 0 0.035937 0.0389 0 0.92022 0.26017 0.070753 0.0098149 4.3616 0.061258 7.3822e-005 0.82882 0.0053826 0.0061214 0.0014717 0.98583 0.99097 3.185e-006 1.274e-005 0.13276 0.81173 0.84228 0.0014416 0.90648 0.51993 0.0019405 0.42392 1.5162 1.5138 16.0094 144.9808 0.00028228 -85.2933 0.29495
1.399 0.98803 5.5169e-005 3.8182 0.012031 1.8406e-005 0.0011543 0.16701 0.00065857 0.16767 0.15325 0 0.035933 0.0389 0 0.92031 0.26021 0.070766 0.0098165 4.3621 0.061268 7.3835e-005 0.82881 0.005383 0.0061218 0.0014711 0.98584 0.99098 3.1835e-006 1.2734e-005 0.13277 0.81226 0.84262 0.0014413 0.90705 0.52009 0.00194 0.42393 1.5175 1.5151 16.0095 144.9808 0.00028173 -85.2959 0.29595
1.4 0.98803 5.5169e-005 3.8182 0.012031 1.8419e-005 0.0011543 0.16707 0.00065857 0.16772 0.1533 0 0.03593 0.0389 0 0.92039 0.26024 0.07078 0.0098182 4.3625 0.061278 7.3848e-005 0.8288 0.0053835 0.0061223 0.0014704 0.98585 0.99098 3.1821e-006 1.2728e-005 0.13277 0.8128 0.84296 0.001441 0.90761 0.52026 0.0019396 0.42394 1.5189 1.5164 16.0095 144.9808 0.00028118 -85.2985 0.29695
1.401 0.98803 5.5169e-005 3.8182 0.012031 1.8433e-005 0.0011543 0.16712 0.00065858 0.16778 0.15335 0 0.035927 0.0389 0 0.92048 0.26028 0.070793 0.0098198 4.363 0.061289 7.3861e-005 0.82879 0.0053839 0.0061228 0.0014698 0.98585 0.99099 3.1806e-006 1.2722e-005 0.13277 0.81333 0.8433 0.0014406 0.90817 0.52042 0.0019392 0.42395 1.5202 1.5177 16.0095 144.9808 0.00028063 -85.3011 0.29795
1.402 0.98803 5.5169e-005 3.8182 0.012031 1.8446e-005 0.0011543 0.16718 0.00065858 0.16783 0.1534 0 0.035923 0.0389 0 0.92056 0.26032 0.070807 0.0098214 4.3634 0.061299 7.3874e-005 0.82878 0.0053844 0.0061232 0.0014692 0.98586 0.991 3.1792e-006 1.2717e-005 0.13278 0.81386 0.84364 0.0014403 0.90873 0.52059 0.0019387 0.42396 1.5215 1.5191 16.0095 144.9808 0.00028009 -85.3037 0.29895
1.403 0.98803 5.5169e-005 3.8182 0.012031 1.8459e-005 0.0011543 0.16723 0.00065858 0.16789 0.15345 0 0.03592 0.0389 0 0.92064 0.26036 0.07082 0.009823 4.3639 0.061309 7.3887e-005 0.82877 0.0053848 0.0061237 0.0014686 0.98587 0.991 3.1777e-006 1.2711e-005 0.13278 0.81439 0.84398 0.00144 0.90929 0.52075 0.0019383 0.42397 1.5228 1.5204 16.0095 144.9809 0.00027955 -85.3062 0.29995
1.404 0.98803 5.5169e-005 3.8182 0.012031 1.8472e-005 0.0011543 0.16729 0.00065858 0.16794 0.1535 0 0.035917 0.0389 0 0.92073 0.26039 0.070834 0.0098247 4.3644 0.061319 7.39e-005 0.82876 0.0053853 0.0061242 0.0014679 0.98588 0.99101 3.1763e-006 1.2705e-005 0.13278 0.81491 0.84431 0.0014397 0.90984 0.52092 0.0019379 0.42398 1.5241 1.5217 16.0095 144.9809 0.00027901 -85.3088 0.30095
1.405 0.98803 5.5169e-005 3.8182 0.012031 1.8485e-005 0.0011543 0.16734 0.00065858 0.168 0.15356 0 0.035913 0.0389 0 0.92081 0.26043 0.070847 0.0098263 4.3648 0.061329 7.3913e-005 0.82875 0.0053857 0.0061246 0.0014673 0.98589 0.99101 3.1749e-006 1.27e-005 0.13279 0.81544 0.84465 0.0014393 0.91039 0.52108 0.0019375 0.424 1.5254 1.523 16.0095 144.9809 0.00027847 -85.3113 0.30195
1.406 0.98803 5.5169e-005 3.8182 0.012031 1.8498e-005 0.0011543 0.1674 0.00065858 0.16805 0.15361 0 0.03591 0.0389 0 0.92089 0.26047 0.07086 0.0098279 4.3653 0.061339 7.3926e-005 0.82874 0.0053862 0.0061251 0.0014667 0.9859 0.99102 3.1735e-006 1.2694e-005 0.13279 0.81596 0.84498 0.001439 0.91093 0.52125 0.0019371 0.42401 1.5267 1.5243 16.0095 144.9809 0.00027793 -85.3138 0.30295
1.407 0.98803 5.5169e-005 3.8182 0.012031 1.8511e-005 0.0011543 0.16745 0.00065858 0.16811 0.15366 0 0.035907 0.0389 0 0.92098 0.26051 0.070874 0.0098295 4.3658 0.061349 7.3939e-005 0.82872 0.0053867 0.0061256 0.0014661 0.9859 0.99102 3.1721e-006 1.2688e-005 0.1328 0.81648 0.84531 0.0014387 0.91147 0.52141 0.0019367 0.42402 1.528 1.5256 16.0096 144.9809 0.0002774 -85.3163 0.30395
1.408 0.98803 5.5169e-005 3.8182 0.012031 1.8524e-005 0.0011543 0.16751 0.00065858 0.16816 0.15371 0 0.035903 0.0389 0 0.92106 0.26054 0.070887 0.0098312 4.3662 0.061359 7.3952e-005 0.82871 0.0053871 0.006126 0.0014655 0.98591 0.99103 3.1707e-006 1.2683e-005 0.1328 0.817 0.84564 0.0014384 0.91201 0.52158 0.0019363 0.42403 1.5293 1.5269 16.0096 144.9809 0.00027687 -85.3187 0.30495
1.409 0.98803 5.5168e-005 3.8182 0.012031 1.8538e-005 0.0011543 0.16756 0.00065858 0.16822 0.15376 0 0.0359 0.0389 0 0.92115 0.26058 0.070901 0.0098328 4.3667 0.061369 7.3965e-005 0.8287 0.0053876 0.0061265 0.0014649 0.98592 0.99103 3.1694e-006 1.2677e-005 0.1328 0.81752 0.84597 0.0014381 0.91255 0.52174 0.0019359 0.42404 1.5306 1.5282 16.0096 144.981 0.00027634 -85.3212 0.30595
1.41 0.98803 5.5168e-005 3.8182 0.012031 1.8551e-005 0.0011543 0.16762 0.00065858 0.16827 0.15381 0 0.035897 0.0389 0 0.92123 0.26062 0.070914 0.0098344 4.3672 0.061379 7.3978e-005 0.82869 0.005388 0.006127 0.0014643 0.98593 0.99104 3.168e-006 1.2672e-005 0.13281 0.81804 0.8463 0.0014378 0.91308 0.52191 0.0019355 0.42405 1.5319 1.5295 16.0096 144.981 0.00027582 -85.3236 0.30695
1.411 0.98803 5.5168e-005 3.8182 0.012031 1.8564e-005 0.0011543 0.16767 0.00065858 0.16832 0.15386 0 0.035893 0.0389 0 0.92131 0.26066 0.070928 0.009836 4.3676 0.061389 7.3991e-005 0.82868 0.0053885 0.0061274 0.0014637 0.98593 0.99104 3.1666e-006 1.2667e-005 0.13281 0.81856 0.84662 0.0014375 0.91361 0.52207 0.0019351 0.42406 1.5332 1.5308 16.0096 144.981 0.00027529 -85.326 0.30795
1.412 0.98803 5.5168e-005 3.8182 0.012031 1.8577e-005 0.0011543 0.16772 0.00065858 0.16838 0.15391 0 0.03589 0.0389 0 0.9214 0.26069 0.070941 0.0098377 4.3681 0.061399 7.4004e-005 0.82867 0.005389 0.0061279 0.0014631 0.98594 0.99105 3.1653e-006 1.2661e-005 0.13281 0.81907 0.84694 0.0014372 0.91413 0.52224 0.0019347 0.42407 1.5345 1.5321 16.0096 144.981 0.00027477 -85.3284 0.30895
1.413 0.98803 5.5168e-005 3.8182 0.012031 1.859e-005 0.0011543 0.16778 0.00065859 0.16843 0.15397 0 0.035887 0.0389 0 0.92148 0.26073 0.070955 0.0098393 4.3686 0.061409 7.4017e-005 0.82866 0.0053894 0.0061284 0.0014626 0.98595 0.99105 3.164e-006 1.2656e-005 0.13282 0.81958 0.84727 0.0014369 0.91466 0.5224 0.0019343 0.42408 1.5357 1.5334 16.0096 144.981 0.00027425 -85.3307 0.30995
1.414 0.98803 5.5168e-005 3.8182 0.012031 1.8603e-005 0.0011543 0.16783 0.00065859 0.16849 0.15402 0 0.035883 0.0389 0 0.92156 0.26077 0.070968 0.0098409 4.369 0.06142 7.403e-005 0.82865 0.0053899 0.0061288 0.001462 0.98596 0.99106 3.1627e-006 1.2651e-005 0.13282 0.82009 0.84759 0.0014366 0.91518 0.52256 0.0019339 0.4241 1.537 1.5347 16.0096 144.981 0.00027374 -85.3331 0.31095
1.415 0.98803 5.5168e-005 3.8182 0.012031 1.8616e-005 0.0011543 0.16789 0.00065859 0.16854 0.15407 0 0.03588 0.0389 0 0.92165 0.26081 0.070982 0.0098426 4.3695 0.06143 7.4043e-005 0.82864 0.0053903 0.0061293 0.0014614 0.98597 0.99106 3.1614e-006 1.2645e-005 0.13283 0.8206 0.84791 0.0014363 0.91569 0.52273 0.0019335 0.42411 1.5383 1.536 16.0097 144.9811 0.00027322 -85.3354 0.31195
1.416 0.98803 5.5168e-005 3.8182 0.012031 1.8629e-005 0.0011543 0.16794 0.00065859 0.1686 0.15412 0 0.035877 0.0389 0 0.92173 0.26084 0.070995 0.0098442 4.37 0.06144 7.4056e-005 0.82863 0.0053908 0.0061298 0.0014609 0.98597 0.99107 3.1601e-006 1.264e-005 0.13283 0.82111 0.84823 0.001436 0.91621 0.52289 0.0019331 0.42412 1.5396 1.5372 16.0097 144.9811 0.00027271 -85.3378 0.31295
1.417 0.98803 5.5168e-005 3.8182 0.012031 1.8643e-005 0.0011543 0.168 0.00065859 0.16865 0.15417 0 0.035873 0.0389 0 0.92182 0.26088 0.071009 0.0098458 4.3704 0.06145 7.4069e-005 0.82862 0.0053913 0.0061302 0.0014603 0.98598 0.99107 3.1588e-006 1.2635e-005 0.13283 0.82161 0.84854 0.0014357 0.91672 0.52306 0.0019328 0.42413 1.5408 1.5385 16.0097 144.9811 0.0002722 -85.3401 0.31395
1.418 0.98803 5.5168e-005 3.8182 0.012031 1.8656e-005 0.0011543 0.16805 0.00065859 0.1687 0.15422 0 0.03587 0.0389 0 0.9219 0.26092 0.071022 0.0098475 4.3709 0.06146 7.4083e-005 0.82861 0.0053917 0.0061307 0.0014598 0.98599 0.99108 3.1575e-006 1.263e-005 0.13284 0.82212 0.84886 0.0014354 0.91722 0.52322 0.0019324 0.42414 1.5421 1.5398 16.0097 144.9811 0.0002717 -85.3424 0.31495
1.419 0.98803 5.5168e-005 3.8182 0.012031 1.8669e-005 0.0011543 0.1681 0.00065859 0.16876 0.15427 0 0.035867 0.0389 0 0.92198 0.26095 0.071036 0.0098491 4.3714 0.06147 7.4096e-005 0.8286 0.0053922 0.0061312 0.0014592 0.98599 0.99108 3.1562e-006 1.2625e-005 0.13284 0.82262 0.84917 0.0014352 0.91773 0.52339 0.001932 0.42415 1.5433 1.541 16.0097 144.9811 0.00027119 -85.3446 0.31595
1.42 0.98803 5.5168e-005 3.8182 0.012031 1.8682e-005 0.0011543 0.16816 0.00065859 0.16881 0.15432 0 0.035864 0.0389 0 0.92207 0.26099 0.071049 0.0098507 4.3719 0.06148 7.4109e-005 0.82859 0.0053926 0.0061317 0.0014586 0.986 0.99109 3.155e-006 1.262e-005 0.13284 0.82312 0.84949 0.0014349 0.91823 0.52355 0.0019316 0.42416 1.5446 1.5423 16.0097 144.9812 0.00027069 -85.3469 0.31695
1.421 0.98803 5.5168e-005 3.8182 0.012031 1.8695e-005 0.0011543 0.16821 0.00065859 0.16887 0.15437 0 0.03586 0.0389 0 0.92215 0.26103 0.071063 0.0098524 4.3723 0.06149 7.4122e-005 0.82858 0.0053931 0.0061321 0.0014581 0.98601 0.99109 3.1537e-006 1.2615e-005 0.13285 0.82362 0.8498 0.0014346 0.91872 0.52371 0.0019313 0.42417 1.5458 1.5436 16.0097 144.9812 0.00027019 -85.3491 0.31795
1.422 0.98803 5.5168e-005 3.8182 0.012031 1.8708e-005 0.0011543 0.16827 0.00065859 0.16892 0.15442 0 0.035857 0.0389 0 0.92224 0.26107 0.071076 0.009854 4.3728 0.0615 7.4135e-005 0.82857 0.0053936 0.0061326 0.0014576 0.98602 0.9911 3.1525e-006 1.261e-005 0.13285 0.82412 0.85011 0.0014343 0.91922 0.52388 0.0019309 0.42419 1.5471 1.5448 16.0097 144.9812 0.00026969 -85.3513 0.31895
1.423 0.98803 5.5168e-005 3.8182 0.012031 1.8721e-005 0.0011543 0.16832 0.00065859 0.16897 0.15447 0 0.035854 0.0389 0 0.92232 0.2611 0.07109 0.0098556 4.3733 0.061511 7.4148e-005 0.82856 0.005394 0.0061331 0.001457 0.98602 0.9911 3.1512e-006 1.2605e-005 0.13286 0.82462 0.85042 0.001434 0.91971 0.52404 0.0019305 0.4242 1.5483 1.5461 16.0097 144.9812 0.00026919 -85.3535 0.31995
1.424 0.98803 5.5167e-005 3.8182 0.012031 1.8734e-005 0.0011543 0.16837 0.00065859 0.16903 0.15452 0 0.035851 0.0389 0 0.9224 0.26114 0.071103 0.0098573 4.3738 0.061521 7.4161e-005 0.82855 0.0053945 0.0061335 0.0014565 0.98603 0.99111 3.15e-006 1.26e-005 0.13286 0.82511 0.85072 0.0014338 0.9202 0.52421 0.0019302 0.42421 1.5496 1.5473 16.0097 144.9812 0.0002687 -85.3557 0.32095
1.425 0.98803 5.5167e-005 3.8182 0.012031 1.8748e-005 0.0011543 0.16843 0.0006586 0.16908 0.15458 0 0.035847 0.0389 0 0.92249 0.26118 0.071117 0.0098589 4.3742 0.061531 7.4174e-005 0.82854 0.005395 0.006134 0.001456 0.98604 0.99111 3.1488e-006 1.2595e-005 0.13286 0.82561 0.85103 0.0014335 0.92069 0.52437 0.0019298 0.42422 1.5508 1.5486 16.0098 144.9812 0.00026821 -85.3579 0.32195
1.426 0.98803 5.5167e-005 3.8182 0.012031 1.8761e-005 0.0011543 0.16848 0.0006586 0.16914 0.15463 0 0.035844 0.0389 0 0.92257 0.26122 0.071131 0.0098605 4.3747 0.061541 7.4187e-005 0.82853 0.0053954 0.0061345 0.0014555 0.98604 0.99112 3.1476e-006 1.259e-005 0.13287 0.8261 0.85134 0.0014332 0.92117 0.52454 0.0019295 0.42423 1.552 1.5498 16.0098 144.9813 0.00026772 -85.3601 0.32295
1.427 0.98803 5.5167e-005 3.8182 0.012031 1.8774e-005 0.0011543 0.16854 0.0006586 0.16919 0.15468 0 0.035841 0.0389 0 0.92266 0.26126 0.071144 0.0098622 4.3752 0.061551 7.42e-005 0.82852 0.0053959 0.006135 0.0014549 0.98605 0.99112 3.1464e-006 1.2586e-005 0.13287 0.82659 0.85164 0.0014329 0.92165 0.5247 0.0019291 0.42424 1.5533 1.551 16.0098 144.9813 0.00026723 -85.3622 0.32395
1.428 0.98803 5.5167e-005 3.8182 0.012031 1.8787e-005 0.0011543 0.16859 0.0006586 0.16924 0.15473 0 0.035837 0.0389 0 0.92274 0.26129 0.071158 0.0098638 4.3757 0.061561 7.4214e-005 0.82851 0.0053963 0.0061354 0.0014544 0.98606 0.99113 3.1452e-006 1.2581e-005 0.13288 0.82708 0.85194 0.0014327 0.92212 0.52486 0.0019288 0.42425 1.5545 1.5523 16.0098 144.9813 0.00026674 -85.3643 0.32495
1.429 0.98803 5.5167e-005 3.8182 0.012031 1.88e-005 0.0011543 0.16864 0.0006586 0.1693 0.15478 0 0.035834 0.0389 0 0.92283 0.26133 0.071171 0.0098654 4.3761 0.061571 7.4227e-005 0.8285 0.0053968 0.0061359 0.0014539 0.98606 0.99113 3.144e-006 1.2576e-005 0.13288 0.82756 0.85224 0.0014324 0.9226 0.52503 0.0019284 0.42427 1.5557 1.5535 16.0098 144.9813 0.00026626 -85.3665 0.32595
1.43 0.98803 5.5167e-005 3.8182 0.012031 1.8813e-005 0.0011543 0.1687 0.0006586 0.16935 0.15483 0 0.035831 0.0389 0 0.92291 0.26137 0.071185 0.0098671 4.3766 0.061581 7.424e-005 0.82849 0.0053973 0.0061364 0.0014534 0.98607 0.99113 3.1429e-006 1.2572e-005 0.13288 0.82805 0.85254 0.0014322 0.92307 0.52519 0.0019281 0.42428 1.5569 1.5547 16.0098 144.9813 0.00026578 -85.3686 0.32695
1.431 0.98803 5.5167e-005 3.8182 0.012031 1.8826e-005 0.0011543 0.16875 0.0006586 0.1694 0.15488 0 0.035828 0.0389 0 0.92299 0.26141 0.071198 0.0098687 4.3771 0.061592 7.4253e-005 0.82848 0.0053977 0.0061369 0.0014529 0.98608 0.99114 3.1417e-006 1.2567e-005 0.13289 0.82853 0.85284 0.0014319 0.92354 0.52535 0.0019277 0.42429 1.5582 1.556 16.0098 144.9814 0.0002653 -85.3706 0.32795
1.432 0.98803 5.5167e-005 3.8182 0.012031 1.8839e-005 0.0011543 0.1688 0.0006586 0.16946 0.15493 0 0.035824 0.0389 0 0.92308 0.26144 0.071212 0.0098703 4.3776 0.061602 7.4266e-005 0.82847 0.0053982 0.0061373 0.0014524 0.98608 0.99114 3.1406e-006 1.2562e-005 0.13289 0.82902 0.85314 0.0014316 0.924 0.52552 0.0019274 0.4243 1.5594 1.5572 16.0098 144.9814 0.00026483 -85.3727 0.32895
1.433 0.98803 5.5167e-005 3.8182 0.012031 1.8853e-005 0.0011543 0.16886 0.0006586 0.16951 0.15498 0 0.035821 0.0389 0 0.92316 0.26148 0.071225 0.009872 4.378 0.061612 7.4279e-005 0.82846 0.0053987 0.0061378 0.0014519 0.98609 0.99115 3.1394e-006 1.2558e-005 0.13289 0.8295 0.85343 0.0014314 0.92447 0.52568 0.0019271 0.42431 1.5606 1.5584 16.0098 144.9814 0.00026435 -85.3748 0.32995
1.434 0.98803 5.5167e-005 3.8182 0.012031 1.8866e-005 0.0011543 0.16891 0.0006586 0.16956 0.15503 0 0.035818 0.0389 0 0.92325 0.26152 0.071239 0.0098736 4.3785 0.061622 7.4292e-005 0.82845 0.0053991 0.0061383 0.0014514 0.9861 0.99115 3.1383e-006 1.2553e-005 0.1329 0.82998 0.85373 0.0014311 0.92493 0.52585 0.0019267 0.42432 1.5618 1.5596 16.0098 144.9814 0.00026388 -85.3768 0.33095
1.435 0.98803 5.5167e-005 3.8182 0.012031 1.8879e-005 0.0011543 0.16896 0.0006586 0.16962 0.15508 0 0.035815 0.0389 0 0.92333 0.26156 0.071253 0.0098752 4.379 0.061632 7.4305e-005 0.82844 0.0053996 0.0061388 0.0014509 0.9861 0.99116 3.1372e-006 1.2549e-005 0.1329 0.83046 0.85402 0.0014309 0.92538 0.52601 0.0019264 0.42433 1.563 1.5608 16.0098 144.9814 0.00026341 -85.3788 0.33195
1.436 0.98803 5.5167e-005 3.8182 0.012031 1.8892e-005 0.0011543 0.16902 0.0006586 0.16967 0.15513 0 0.035812 0.0389 0 0.92342 0.26159 0.071266 0.0098769 4.3795 0.061642 7.4319e-005 0.82843 0.0054001 0.0061392 0.0014504 0.98611 0.99116 3.1361e-006 1.2544e-005 0.13291 0.83093 0.85431 0.0014306 0.92584 0.52617 0.0019261 0.42435 1.5642 1.562 16.0098 144.9814 0.00026294 -85.3808 0.33295
1.437 0.98803 5.5167e-005 3.8182 0.012031 1.8905e-005 0.0011543 0.16907 0.00065861 0.16972 0.15518 0 0.035808 0.0389 0 0.9235 0.26163 0.07128 0.0098785 4.38 0.061652 7.4332e-005 0.82842 0.0054005 0.0061397 0.0014499 0.98612 0.99116 3.135e-006 1.254e-005 0.13291 0.83141 0.85461 0.0014304 0.92629 0.52634 0.0019257 0.42436 1.5654 1.5632 16.0098 144.9815 0.00026247 -85.3828 0.33395
1.438 0.98803 5.5167e-005 3.8182 0.012031 1.8918e-005 0.0011543 0.16912 0.00065861 0.16978 0.15523 0 0.035805 0.0389 0 0.92359 0.26167 0.071293 0.0098802 4.3804 0.061663 7.4345e-005 0.82841 0.005401 0.0061402 0.0014495 0.98612 0.99117 3.1339e-006 1.2535e-005 0.13291 0.83188 0.85489 0.0014301 0.92674 0.5265 0.0019254 0.42437 1.5666 1.5644 16.0099 144.9815 0.00026201 -85.3848 0.33495
1.439 0.98803 5.5167e-005 3.8182 0.012031 1.8931e-005 0.0011543 0.16918 0.00065861 0.16983 0.15528 0 0.035802 0.0389 0 0.92367 0.26171 0.071307 0.0098818 4.3809 0.061673 7.4358e-005 0.8284 0.0054015 0.0061407 0.001449 0.98613 0.99117 3.1328e-006 1.2531e-005 0.13292 0.83236 0.85518 0.0014299 0.92718 0.52666 0.0019251 0.42438 1.5678 1.5656 16.0099 144.9815 0.00026155 -85.3868 0.33595
1.44 0.98803 5.5166e-005 3.8182 0.012031 1.8944e-005 0.0011543 0.16923 0.00065861 0.16988 0.15533 0 0.035799 0.0389 0 0.92375 0.26174 0.07132 0.0098834 4.3814 0.061683 7.4371e-005 0.82839 0.0054019 0.0061411 0.0014485 0.98614 0.99118 3.1317e-006 1.2527e-005 0.13292 0.83283 0.85547 0.0014296 0.92762 0.52683 0.0019248 0.42439 1.569 1.5668 16.0099 144.9815 0.00026109 -85.3887 0.33695
1.441 0.98803 5.5166e-005 3.8182 0.012031 1.8958e-005 0.0011543 0.16928 0.00065861 0.16994 0.15538 0 0.035795 0.0389 0 0.92384 0.26178 0.071334 0.0098851 4.3819 0.061693 7.4384e-005 0.82838 0.0054024 0.0061416 0.001448 0.98614 0.99118 3.1306e-006 1.2522e-005 0.13293 0.8333 0.85576 0.0014294 0.92807 0.52699 0.0019245 0.4244 1.5701 1.568 16.0099 144.9815 0.00026063 -85.3907 0.33795
1.442 0.98803 5.5166e-005 3.8182 0.012031 1.8971e-005 0.0011543 0.16934 0.00065861 0.16999 0.15543 0 0.035792 0.0389 0 0.92392 0.26182 0.071348 0.0098867 4.3824 0.061703 7.4398e-005 0.82837 0.0054029 0.0061421 0.0014476 0.98615 0.99118 3.1295e-006 1.2518e-005 0.13293 0.83376 0.85604 0.0014291 0.9285 0.52715 0.0019242 0.42442 1.5713 1.5692 16.0099 144.9816 0.00026017 -85.3926 0.33895
1.443 0.98803 5.5166e-005 3.8182 0.012031 1.8984e-005 0.0011543 0.16939 0.00065861 0.17004 0.15548 0 0.035789 0.0389 0 0.92401 0.26186 0.071361 0.0098884 4.3828 0.061713 7.4411e-005 0.82836 0.0054034 0.0061426 0.0014471 0.98615 0.99119 3.1285e-006 1.2514e-005 0.13293 0.83423 0.85632 0.0014289 0.92894 0.52732 0.0019238 0.42443 1.5725 1.5704 16.0099 144.9816 0.00025972 -85.3945 0.33995
1.444 0.98803 5.5166e-005 3.8182 0.012031 1.8997e-005 0.0011543 0.16944 0.00065861 0.1701 0.15553 0 0.035786 0.0389 0 0.92409 0.2619 0.071375 0.00989 4.3833 0.061724 7.4424e-005 0.82835 0.0054038 0.006143 0.0014466 0.98616 0.99119 3.1274e-006 1.251e-005 0.13294 0.8347 0.85661 0.0014287 0.92937 0.52748 0.0019235 0.42444 1.5737 1.5716 16.0099 144.9816 0.00025926 -85.3964 0.34095
1.445 0.98803 5.5166e-005 3.8182 0.012031 1.901e-005 0.0011543 0.1695 0.00065861 0.17015 0.15558 0 0.035783 0.0389 0 0.92418 0.26193 0.071388 0.0098916 4.3838 0.061734 7.4437e-005 0.82834 0.0054043 0.0061435 0.0014462 0.98617 0.9912 3.1264e-006 1.2506e-005 0.13294 0.83516 0.85689 0.0014284 0.9298 0.52764 0.0019232 0.42445 1.5748 1.5727 16.0099 144.9816 0.00025881 -85.3983 0.34195
1.446 0.98803 5.5166e-005 3.8182 0.012031 1.9023e-005 0.0011543 0.16955 0.00065861 0.1702 0.15563 0 0.035779 0.0389 0 0.92426 0.26197 0.071402 0.0098933 4.3843 0.061744 7.445e-005 0.82833 0.0054048 0.006144 0.0014457 0.98617 0.9912 3.1253e-006 1.2501e-005 0.13295 0.83562 0.85717 0.0014282 0.93023 0.52781 0.0019229 0.42446 1.576 1.5739 16.0099 144.9816 0.00025837 -85.4002 0.34295
1.447 0.98803 5.5166e-005 3.8182 0.012031 1.9036e-005 0.0011543 0.1696 0.00065861 0.17026 0.15568 0 0.035776 0.0389 0 0.92435 0.26201 0.071416 0.0098949 4.3848 0.061754 7.4463e-005 0.82832 0.0054052 0.0061445 0.0014453 0.98618 0.9912 3.1243e-006 1.2497e-005 0.13295 0.83608 0.85745 0.001428 0.93065 0.52797 0.0019226 0.42447 1.5772 1.5751 16.0099 144.9816 0.00025792 -85.402 0.34395
1.448 0.98803 5.5166e-005 3.8182 0.012031 1.9049e-005 0.0011543 0.16965 0.00065861 0.17031 0.15573 0 0.035773 0.0389 0 0.92443 0.26205 0.071429 0.0098966 4.3853 0.061764 7.4477e-005 0.82831 0.0054057 0.006145 0.0014448 0.98618 0.99121 3.1233e-006 1.2493e-005 0.13295 0.83654 0.85773 0.0014277 0.93107 0.52813 0.0019223 0.42449 1.5783 1.5763 16.0099 144.9817 0.00025747 -85.4039 0.34495
1.449 0.98803 5.5166e-005 3.8182 0.012031 1.9063e-005 0.0011543 0.16971 0.00065862 0.17036 0.15578 0 0.03577 0.0389 0 0.92452 0.26208 0.071443 0.0098982 4.3857 0.061774 7.449e-005 0.8283 0.0054062 0.0061454 0.0014444 0.98619 0.99121 3.1223e-006 1.2489e-005 0.13296 0.837 0.858 0.0014275 0.93149 0.52829 0.001922 0.4245 1.5795 1.5774 16.0099 144.9817 0.00025703 -85.4057 0.34595
1.45 0.98803 5.5166e-005 3.8182 0.012031 1.9076e-005 0.0011543 0.16976 0.00065862 0.17041 0.15583 0 0.035767 0.0389 0 0.9246 0.26212 0.071457 0.0098998 4.3862 0.061785 7.4503e-005 0.82829 0.0054066 0.0061459 0.001444 0.98619 0.99122 3.1213e-006 1.2485e-005 0.13296 0.83746 0.85828 0.0014273 0.93191 0.52846 0.0019217 0.42451 1.5806 1.5786 16.0099 144.9817 0.00025659 -85.4075 0.34695
1.451 0.98803 5.5166e-005 3.8182 0.012031 1.9089e-005 0.0011543 0.16981 0.00065862 0.17047 0.15588 0 0.035763 0.0389 0 0.92468 0.26216 0.07147 0.0099015 4.3867 0.061795 7.4516e-005 0.82828 0.0054071 0.0061464 0.0014435 0.9862 0.99122 3.1203e-006 1.2481e-005 0.13296 0.83791 0.85855 0.0014271 0.93232 0.52862 0.0019214 0.42452 1.5818 1.5797 16.0099 144.9817 0.00025615 -85.4093 0.34795
1.452 0.98803 5.5166e-005 3.8182 0.012031 1.9102e-005 0.0011543 0.16987 0.00065862 0.17052 0.15593 0 0.03576 0.0389 0 0.92477 0.2622 0.071484 0.0099031 4.3872 0.061805 7.4529e-005 0.82827 0.0054076 0.0061469 0.0014431 0.98621 0.99122 3.1193e-006 1.2477e-005 0.13297 0.83837 0.85882 0.0014268 0.93274 0.52878 0.0019211 0.42453 1.5829 1.5809 16.0099 144.9817 0.00025571 -85.4111 0.34895
1.453 0.98803 5.5166e-005 3.8182 0.012031 1.9115e-005 0.0011543 0.16992 0.00065862 0.17057 0.15597 0 0.035757 0.0389 0 0.92485 0.26224 0.071497 0.0099048 4.3877 0.061815 7.4543e-005 0.82826 0.0054081 0.0061474 0.0014427 0.98621 0.99123 3.1183e-006 1.2473e-005 0.13297 0.83882 0.8591 0.0014266 0.93314 0.52895 0.0019208 0.42455 1.5841 1.5821 16.0099 144.9818 0.00025528 -85.4129 0.34995
1.454 0.98803 5.5166e-005 3.8182 0.012031 1.9128e-005 0.0011543 0.16997 0.00065862 0.17062 0.15602 0 0.035754 0.0389 0 0.92494 0.26227 0.071511 0.0099064 4.3882 0.061825 7.4556e-005 0.82825 0.0054085 0.0061479 0.0014422 0.98622 0.99123 3.1173e-006 1.2469e-005 0.13298 0.83927 0.85937 0.0014264 0.93355 0.52911 0.0019205 0.42456 1.5852 1.5832 16.0099 144.9818 0.00025485 -85.4147 0.35095
1.455 0.98803 5.5166e-005 3.8182 0.012031 1.9141e-005 0.0011543 0.17002 0.00065862 0.17068 0.15607 0 0.035751 0.0389 0 0.92502 0.26231 0.071525 0.0099081 4.3887 0.061836 7.4569e-005 0.82824 0.005409 0.0061483 0.0014418 0.98622 0.99123 3.1164e-006 1.2465e-005 0.13298 0.83972 0.85964 0.0014262 0.93395 0.52927 0.0019203 0.42457 1.5864 1.5843 16.0099 144.9818 0.00025441 -85.4164 0.35195
1.456 0.98803 5.5165e-005 3.8182 0.012031 1.9154e-005 0.0011543 0.17008 0.00065862 0.17073 0.15612 0 0.035747 0.0389 0 0.92511 0.26235 0.071538 0.0099097 4.3891 0.061846 7.4582e-005 0.82823 0.0054095 0.0061488 0.0014414 0.98623 0.99124 3.1154e-006 1.2462e-005 0.13298 0.84017 0.8599 0.0014259 0.93436 0.52943 0.00192 0.42458 1.5875 1.5855 16.01 144.9818 0.00025399 -85.4182 0.35295
1.457 0.98803 5.5165e-005 3.8182 0.012031 1.9168e-005 0.0011543 0.17013 0.00065862 0.17078 0.15617 0 0.035744 0.0389 0 0.92519 0.26239 0.071552 0.0099113 4.3896 0.061856 7.4595e-005 0.82822 0.00541 0.0061493 0.001441 0.98623 0.99124 3.1144e-006 1.2458e-005 0.13299 0.84061 0.86017 0.0014257 0.93476 0.5296 0.0019197 0.42459 1.5886 1.5866 16.01 144.9818 0.00025356 -85.4199 0.35395
1.458 0.98803 5.5165e-005 3.8182 0.012031 1.9181e-005 0.0011543 0.17018 0.00065862 0.17083 0.15622 0 0.035741 0.0389 0 0.92528 0.26242 0.071566 0.009913 4.3901 0.061866 7.4609e-005 0.82821 0.0054104 0.0061498 0.0014406 0.98624 0.99124 3.1135e-006 1.2454e-005 0.13299 0.84106 0.86044 0.0014255 0.93515 0.52976 0.0019194 0.42461 1.5898 1.5878 16.01 144.9819 0.00025313 -85.4216 0.35495
1.459 0.98803 5.5165e-005 3.8182 0.01203 1.9194e-005 0.0011543 0.17023 0.00065862 0.17089 0.15627 0 0.035738 0.0389 0 0.92536 0.26246 0.071579 0.0099146 4.3906 0.061876 7.4622e-005 0.8282 0.0054109 0.0061503 0.0014402 0.98624 0.99125 3.1126e-006 1.245e-005 0.133 0.8415 0.8607 0.0014253 0.93555 0.52992 0.0019191 0.42462 1.5909 1.5889 16.01 144.9819 0.00025271 -85.4233 0.35595
1.46 0.98803 5.5165e-005 3.8182 0.01203 1.9207e-005 0.0011543 0.17029 0.00065862 0.17094 0.15632 0 0.035735 0.0389 0 0.92545 0.2625 0.071593 0.0099163 4.3911 0.061887 7.4635e-005 0.82819 0.0054114 0.0061508 0.0014398 0.98625 0.99125 3.1116e-006 1.2447e-005 0.133 0.84195 0.86097 0.0014251 0.93594 0.53008 0.0019189 0.42463 1.592 1.59 16.01 144.9819 0.00025229 -85.425 0.35695
1.461 0.98803 5.5165e-005 3.8182 0.01203 1.922e-005 0.0011543 0.17034 0.00065862 0.17099 0.15637 0 0.035732 0.0389 0 0.92553 0.26254 0.071607 0.0099179 4.3916 0.061897 7.4648e-005 0.82818 0.0054119 0.0061512 0.0014394 0.98625 0.99126 3.1107e-006 1.2443e-005 0.133 0.84239 0.86123 0.0014249 0.93633 0.53025 0.0019186 0.42464 1.5932 1.5912 16.01 144.9819 0.00025187 -85.4267 0.35795
1.462 0.98803 5.5165e-005 3.8182 0.01203 1.9233e-005 0.0011543 0.17039 0.00065863 0.17104 0.15642 0 0.035729 0.0389 0 0.92562 0.26258 0.07162 0.0099196 4.3921 0.061907 7.4662e-005 0.82817 0.0054123 0.0061517 0.0014389 0.98626 0.99126 3.1098e-006 1.2439e-005 0.13301 0.84283 0.86149 0.0014247 0.93671 0.53041 0.0019183 0.42465 1.5943 1.5923 16.01 144.9819 0.00025145 -85.4284 0.35895
1.463 0.98803 5.5165e-005 3.8182 0.01203 1.9246e-005 0.0011543 0.17044 0.00065863 0.1711 0.15647 0 0.035725 0.0389 0 0.9257 0.26261 0.071634 0.0099212 4.3926 0.061917 7.4675e-005 0.82816 0.0054128 0.0061522 0.0014386 0.98627 0.99126 3.1089e-006 1.2435e-005 0.13301 0.84327 0.86175 0.0014245 0.9371 0.53057 0.001918 0.42467 1.5954 1.5934 16.01 144.9819 0.00025103 -85.43 0.35995
1.464 0.98803 5.5165e-005 3.8182 0.01203 1.9259e-005 0.0011543 0.17049 0.00065863 0.17115 0.15652 0 0.035722 0.0389 0 0.92579 0.26265 0.071648 0.0099229 4.3931 0.061927 7.4688e-005 0.82815 0.0054133 0.0061527 0.0014382 0.98627 0.99127 3.108e-006 1.2432e-005 0.13302 0.8437 0.86201 0.0014243 0.93748 0.53073 0.0019178 0.42468 1.5965 1.5945 16.01 144.982 0.00025062 -85.4317 0.36095
1.465 0.98803 5.5165e-005 3.8182 0.01203 1.9273e-005 0.0011543 0.17055 0.00065863 0.1712 0.15657 0 0.035719 0.0389 0 0.92587 0.26269 0.071661 0.0099245 4.3936 0.061938 7.4701e-005 0.82814 0.0054138 0.0061532 0.0014378 0.98628 0.99127 3.1071e-006 1.2428e-005 0.13302 0.84414 0.86227 0.0014241 0.93786 0.5309 0.0019175 0.42469 1.5976 1.5956 16.01 144.982 0.0002502 -85.4333 0.36195
1.466 0.98803 5.5165e-005 3.8182 0.01203 1.9286e-005 0.0011543 0.1706 0.00065863 0.17125 0.15661 0 0.035716 0.0389 0 0.92596 0.26273 0.071675 0.0099262 4.3941 0.061948 7.4715e-005 0.82813 0.0054142 0.0061537 0.0014374 0.98628 0.99127 3.1062e-006 1.2425e-005 0.13302 0.84457 0.86253 0.0014239 0.93824 0.53106 0.0019172 0.4247 1.5987 1.5968 16.01 144.982 0.00024979 -85.435 0.36295
1.467 0.98803 5.5165e-005 3.8182 0.01203 1.9299e-005 0.0011543 0.17065 0.00065863 0.1713 0.15666 0 0.035713 0.0389 0 0.92604 0.26277 0.071689 0.0099278 4.3945 0.061958 7.4728e-005 0.82812 0.0054147 0.0061542 0.001437 0.98629 0.99128 3.1053e-006 1.2421e-005 0.13303 0.84501 0.86279 0.0014237 0.93861 0.53122 0.001917 0.42471 1.5998 1.5979 16.01 144.982 0.00024938 -85.4366 0.36395
1.468 0.98803 5.5165e-005 3.8182 0.01203 1.9312e-005 0.0011543 0.1707 0.00065863 0.17136 0.15671 0 0.03571 0.0389 0 0.92613 0.2628 0.071702 0.0099295 4.395 0.061968 7.4741e-005 0.82811 0.0054152 0.0061546 0.0014366 0.98629 0.99128 3.1044e-006 1.2418e-005 0.13303 0.84544 0.86304 0.0014235 0.93899 0.53138 0.0019167 0.42473 1.6009 1.599 16.01 144.982 0.00024897 -85.4382 0.36495
1.469 0.98803 5.5165e-005 3.8182 0.01203 1.9325e-005 0.0011543 0.17075 0.00065863 0.17141 0.15676 0 0.035707 0.0389 0 0.92621 0.26284 0.071716 0.0099311 4.3955 0.061978 7.4754e-005 0.8281 0.0054157 0.0061551 0.0014362 0.9863 0.99128 3.1035e-006 1.2414e-005 0.13304 0.84587 0.8633 0.0014233 0.93936 0.53154 0.0019165 0.42474 1.602 1.6001 16.01 144.9821 0.00024857 -85.4398 0.36595
1.47 0.98803 5.5165e-005 3.8182 0.01203 1.9338e-005 0.0011543 0.17081 0.00065863 0.17146 0.15681 0 0.035703 0.0389 0 0.9263 0.26288 0.07173 0.0099328 4.396 0.061989 7.4768e-005 0.82809 0.0054161 0.0061556 0.0014358 0.9863 0.99129 3.1027e-006 1.2411e-005 0.13304 0.8463 0.86355 0.0014231 0.93972 0.53171 0.0019162 0.42475 1.6031 1.6012 16.01 144.9821 0.00024816 -85.4413 0.36695
1.471 0.98803 5.5165e-005 3.8182 0.01203 1.9351e-005 0.0011543 0.17086 0.00065863 0.17151 0.15686 0 0.0357 0.0389 0 0.92638 0.26292 0.071743 0.0099344 4.3965 0.061999 7.4781e-005 0.82808 0.0054166 0.0061561 0.0014355 0.98631 0.99129 3.1018e-006 1.2407e-005 0.13304 0.84673 0.8638 0.0014229 0.94009 0.53187 0.0019159 0.42476 1.6042 1.6023 16.01 144.9821 0.00024776 -85.4429 0.36795
1.472 0.98803 5.5164e-005 3.8182 0.01203 1.9364e-005 0.0011543 0.17091 0.00065863 0.17156 0.15691 0 0.035697 0.0389 0 0.92647 0.26296 0.071757 0.0099361 4.397 0.062009 7.4794e-005 0.82807 0.0054171 0.0061566 0.0014351 0.98631 0.99129 3.1009e-006 1.2404e-005 0.13305 0.84715 0.86405 0.0014227 0.94045 0.53203 0.0019157 0.42477 1.6053 1.6034 16.01 144.9821 0.00024736 -85.4445 0.36895
1.473 0.98803 5.5164e-005 3.8182 0.01203 1.9378e-005 0.0011543 0.17096 0.00065863 0.17162 0.15696 0 0.035694 0.0389 0 0.92655 0.26299 0.071771 0.0099377 4.3975 0.062019 7.4807e-005 0.82806 0.0054176 0.0061571 0.0014347 0.98632 0.99129 3.1001e-006 1.24e-005 0.13305 0.84758 0.8643 0.0014225 0.94081 0.53219 0.0019154 0.42479 1.6064 1.6045 16.01 144.9821 0.00024696 -85.446 0.36995
1.474 0.98803 5.5164e-005 3.8182 0.01203 1.9391e-005 0.0011543 0.17101 0.00065863 0.17167 0.157 0 0.035691 0.0389 0 0.92664 0.26303 0.071785 0.0099394 4.398 0.06203 7.4821e-005 0.82805 0.0054181 0.0061576 0.0014344 0.98632 0.9913 3.0993e-006 1.2397e-005 0.13306 0.848 0.86455 0.0014223 0.94117 0.53235 0.0019152 0.4248 1.6075 1.6055 16.01 144.9822 0.00024656 -85.4475 0.37095
1.475 0.98803 5.5164e-005 3.8182 0.01203 1.9404e-005 0.0011543 0.17107 0.00065864 0.17172 0.15705 0 0.035688 0.0389 0 0.92672 0.26307 0.071798 0.009941 4.3985 0.06204 7.4834e-005 0.82803 0.0054185 0.0061581 0.001434 0.98632 0.9913 3.0984e-006 1.2394e-005 0.13306 0.84842 0.8648 0.0014221 0.94153 0.53251 0.0019149 0.42481 1.6085 1.6066 16.01 144.9822 0.00024617 -85.4491 0.37195
1.476 0.98803 5.5164e-005 3.8182 0.01203 1.9417e-005 0.0011543 0.17112 0.00065864 0.17177 0.1571 0 0.035685 0.0389 0 0.92681 0.26311 0.071812 0.0099427 4.399 0.06205 7.4847e-005 0.82802 0.005419 0.0061585 0.0014336 0.98633 0.9913 3.0976e-006 1.239e-005 0.13306 0.84885 0.86505 0.0014219 0.94189 0.53268 0.0019147 0.42482 1.6096 1.6077 16.01 144.9822 0.00024577 -85.4506 0.37295
1.477 0.98803 5.5164e-005 3.8182 0.01203 1.943e-005 0.0011543 0.17117 0.00065864 0.17182 0.15715 0 0.035682 0.0389 0 0.92689 0.26315 0.071826 0.0099443 4.3995 0.06206 7.486e-005 0.82801 0.0054195 0.006159 0.0014333 0.98633 0.99131 3.0968e-006 1.2387e-005 0.13307 0.84926 0.86529 0.0014217 0.94224 0.53284 0.0019144 0.42484 1.6107 1.6088 16.01 144.9822 0.00024538 -85.4521 0.37395
1.478 0.98803 5.5164e-005 3.8182 0.01203 1.9443e-005 0.0011543 0.17122 0.00065864 0.17187 0.1572 0 0.035678 0.0389 0 0.92698 0.26318 0.071839 0.009946 4.4 0.062071 7.4874e-005 0.828 0.00542 0.0061595 0.0014329 0.98634 0.99131 3.0959e-006 1.2384e-005 0.13307 0.84968 0.86554 0.0014215 0.94259 0.533 0.0019142 0.42485 1.6118 1.6099 16.01 144.9822 0.00024499 -85.4536 0.37495
1.479 0.98803 5.5164e-005 3.8182 0.01203 1.9456e-005 0.0011543 0.17127 0.00065864 0.17193 0.15725 0 0.035675 0.0389 0 0.92707 0.26322 0.071853 0.0099476 4.4005 0.062081 7.4887e-005 0.82799 0.0054205 0.00616 0.0014326 0.98634 0.99131 3.0951e-006 1.2381e-005 0.13308 0.8501 0.86578 0.0014214 0.94294 0.53316 0.001914 0.42486 1.6128 1.6109 16.01 144.9822 0.0002446 -85.4551 0.37595
1.48 0.98803 5.5164e-005 3.8182 0.01203 1.9469e-005 0.0011543 0.17132 0.00065864 0.17198 0.1573 0 0.035672 0.0389 0 0.92715 0.26326 0.071867 0.0099493 4.401 0.062091 7.49e-005 0.82798 0.0054209 0.0061605 0.0014322 0.98635 0.99132 3.0943e-006 1.2377e-005 0.13308 0.85052 0.86603 0.0014212 0.94328 0.53332 0.0019137 0.42487 1.6139 1.612 16.01 144.9823 0.00024421 -85.4565 0.37695
1.481 0.98803 5.5164e-005 3.8182 0.01203 1.9483e-005 0.0011543 0.17137 0.00065864 0.17203 0.15734 0 0.035669 0.0389 0 0.92724 0.2633 0.071881 0.0099509 4.4015 0.062101 7.4914e-005 0.82797 0.0054214 0.006161 0.0014319 0.98635 0.99132 3.0935e-006 1.2374e-005 0.13308 0.85093 0.86627 0.001421 0.94363 0.53348 0.0019135 0.42488 1.6149 1.6131 16.01 144.9823 0.00024383 -85.458 0.37795
1.482 0.98803 5.5164e-005 3.8182 0.01203 1.9496e-005 0.0011543 0.17143 0.00065864 0.17208 0.15739 0 0.035666 0.0389 0 0.92732 0.26334 0.071894 0.0099526 4.402 0.062112 7.4927e-005 0.82796 0.0054219 0.0061615 0.0014315 0.98636 0.99132 3.0927e-006 1.2371e-005 0.13309 0.85134 0.86651 0.0014208 0.94397 0.53365 0.0019133 0.4249 1.616 1.6142 16.01 144.9823 0.00024344 -85.4594 0.37895
1.483 0.98803 5.5164e-005 3.8182 0.01203 1.9509e-005 0.0011543 0.17148 0.00065864 0.17213 0.15744 0 0.035663 0.0389 0 0.92741 0.26337 0.071908 0.0099542 4.4025 0.062122 7.494e-005 0.82795 0.0054224 0.006162 0.0014312 0.98636 0.99133 3.0919e-006 1.2368e-005 0.13309 0.85176 0.86675 0.0014206 0.94431 0.53381 0.001913 0.42491 1.6171 1.6152 16.01 144.9823 0.00024306 -85.4609 0.37995
1.484 0.98803 5.5164e-005 3.8182 0.01203 1.9522e-005 0.0011543 0.17153 0.00065864 0.17218 0.15749 0 0.03566 0.0389 0 0.92749 0.26341 0.071922 0.0099559 4.403 0.062132 7.4954e-005 0.82794 0.0054229 0.0061625 0.0014308 0.98637 0.99133 3.0912e-006 1.2365e-005 0.1331 0.85217 0.86699 0.0014205 0.94464 0.53397 0.0019128 0.42492 1.6181 1.6163 16.01 144.9823 0.00024268 -85.4623 0.38095
1.485 0.98803 5.5164e-005 3.8182 0.01203 1.9535e-005 0.0011543 0.17158 0.00065864 0.17223 0.15754 0 0.035657 0.0389 0 0.92758 0.26345 0.071936 0.0099575 4.4035 0.062142 7.4967e-005 0.82793 0.0054233 0.006163 0.0014305 0.98637 0.99133 3.0904e-006 1.2362e-005 0.1331 0.85258 0.86723 0.0014203 0.94498 0.53413 0.0019126 0.42493 1.6192 1.6173 16.01 144.9824 0.0002423 -85.4637 0.38195
1.486 0.98803 5.5164e-005 3.8182 0.01203 1.9548e-005 0.0011543 0.17163 0.00065864 0.17229 0.15758 0 0.035654 0.0389 0 0.92766 0.26349 0.071949 0.0099592 4.404 0.062153 7.498e-005 0.82792 0.0054238 0.0061635 0.0014302 0.98638 0.99133 3.0896e-006 1.2358e-005 0.1331 0.85299 0.86746 0.0014201 0.94531 0.53429 0.0019123 0.42495 1.6202 1.6184 16.01 144.9824 0.00024192 -85.4651 0.38295
1.487 0.98803 5.5163e-005 3.8182 0.01203 1.9561e-005 0.0011543 0.17168 0.00065864 0.17234 0.15763 0 0.035651 0.0389 0 0.92775 0.26353 0.071963 0.0099608 4.4045 0.062163 7.4993e-005 0.82791 0.0054243 0.006164 0.0014298 0.98638 0.99134 3.0889e-006 1.2355e-005 0.13311 0.85339 0.8677 0.0014199 0.94564 0.53445 0.0019121 0.42496 1.6213 1.6194 16.01 144.9824 0.00024154 -85.4665 0.38395
1.488 0.98803 5.5163e-005 3.8182 0.01203 1.9574e-005 0.0011543 0.17173 0.00065864 0.17239 0.15768 0 0.035648 0.0389 0 0.92783 0.26357 0.071977 0.0099625 4.405 0.062173 7.5007e-005 0.8279 0.0054248 0.0061644 0.0014295 0.98638 0.99134 3.0881e-006 1.2352e-005 0.13311 0.8538 0.86793 0.0014198 0.94597 0.53461 0.0019119 0.42497 1.6223 1.6205 16.01 144.9824 0.00024117 -85.4679 0.38495
1.489 0.98803 5.5163e-005 3.8182 0.01203 1.9587e-005 0.0011543 0.17178 0.00065865 0.17244 0.15773 0 0.035645 0.0389 0 0.92792 0.2636 0.071991 0.0099642 4.4055 0.062184 7.502e-005 0.82789 0.0054253 0.0061649 0.0014292 0.98639 0.99134 3.0873e-006 1.2349e-005 0.13312 0.8542 0.86817 0.0014196 0.9463 0.53477 0.0019116 0.42498 1.6233 1.6215 16.01 144.9824 0.0002408 -85.4693 0.38595
1.49 0.98803 5.5163e-005 3.8182 0.01203 1.9601e-005 0.0011543 0.17184 0.00065865 0.17249 0.15778 0 0.035641 0.0389 0 0.92801 0.26364 0.072004 0.0099658 4.406 0.062194 7.5033e-005 0.82788 0.0054258 0.0061654 0.0014288 0.98639 0.99135 3.0866e-006 1.2346e-005 0.13312 0.85461 0.8684 0.0014194 0.94662 0.53493 0.0019114 0.42499 1.6244 1.6226 16.01 144.9825 0.00024042 -85.4707 0.38695
1.491 0.98803 5.5163e-005 3.8182 0.01203 1.9614e-005 0.0011543 0.17189 0.00065865 0.17254 0.15783 0 0.035638 0.0389 0 0.92809 0.26368 0.072018 0.0099675 4.4065 0.062204 7.5047e-005 0.82787 0.0054263 0.0061659 0.0014285 0.9864 0.99135 3.0858e-006 1.2343e-005 0.13312 0.85501 0.86863 0.0014192 0.94695 0.5351 0.0019112 0.42501 1.6254 1.6236 16.01 144.9825 0.00024005 -85.4721 0.38795
1.492 0.98803 5.5163e-005 3.8182 0.01203 1.9627e-005 0.0011543 0.17194 0.00065865 0.17259 0.15787 0 0.035635 0.0389 0 0.92818 0.26372 0.072032 0.0099691 4.407 0.062214 7.506e-005 0.82786 0.0054267 0.0061664 0.0014282 0.9864 0.99135 3.0851e-006 1.234e-005 0.13313 0.85541 0.86887 0.0014191 0.94727 0.53526 0.001911 0.42502 1.6264 1.6246 16.01 144.9825 0.00023968 -85.4734 0.38895
1.493 0.98803 5.5163e-005 3.8182 0.01203 1.964e-005 0.0011543 0.17199 0.00065865 0.17264 0.15792 0 0.035632 0.0389 0 0.92826 0.26376 0.072046 0.0099708 4.4075 0.062225 7.5073e-005 0.82785 0.0054272 0.0061669 0.0014279 0.9864 0.99135 3.0844e-006 1.2337e-005 0.13313 0.85581 0.8691 0.0014189 0.94759 0.53542 0.0019108 0.42503 1.6275 1.6257 16.01 144.9825 0.00023932 -85.4747 0.38995
1.494 0.98803 5.5163e-005 3.8182 0.01203 1.9653e-005 0.0011543 0.17204 0.00065865 0.17269 0.15797 0 0.035629 0.0389 0 0.92835 0.26379 0.07206 0.0099724 4.408 0.062235 7.5087e-005 0.82784 0.0054277 0.0061674 0.0014276 0.98641 0.99136 3.0836e-006 1.2335e-005 0.13314 0.85621 0.86933 0.0014187 0.9479 0.53558 0.0019105 0.42504 1.6285 1.6267 16.01 144.9825 0.00023895 -85.4761 0.39095
1.495 0.98803 5.5163e-005 3.8182 0.01203 1.9666e-005 0.0011543 0.17209 0.00065865 0.17274 0.15802 0 0.035626 0.0389 0 0.92843 0.26383 0.072073 0.0099741 4.4085 0.062245 7.51e-005 0.82783 0.0054282 0.0061679 0.0014272 0.98641 0.99136 3.0829e-006 1.2332e-005 0.13314 0.8566 0.86955 0.0014186 0.94822 0.53574 0.0019103 0.42506 1.6295 1.6277 16.01 144.9826 0.00023859 -85.4774 0.39195
1.496 0.98803 5.5163e-005 3.8182 0.01203 1.9679e-005 0.0011543 0.17214 0.00065865 0.1728 0.15806 0 0.035623 0.0389 0 0.92852 0.26387 0.072087 0.0099757 4.409 0.062255 7.5113e-005 0.82782 0.0054287 0.0061684 0.0014269 0.98642 0.99136 3.0822e-006 1.2329e-005 0.13314 0.857 0.86978 0.0014184 0.94853 0.5359 0.0019101 0.42507 1.6305 1.6288 16.01 144.9826 0.00023823 -85.4787 0.39295
1.497 0.98803 5.5163e-005 3.8182 0.01203 1.9692e-005 0.0011543 0.17219 0.00065865 0.17285 0.15811 0 0.03562 0.0389 0 0.9286 0.26391 0.072101 0.0099774 4.4096 0.062266 7.5127e-005 0.82781 0.0054292 0.0061689 0.0014266 0.98642 0.99136 3.0815e-006 1.2326e-005 0.13315 0.85739 0.87001 0.0014183 0.94884 0.53606 0.0019099 0.42508 1.6316 1.6298 16.01 144.9826 0.00023787 -85.48 0.39395
1.498 0.98803 5.5163e-005 3.8182 0.01203 1.9706e-005 0.0011543 0.17224 0.00065865 0.1729 0.15816 0 0.035617 0.0389 0 0.92869 0.26395 0.072115 0.0099791 4.4101 0.062276 7.514e-005 0.8278 0.0054297 0.0061694 0.0014263 0.98643 0.99137 3.0808e-006 1.2323e-005 0.13315 0.85779 0.87024 0.0014181 0.94915 0.53622 0.0019097 0.42509 1.6326 1.6308 16.01 144.9826 0.00023751 -85.4813 0.39495
1.499 0.98803 5.5163e-005 3.8182 0.01203 1.9719e-005 0.0011543 0.17229 0.00065865 0.17295 0.15821 0 0.035614 0.0389 0 0.92878 0.26399 0.072128 0.0099807 4.4106 0.062286 7.5153e-005 0.82779 0.0054301 0.0061699 0.001426 0.98643 0.99137 3.0801e-006 1.232e-005 0.13316 0.85818 0.87046 0.0014179 0.94946 0.53638 0.0019095 0.42511 1.6336 1.6318 16.01 144.9826 0.00023715 -85.4826 0.39595
1.5 0.98803 5.5163e-005 3.8182 0.01203 1.9732e-005 0.0011543 0.17234 0.00065865 0.173 0.15826 0 0.035611 0.0389 0 0.92886 0.26402 0.072142 0.0099824 4.4111 0.062297 7.5167e-005 0.82778 0.0054306 0.0061704 0.0014257 0.98643 0.99137 3.0794e-006 1.2318e-005 0.13316 0.85857 0.87068 0.0014178 0.94976 0.53654 0.0019093 0.42512 1.6346 1.6328 16.01 144.9826 0.00023679 -85.4839 0.39695
1.501 0.98803 5.5163e-005 3.8182 0.01203 1.9745e-005 0.0011543 0.1724 0.00065865 0.17305 0.1583 0 0.035608 0.0389 0 0.92895 0.26406 0.072156 0.009984 4.4116 0.062307 7.518e-005 0.82777 0.0054311 0.0061709 0.0014254 0.98644 0.99137 3.0787e-006 1.2315e-005 0.13316 0.85896 0.87091 0.0014176 0.95007 0.5367 0.0019091 0.42513 1.6356 1.6339 16.01 144.9827 0.00023644 -85.4852 0.39795
1.502 0.98803 5.5163e-005 3.8182 0.01203 1.9758e-005 0.0011543 0.17245 0.00065866 0.1731 0.15835 0 0.035605 0.0389 0 0.92903 0.2641 0.07217 0.0099857 4.4121 0.062317 7.5194e-005 0.82776 0.0054316 0.0061714 0.0014251 0.98644 0.99138 3.078e-006 1.2312e-005 0.13317 0.85935 0.87113 0.0014175 0.95037 0.53686 0.0019089 0.42514 1.6366 1.6349 16.01 144.9827 0.00023608 -85.4864 0.39895
1.503 0.98803 5.5162e-005 3.8182 0.01203 1.9771e-005 0.0011543 0.1725 0.00065866 0.17315 0.1584 0 0.035602 0.0389 0 0.92912 0.26414 0.072184 0.0099874 4.4126 0.062328 7.5207e-005 0.82775 0.0054321 0.0061719 0.0014248 0.98644 0.99138 3.0773e-006 1.2309e-005 0.13317 0.85974 0.87135 0.0014173 0.95067 0.53702 0.0019087 0.42516 1.6376 1.6359 16.01 144.9827 0.00023573 -85.4877 0.39995
1.504 0.98803 5.5162e-005 3.8182 0.01203 1.9784e-005 0.0011543 0.17255 0.00065866 0.1732 0.15845 0 0.035599 0.0389 0 0.9292 0.26418 0.072197 0.009989 4.4131 0.062338 7.522e-005 0.82774 0.0054326 0.0061724 0.0014245 0.98645 0.99138 3.0766e-006 1.2307e-005 0.13318 0.86012 0.87157 0.0014171 0.95096 0.53718 0.0019085 0.42517 1.6386 1.6369 16.01 144.9827 0.00023538 -85.4889 0.40095
1.505 0.98803 5.5162e-005 3.8182 0.01203 1.9797e-005 0.0011543 0.1726 0.00065866 0.17325 0.15849 0 0.035596 0.0389 0 0.92929 0.26422 0.072211 0.0099907 4.4136 0.062348 7.5234e-005 0.82773 0.0054331 0.0061729 0.0014242 0.98645 0.99138 3.076e-006 1.2304e-005 0.13318 0.86051 0.87179 0.001417 0.95126 0.53734 0.0019083 0.42518 1.6396 1.6379 16.01 144.9827 0.00023503 -85.4902 0.40195
1.506 0.98803 5.5162e-005 3.8182 0.01203 1.9811e-005 0.0011543 0.17265 0.00065866 0.1733 0.15854 0 0.035593 0.0389 0 0.92938 0.26425 0.072225 0.0099923 4.4141 0.062358 7.5247e-005 0.82772 0.0054336 0.0061734 0.0014239 0.98646 0.99139 3.0753e-006 1.2301e-005 0.13318 0.86089 0.87201 0.0014168 0.95155 0.5375 0.0019081 0.42519 1.6406 1.6389 16.01 144.9828 0.00023468 -85.4914 0.40295
1.507 0.98803 5.5162e-005 3.8182 0.01203 1.9824e-005 0.0011543 0.1727 0.00065866 0.17335 0.15859 0 0.03559 0.0389 0 0.92946 0.26429 0.072239 0.009994 4.4146 0.062369 7.526e-005 0.82771 0.005434 0.0061739 0.0014236 0.98646 0.99139 3.0746e-006 1.2299e-005 0.13319 0.86127 0.87223 0.0014167 0.95185 0.53766 0.0019079 0.42521 1.6416 1.6399 16.01 144.9828 0.00023434 -85.4926 0.40395
1.508 0.98803 5.5162e-005 3.8182 0.01203 1.9837e-005 0.0011543 0.17275 0.00065866 0.1734 0.15864 0 0.035587 0.0389 0 0.92955 0.26433 0.072253 0.0099957 4.4152 0.062379 7.5274e-005 0.8277 0.0054345 0.0061744 0.0014233 0.98646 0.99139 3.074e-006 1.2296e-005 0.13319 0.86165 0.87244 0.0014165 0.95214 0.53782 0.0019077 0.42522 1.6426 1.6409 16.01 144.9828 0.00023399 -85.4938 0.40495
1.509 0.98803 5.5162e-005 3.8182 0.01203 1.985e-005 0.0011543 0.1728 0.00065866 0.17345 0.15868 0 0.035584 0.0389 0 0.92963 0.26437 0.072267 0.0099973 4.4157 0.062389 7.5287e-005 0.82769 0.005435 0.0061749 0.0014231 0.98647 0.99139 3.0733e-006 1.2293e-005 0.1332 0.86203 0.87266 0.0014164 0.95242 0.53798 0.0019075 0.42523 1.6436 1.6419 16.01 144.9828 0.00023365 -85.495 0.40595
1.51 0.98803 5.5162e-005 3.8182 0.01203 1.9863e-005 0.0011543 0.17285 0.00065866 0.1735 0.15873 0 0.035581 0.0389 0 0.92972 0.26441 0.07228 0.009999 4.4162 0.0624 7.5301e-005 0.82768 0.0054355 0.0061754 0.0014228 0.98647 0.9914 3.0727e-006 1.2291e-005 0.1332 0.86241 0.87288 0.0014162 0.95271 0.53814 0.0019073 0.42524 1.6445 1.6428 16.01 144.9828 0.00023331 -85.4962 0.40695
1.511 0.98803 5.5162e-005 3.8182 0.01203 1.9876e-005 0.0011543 0.1729 0.00065866 0.17355 0.15878 0 0.035578 0.0389 0 0.92981 0.26445 0.072294 0.010001 4.4167 0.06241 7.5314e-005 0.82767 0.005436 0.0061759 0.0014225 0.98647 0.9914 3.072e-006 1.2288e-005 0.1332 0.86279 0.87309 0.0014161 0.953 0.5383 0.0019071 0.42526 1.6455 1.6438 16.0099 144.9829 0.00023297 -85.4974 0.40795
1.512 0.98803 5.5162e-005 3.8182 0.01203 1.9889e-005 0.0011543 0.17295 0.00065866 0.1736 0.15882 0 0.035575 0.0389 0 0.92989 0.26448 0.072308 0.010002 4.4172 0.06242 7.5327e-005 0.82765 0.0054365 0.0061764 0.0014222 0.98648 0.9914 3.0714e-006 1.2286e-005 0.13321 0.86317 0.8733 0.001416 0.95328 0.53846 0.0019069 0.42527 1.6465 1.6448 16.0099 144.9829 0.00023263 -85.4986 0.40895
1.513 0.98803 5.5162e-005 3.8182 0.01203 1.9902e-005 0.0011543 0.173 0.00065866 0.17365 0.15887 0 0.035572 0.0389 0 0.92998 0.26452 0.072322 0.010004 4.4177 0.062431 7.5341e-005 0.82764 0.005437 0.0061769 0.0014219 0.98648 0.9914 3.0708e-006 1.2283e-005 0.13321 0.86354 0.87352 0.0014158 0.95356 0.53862 0.0019067 0.42528 1.6475 1.6458 16.0099 144.9829 0.00023229 -85.4997 0.40995
1.514 0.98803 5.5162e-005 3.8182 0.01203 1.9916e-005 0.0011544 0.17305 0.00065866 0.1737 0.15892 0 0.035569 0.0389 0 0.93006 0.26456 0.072336 0.010006 4.4182 0.062441 7.5354e-005 0.82763 0.0054375 0.0061774 0.0014217 0.98649 0.99141 3.0701e-006 1.228e-005 0.13322 0.86392 0.87373 0.0014157 0.95384 0.53878 0.0019065 0.42529 1.6484 1.6468 16.0099 144.9829 0.00023195 -85.5009 0.41095
1.515 0.98803 5.5162e-005 3.8182 0.01203 1.9929e-005 0.0011544 0.1731 0.00065866 0.17375 0.15897 0 0.035566 0.0389 0 0.93015 0.2646 0.07235 0.010007 4.4188 0.062451 7.5368e-005 0.82762 0.005438 0.0061779 0.0014214 0.98649 0.99141 3.0695e-006 1.2278e-005 0.13322 0.86429 0.87394 0.0014155 0.95412 0.53894 0.0019063 0.42531 1.6494 1.6477 16.0099 144.9829 0.00023162 -85.5021 0.41195
1.516 0.98803 5.5162e-005 3.8182 0.01203 1.9942e-005 0.0011544 0.17315 0.00065867 0.1738 0.15901 0 0.035563 0.0389 0 0.93024 0.26464 0.072363 0.010009 4.4193 0.062462 7.5381e-005 0.82761 0.0054385 0.0061784 0.0014211 0.98649 0.99141 3.0689e-006 1.2275e-005 0.13322 0.86466 0.87415 0.0014154 0.95439 0.5391 0.0019062 0.42532 1.6504 1.6487 16.0099 144.983 0.00023128 -85.5032 0.41295
1.517 0.98803 5.5162e-005 3.8182 0.01203 1.9955e-005 0.0011544 0.1732 0.00065867 0.17385 0.15906 0 0.03556 0.0389 0 0.93032 0.26468 0.072377 0.010011 4.4198 0.062472 7.5394e-005 0.8276 0.005439 0.0061789 0.0014208 0.9865 0.99141 3.0683e-006 1.2273e-005 0.13323 0.86503 0.87436 0.0014152 0.95467 0.53926 0.001906 0.42533 1.6513 1.6497 16.0099 144.983 0.00023095 -85.5043 0.41395
1.518 0.98803 5.5162e-005 3.8182 0.01203 1.9968e-005 0.0011544 0.17325 0.00065867 0.1739 0.15911 0 0.035557 0.0389 0 0.93041 0.26471 0.072391 0.010012 4.4203 0.062482 7.5408e-005 0.82759 0.0054394 0.0061794 0.0014206 0.9865 0.99142 3.0677e-006 1.2271e-005 0.13323 0.8654 0.87457 0.0014151 0.95494 0.53942 0.0019058 0.42534 1.6523 1.6506 16.0099 144.983 0.00023062 -85.5055 0.41495
1.519 0.98803 5.5161e-005 3.8182 0.01203 1.9981e-005 0.0011544 0.1733 0.00065867 0.17395 0.15915 0 0.035554 0.0389 0 0.93049 0.26475 0.072405 0.010014 4.4208 0.062493 7.5421e-005 0.82758 0.0054399 0.0061799 0.0014203 0.9865 0.99142 3.067e-006 1.2268e-005 0.13324 0.86577 0.87477 0.001415 0.95521 0.53958 0.0019056 0.42536 1.6533 1.6516 16.0099 144.983 0.00023029 -85.5066 0.41595
1.52 0.98803 5.5161e-005 3.8182 0.01203 1.9994e-005 0.0011544 0.17335 0.00065867 0.174 0.1592 0 0.035551 0.0389 0 0.93058 0.26479 0.072419 0.010016 4.4213 0.062503 7.5435e-005 0.82757 0.0054404 0.0061804 0.00142 0.98651 0.99142 3.0664e-006 1.2266e-005 0.13324 0.86614 0.87498 0.0014148 0.95548 0.53974 0.0019054 0.42537 1.6542 1.6526 16.0099 144.983 0.00022996 -85.5077 0.41695
1.521 0.98803 5.5161e-005 3.8182 0.01203 2.0007e-005 0.0011544 0.1734 0.00065867 0.17405 0.15925 0 0.035548 0.0389 0 0.93067 0.26483 0.072433 0.010017 4.4219 0.062513 7.5448e-005 0.82756 0.0054409 0.0061809 0.0014198 0.98651 0.99142 3.0658e-006 1.2263e-005 0.13324 0.8665 0.87519 0.0014147 0.95575 0.5399 0.0019052 0.42538 1.6552 1.6535 16.0099 144.983 0.00022964 -85.5088 0.41795
1.522 0.98803 5.5161e-005 3.8182 0.01203 2.002e-005 0.0011544 0.17345 0.00065867 0.1741 0.15929 0 0.035545 0.0389 0 0.93075 0.26487 0.072447 0.010019 4.4224 0.062524 7.5461e-005 0.82755 0.0054414 0.0061814 0.0014195 0.98651 0.99142 3.0652e-006 1.2261e-005 0.13325 0.86687 0.87539 0.0014146 0.95601 0.54006 0.0019051 0.42539 1.6561 1.6545 16.0099 144.9831 0.00022931 -85.5099 0.41895
1.523 0.98803 5.5161e-005 3.8182 0.01203 2.0034e-005 0.0011544 0.1735 0.00065867 0.17415 0.15934 0 0.035542 0.0389 0 0.93084 0.26491 0.072461 0.010021 4.4229 0.062534 7.5475e-005 0.82754 0.0054419 0.0061819 0.0014193 0.98652 0.99143 3.0647e-006 1.2259e-005 0.13325 0.86723 0.8756 0.0014144 0.95628 0.54022 0.0019049 0.42541 1.6571 1.6554 16.0099 144.9831 0.00022899 -85.511 0.41995
1.524 0.98803 5.5161e-005 3.8182 0.01203 2.0047e-005 0.0011544 0.17355 0.00065867 0.1742 0.15939 0 0.035539 0.0389 0 0.93092 0.26495 0.072474 0.010022 4.4234 0.062544 7.5488e-005 0.82753 0.0054424 0.0061824 0.001419 0.98652 0.99143 3.0641e-006 1.2256e-005 0.13326 0.8676 0.8758 0.0014143 0.95654 0.54038 0.0019047 0.42542 1.658 1.6564 16.0099 144.9831 0.00022866 -85.5121 0.42095
1.525 0.98803 5.5161e-005 3.8182 0.01203 2.006e-005 0.0011544 0.1736 0.00065867 0.17425 0.15943 0 0.035536 0.0389 0 0.93101 0.26498 0.072488 0.010024 4.4239 0.062555 7.5502e-005 0.82752 0.0054429 0.0061829 0.0014188 0.98652 0.99143 3.0635e-006 1.2254e-005 0.13326 0.86796 0.876 0.0014141 0.9568 0.54054 0.0019045 0.42543 1.659 1.6573 16.0099 144.9831 0.00022834 -85.5131 0.42195
1.526 0.98803 5.5161e-005 3.8182 0.01203 2.0073e-005 0.0011544 0.17365 0.00065867 0.1743 0.15948 0 0.035533 0.0389 0 0.9311 0.26502 0.072502 0.010026 4.4245 0.062565 7.5515e-005 0.82751 0.0054434 0.0061834 0.0014185 0.98653 0.99143 3.0629e-006 1.2252e-005 0.13327 0.86832 0.8762 0.001414 0.95706 0.5407 0.0019044 0.42544 1.6599 1.6583 16.0099 144.9831 0.00022802 -85.5142 0.42295
1.527 0.98803 5.5161e-005 3.8182 0.01203 2.0086e-005 0.0011544 0.1737 0.00065867 0.17435 0.15953 0 0.03553 0.0389 0 0.93118 0.26506 0.072516 0.010027 4.425 0.062575 7.5529e-005 0.8275 0.0054439 0.006184 0.0014182 0.98653 0.99144 3.0623e-006 1.2249e-005 0.13327 0.86868 0.87641 0.0014139 0.95732 0.54086 0.0019042 0.42546 1.6608 1.6592 16.0099 144.9832 0.0002277 -85.5153 0.42395
1.528 0.98803 5.5161e-005 3.8182 0.01203 2.0099e-005 0.0011544 0.17375 0.00065867 0.1744 0.15957 0 0.035527 0.0389 0 0.93127 0.2651 0.07253 0.010029 4.4255 0.062586 7.5542e-005 0.82749 0.0054444 0.0061845 0.001418 0.98653 0.99144 3.0618e-006 1.2247e-005 0.13327 0.86904 0.87661 0.0014138 0.95757 0.54102 0.001904 0.42547 1.6618 1.6602 16.0099 144.9832 0.00022739 -85.5163 0.42495
1.529 0.98803 5.5161e-005 3.8182 0.01203 2.0112e-005 0.0011544 0.1738 0.00065867 0.17445 0.15962 0 0.035524 0.0389 0 0.93136 0.26514 0.072544 0.010031 4.426 0.062596 7.5555e-005 0.82748 0.0054449 0.006185 0.0014178 0.98654 0.99144 3.0612e-006 1.2245e-005 0.13328 0.86939 0.87681 0.0014136 0.95783 0.54118 0.0019039 0.42548 1.6627 1.6611 16.0099 144.9832 0.00022707 -85.5174 0.42595
1.53 0.98803 5.5161e-005 3.8182 0.01203 2.0125e-005 0.0011544 0.17385 0.00065868 0.1745 0.15967 0 0.035521 0.0389 0 0.93144 0.26518 0.072558 0.010032 4.4265 0.062606 7.5569e-005 0.82747 0.0054454 0.0061855 0.0014175 0.98654 0.99144 3.0606e-006 1.2242e-005 0.13328 0.86975 0.877 0.0014135 0.95808 0.54133 0.0019037 0.42549 1.6636 1.662 16.0099 144.9832 0.00022675 -85.5184 0.42695
1.531 0.98803 5.5161e-005 3.8182 0.01203 2.0139e-005 0.0011544 0.1739 0.00065868 0.17455 0.15971 0 0.035518 0.0389 0 0.93153 0.26522 0.072572 0.010034 4.4271 0.062617 7.5582e-005 0.82746 0.0054459 0.006186 0.0014173 0.98654 0.99144 3.0601e-006 1.224e-005 0.13329 0.8701 0.8772 0.0014134 0.95833 0.54149 0.0019035 0.42551 1.6646 1.663 16.0098 144.9832 0.00022644 -85.5194 0.42795
1.532 0.98803 5.5161e-005 3.8182 0.012029 2.0152e-005 0.0011544 0.17394 0.00065868 0.1746 0.15976 0 0.035515 0.0389 0 0.93161 0.26525 0.072586 0.010036 4.4276 0.062627 7.5596e-005 0.82745 0.0054464 0.0061865 0.001417 0.98655 0.99145 3.0595e-006 1.2238e-005 0.13329 0.87046 0.8774 0.0014132 0.95858 0.54165 0.0019034 0.42552 1.6655 1.6639 16.0098 144.9833 0.00022613 -85.5205 0.42895
1.533 0.98803 5.5161e-005 3.8182 0.012029 2.0165e-005 0.0011544 0.17399 0.00065868 0.17465 0.15981 0 0.035512 0.0389 0 0.9317 0.26529 0.072599 0.010037 4.4281 0.062638 7.5609e-005 0.82744 0.0054469 0.006187 0.0014168 0.98655 0.99145 3.059e-006 1.2236e-005 0.13329 0.87081 0.8776 0.0014131 0.95883 0.54181 0.0019032 0.42553 1.6664 1.6648 16.0098 144.9833 0.00022582 -85.5215 0.42995
1.534 0.98803 5.516e-005 3.8182 0.012029 2.0178e-005 0.0011544 0.17404 0.00065868 0.1747 0.15985 0 0.035509 0.0389 0 0.93179 0.26533 0.072613 0.010039 4.4286 0.062648 7.5623e-005 0.82743 0.0054474 0.0061875 0.0014165 0.98655 0.99145 3.0584e-006 1.2234e-005 0.1333 0.87116 0.87779 0.001413 0.95907 0.54197 0.001903 0.42555 1.6673 1.6658 16.0098 144.9833 0.00022551 -85.5225 0.43095
1.535 0.98803 5.516e-005 3.8182 0.012029 2.0191e-005 0.0011544 0.17409 0.00065868 0.17475 0.1599 0 0.035506 0.0389 0 0.93187 0.26537 0.072627 0.010041 4.4292 0.062658 7.5636e-005 0.82742 0.0054479 0.006188 0.0014163 0.98656 0.99145 3.0579e-006 1.2231e-005 0.1333 0.87151 0.87799 0.0014129 0.95932 0.54213 0.0019029 0.42556 1.6683 1.6667 16.0098 144.9833 0.0002252 -85.5235 0.43195
1.536 0.98803 5.516e-005 3.8182 0.012029 2.0204e-005 0.0011544 0.17414 0.00065868 0.1748 0.15995 0 0.035503 0.0389 0 0.93196 0.26541 0.072641 0.010042 4.4297 0.062669 7.565e-005 0.82741 0.0054484 0.0061885 0.0014161 0.98656 0.99145 3.0573e-006 1.2229e-005 0.13331 0.87186 0.87818 0.0014127 0.95956 0.54229 0.0019027 0.42557 1.6692 1.6676 16.0098 144.9833 0.00022489 -85.5245 0.43295
1.537 0.98803 5.516e-005 3.8182 0.012029 2.0217e-005 0.0011544 0.17419 0.00065868 0.17485 0.15999 0 0.035501 0.0389 0 0.93205 0.26545 0.072655 0.010044 4.4302 0.062679 7.5663e-005 0.8274 0.0054489 0.006189 0.0014158 0.98656 0.99146 3.0568e-006 1.2227e-005 0.13331 0.87221 0.87837 0.0014126 0.9598 0.54245 0.0019025 0.42558 1.6701 1.6685 16.0098 144.9834 0.00022458 -85.5255 0.43395
1.538 0.98803 5.516e-005 3.8182 0.012029 2.023e-005 0.0011544 0.17424 0.00065868 0.17489 0.16004 0 0.035498 0.0389 0 0.93213 0.26549 0.072669 0.010046 4.4307 0.062689 7.5677e-005 0.82739 0.0054494 0.0061895 0.0014156 0.98656 0.99146 3.0563e-006 1.2225e-005 0.13331 0.87256 0.87857 0.0014125 0.96004 0.5426 0.0019024 0.4256 1.671 1.6695 16.0098 144.9834 0.00022428 -85.5265 0.43495
1.539 0.98803 5.516e-005 3.8182 0.012029 2.0244e-005 0.0011544 0.17429 0.00065868 0.17494 0.16008 0 0.035495 0.0389 0 0.93222 0.26552 0.072683 0.010047 4.4313 0.0627 7.569e-005 0.82738 0.0054499 0.0061901 0.0014154 0.98657 0.99146 3.0557e-006 1.2223e-005 0.13332 0.8729 0.87876 0.0014124 0.96028 0.54276 0.0019022 0.42561 1.6719 1.6704 16.0098 144.9834 0.00022398 -85.5274 0.43595
1.54 0.98803 5.516e-005 3.8182 0.012029 2.0257e-005 0.0011544 0.17434 0.00065868 0.17499 0.16013 0 0.035492 0.0389 0 0.93231 0.26556 0.072697 0.010049 4.4318 0.06271 7.5704e-005 0.82737 0.0054504 0.0061906 0.0014151 0.98657 0.99146 3.0552e-006 1.2221e-005 0.13332 0.87325 0.87895 0.0014123 0.96052 0.54292 0.0019021 0.42562 1.6728 1.6713 16.0098 144.9834 0.00022367 -85.5284 0.43695
1.541 0.98803 5.516e-005 3.8182 0.012029 2.027e-005 0.0011544 0.17439 0.00065868 0.17504 0.16018 0 0.035489 0.0389 0 0.93239 0.2656 0.072711 0.010051 4.4323 0.062721 7.5717e-005 0.82736 0.0054509 0.0061911 0.0014149 0.98657 0.99146 3.0547e-006 1.2219e-005 0.13333 0.87359 0.87914 0.0014121 0.96075 0.54308 0.0019019 0.42563 1.6737 1.6722 16.0098 144.9834 0.00022337 -85.5294 0.43795
1.542 0.98803 5.516e-005 3.8182 0.012029 2.0283e-005 0.0011544 0.17444 0.00065868 0.17509 0.16022 0 0.035486 0.0389 0 0.93248 0.26564 0.072725 0.010052 4.4328 0.062731 7.5731e-005 0.82734 0.0054514 0.0061916 0.0014147 0.98658 0.99147 3.0542e-006 1.2217e-005 0.13333 0.87394 0.87933 0.001412 0.96099 0.54324 0.0019018 0.42565 1.6746 1.6731 16.0098 144.9835 0.00022307 -85.5303 0.43895
1.543 0.98803 5.516e-005 3.8182 0.012029 2.0296e-005 0.0011544 0.17449 0.00065868 0.17514 0.16027 0 0.035483 0.0389 0 0.93257 0.26568 0.072739 0.010054 4.4334 0.062741 7.5744e-005 0.82733 0.0054519 0.0061921 0.0014145 0.98658 0.99147 3.0537e-006 1.2215e-005 0.13334 0.87428 0.87952 0.0014119 0.96122 0.5434 0.0019016 0.42566 1.6755 1.674 16.0098 144.9835 0.00022277 -85.5313 0.43995
1.544 0.98803 5.516e-005 3.8182 0.012029 2.0309e-005 0.0011544 0.17453 0.00065869 0.17519 0.16031 0 0.03548 0.0389 0 0.93265 0.26572 0.072753 0.010056 4.4339 0.062752 7.5757e-005 0.82732 0.0054524 0.0061926 0.0014142 0.98658 0.99147 3.0532e-006 1.2213e-005 0.13334 0.87462 0.8797 0.0014118 0.96145 0.54356 0.0019015 0.42567 1.6764 1.6749 16.0098 144.9835 0.00022248 -85.5322 0.44095
1.545 0.98803 5.516e-005 3.8182 0.012029 2.0322e-005 0.0011544 0.17458 0.00065869 0.17524 0.16036 0 0.035477 0.0389 0 0.93274 0.26576 0.072767 0.010057 4.4344 0.062762 7.5771e-005 0.82731 0.0054529 0.0061931 0.001414 0.98658 0.99147 3.0526e-006 1.2211e-005 0.13334 0.87496 0.87989 0.0014117 0.96168 0.54371 0.0019013 0.42569 1.6773 1.6758 16.0097 144.9835 0.00022218 -85.5332 0.44195
1.546 0.98803 5.516e-005 3.8182 0.012029 2.0335e-005 0.0011544 0.17463 0.00065869 0.17529 0.16041 0 0.035474 0.0389 0 0.93283 0.26579 0.072781 0.010059 4.435 0.062773 7.5784e-005 0.8273 0.0054534 0.0061936 0.0014138 0.98659 0.99147 3.0521e-006 1.2209e-005 0.13335 0.8753 0.88008 0.0014116 0.96191 0.54387 0.0019012 0.4257 1.6782 1.6767 16.0097 144.9835 0.00022188 -85.5341 0.44295
1.547 0.98803 5.516e-005 3.8182 0.012029 2.0349e-005 0.0011544 0.17468 0.00065869 0.17534 0.16045 0 0.035471 0.0389 0 0.93291 0.26583 0.072794 0.010061 4.4355 0.062783 7.5798e-005 0.82729 0.0054539 0.0061942 0.0014136 0.98659 0.99147 3.0516e-006 1.2207e-005 0.13335 0.87563 0.88026 0.0014114 0.96214 0.54403 0.001901 0.42571 1.6791 1.6776 16.0097 144.9836 0.00022159 -85.535 0.44395
1.548 0.98803 5.516e-005 3.8182 0.012029 2.0362e-005 0.0011544 0.17473 0.00065869 0.17538 0.1605 0 0.035468 0.0389 0 0.933 0.26587 0.072808 0.010062 4.436 0.062793 7.5811e-005 0.82728 0.0054544 0.0061947 0.0014134 0.98659 0.99148 3.0512e-006 1.2205e-005 0.13336 0.87597 0.88045 0.0014113 0.96236 0.54419 0.0019009 0.42572 1.68 1.6785 16.0097 144.9836 0.0002213 -85.5359 0.44495
1.549 0.98803 5.516e-005 3.8182 0.012029 2.0375e-005 0.0011544 0.17478 0.00065869 0.17543 0.16054 0 0.035466 0.0389 0 0.93309 0.26591 0.072822 0.010064 4.4365 0.062804 7.5825e-005 0.82727 0.0054549 0.0061952 0.0014132 0.9866 0.99148 3.0507e-006 1.2203e-005 0.13336 0.87631 0.88063 0.0014112 0.96259 0.54435 0.0019007 0.42574 1.6809 1.6794 16.0097 144.9836 0.000221 -85.5368 0.44595
1.55 0.98803 5.5159e-005 3.8182 0.012029 2.0388e-005 0.0011544 0.17483 0.00065869 0.17548 0.16059 0 0.035463 0.0389 0 0.93317 0.26595 0.072836 0.010066 4.4371 0.062814 7.5838e-005 0.82726 0.0054554 0.0061957 0.0014129 0.9866 0.99148 3.0502e-006 1.2201e-005 0.13336 0.87664 0.88082 0.0014111 0.96281 0.5445 0.0019006 0.42575 1.6818 1.6803 16.0097 144.9836 0.00022071 -85.5378 0.44695
1.551 0.98803 5.5159e-005 3.8182 0.012029 2.0401e-005 0.0011544 0.17488 0.00065869 0.17553 0.16064 0 0.03546 0.0389 0 0.93326 0.26599 0.07285 0.010067 4.4376 0.062825 7.5852e-005 0.82725 0.0054559 0.0061962 0.0014127 0.9866 0.99148 3.0497e-006 1.2199e-005 0.13337 0.87698 0.881 0.001411 0.96303 0.54466 0.0019004 0.42576 1.6826 1.6811 16.0097 144.9836 0.00022042 -85.5387 0.44795
1.552 0.98803 5.5159e-005 3.8182 0.012029 2.0414e-005 0.0011544 0.17492 0.00065869 0.17558 0.16068 0 0.035457 0.0389 0 0.93335 0.26603 0.072864 0.010069 4.4381 0.062835 7.5866e-005 0.82724 0.0054564 0.0061967 0.0014125 0.9866 0.99148 3.0492e-006 1.2197e-005 0.13337 0.87731 0.88118 0.0014109 0.96325 0.54482 0.0019003 0.42577 1.6835 1.682 16.0097 144.9837 0.00022014 -85.5395 0.44895
1.553 0.98803 5.5159e-005 3.8182 0.012029 2.0427e-005 0.0011544 0.17497 0.00065869 0.17563 0.16073 0 0.035454 0.0389 0 0.93343 0.26607 0.072878 0.010071 4.4387 0.062845 7.5879e-005 0.82723 0.0054569 0.0061972 0.0014123 0.98661 0.99149 3.0487e-006 1.2195e-005 0.13338 0.87764 0.88136 0.0014108 0.96347 0.54498 0.0019001 0.42579 1.6844 1.6829 16.0097 144.9837 0.00021985 -85.5404 0.44995
1.554 0.98803 5.5159e-005 3.8182 0.012029 2.044e-005 0.0011544 0.17502 0.00065869 0.17568 0.16077 0 0.035451 0.0389 0 0.93352 0.2661 0.072892 0.010072 4.4392 0.062856 7.5893e-005 0.82722 0.0054574 0.0061978 0.0014121 0.98661 0.99149 3.0483e-006 1.2193e-005 0.13338 0.87797 0.88155 0.0014107 0.96369 0.54514 0.0019 0.4258 1.6853 1.6838 16.0097 144.9837 0.00021956 -85.5413 0.45095
1.555 0.98803 5.5159e-005 3.8182 0.012029 2.0453e-005 0.0011544 0.17507 0.00065869 0.17572 0.16082 0 0.035448 0.0389 0 0.93361 0.26614 0.072906 0.010074 4.4397 0.062866 7.5906e-005 0.82721 0.0054579 0.0061983 0.0014119 0.98661 0.99149 3.0478e-006 1.2191e-005 0.13339 0.8783 0.88173 0.0014106 0.9639 0.54529 0.0018998 0.42581 1.6861 1.6847 16.0097 144.9837 0.00021928 -85.5422 0.45195
1.556 0.98803 5.5159e-005 3.8182 0.012029 2.0467e-005 0.0011544 0.17512 0.00065869 0.17577 0.16086 0 0.035445 0.0389 0 0.93369 0.26618 0.07292 0.010076 4.4403 0.062877 7.592e-005 0.8272 0.0054584 0.0061988 0.0014117 0.98662 0.99149 3.0473e-006 1.2189e-005 0.13339 0.87863 0.8819 0.0014105 0.96411 0.54545 0.0018997 0.42583 1.687 1.6855 16.0097 144.9837 0.00021899 -85.5431 0.45295
1.557 0.98803 5.5159e-005 3.8182 0.012029 2.048e-005 0.0011544 0.17517 0.00065869 0.17582 0.16091 0 0.035442 0.0389 0 0.93378 0.26622 0.072934 0.010077 4.4408 0.062887 7.5933e-005 0.82719 0.0054589 0.0061993 0.0014115 0.98662 0.99149 3.0468e-006 1.2187e-005 0.13339 0.87895 0.88208 0.0014103 0.96433 0.54561 0.0018996 0.42584 1.6879 1.6864 16.0096 144.9837 0.00021871 -85.5439 0.45395
1.558 0.98803 5.5159e-005 3.8182 0.012029 2.0493e-005 0.0011544 0.17522 0.00065869 0.17587 0.16095 0 0.03544 0.0389 0 0.93387 0.26626 0.072948 0.010079 4.4413 0.062897 7.5947e-005 0.82718 0.0054594 0.0061998 0.0014113 0.98662 0.99149 3.0464e-006 1.2185e-005 0.1334 0.87928 0.88226 0.0014102 0.96454 0.54577 0.0018994 0.42585 1.6887 1.6873 16.0096 144.9838 0.00021843 -85.5448 0.45495
1.559 0.98803 5.5159e-005 3.8182 0.012029 2.0506e-005 0.0011544 0.17526 0.0006587 0.17592 0.161 0 0.035437 0.0389 0 0.93395 0.2663 0.072962 0.010081 4.4419 0.062908 7.596e-005 0.82717 0.0054599 0.0062003 0.0014111 0.98662 0.9915 3.0459e-006 1.2184e-005 0.1334 0.87961 0.88244 0.0014101 0.96475 0.54592 0.0018993 0.42586 1.6896 1.6881 16.0096 144.9838 0.00021815 -85.5456 0.45595
1.56 0.98803 5.5159e-005 3.8182 0.012029 2.0519e-005 0.0011544 0.17531 0.0006587 0.17597 0.16105 0 0.035434 0.0389 0 0.93404 0.26634 0.072976 0.010082 4.4424 0.062918 7.5974e-005 0.82716 0.0054604 0.0062008 0.0014109 0.98663 0.9915 3.0455e-006 1.2182e-005 0.13341 0.87993 0.88262 0.00141 0.96496 0.54608 0.0018992 0.42588 1.6905 1.689 16.0096 144.9838 0.00021787 -85.5465 0.45695
1.561 0.98803 5.5159e-005 3.8182 0.012029 2.0532e-005 0.0011544 0.17536 0.0006587 0.17601 0.16109 0 0.035431 0.0389 0 0.93413 0.26638 0.07299 0.010084 4.4429 0.062929 7.5987e-005 0.82715 0.0054609 0.0062014 0.0014107 0.98663 0.9915 3.045e-006 1.218e-005 0.13341 0.88025 0.88279 0.0014099 0.96517 0.54624 0.001899 0.42589 1.6913 1.6899 16.0096 144.9838 0.00021759 -85.5473 0.45795
1.562 0.98803 5.5159e-005 3.8182 0.012029 2.0545e-005 0.0011544 0.17541 0.0006587 0.17606 0.16114 0 0.035428 0.0389 0 0.93421 0.26642 0.073004 0.010086 4.4435 0.062939 7.6001e-005 0.82714 0.0054614 0.0062019 0.0014105 0.98663 0.9915 3.0446e-006 1.2178e-005 0.13341 0.88058 0.88297 0.0014098 0.96537 0.5464 0.0018989 0.4259 1.6922 1.6907 16.0096 144.9838 0.00021732 -85.5481 0.45895
1.563 0.98803 5.5159e-005 3.8182 0.012029 2.0558e-005 0.0011544 0.17546 0.0006587 0.17611 0.16118 0 0.035425 0.0389 0 0.9343 0.26645 0.073018 0.010088 4.444 0.062949 7.6014e-005 0.82713 0.0054619 0.0062024 0.0014103 0.98663 0.9915 3.0441e-006 1.2176e-005 0.13342 0.8809 0.88314 0.0014097 0.96558 0.54655 0.0018988 0.42591 1.693 1.6916 16.0096 144.9839 0.00021704 -85.549 0.45995
1.564 0.98803 5.5159e-005 3.8182 0.012029 2.0572e-005 0.0011544 0.1755 0.0006587 0.17616 0.16123 0 0.035422 0.0389 0 0.93439 0.26649 0.073032 0.010089 4.4446 0.06296 7.6028e-005 0.82712 0.0054624 0.0062029 0.0014101 0.98664 0.9915 3.0437e-006 1.2175e-005 0.13342 0.88122 0.88331 0.0014096 0.96578 0.54671 0.0018986 0.42593 1.6939 1.6924 16.0096 144.9839 0.00021676 -85.5498 0.46095
1.565 0.98803 5.5159e-005 3.8182 0.012029 2.0585e-005 0.0011544 0.17555 0.0006587 0.17621 0.16127 0 0.03542 0.0389 0 0.93447 0.26653 0.073046 0.010091 4.4451 0.06297 7.6041e-005 0.82711 0.0054629 0.0062034 0.0014099 0.98664 0.99151 3.0432e-006 1.2173e-005 0.13343 0.88154 0.88349 0.0014095 0.96598 0.54687 0.0018985 0.42594 1.6947 1.6933 16.0096 144.9839 0.00021649 -85.5506 0.46195
1.566 0.98803 5.5158e-005 3.8182 0.012029 2.0598e-005 0.0011544 0.1756 0.0006587 0.17625 0.16132 0 0.035417 0.0389 0 0.93456 0.26657 0.07306 0.010093 4.4456 0.062981 7.6055e-005 0.8271 0.0054635 0.006204 0.0014097 0.98664 0.99151 3.0428e-006 1.2171e-005 0.13343 0.88185 0.88366 0.0014094 0.96618 0.54703 0.0018984 0.42595 1.6956 1.6942 16.0096 144.9839 0.00021622 -85.5514 0.46295
1.567 0.98803 5.5158e-005 3.8182 0.012029 2.0611e-005 0.0011544 0.17565 0.0006587 0.1763 0.16136 0 0.035414 0.0389 0 0.93465 0.26661 0.073074 0.010094 4.4462 0.062991 7.6069e-005 0.82708 0.005464 0.0062045 0.0014095 0.98664 0.99151 3.0424e-006 1.2169e-005 0.13344 0.88217 0.88383 0.0014093 0.96638 0.54718 0.0018982 0.42597 1.6964 1.695 16.0096 144.9839 0.00021595 -85.5522 0.46395
1.568 0.98803 5.5158e-005 3.8182 0.012029 2.0624e-005 0.0011544 0.1757 0.0006587 0.17635 0.16141 0 0.035411 0.0389 0 0.93474 0.26665 0.073088 0.010096 4.4467 0.063002 7.6082e-005 0.82707 0.0054645 0.006205 0.0014093 0.98665 0.99151 3.0419e-006 1.2168e-005 0.13344 0.88249 0.884 0.0014092 0.96658 0.54734 0.0018981 0.42598 1.6973 1.6958 16.0095 144.984 0.00021568 -85.553 0.46495
1.569 0.98803 5.5158e-005 3.8182 0.012029 2.0637e-005 0.0011544 0.17574 0.0006587 0.1764 0.16145 0 0.035408 0.0389 0 0.93482 0.26669 0.073102 0.010098 4.4472 0.063012 7.6096e-005 0.82706 0.005465 0.0062055 0.0014092 0.98665 0.99151 3.0415e-006 1.2166e-005 0.13344 0.8828 0.88417 0.0014091 0.96678 0.5475 0.001898 0.42599 1.6981 1.6967 16.0095 144.984 0.00021541 -85.5538 0.46595
1.57 0.98803 5.5158e-005 3.8182 0.012029 2.065e-005 0.0011544 0.17579 0.0006587 0.17645 0.1615 0 0.035405 0.0389 0 0.93491 0.26673 0.073116 0.010099 4.4478 0.063023 7.6109e-005 0.82705 0.0054655 0.006206 0.001409 0.98665 0.99151 3.0411e-006 1.2164e-005 0.13345 0.88312 0.88434 0.001409 0.96697 0.54765 0.0018978 0.426 1.6989 1.6975 16.0095 144.984 0.00021514 -85.5546 0.46695
1.571 0.98803 5.5158e-005 3.8182 0.012029 2.0663e-005 0.0011544 0.17584 0.0006587 0.17649 0.16154 0 0.035402 0.0389 0 0.935 0.26677 0.07313 0.010101 4.4483 0.063033 7.6123e-005 0.82704 0.005466 0.0062066 0.0014088 0.98665 0.99152 3.0407e-006 1.2163e-005 0.13345 0.88343 0.88451 0.0014089 0.96717 0.54781 0.0018977 0.42602 1.6998 1.6984 16.0095 144.984 0.00021487 -85.5554 0.46795
1.572 0.98803 5.5158e-005 3.8182 0.012029 2.0676e-005 0.0011544 0.17589 0.0006587 0.17654 0.16159 0 0.0354 0.0389 0 0.93508 0.2668 0.073144 0.010103 4.4489 0.063043 7.6136e-005 0.82703 0.0054665 0.0062071 0.0014086 0.98666 0.99152 3.0403e-006 1.2161e-005 0.13346 0.88374 0.88468 0.0014088 0.96736 0.54797 0.0018976 0.42603 1.7006 1.6992 16.0095 144.984 0.00021461 -85.5562 0.46895
1.573 0.98803 5.5158e-005 3.8182 0.012029 2.069e-005 0.0011544 0.17594 0.0006587 0.17659 0.16163 0 0.035397 0.0389 0 0.93517 0.26684 0.073158 0.010104 4.4494 0.063054 7.615e-005 0.82702 0.005467 0.0062076 0.0014084 0.98666 0.99152 3.0398e-006 1.2159e-005 0.13346 0.88406 0.88485 0.0014087 0.96755 0.54813 0.0018975 0.42604 1.7014 1.7001 16.0095 144.9841 0.00021434 -85.5569 0.46995
1.574 0.98803 5.5158e-005 3.8182 0.012029 2.0703e-005 0.0011544 0.17598 0.00065871 0.17664 0.16168 0 0.035394 0.0389 0 0.93526 0.26688 0.073172 0.010106 4.45 0.063064 7.6164e-005 0.82701 0.0054675 0.0062081 0.0014082 0.98666 0.99152 3.0394e-006 1.2158e-005 0.13347 0.88437 0.88502 0.0014086 0.96774 0.54828 0.0018973 0.42606 1.7023 1.7009 16.0095 144.9841 0.00021408 -85.5577 0.47095
1.575 0.98803 5.5158e-005 3.8182 0.012029 2.0716e-005 0.0011544 0.17603 0.00065871 0.17669 0.16172 0 0.035391 0.0389 0 0.93535 0.26692 0.073186 0.010108 4.4505 0.063075 7.6177e-005 0.827 0.005468 0.0062086 0.0014081 0.98666 0.99152 3.039e-006 1.2156e-005 0.13347 0.88468 0.88518 0.0014086 0.96793 0.54844 0.0018972 0.42607 1.7031 1.7017 16.0095 144.9841 0.00021381 -85.5585 0.47195
1.576 0.98803 5.5158e-005 3.8182 0.012029 2.0729e-005 0.0011544 0.17608 0.00065871 0.17673 0.16177 0 0.035388 0.0389 0 0.93543 0.26696 0.0732 0.010109 4.451 0.063085 7.6191e-005 0.82699 0.0054685 0.0062092 0.0014079 0.98666 0.99152 3.0386e-006 1.2154e-005 0.13347 0.88498 0.88535 0.0014085 0.96812 0.5486 0.0018971 0.42608 1.7039 1.7025 16.0095 144.9841 0.00021355 -85.5592 0.47295
1.577 0.98803 5.5158e-005 3.8182 0.012029 2.0742e-005 0.0011544 0.17613 0.00065871 0.17678 0.16181 0 0.035385 0.0389 0 0.93552 0.267 0.073214 0.010111 4.4516 0.063096 7.6204e-005 0.82698 0.0054691 0.0062097 0.0014077 0.98667 0.99152 3.0382e-006 1.2153e-005 0.13348 0.88529 0.88552 0.0014084 0.96831 0.54875 0.001897 0.42609 1.7047 1.7034 16.0094 144.9841 0.00021329 -85.56 0.47395
1.578 0.98803 5.5158e-005 3.8182 0.012029 2.0755e-005 0.0011544 0.17617 0.00065871 0.17683 0.16186 0 0.035383 0.0389 0 0.93561 0.26704 0.073229 0.010113 4.4521 0.063106 7.6218e-005 0.82697 0.0054696 0.0062102 0.0014075 0.98667 0.99153 3.0378e-006 1.2151e-005 0.13348 0.8856 0.88568 0.0014083 0.9685 0.54891 0.0018969 0.42611 1.7056 1.7042 16.0094 144.9842 0.00021303 -85.5607 0.47495
1.579 0.98803 5.5158e-005 3.8182 0.012029 2.0768e-005 0.0011544 0.17622 0.00065871 0.17688 0.1619 0 0.03538 0.0389 0 0.93569 0.26708 0.073243 0.010114 4.4527 0.063117 7.6231e-005 0.82696 0.0054701 0.0062107 0.0014074 0.98667 0.99153 3.0374e-006 1.215e-005 0.13349 0.8859 0.88584 0.0014082 0.96868 0.54907 0.0018967 0.42612 1.7064 1.705 16.0094 144.9842 0.00021277 -85.5615 0.47595
1.58 0.98803 5.5158e-005 3.8182 0.012029 2.0781e-005 0.0011544 0.17627 0.00065871 0.17692 0.16195 0 0.035377 0.0389 0 0.93578 0.26712 0.073257 0.010116 4.4532 0.063127 7.6245e-005 0.82695 0.0054706 0.0062113 0.0014072 0.98667 0.99153 3.037e-006 1.2148e-005 0.13349 0.88621 0.88601 0.0014081 0.96886 0.54922 0.0018966 0.42613 1.7072 1.7058 16.0094 144.9842 0.00021251 -85.5622 0.47695
1.581 0.98803 5.5157e-005 3.8182 0.012029 2.0795e-005 0.0011544 0.17632 0.00065871 0.17697 0.16199 0 0.035374 0.0389 0 0.93587 0.26716 0.073271 0.010118 4.4538 0.063137 7.6259e-005 0.82694 0.0054711 0.0062118 0.001407 0.98668 0.99153 3.0366e-006 1.2146e-005 0.13349 0.88651 0.88617 0.001408 0.96905 0.54938 0.0018965 0.42615 1.708 1.7067 16.0094 144.9842 0.00021226 -85.5629 0.47795
1.582 0.98803 5.5157e-005 3.8182 0.012029 2.0808e-005 0.0011544 0.17636 0.00065871 0.17702 0.16204 0 0.035371 0.0389 0 0.93596 0.26719 0.073285 0.010119 4.4543 0.063148 7.6272e-005 0.82693 0.0054716 0.0062123 0.0014068 0.98668 0.99153 3.0362e-006 1.2145e-005 0.1335 0.88681 0.88633 0.0014079 0.96923 0.54953 0.0018964 0.42616 1.7088 1.7075 16.0094 144.9842 0.000212 -85.5637 0.47895
1.583 0.98803 5.5157e-005 3.8182 0.012029 2.0821e-005 0.0011544 0.17641 0.00065871 0.17707 0.16208 0 0.035369 0.0389 0 0.93604 0.26723 0.073299 0.010121 4.4549 0.063158 7.6286e-005 0.82692 0.0054721 0.0062128 0.0014067 0.98668 0.99153 3.0358e-006 1.2143e-005 0.1335 0.88712 0.88649 0.0014078 0.96941 0.54969 0.0018963 0.42617 1.7096 1.7083 16.0094 144.9843 0.00021174 -85.5644 0.47995
1.584 0.98803 5.5157e-005 3.8182 0.012029 2.0834e-005 0.0011544 0.17646 0.00065871 0.17711 0.16213 0 0.035366 0.0389 0 0.93613 0.26727 0.073313 0.010123 4.4554 0.063169 7.6299e-005 0.82691 0.0054726 0.0062134 0.0014065 0.98668 0.99153 3.0354e-006 1.2142e-005 0.13351 0.88742 0.88666 0.0014077 0.96959 0.54985 0.0018962 0.42618 1.7104 1.7091 16.0094 144.9843 0.00021149 -85.5651 0.48095
1.585 0.98803 5.5157e-005 3.8182 0.012029 2.0847e-005 0.0011544 0.17651 0.00065871 0.17716 0.16217 0 0.035363 0.0389 0 0.93622 0.26731 0.073327 0.010124 4.4559 0.063179 7.6313e-005 0.8269 0.0054731 0.0062139 0.0014063 0.98668 0.99154 3.0351e-006 1.214e-005 0.13351 0.88772 0.88682 0.0014076 0.96977 0.55 0.001896 0.4262 1.7113 1.7099 16.0094 144.9843 0.00021124 -85.5658 0.48195
1.586 0.98803 5.5157e-005 3.8182 0.012029 2.086e-005 0.0011544 0.17655 0.00065871 0.17721 0.16221 0 0.03536 0.0389 0 0.93631 0.26735 0.073341 0.010126 4.4565 0.06319 7.6327e-005 0.82689 0.0054737 0.0062144 0.0014062 0.98669 0.99154 3.0347e-006 1.2139e-005 0.13352 0.88802 0.88698 0.0014076 0.96994 0.55016 0.0018959 0.42621 1.7121 1.7107 16.0093 144.9843 0.00021099 -85.5665 0.48295
1.587 0.98803 5.5157e-005 3.8182 0.012029 2.0873e-005 0.0011544 0.1766 0.00065871 0.17726 0.16226 0 0.035357 0.0389 0 0.93639 0.26739 0.073355 0.010128 4.457 0.0632 7.634e-005 0.82688 0.0054742 0.0062149 0.001406 0.98669 0.99154 3.0343e-006 1.2137e-005 0.13352 0.88831 0.88713 0.0014075 0.97012 0.55032 0.0018958 0.42622 1.7129 1.7115 16.0093 144.9843 0.00021073 -85.5672 0.48395
1.588 0.98803 5.5157e-005 3.8182 0.012029 2.0886e-005 0.0011544 0.17665 0.00065871 0.1773 0.1623 0 0.035355 0.0389 0 0.93648 0.26743 0.073369 0.01013 4.4576 0.063211 7.6354e-005 0.82687 0.0054747 0.0062155 0.0014058 0.98669 0.99154 3.0339e-006 1.2136e-005 0.13352 0.88861 0.88729 0.0014074 0.97029 0.55047 0.0018957 0.42624 1.7137 1.7123 16.0093 144.9844 0.00021048 -85.5679 0.48495
1.589 0.98803 5.5157e-005 3.8182 0.012029 2.0899e-005 0.0011544 0.1767 0.00065872 0.17735 0.16235 0 0.035352 0.0389 0 0.93657 0.26747 0.073383 0.010131 4.4581 0.063221 7.6368e-005 0.82686 0.0054752 0.006216 0.0014057 0.98669 0.99154 3.0336e-006 1.2134e-005 0.13353 0.88891 0.88745 0.0014073 0.97047 0.55063 0.0018956 0.42625 1.7145 1.7131 16.0093 144.9844 0.00021023 -85.5686 0.48595
1.59 0.98803 5.5157e-005 3.8182 0.012029 2.0913e-005 0.0011544 0.17674 0.00065872 0.1774 0.16239 0 0.035349 0.0389 0 0.93665 0.26751 0.073397 0.010133 4.4587 0.063232 7.6381e-005 0.82684 0.0054757 0.0062165 0.0014055 0.9867 0.99154 3.0332e-006 1.2133e-005 0.13353 0.8892 0.88761 0.0014072 0.97064 0.55078 0.0018955 0.42626 1.7153 1.7139 16.0093 144.9844 0.00020999 -85.5693 0.48695
1.591 0.98803 5.5157e-005 3.8182 0.012029 2.0926e-005 0.0011544 0.17679 0.00065872 0.17744 0.16244 0 0.035346 0.0389 0 0.93674 0.26755 0.073411 0.010135 4.4592 0.063242 7.6395e-005 0.82683 0.0054762 0.006217 0.0014054 0.9867 0.99154 3.0328e-006 1.2131e-005 0.13354 0.8895 0.88776 0.0014071 0.97081 0.55094 0.0018954 0.42627 1.716 1.7147 16.0093 144.9844 0.00020974 -85.57 0.48795
1.592 0.98803 5.5157e-005 3.8182 0.012029 2.0939e-005 0.0011544 0.17684 0.00065872 0.17749 0.16248 0 0.035343 0.0389 0 0.93683 0.26758 0.073426 0.010136 4.4598 0.063253 7.6408e-005 0.82682 0.0054767 0.0062176 0.0014052 0.9867 0.99155 3.0325e-006 1.213e-005 0.13354 0.88979 0.88792 0.0014071 0.97098 0.5511 0.0018953 0.42629 1.7168 1.7155 16.0093 144.9844 0.00020949 -85.5707 0.48895
1.593 0.98803 5.5157e-005 3.8182 0.012029 2.0952e-005 0.0011544 0.17688 0.00065872 0.17754 0.16252 0 0.035341 0.0389 0 0.93692 0.26762 0.07344 0.010138 4.4603 0.063263 7.6422e-005 0.82681 0.0054773 0.0062181 0.001405 0.9867 0.99155 3.0321e-006 1.2128e-005 0.13355 0.89008 0.88808 0.001407 0.97115 0.55125 0.0018951 0.4263 1.7176 1.7163 16.0093 144.9845 0.00020925 -85.5713 0.48995
1.594 0.98803 5.5157e-005 3.8182 0.012029 2.0965e-005 0.0011544 0.17693 0.00065872 0.17759 0.16257 0 0.035338 0.0389 0 0.937 0.26766 0.073454 0.01014 4.4609 0.063274 7.6436e-005 0.8268 0.0054778 0.0062186 0.0014049 0.9867 0.99155 3.0317e-006 1.2127e-005 0.13355 0.89038 0.88823 0.0014069 0.97132 0.55141 0.001895 0.42631 1.7184 1.7171 16.0092 144.9845 0.000209 -85.572 0.49095
1.595 0.98803 5.5157e-005 3.8182 0.012029 2.0978e-005 0.0011544 0.17698 0.00065872 0.17763 0.16261 0 0.035335 0.0389 0 0.93709 0.2677 0.073468 0.010141 4.4614 0.063284 7.6449e-005 0.82679 0.0054783 0.0062191 0.0014047 0.98671 0.99155 3.0314e-006 1.2125e-005 0.13355 0.89067 0.88839 0.0014068 0.97148 0.55156 0.0018949 0.42633 1.7192 1.7179 16.0092 144.9845 0.00020876 -85.5727 0.49195
1.596 0.98803 5.5157e-005 3.8182 0.012029 2.0991e-005 0.0011544 0.17702 0.00065872 0.17768 0.16266 0 0.035332 0.0389 0 0.93718 0.26774 0.073482 0.010143 4.462 0.063295 7.6463e-005 0.82678 0.0054788 0.0062197 0.0014046 0.98671 0.99155 3.031e-006 1.2124e-005 0.13356 0.89096 0.88854 0.0014067 0.97165 0.55172 0.0018948 0.42634 1.72 1.7187 16.0092 144.9845 0.00020852 -85.5733 0.49295
1.597 0.98803 5.5156e-005 3.8182 0.012029 2.1004e-005 0.0011544 0.17707 0.00065872 0.17773 0.1627 0 0.03533 0.0389 0 0.93727 0.26778 0.073496 0.010145 4.4625 0.063305 7.6477e-005 0.82677 0.0054793 0.0062202 0.0014044 0.98671 0.99155 3.0307e-006 1.2123e-005 0.13356 0.89124 0.88869 0.0014066 0.97182 0.55188 0.0018947 0.42635 1.7208 1.7195 16.0092 144.9845 0.00020828 -85.574 0.49395
1.598 0.98803 5.5156e-005 3.8182 0.012029 2.1018e-005 0.0011544 0.17712 0.00065872 0.17777 0.16275 0 0.035327 0.0389 0 0.93735 0.26782 0.07351 0.010146 4.4631 0.063316 7.649e-005 0.82676 0.0054798 0.0062207 0.0014043 0.98671 0.99155 3.0303e-006 1.2121e-005 0.13357 0.89153 0.88885 0.0014066 0.97198 0.55203 0.0018946 0.42636 1.7215 1.7203 16.0092 144.9846 0.00020804 -85.5746 0.49495
1.599 0.98803 5.5156e-005 3.8182 0.012029 2.1031e-005 0.0011544 0.17717 0.00065872 0.17782 0.16279 0 0.035324 0.0389 0 0.93744 0.26786 0.073524 0.010148 4.4637 0.063326 7.6504e-005 0.82675 0.0054804 0.0062213 0.0014041 0.98671 0.99155 3.03e-006 1.212e-005 0.13357 0.89182 0.889 0.0014065 0.97214 0.55219 0.0018945 0.42638 1.7223 1.721 16.0092 144.9846 0.0002078 -85.5753 0.49595
1.6 0.98803 5.5156e-005 3.8182 0.012029 2.1044e-005 0.0011544 0.17721 0.00065872 0.17787 0.16283 0 0.035321 0.0389 0 0.93753 0.2679 0.073538 0.01015 4.4642 0.063337 7.6518e-005 0.82674 0.0054809 0.0062218 0.001404 0.98672 0.99156 3.0296e-006 1.2118e-005 0.13358 0.89211 0.88915 0.0014064 0.9723 0.55234 0.0018944 0.42639 1.7231 1.7218 16.0092 144.9846 0.00020756 -85.5759 0.49695
1.601 0.98803 5.5156e-005 3.8182 0.012029 2.1057e-005 0.0011544 0.17726 0.00065872 0.17791 0.16288 0 0.035319 0.0389 0 0.93762 0.26794 0.073552 0.010151 4.4648 0.063347 7.6531e-005 0.82673 0.0054814 0.0062223 0.0014038 0.98672 0.99156 3.0293e-006 1.2117e-005 0.13358 0.89239 0.8893 0.0014063 0.97246 0.5525 0.0018943 0.4264 1.7239 1.7226 16.0091 144.9846 0.00020732 -85.5766 0.49795
1.602 0.98803 5.5156e-005 3.8182 0.012029 2.107e-005 0.0011544 0.17731 0.00065872 0.17796 0.16292 0 0.035316 0.0389 0 0.93771 0.26798 0.073567 0.010153 4.4653 0.063358 7.6545e-005 0.82672 0.0054819 0.0062229 0.0014037 0.98672 0.99156 3.0289e-006 1.2116e-005 0.13358 0.89268 0.88945 0.0014062 0.97262 0.55265 0.0018942 0.42642 1.7246 1.7234 16.0091 144.9846 0.00020708 -85.5772 0.49895
1.603 0.98803 5.5156e-005 3.8182 0.012029 2.1083e-005 0.0011544 0.17735 0.00065872 0.17801 0.16297 0 0.035313 0.0389 0 0.93779 0.26802 0.073581 0.010155 4.4659 0.063368 7.6558e-005 0.82671 0.0054824 0.0062234 0.0014035 0.98672 0.99156 3.0286e-006 1.2114e-005 0.13359 0.89296 0.8896 0.0014062 0.97278 0.55281 0.0018941 0.42643 1.7254 1.7241 16.0091 144.9847 0.00020685 -85.5778 0.49995
1.604 0.98803 5.5156e-005 3.8182 0.012028 2.1096e-005 0.0011544 0.1774 0.00065873 0.17805 0.16301 0 0.03531 0.0389 0 0.93788 0.26805 0.073595 0.010157 4.4664 0.063379 7.6572e-005 0.8267 0.0054829 0.0062239 0.0014034 0.98672 0.99156 3.0283e-006 1.2113e-005 0.13359 0.89324 0.88975 0.0014061 0.97294 0.55296 0.001894 0.42644 1.7262 1.7249 16.0091 144.9847 0.00020661 -85.5785 0.50095
1.605 0.98803 5.5156e-005 3.8182 0.012028 2.1109e-005 0.0011544 0.17745 0.00065873 0.1781 0.16305 0 0.035308 0.0389 0 0.93797 0.26809 0.073609 0.010158 4.467 0.063389 7.6586e-005 0.82669 0.0054835 0.0062244 0.0014032 0.98672 0.99156 3.0279e-006 1.2112e-005 0.1336 0.89352 0.8899 0.001406 0.9731 0.55312 0.0018939 0.42645 1.727 1.7257 16.0091 144.9847 0.00020638 -85.5791 0.50195
1.606 0.98803 5.5156e-005 3.8182 0.012028 2.1122e-005 0.0011544 0.17749 0.00065873 0.17815 0.1631 0 0.035305 0.0389 0 0.93806 0.26813 0.073623 0.01016 4.4675 0.0634 7.6599e-005 0.82668 0.005484 0.006225 0.0014031 0.98673 0.99156 3.0276e-006 1.211e-005 0.1336 0.89381 0.89004 0.0014059 0.97325 0.55327 0.0018938 0.42647 1.7277 1.7265 16.0091 144.9847 0.00020614 -85.5797 0.50295
1.607 0.98803 5.5156e-005 3.8182 0.012028 2.1136e-005 0.0011544 0.17754 0.00065873 0.17819 0.16314 0 0.035302 0.0389 0 0.93814 0.26817 0.073637 0.010162 4.4681 0.06341 7.6613e-005 0.82667 0.0054845 0.0062255 0.0014029 0.98673 0.99156 3.0273e-006 1.2109e-005 0.13361 0.89409 0.89019 0.0014059 0.97341 0.55343 0.0018937 0.42648 1.7285 1.7272 16.0091 144.9847 0.00020591 -85.5803 0.50395
1.608 0.98803 5.5156e-005 3.8182 0.012028 2.1149e-005 0.0011544 0.17758 0.00065873 0.17824 0.16318 0 0.035299 0.0389 0 0.93823 0.26821 0.073651 0.010163 4.4687 0.063421 7.6627e-005 0.82666 0.005485 0.006226 0.0014028 0.98673 0.99157 3.027e-006 1.2108e-005 0.13361 0.89436 0.89034 0.0014058 0.97356 0.55358 0.0018936 0.42649 1.7292 1.728 16.0091 144.9848 0.00020568 -85.5809 0.50495
1.609 0.98803 5.5156e-005 3.8182 0.012028 2.1162e-005 0.0011544 0.17763 0.00065873 0.17829 0.16323 0 0.035297 0.0389 0 0.93832 0.26825 0.073666 0.010165 4.4692 0.063431 7.664e-005 0.82665 0.0054855 0.0062266 0.0014027 0.98673 0.99157 3.0266e-006 1.2106e-005 0.13361 0.89464 0.89049 0.0014057 0.97371 0.55374 0.0018935 0.42651 1.73 1.7287 16.009 144.9848 0.00020545 -85.5815 0.50595
1.61 0.98803 5.5156e-005 3.8182 0.012028 2.1175e-005 0.0011544 0.17768 0.00065873 0.17833 0.16327 0 0.035294 0.0389 0 0.93841 0.26829 0.07368 0.010167 4.4698 0.063442 7.6654e-005 0.82663 0.0054861 0.0062271 0.0014025 0.98673 0.99157 3.0263e-006 1.2105e-005 0.13362 0.89492 0.89063 0.0014056 0.97386 0.55389 0.0018934 0.42652 1.7308 1.7295 16.009 144.9848 0.00020522 -85.5821 0.50695
1.611 0.98803 5.5156e-005 3.8182 0.012028 2.1188e-005 0.0011544 0.17772 0.00065873 0.17838 0.16332 0 0.035291 0.0389 0 0.93849 0.26833 0.073694 0.010168 4.4703 0.063452 7.6668e-005 0.82662 0.0054866 0.0062276 0.0014024 0.98674 0.99157 3.026e-006 1.2104e-005 0.13362 0.8952 0.89078 0.0014056 0.97402 0.55405 0.0018933 0.42653 1.7315 1.7303 16.009 144.9848 0.00020499 -85.5827 0.50795
1.612 0.98803 5.5155e-005 3.8182 0.012028 2.1201e-005 0.0011544 0.17777 0.00065873 0.17842 0.16336 0 0.035288 0.0389 0 0.93858 0.26837 0.073708 0.01017 4.4709 0.063463 7.6682e-005 0.82661 0.0054871 0.0062282 0.0014022 0.98674 0.99157 3.0257e-006 1.2103e-005 0.13363 0.89547 0.89092 0.0014055 0.97417 0.5542 0.0018932 0.42654 1.7323 1.731 16.009 144.9848 0.00020476 -85.5833 0.50895
1.613 0.98803 5.5155e-005 3.8182 0.012028 2.1214e-005 0.0011544 0.17782 0.00065873 0.17847 0.1634 0 0.035286 0.0389 0 0.93867 0.26841 0.073722 0.010172 4.4714 0.063473 7.6695e-005 0.8266 0.0054876 0.0062287 0.0014021 0.98674 0.99157 3.0254e-006 1.2101e-005 0.13363 0.89575 0.89107 0.0014054 0.97431 0.55436 0.0018931 0.42656 1.733 1.7318 16.009 144.9849 0.00020454 -85.5839 0.50995
1.614 0.98803 5.5155e-005 3.8182 0.012028 2.1227e-005 0.0011544 0.17786 0.00065873 0.17852 0.16345 0 0.035283 0.0389 0 0.93876 0.26845 0.073736 0.010173 4.472 0.063484 7.6709e-005 0.82659 0.0054881 0.0062292 0.001402 0.98674 0.99157 3.025e-006 1.21e-005 0.13364 0.89602 0.89121 0.0014053 0.97446 0.55451 0.001893 0.42657 1.7338 1.7325 16.009 144.9849 0.00020431 -85.5845 0.51095
1.615 0.98803 5.5155e-005 3.8182 0.012028 2.1241e-005 0.0011544 0.17791 0.00065873 0.17856 0.16349 0 0.03528 0.0389 0 0.93885 0.26849 0.07375 0.010175 4.4726 0.063494 7.6723e-005 0.82658 0.0054887 0.0062298 0.0014018 0.98674 0.99157 3.0247e-006 1.2099e-005 0.13364 0.8963 0.89135 0.0014053 0.97461 0.55467 0.0018929 0.42658 1.7345 1.7333 16.009 144.9849 0.00020409 -85.5851 0.51195
1.616 0.98803 5.5155e-005 3.8182 0.012028 2.1254e-005 0.0011544 0.17796 0.00065873 0.17861 0.16353 0 0.035277 0.0389 0 0.93893 0.26853 0.073765 0.010177 4.4731 0.063505 7.6736e-005 0.82657 0.0054892 0.0062303 0.0014017 0.98674 0.99157 3.0244e-006 1.2098e-005 0.13364 0.89657 0.89149 0.0014052 0.97475 0.55482 0.0018928 0.4266 1.7352 1.734 16.0089 144.9849 0.00020386 -85.5857 0.51295
1.617 0.98803 5.5155e-005 3.8182 0.012028 2.1267e-005 0.0011544 0.178 0.00065873 0.17866 0.16358 0 0.035275 0.0389 0 0.93902 0.26857 0.073779 0.010179 4.4737 0.063515 7.675e-005 0.82656 0.0054897 0.0062308 0.0014016 0.98675 0.99158 3.0241e-006 1.2096e-005 0.13365 0.89684 0.89164 0.0014051 0.9749 0.55498 0.0018928 0.42661 1.736 1.7348 16.0089 144.9849 0.00020364 -85.5862 0.51395
1.618 0.98803 5.5155e-005 3.8182 0.012028 2.128e-005 0.0011544 0.17805 0.00065873 0.1787 0.16362 0 0.035272 0.0389 0 0.93911 0.2686 0.073793 0.01018 4.4743 0.063526 7.6764e-005 0.82655 0.0054902 0.0062314 0.0014014 0.98675 0.99158 3.0238e-006 1.2095e-005 0.13365 0.89711 0.89178 0.0014051 0.97504 0.55513 0.0018927 0.42662 1.7367 1.7355 16.0089 144.985 0.00020341 -85.5868 0.51495
1.619 0.98803 5.5155e-005 3.8182 0.012028 2.1293e-005 0.0011544 0.17809 0.00065873 0.17875 0.16366 0 0.035269 0.0389 0 0.9392 0.26864 0.073807 0.010182 4.4748 0.063536 7.6777e-005 0.82654 0.0054907 0.0062319 0.0014013 0.98675 0.99158 3.0235e-006 1.2094e-005 0.13366 0.89738 0.89192 0.001405 0.97519 0.55529 0.0018926 0.42664 1.7375 1.7363 16.0089 144.985 0.00020319 -85.5874 0.51595
1.62 0.98803 5.5155e-005 3.8182 0.012028 2.1306e-005 0.0011544 0.17814 0.00065874 0.17879 0.16371 0 0.035267 0.0389 0 0.93929 0.26868 0.073821 0.010184 4.4754 0.063547 7.6791e-005 0.82653 0.0054913 0.0062325 0.0014012 0.98675 0.99158 3.0232e-006 1.2093e-005 0.13366 0.89765 0.89206 0.0014049 0.97533 0.55544 0.0018925 0.42665 1.7382 1.737 16.0089 144.985 0.00020297 -85.5879 0.51695
1.621 0.98803 5.5155e-005 3.8182 0.012028 2.1319e-005 0.0011544 0.17819 0.00065874 0.17884 0.16375 0 0.035264 0.0389 0 0.93937 0.26872 0.073835 0.010185 4.4759 0.063557 7.6805e-005 0.82652 0.0054918 0.006233 0.001401 0.98675 0.99158 3.0229e-006 1.2092e-005 0.13367 0.89792 0.8922 0.0014049 0.97547 0.5556 0.0018924 0.42666 1.7389 1.7377 16.0089 144.985 0.00020275 -85.5885 0.51795
1.622 0.98803 5.5155e-005 3.8182 0.012028 2.1332e-005 0.0011544 0.17823 0.00065874 0.17889 0.16379 0 0.035261 0.0389 0 0.93946 0.26876 0.07385 0.010187 4.4765 0.063568 7.6818e-005 0.82651 0.0054923 0.0062335 0.0014009 0.98675 0.99158 3.0226e-006 1.209e-005 0.13367 0.89818 0.89234 0.0014048 0.97561 0.55575 0.0018923 0.42667 1.7397 1.7385 16.0088 144.985 0.00020253 -85.589 0.51895
1.623 0.98803 5.5155e-005 3.8182 0.012028 2.1345e-005 0.0011544 0.17828 0.00065874 0.17893 0.16384 0 0.035258 0.0389 0 0.93955 0.2688 0.073864 0.010189 4.4771 0.063579 7.6832e-005 0.8265 0.0054928 0.0062341 0.0014008 0.98676 0.99158 3.0223e-006 1.2089e-005 0.13367 0.89845 0.89248 0.0014047 0.97575 0.5559 0.0018922 0.42669 1.7404 1.7392 16.0088 144.9851 0.00020231 -85.5896 0.51995
1.624 0.98803 5.5155e-005 3.8182 0.012028 2.1359e-005 0.0011544 0.17832 0.00065874 0.17898 0.16388 0 0.035256 0.0389 0 0.93964 0.26884 0.073878 0.01019 4.4776 0.063589 7.6846e-005 0.82649 0.0054934 0.0062346 0.0014006 0.98676 0.99158 3.022e-006 1.2088e-005 0.13368 0.89872 0.89262 0.0014047 0.97589 0.55606 0.0018921 0.4267 1.7411 1.7399 16.0088 144.9851 0.0002021 -85.5901 0.52095
1.625 0.98803 5.5155e-005 3.8182 0.012028 2.1372e-005 0.0011544 0.17837 0.00065874 0.17902 0.16392 0 0.035253 0.0389 0 0.93973 0.26888 0.073892 0.010192 4.4782 0.0636 7.686e-005 0.82648 0.0054939 0.0062351 0.0014005 0.98676 0.99158 3.0217e-006 1.2087e-005 0.13368 0.89898 0.89275 0.0014046 0.97603 0.55621 0.001892 0.42671 1.7419 1.7407 16.0088 144.9851 0.00020188 -85.5907 0.52195
1.626 0.98803 5.5155e-005 3.8182 0.012028 2.1385e-005 0.0011544 0.17841 0.00065874 0.17907 0.16397 0 0.03525 0.0389 0 0.93981 0.26892 0.073906 0.010194 4.4788 0.06361 7.6873e-005 0.82647 0.0054944 0.0062357 0.0014004 0.98676 0.99159 3.0215e-006 1.2086e-005 0.13369 0.89924 0.89289 0.0014045 0.97616 0.55637 0.001892 0.42673 1.7426 1.7414 16.0088 144.9851 0.00020166 -85.5912 0.52295
1.627 0.98803 5.5155e-005 3.8182 0.012028 2.1398e-005 0.0011544 0.17846 0.00065874 0.17911 0.16401 0 0.035248 0.0389 0 0.9399 0.26896 0.073921 0.010195 4.4793 0.063621 7.6887e-005 0.82646 0.0054949 0.0062362 0.0014003 0.98676 0.99159 3.0212e-006 1.2085e-005 0.13369 0.89951 0.89303 0.0014045 0.9763 0.55652 0.0018919 0.42674 1.7433 1.7421 16.0088 144.9851 0.00020145 -85.5917 0.52395
1.628 0.98803 5.5154e-005 3.8182 0.012028 2.1411e-005 0.0011544 0.17851 0.00065874 0.17916 0.16405 0 0.035245 0.0389 0 0.93999 0.269 0.073935 0.010197 4.4799 0.063631 7.6901e-005 0.82645 0.0054955 0.0062367 0.0014001 0.98676 0.99159 3.0209e-006 1.2083e-005 0.1337 0.89977 0.89316 0.0014044 0.97643 0.55668 0.0018918 0.42675 1.744 1.7429 16.0088 144.9852 0.00020123 -85.5923 0.52495
1.629 0.98803 5.5154e-005 3.8182 0.012028 2.1424e-005 0.0011544 0.17855 0.00065874 0.17921 0.16409 0 0.035242 0.0389 0 0.94008 0.26904 0.073949 0.010199 4.4805 0.063642 7.6915e-005 0.82644 0.005496 0.0062373 0.0014 0.98677 0.99159 3.0206e-006 1.2082e-005 0.1337 0.90003 0.8933 0.0014043 0.97657 0.55683 0.0018917 0.42676 1.7448 1.7436 16.0087 144.9852 0.00020102 -85.5928 0.52595
1.63 0.98803 5.5154e-005 3.8182 0.012028 2.1437e-005 0.0011544 0.1786 0.00065874 0.17925 0.16414 0 0.03524 0.0389 0 0.94017 0.26908 0.073963 0.010201 4.481 0.063652 7.6928e-005 0.82642 0.0054965 0.0062378 0.0013999 0.98677 0.99159 3.0203e-006 1.2081e-005 0.1337 0.90029 0.89343 0.0014043 0.9767 0.55698 0.0018916 0.42678 1.7455 1.7443 16.0087 144.9852 0.00020081 -85.5933 0.52695
1.631 0.98803 5.5154e-005 3.8182 0.012028 2.145e-005 0.0011544 0.17864 0.00065874 0.1793 0.16418 0 0.035237 0.0389 0 0.94025 0.26912 0.073977 0.010202 4.4816 0.063663 7.6942e-005 0.82641 0.005497 0.0062384 0.0013998 0.98677 0.99159 3.02e-006 1.208e-005 0.13371 0.90055 0.89357 0.0014042 0.97683 0.55714 0.0018915 0.42679 1.7462 1.745 16.0087 144.9852 0.0002006 -85.5939 0.52795
1.632 0.98803 5.5154e-005 3.8182 0.012028 2.1464e-005 0.0011544 0.17869 0.00065874 0.17934 0.16422 0 0.035234 0.0389 0 0.94034 0.26916 0.073992 0.010204 4.4822 0.063673 7.6956e-005 0.8264 0.0054976 0.0062389 0.0013997 0.98677 0.99159 3.0198e-006 1.2079e-005 0.13371 0.90081 0.8937 0.0014041 0.97697 0.55729 0.0018914 0.4268 1.7469 1.7458 16.0087 144.9852 0.00020038 -85.5944 0.52895
1.633 0.98803 5.5154e-005 3.8182 0.012028 2.1477e-005 0.0011544 0.17873 0.00065874 0.17939 0.16427 0 0.035232 0.0389 0 0.94043 0.2692 0.074006 0.010206 4.4827 0.063684 7.6969e-005 0.82639 0.0054981 0.0062394 0.0013995 0.98677 0.99159 3.0195e-006 1.2078e-005 0.13372 0.90107 0.89384 0.0014041 0.9771 0.55744 0.0018914 0.42682 1.7476 1.7465 16.0087 144.9853 0.00020017 -85.5949 0.52995
1.634 0.98803 5.5154e-005 3.8182 0.012028 2.149e-005 0.0011544 0.17878 0.00065874 0.17943 0.16431 0 0.035229 0.0389 0 0.94052 0.26924 0.07402 0.010207 4.4833 0.063695 7.6983e-005 0.82638 0.0054986 0.00624 0.0013994 0.98677 0.99159 3.0192e-006 1.2077e-005 0.13372 0.90133 0.89397 0.001404 0.97723 0.5576 0.0018913 0.42683 1.7483 1.7472 16.0087 144.9853 0.00019996 -85.5954 0.53095
1.635 0.98803 5.5154e-005 3.8182 0.012028 2.1503e-005 0.0011544 0.17883 0.00065874 0.17948 0.16435 0 0.035226 0.0389 0 0.94061 0.26927 0.074034 0.010209 4.4839 0.063705 7.6997e-005 0.82637 0.0054991 0.0062405 0.0013993 0.98678 0.99159 3.0189e-006 1.2076e-005 0.13373 0.90158 0.8941 0.0014039 0.97736 0.55775 0.0018912 0.42684 1.7491 1.7479 16.0086 144.9853 0.00019976 -85.5959 0.53195
1.636 0.98803 5.5154e-005 3.8182 0.012028 2.1516e-005 0.0011544 0.17887 0.00065875 0.17952 0.16439 0 0.035224 0.0389 0 0.94069 0.26931 0.074048 0.010211 4.4844 0.063716 7.7011e-005 0.82636 0.0054997 0.0062411 0.0013992 0.98678 0.9916 3.0187e-006 1.2075e-005 0.13373 0.90184 0.89424 0.0014039 0.97748 0.55791 0.0018911 0.42685 1.7498 1.7486 16.0086 144.9853 0.00019955 -85.5964 0.53295
1.637 0.98803 5.5154e-005 3.8182 0.012028 2.1529e-005 0.0011544 0.17892 0.00065875 0.17957 0.16444 0 0.035221 0.0389 0 0.94078 0.26935 0.074063 0.010212 4.485 0.063726 7.7024e-005 0.82635 0.0055002 0.0062416 0.0013991 0.98678 0.9916 3.0184e-006 1.2074e-005 0.13374 0.90209 0.89437 0.0014038 0.97761 0.55806 0.001891 0.42687 1.7505 1.7493 16.0086 144.9853 0.00019934 -85.5969 0.53395
1.638 0.98803 5.5154e-005 3.8182 0.012028 2.1542e-005 0.0011544 0.17896 0.00065875 0.17962 0.16448 0 0.035218 0.0389 0 0.94087 0.26939 0.074077 0.010214 4.4856 0.063737 7.7038e-005 0.82634 0.0055007 0.0062421 0.0013989 0.98678 0.9916 3.0181e-006 1.2072e-005 0.13374 0.90235 0.8945 0.0014038 0.97774 0.55821 0.001891 0.42688 1.7512 1.75 16.0086 144.9854 0.00019913 -85.5974 0.53495
1.639 0.98803 5.5154e-005 3.8182 0.012028 2.1555e-005 0.0011544 0.17901 0.00065875 0.17966 0.16452 0 0.035216 0.0389 0 0.94096 0.26943 0.074091 0.010216 4.4862 0.063747 7.7052e-005 0.82633 0.0055013 0.0062427 0.0013988 0.98678 0.9916 3.0179e-006 1.2071e-005 0.13374 0.9026 0.89463 0.0014037 0.97786 0.55837 0.0018909 0.42689 1.7519 1.7507 16.0086 144.9854 0.00019893 -85.5979 0.53595
1.64 0.98803 5.5154e-005 3.8182 0.012028 2.1568e-005 0.0011544 0.17905 0.00065875 0.17971 0.16457 0 0.035213 0.0389 0 0.94105 0.26947 0.074105 0.010218 4.4867 0.063758 7.7066e-005 0.82632 0.0055018 0.0062432 0.0013987 0.98678 0.9916 3.0176e-006 1.207e-005 0.13375 0.90286 0.89476 0.0014036 0.97799 0.55852 0.0018908 0.42691 1.7526 1.7514 16.0086 144.9854 0.00019872 -85.5984 0.53695
1.641 0.98803 5.5154e-005 3.8182 0.012028 2.1582e-005 0.0011544 0.1791 0.00065875 0.17975 0.16461 0 0.03521 0.0389 0 0.94114 0.26951 0.07412 0.010219 4.4873 0.063768 7.7079e-005 0.82631 0.0055023 0.0062438 0.0013986 0.98678 0.9916 3.0174e-006 1.2069e-005 0.13375 0.90311 0.89489 0.0014036 0.97811 0.55867 0.0018907 0.42692 1.7533 1.7521 16.0085 144.9854 0.00019852 -85.5989 0.53795
1.642 0.98803 5.5154e-005 3.8182 0.012028 2.1595e-005 0.0011544 0.17914 0.00065875 0.1798 0.16465 0 0.035208 0.0389 0 0.94122 0.26955 0.074134 0.010221 4.4879 0.063779 7.7093e-005 0.8263 0.0055028 0.0062443 0.0013985 0.98679 0.9916 3.0171e-006 1.2068e-005 0.13376 0.90336 0.89502 0.0014035 0.97824 0.55883 0.0018906 0.42693 1.754 1.7528 16.0085 144.9854 0.00019832 -85.5994 0.53895
1.643 0.98803 5.5154e-005 3.8182 0.012028 2.1608e-005 0.0011544 0.17919 0.00065875 0.17984 0.16469 0 0.035205 0.0389 0 0.94131 0.26959 0.074148 0.010223 4.4885 0.06379 7.7107e-005 0.82629 0.0055034 0.0062449 0.0013984 0.98679 0.9916 3.0168e-006 1.2067e-005 0.13376 0.90361 0.89515 0.0014035 0.97836 0.55898 0.0018906 0.42694 1.7547 1.7535 16.0085 144.9855 0.00019811 -85.5998 0.53995
1.644 0.98803 5.5153e-005 3.8182 0.012028 2.1621e-005 0.0011544 0.17923 0.00065875 0.17989 0.16474 0 0.035202 0.0389 0 0.9414 0.26963 0.074162 0.010224 4.489 0.0638 7.7121e-005 0.82628 0.0055039 0.0062454 0.0013983 0.98679 0.9916 3.0166e-006 1.2066e-005 0.13377 0.90386 0.89528 0.0014034 0.97848 0.55913 0.0018905 0.42696 1.7554 1.7542 16.0085 144.9855 0.00019791 -85.6003 0.54095
1.645 0.98803 5.5153e-005 3.8182 0.012028 2.1634e-005 0.0011544 0.17928 0.00065875 0.17993 0.16478 0 0.0352 0.0389 0 0.94149 0.26967 0.074177 0.010226 4.4896 0.063811 7.7135e-005 0.82627 0.0055044 0.0062459 0.0013982 0.98679 0.9916 3.0163e-006 1.2065e-005 0.13377 0.90411 0.8954 0.0014033 0.9786 0.55929 0.0018904 0.42697 1.7561 1.7549 16.0085 144.9855 0.00019771 -85.6008 0.54195
1.646 0.98803 5.5153e-005 3.8182 0.012028 2.1647e-005 0.0011544 0.17932 0.00065875 0.17998 0.16482 0 0.035197 0.0389 0 0.94158 0.26971 0.074191 0.010228 4.4902 0.063821 7.7148e-005 0.82626 0.005505 0.0062465 0.001398 0.98679 0.99161 3.0161e-006 1.2064e-005 0.13377 0.90435 0.89553 0.0014033 0.97872 0.55944 0.0018903 0.42698 1.7568 1.7556 16.0085 144.9855 0.00019751 -85.6013 0.54295
1.647 0.98803 5.5153e-005 3.8182 0.012028 2.166e-005 0.0011544 0.17937 0.00065875 0.18002 0.16486 0 0.035194 0.0389 0 0.94167 0.26975 0.074205 0.010229 4.4907 0.063832 7.7162e-005 0.82625 0.0055055 0.006247 0.0013979 0.98679 0.99161 3.0158e-006 1.2063e-005 0.13378 0.9046 0.89566 0.0014032 0.97884 0.55959 0.0018903 0.427 1.7574 1.7563 16.0084 144.9855 0.00019731 -85.6017 0.54395
1.648 0.98803 5.5153e-005 3.8182 0.012028 2.1673e-005 0.0011544 0.17941 0.00065875 0.18007 0.1649 0 0.035192 0.0389 0 0.94175 0.26979 0.074219 0.010231 4.4913 0.063843 7.7176e-005 0.82623 0.005506 0.0062476 0.0013978 0.98679 0.99161 3.0156e-006 1.2062e-005 0.13378 0.90485 0.89578 0.0014032 0.97896 0.55975 0.0018902 0.42701 1.7581 1.757 16.0084 144.9856 0.00019711 -85.6022 0.54495
1.649 0.98803 5.5153e-005 3.8182 0.012028 2.1686e-005 0.0011544 0.17946 0.00065875 0.18011 0.16495 0 0.035189 0.0389 0 0.94184 0.26983 0.074234 0.010233 4.4919 0.063853 7.719e-005 0.82622 0.0055066 0.0062481 0.0013977 0.9868 0.99161 3.0153e-006 1.2061e-005 0.13379 0.90509 0.89591 0.0014031 0.97908 0.5599 0.0018901 0.42702 1.7588 1.7577 16.0084 144.9856 0.00019691 -85.6027 0.54595
1.65 0.98803 5.5153e-005 3.8182 0.012028 2.17e-005 0.0011544 0.1795 0.00065875 0.18016 0.16499 0 0.035186 0.0389 0 0.94193 0.26987 0.074248 0.010234 4.4925 0.063864 7.7203e-005 0.82621 0.0055071 0.0062487 0.0013976 0.9868 0.99161 3.0151e-006 1.206e-005 0.13379 0.90534 0.89603 0.0014031 0.9792 0.56005 0.00189 0.42703 1.7595 1.7584 16.0084 144.9856 0.00019672 -85.6031 0.54695
1.651 0.98803 5.5153e-005 3.8182 0.012028 2.1713e-005 0.0011544 0.17955 0.00065875 0.1802 0.16503 0 0.035184 0.0389 0 0.94202 0.26991 0.074262 0.010236 4.4931 0.063874 7.7217e-005 0.8262 0.0055076 0.0062492 0.0013975 0.9868 0.99161 3.0148e-006 1.2059e-005 0.1338 0.90558 0.89616 0.001403 0.97931 0.56021 0.00189 0.42705 1.7602 1.7591 16.0084 144.9856 0.00019652 -85.6036 0.54795
1.652 0.98803 5.5153e-005 3.8182 0.012028 2.1726e-005 0.0011544 0.17959 0.00065875 0.18025 0.16507 0 0.035181 0.0389 0 0.94211 0.26995 0.074276 0.010238 4.4936 0.063885 7.7231e-005 0.82619 0.0055081 0.0062498 0.0013974 0.9868 0.99161 3.0146e-006 1.2058e-005 0.1338 0.90583 0.89628 0.0014029 0.97943 0.56036 0.0018899 0.42706 1.7609 1.7598 16.0084 144.9856 0.00019632 -85.604 0.54895
1.653 0.98803 5.5153e-005 3.8182 0.012028 2.1739e-005 0.0011544 0.17964 0.00065876 0.18029 0.16512 0 0.035179 0.0389 0 0.9422 0.26999 0.074291 0.01024 4.4942 0.063895 7.7245e-005 0.82618 0.0055087 0.0062503 0.0013973 0.9868 0.99161 3.0144e-006 1.2057e-005 0.13381 0.90607 0.89641 0.0014029 0.97954 0.56051 0.0018898 0.42707 1.7615 1.7604 16.0083 144.9857 0.00019613 -85.6045 0.54995
1.654 0.98803 5.5153e-005 3.8182 0.012028 2.1752e-005 0.0011544 0.17968 0.00065876 0.18034 0.16516 0 0.035176 0.0389 0 0.94229 0.27003 0.074305 0.010241 4.4948 0.063906 7.7259e-005 0.82617 0.0055092 0.0062509 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.13381 0.90631 0.89653 0.0014028 0.97966 0.56066 0.0018897 0.42709 1.7622 1.7611 16.0083 144.9857 0.00019593 -85.6049 0.55095
1.655 0.98803 5.5153e-005 3.8182 0.012028 2.1765e-005 0.0011544 0.17973 0.00065876 0.18038 0.1652 0 0.035173 0.0389 0 0.94237 0.27007 0.074319 0.010243 4.4954 0.063917 7.7272e-005 0.82616 0.0055097 0.0062514 0.0013971 0.9868 0.99161 3.0139e-006 1.2055e-005 0.13381 0.90655 0.89666 0.0014028 0.97977 0.56082 0.0018897 0.4271 1.7629 1.7618 16.0083 144.9857 0.00019574 -85.6054 0.55195
1.656 0.98803 5.5153e-005 3.8182 0.012028 2.1778e-005 0.0011544 0.17977 0.00065876 0.18043 0.16524 0 0.035171 0.0389 0 0.94246 0.27011 0.074334 0.010245 4.4959 0.063927 7.7286e-005 0.82615 0.0055103 0.0062519 0.001397 0.98681 0.99161 3.0137e-006 1.2055e-005 0.13382 0.90679 0.89678 0.0014027 0.97988 0.56097 0.0018896 0.42711 1.7636 1.7625 16.0083 144.9857 0.00019555 -85.6058 0.55295
1.657 0.98803 5.5153e-005 3.8182 0.012028 2.1791e-005 0.0011544 0.17982 0.00065876 0.18047 0.16528 0 0.035168 0.0389 0 0.94255 0.27015 0.074348 0.010246 4.4965 0.063938 7.73e-005 0.82614 0.0055108 0.0062525 0.0013969 0.98681 0.99162 3.0134e-006 1.2054e-005 0.13382 0.90703 0.8969 0.0014027 0.98 0.56112 0.0018895 0.42712 1.7642 1.7632 16.0083 144.9857 0.00019536 -85.6062 0.55395
1.658 0.98803 5.5153e-005 3.8182 0.012028 2.1805e-005 0.0011544 0.17986 0.00065876 0.18052 0.16533 0 0.035166 0.0389 0 0.94264 0.27019 0.074362 0.010248 4.4971 0.063948 7.7314e-005 0.82613 0.0055113 0.006253 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.13383 0.90727 0.89702 0.0014026 0.98011 0.56127 0.0018895 0.42714 1.7649 1.7638 16.0083 144.9858 0.00019516 -85.6067 0.55495
1.659 0.98803 5.5152e-005 3.8182 0.012028 2.1818e-005 0.0011544 0.17991 0.00065876 0.18056 0.16537 0 0.035163 0.0389 0 0.94273 0.27022 0.074376 0.01025 4.4977 0.063959 7.7328e-005 0.82612 0.0055119 0.0062536 0.0013967 0.98681 0.99162 3.013e-006 1.2052e-005 0.13383 0.90751 0.89714 0.0014026 0.98022 0.56143 0.0018894 0.42715 1.7656 1.7645 16.0082 144.9858 0.00019497 -85.6071 0.55595
1.66 0.98803 5.5152e-005 3.8182 0.012028 2.1831e-005 0.0011544 0.17995 0.00065876 0.1806 0.16541 0 0.03516 0.0389 0 0.94282 0.27026 0.074391 0.010252 4.4983 0.06397 7.7341e-005 0.82611 0.0055124 0.0062541 0.0013966 0.98681 0.99162 3.0127e-006 1.2051e-005 0.13384 0.90775 0.89726 0.0014025 0.98033 0.56158 0.0018893 0.42716 1.7663 1.7652 16.0082 144.9858 0.00019478 -85.6075 0.55695
1.661 0.98803 5.5152e-005 3.8182 0.012028 2.1844e-005 0.0011544 0.17999 0.00065876 0.18065 0.16545 0 0.035158 0.0389 0 0.94291 0.2703 0.074405 0.010253 4.4989 0.06398 7.7355e-005 0.8261 0.0055129 0.0062547 0.0013965 0.98681 0.99162 3.0125e-006 1.205e-005 0.13384 0.90798 0.89738 0.0014025 0.98044 0.56173 0.0018893 0.42718 1.7669 1.7658 16.0082 144.9858 0.00019459 -85.608 0.55795
1.662 0.98803 5.5152e-005 3.8182 0.012028 2.1857e-005 0.0011544 0.18004 0.00065876 0.18069 0.16549 0 0.035155 0.0389 0 0.94299 0.27034 0.074419 0.010255 4.4994 0.063991 7.7369e-005 0.82609 0.0055135 0.0062552 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.13385 0.90822 0.8975 0.0014024 0.98054 0.56188 0.0018892 0.42719 1.7676 1.7665 16.0082 144.9858 0.0001944 -85.6084 0.55895
1.663 0.98803 5.5152e-005 3.8182 0.012028 2.187e-005 0.0011544 0.18008 0.00065876 0.18074 0.16554 0 0.035152 0.0389 0 0.94308 0.27038 0.074434 0.010257 4.5 0.064001 7.7383e-005 0.82608 0.005514 0.0062558 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.13385 0.90845 0.89762 0.0014024 0.98065 0.56204 0.0018891 0.4272 1.7683 1.7672 16.0082 144.9859 0.00019422 -85.6088 0.55995
1.664 0.98803 5.5152e-005 3.8182 0.012028 2.1883e-005 0.0011544 0.18013 0.00065876 0.18078 0.16558 0 0.03515 0.0389 0 0.94317 0.27042 0.074448 0.010258 4.5006 0.064012 7.7397e-005 0.82607 0.0055145 0.0062563 0.0013962 0.98682 0.99162 3.0118e-006 1.2047e-005 0.13385 0.90869 0.89774 0.0014023 0.98076 0.56219 0.0018891 0.42721 1.7689 1.7678 16.0081 144.9859 0.00019403 -85.6092 0.56095
1.665 0.98803 5.5152e-005 3.8182 0.012028 2.1896e-005 0.0011544 0.18017 0.00065876 0.18083 0.16562 0 0.035147 0.0389 0 0.94326 0.27046 0.074462 0.01026 4.5012 0.064023 7.741e-005 0.82605 0.0055151 0.0062569 0.0013961 0.98682 0.99162 3.0116e-006 1.2046e-005 0.13386 0.90892 0.89786 0.0014023 0.98087 0.56234 0.001889 0.42723 1.7696 1.7685 16.0081 144.9859 0.00019384 -85.6096 0.56195
1.666 0.98803 5.5152e-005 3.8182 0.012028 2.1909e-005 0.0011544 0.18022 0.00065876 0.18087 0.16566 0 0.035145 0.0389 0 0.94335 0.2705 0.074476 0.010262 4.5018 0.064033 7.7424e-005 0.82604 0.0055156 0.0062574 0.001396 0.98682 0.99162 3.0114e-006 1.2046e-005 0.13386 0.90916 0.89798 0.0014022 0.98097 0.56249 0.0018889 0.42724 1.7702 1.7692 16.0081 144.9859 0.00019366 -85.6101 0.56295
1.667 0.98803 5.5152e-005 3.8182 0.012028 2.1923e-005 0.0011544 0.18026 0.00065876 0.18092 0.1657 0 0.035142 0.0389 0 0.94344 0.27054 0.074491 0.010263 4.5024 0.064044 7.7438e-005 0.82603 0.0055162 0.006258 0.0013959 0.98682 0.99162 3.0112e-006 1.2045e-005 0.13387 0.90939 0.8981 0.0014022 0.98108 0.56264 0.0018889 0.42725 1.7709 1.7698 16.0081 144.9859 0.00019347 -85.6105 0.56395
1.668 0.98803 5.5152e-005 3.8182 0.012028 2.1936e-005 0.0011544 0.18031 0.00065876 0.18096 0.16574 0 0.03514 0.0389 0 0.94353 0.27058 0.074505 0.010265 4.5029 0.064054 7.7452e-005 0.82602 0.0055167 0.0062585 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.13387 0.90962 0.89822 0.0014021 0.98118 0.5628 0.0018888 0.42727 1.7715 1.7705 16.0081 144.986 0.00019329 -85.6109 0.56495
1.669 0.98803 5.5152e-005 3.8182 0.012028 2.1949e-005 0.0011544 0.18035 0.00065876 0.181 0.16579 0 0.035137 0.0389 0 0.94362 0.27062 0.074519 0.010267 4.5035 0.064065 7.7466e-005 0.82601 0.0055172 0.0062591 0.0013957 0.98682 0.99162 3.0107e-006 1.2043e-005 0.13388 0.90985 0.89833 0.0014021 0.98128 0.56295 0.0018887 0.42728 1.7722 1.7711 16.0081 144.986 0.0001931 -85.6113 0.56595
1.67 0.98803 5.5152e-005 3.8182 0.012028 2.1962e-005 0.0011545 0.18039 0.00065877 0.18105 0.16583 0 0.035134 0.0389 0 0.9437 0.27066 0.074534 0.010269 4.5041 0.064076 7.748e-005 0.826 0.0055178 0.0062596 0.0013956 0.98682 0.99163 3.0105e-006 1.2042e-005 0.13388 0.91008 0.89845 0.001402 0.98139 0.5631 0.0018887 0.42729 1.7728 1.7718 16.008 144.986 0.00019292 -85.6117 0.56695
1.671 0.98803 5.5152e-005 3.8182 0.012028 2.1975e-005 0.0011545 0.18044 0.00065877 0.18109 0.16587 0 0.035132 0.0389 0 0.94379 0.2707 0.074548 0.01027 4.5047 0.064086 7.7493e-005 0.82599 0.0055183 0.0062602 0.0013955 0.98682 0.99163 3.0103e-006 1.2041e-005 0.13389 0.91031 0.89857 0.001402 0.98149 0.56325 0.0018886 0.4273 1.7735 1.7725 16.008 144.986 0.00019274 -85.6121 0.56795
1.672 0.98803 5.5152e-005 3.8182 0.012028 2.1988e-005 0.0011545 0.18048 0.00065877 0.18114 0.16591 0 0.035129 0.0389 0 0.94388 0.27074 0.074562 0.010272 4.5053 0.064097 7.7507e-005 0.82598 0.0055188 0.0062607 0.0013954 0.98683 0.99163 3.0101e-006 1.204e-005 0.13389 0.91054 0.89868 0.0014019 0.98159 0.5634 0.0018885 0.42732 1.7741 1.7731 16.008 144.986 0.00019256 -85.6125 0.56895
1.673 0.98803 5.5152e-005 3.8182 0.012028 2.2001e-005 0.0011545 0.18053 0.00065877 0.18118 0.16595 0 0.035127 0.0389 0 0.94397 0.27078 0.074577 0.010274 4.5059 0.064108 7.7521e-005 0.82597 0.0055194 0.0062613 0.0013953 0.98683 0.99163 3.0099e-006 1.204e-005 0.13389 0.91077 0.8988 0.0014019 0.98169 0.56356 0.0018885 0.42733 1.7748 1.7738 16.008 144.9861 0.00019237 -85.6129 0.56995
1.674 0.98803 5.5152e-005 3.8182 0.012028 2.2014e-005 0.0011545 0.18057 0.00065877 0.18122 0.16599 0 0.035124 0.0389 0 0.94406 0.27082 0.074591 0.010275 4.5065 0.064118 7.7535e-005 0.82596 0.0055199 0.0062618 0.0013953 0.98683 0.99163 3.0097e-006 1.2039e-005 0.1339 0.91099 0.89891 0.0014018 0.98179 0.56371 0.0018884 0.42734 1.7754 1.7744 16.008 144.9861 0.00019219 -85.6133 0.57095
1.675 0.98803 5.5151e-005 3.8182 0.012028 2.2027e-005 0.0011545 0.18061 0.00065877 0.18127 0.16604 0 0.035121 0.0389 0 0.94415 0.27086 0.074605 0.010277 4.507 0.064129 7.7549e-005 0.82595 0.0055204 0.0062624 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.1339 0.91122 0.89903 0.0014018 0.98189 0.56386 0.0018884 0.42736 1.7761 1.7751 16.0079 144.9861 0.00019201 -85.6136 0.57195
1.676 0.98803 5.5151e-005 3.8182 0.012028 2.2041e-005 0.0011545 0.18066 0.00065877 0.18131 0.16608 0 0.035119 0.0389 0 0.94424 0.2709 0.07462 0.010279 4.5076 0.064139 7.7563e-005 0.82594 0.005521 0.0062629 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.13391 0.91145 0.89914 0.0014017 0.98199 0.56401 0.0018883 0.42737 1.7767 1.7757 16.0079 144.9861 0.00019184 -85.614 0.57295
1.677 0.98803 5.5151e-005 3.8182 0.012027 2.2054e-005 0.0011545 0.1807 0.00065877 0.18136 0.16612 0 0.035116 0.0389 0 0.94433 0.27094 0.074634 0.010281 4.5082 0.06415 7.7576e-005 0.82593 0.0055215 0.0062635 0.001395 0.98683 0.99163 3.0091e-006 1.2036e-005 0.13391 0.91167 0.89925 0.0014017 0.98209 0.56416 0.0018882 0.42738 1.7774 1.7763 16.0079 144.9861 0.00019166 -85.6144 0.57395
1.678 0.98803 5.5151e-005 3.8182 0.012027 2.2067e-005 0.0011545 0.18075 0.00065877 0.1814 0.16616 0 0.035114 0.0389 0 0.94441 0.27098 0.074648 0.010282 4.5088 0.064161 7.759e-005 0.82592 0.0055221 0.006264 0.0013949 0.98683 0.99163 3.0089e-006 1.2035e-005 0.13392 0.9119 0.89937 0.0014016 0.98219 0.56431 0.0018882 0.42739 1.778 1.777 16.0079 144.9862 0.00019148 -85.6148 0.57495
1.679 0.98803 5.5151e-005 3.8182 0.012027 2.208e-005 0.0011545 0.18079 0.00065877 0.18144 0.1662 0 0.035111 0.0389 0 0.9445 0.27102 0.074663 0.010284 4.5094 0.064171 7.7604e-005 0.82591 0.0055226 0.0062646 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.13392 0.91212 0.89948 0.0014016 0.98229 0.56447 0.0018881 0.42741 1.7786 1.7776 16.0079 144.9862 0.0001913 -85.6152 0.57595
1.68 0.98803 5.5151e-005 3.8182 0.012027 2.2093e-005 0.0011545 0.18083 0.00065877 0.18149 0.16624 0 0.035109 0.0389 0 0.94459 0.27106 0.074677 0.010286 4.51 0.064182 7.7618e-005 0.8259 0.0055231 0.0062652 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.13393 0.91234 0.89959 0.0014015 0.98238 0.56462 0.001888 0.42742 1.7793 1.7783 16.0078 144.9862 0.00019113 -85.6155 0.57695
1.681 0.98803 5.5151e-005 3.8182 0.012027 2.2106e-005 0.0011545 0.18088 0.00065877 0.18153 0.16628 0 0.035106 0.0389 0 0.94468 0.2711 0.074691 0.010287 4.5106 0.064193 7.7632e-005 0.82589 0.0055237 0.0062657 0.0013946 0.98684 0.99163 3.0083e-006 1.2033e-005 0.13393 0.91256 0.8997 0.0014015 0.98248 0.56477 0.001888 0.42743 1.7799 1.7789 16.0078 144.9862 0.00019095 -85.6159 0.57795
1.682 0.98803 5.5151e-005 3.8182 0.012027 2.2119e-005 0.0011545 0.18092 0.00065877 0.18158 0.16633 0 0.035104 0.0389 0 0.94477 0.27114 0.074706 0.010289 4.5112 0.064203 7.7646e-005 0.82587 0.0055242 0.0062663 0.0013945 0.98684 0.99163 3.0081e-006 1.2032e-005 0.13393 0.91279 0.89982 0.0014014 0.98257 0.56492 0.0018879 0.42745 1.7806 1.7795 16.0078 144.9862 0.00019077 -85.6163 0.57895
1.683 0.98803 5.5151e-005 3.8182 0.012027 2.2132e-005 0.0011545 0.18097 0.00065877 0.18162 0.16637 0 0.035101 0.0389 0 0.94486 0.27118 0.07472 0.010291 4.5118 0.064214 7.766e-005 0.82586 0.0055248 0.0062668 0.0013945 0.98684 0.99164 3.0079e-006 1.2031e-005 0.13394 0.91301 0.89993 0.0014014 0.98267 0.56507 0.0018879 0.42746 1.7812 1.7802 16.0078 144.9863 0.0001906 -85.6166 0.57995
1.684 0.98803 5.5151e-005 3.8182 0.012027 2.2145e-005 0.0011545 0.18101 0.00065877 0.18166 0.16641 0 0.035098 0.0389 0 0.94495 0.27122 0.074734 0.010292 4.5124 0.064225 7.7673e-005 0.82585 0.0055253 0.0062674 0.0013944 0.98684 0.99164 3.0077e-006 1.2031e-005 0.13394 0.91323 0.90004 0.0014014 0.98276 0.56522 0.0018878 0.42747 1.7818 1.7808 16.0078 144.9863 0.00019043 -85.617 0.58095
1.685 0.98803 5.5151e-005 3.8182 0.012027 2.2159e-005 0.0011545 0.18105 0.00065877 0.18171 0.16645 0 0.035096 0.0389 0 0.94504 0.27126 0.074749 0.010294 4.5129 0.064235 7.7687e-005 0.82584 0.0055258 0.0062679 0.0013943 0.98684 0.99164 3.0075e-006 1.203e-005 0.13395 0.91345 0.90015 0.0014013 0.98286 0.56537 0.0018878 0.42748 1.7824 1.7814 16.0077 144.9863 0.00019025 -85.6174 0.58195
1.686 0.98803 5.5151e-005 3.8182 0.012027 2.2172e-005 0.0011545 0.1811 0.00065877 0.18175 0.16649 0 0.035093 0.0389 0 0.94513 0.2713 0.074763 0.010296 4.5135 0.064246 7.7701e-005 0.82583 0.0055264 0.0062685 0.0013942 0.98684 0.99164 3.0073e-006 1.2029e-005 0.13395 0.91367 0.90026 0.0014013 0.98295 0.56552 0.0018877 0.4275 1.7831 1.7821 16.0077 144.9863 0.00019008 -85.6177 0.58295
1.687 0.98803 5.5151e-005 3.8182 0.012027 2.2185e-005 0.0011545 0.18114 0.00065878 0.18179 0.16653 0 0.035091 0.0389 0 0.94522 0.27134 0.074777 0.010298 4.5141 0.064256 7.7715e-005 0.82582 0.0055269 0.006269 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.13396 0.91388 0.90037 0.0014012 0.98304 0.56568 0.0018876 0.42751 1.7837 1.7827 16.0077 144.9863 0.00018991 -85.6181 0.58395
1.688 0.98803 5.5151e-005 3.8182 0.012027 2.2198e-005 0.0011545 0.18118 0.00065878 0.18184 0.16657 0 0.035088 0.0389 0 0.9453 0.27138 0.074792 0.010299 4.5147 0.064267 7.7729e-005 0.82581 0.0055275 0.0062696 0.001394 0.98684 0.99164 3.0069e-006 1.2028e-005 0.13396 0.9141 0.90048 0.0014012 0.98313 0.56583 0.0018876 0.42752 1.7843 1.7833 16.0077 144.9864 0.00018974 -85.6184 0.58495
1.689 0.98803 5.5151e-005 3.8182 0.012027 2.2211e-005 0.0011545 0.18123 0.00065878 0.18188 0.16661 0 0.035086 0.0389 0 0.94539 0.27142 0.074806 0.010301 4.5153 0.064278 7.7743e-005 0.8258 0.005528 0.0062702 0.001394 0.98684 0.99164 3.0067e-006 1.2027e-005 0.13397 0.91432 0.90058 0.0014011 0.98322 0.56598 0.0018875 0.42754 1.7849 1.7839 16.0077 144.9864 0.00018957 -85.6188 0.58595
1.69 0.98803 5.515e-005 3.8182 0.012027 2.2224e-005 0.0011545 0.18127 0.00065878 0.18192 0.16665 0 0.035083 0.0389 0 0.94548 0.27146 0.074821 0.010303 4.5159 0.064288 7.7757e-005 0.82579 0.0055286 0.0062707 0.0013939 0.98685 0.99164 3.0066e-006 1.2026e-005 0.13397 0.91453 0.90069 0.0014011 0.98331 0.56613 0.0018875 0.42755 1.7856 1.7846 16.0076 144.9864 0.0001894 -85.6192 0.58695
1.691 0.98803 5.515e-005 3.8182 0.012027 2.2237e-005 0.0011545 0.18131 0.00065878 0.18197 0.16669 0 0.035081 0.0389 0 0.94557 0.2715 0.074835 0.010304 4.5165 0.064299 7.7771e-005 0.82578 0.0055291 0.0062713 0.0013938 0.98685 0.99164 3.0064e-006 1.2025e-005 0.13397 0.91475 0.9008 0.0014011 0.9834 0.56628 0.0018874 0.42756 1.7862 1.7852 16.0076 144.9864 0.00018923 -85.6195 0.58795
1.692 0.98803 5.515e-005 3.8182 0.012027 2.225e-005 0.0011545 0.18136 0.00065878 0.18201 0.16674 0 0.035078 0.0389 0 0.94566 0.27154 0.074849 0.010306 4.5171 0.06431 7.7784e-005 0.82577 0.0055296 0.0062718 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.13398 0.91496 0.90091 0.001401 0.98349 0.56643 0.0018874 0.42757 1.7868 1.7858 16.0076 144.9864 0.00018906 -85.6198 0.58895
1.693 0.98803 5.515e-005 3.8182 0.012027 2.2264e-005 0.0011545 0.1814 0.00065878 0.18205 0.16678 0 0.035076 0.0389 0 0.94575 0.27158 0.074864 0.010308 4.5177 0.06432 7.7798e-005 0.82576 0.0055302 0.0062724 0.0013936 0.98685 0.99164 3.006e-006 1.2024e-005 0.13398 0.91518 0.90102 0.001401 0.98358 0.56658 0.0018873 0.42759 1.7874 1.7864 16.0076 144.9865 0.00018889 -85.6202 0.58995
1.694 0.98803 5.515e-005 3.8182 0.012027 2.2277e-005 0.0011545 0.18144 0.00065878 0.1821 0.16682 0 0.035073 0.0389 0 0.94584 0.27162 0.074878 0.01031 4.5183 0.064331 7.7812e-005 0.82575 0.0055307 0.0062729 0.0013936 0.98685 0.99164 3.0058e-006 1.2023e-005 0.13399 0.91539 0.90112 0.0014009 0.98367 0.56673 0.0018872 0.4276 1.788 1.7871 16.0076 144.9865 0.00018872 -85.6205 0.59095
1.695 0.98803 5.515e-005 3.8182 0.012027 2.229e-005 0.0011545 0.18149 0.00065878 0.18214 0.16686 0 0.035071 0.0389 0 0.94593 0.27166 0.074893 0.010311 4.5189 0.064342 7.7826e-005 0.82574 0.0055313 0.0062735 0.0013935 0.98685 0.99164 3.0056e-006 1.2022e-005 0.13399 0.91561 0.90123 0.0014009 0.98376 0.56688 0.0018872 0.42761 1.7887 1.7877 16.0075 144.9865 0.00018855 -85.6209 0.59195
1.696 0.98803 5.515e-005 3.8182 0.012027 2.2303e-005 0.0011545 0.18153 0.00065878 0.18218 0.1669 0 0.035068 0.0389 0 0.94602 0.2717 0.074907 0.010313 4.5195 0.064352 7.784e-005 0.82573 0.0055318 0.0062741 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.134 0.91582 0.90133 0.0014008 0.98384 0.56703 0.0018871 0.42763 1.7893 1.7883 16.0075 144.9865 0.00018839 -85.6212 0.59295
1.697 0.98803 5.515e-005 3.8182 0.012027 2.2316e-005 0.0011545 0.18157 0.00065878 0.18223 0.16694 0 0.035065 0.0389 0 0.94611 0.27174 0.074921 0.010315 4.5201 0.064363 7.7854e-005 0.82571 0.0055324 0.0062746 0.0013933 0.98685 0.99164 3.0053e-006 1.2021e-005 0.134 0.91603 0.90144 0.0014008 0.98393 0.56718 0.0018871 0.42764 1.7899 1.7889 16.0075 144.9865 0.00018822 -85.6215 0.59395
1.698 0.98803 5.515e-005 3.8182 0.012027 2.2329e-005 0.0011545 0.18162 0.00065878 0.18227 0.16698 0 0.035063 0.0389 0 0.9462 0.27178 0.074936 0.010316 4.5207 0.064374 7.7868e-005 0.8257 0.0055329 0.0062752 0.0013932 0.98685 0.99165 3.0051e-006 1.202e-005 0.13401 0.91624 0.90155 0.0014008 0.98402 0.56733 0.001887 0.42765 1.7905 1.7895 16.0075 144.9866 0.00018806 -85.6219 0.59495
1.699 0.98803 5.515e-005 3.8182 0.012027 2.2342e-005 0.0011545 0.18166 0.00065878 0.18231 0.16702 0 0.03506 0.0389 0 0.94629 0.27182 0.07495 0.010318 4.5213 0.064384 7.7882e-005 0.82569 0.0055334 0.0062757 0.0013932 0.98685 0.99165 3.0049e-006 1.202e-005 0.13401 0.91645 0.90165 0.0014007 0.9841 0.56748 0.001887 0.42766 1.7911 1.7901 16.0075 144.9866 0.00018789 -85.6222 0.59595
1.7 0.98803 5.515e-005 3.8182 0.012027 2.2355e-005 0.0011545 0.1817 0.00065878 0.18236 0.16706 0 0.035058 0.0389 0 0.94637 0.27186 0.074964 0.01032 4.5219 0.064395 7.7896e-005 0.82568 0.005534 0.0062763 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.13401 0.91666 0.90175 0.0014007 0.98419 0.56763 0.0018869 0.42768 1.7917 1.7907 16.0074 144.9866 0.00018773 -85.6225 0.59695
1.701 0.98803 5.515e-005 3.8182 0.012027 2.2368e-005 0.0011545 0.18175 0.00065878 0.1824 0.1671 0 0.035055 0.0389 0 0.94646 0.2719 0.074979 0.010322 4.5225 0.064406 7.791e-005 0.82567 0.0055345 0.0062769 0.001393 0.98686 0.99165 3.0046e-006 1.2018e-005 0.13402 0.91687 0.90186 0.0014006 0.98427 0.56779 0.0018869 0.42769 1.7923 1.7913 16.0074 144.9866 0.00018756 -85.6229 0.59795
1.702 0.98803 5.515e-005 3.8182 0.012027 2.2382e-005 0.0011545 0.18179 0.00065878 0.18244 0.16714 0 0.035053 0.0389 0 0.94655 0.27194 0.074993 0.010323 4.5231 0.064416 7.7923e-005 0.82566 0.0055351 0.0062774 0.0013929 0.98686 0.99165 3.0044e-006 1.2018e-005 0.13402 0.91708 0.90196 0.0014006 0.98436 0.56794 0.0018868 0.4277 1.7929 1.792 16.0074 144.9866 0.0001874 -85.6232 0.59895
1.703 0.98803 5.515e-005 3.8182 0.012027 2.2395e-005 0.0011545 0.18183 0.00065878 0.18249 0.16718 0 0.03505 0.0389 0 0.94664 0.27198 0.075008 0.010325 4.5237 0.064427 7.7937e-005 0.82565 0.0055356 0.006278 0.0013929 0.98686 0.99165 3.0042e-006 1.2017e-005 0.13403 0.91728 0.90207 0.0014006 0.98444 0.56809 0.0018868 0.42772 1.7935 1.7926 16.0074 144.9867 0.00018724 -85.6235 0.59995
1.704 0.98803 5.515e-005 3.8182 0.012027 2.2408e-005 0.0011545 0.18188 0.00065878 0.18253 0.16722 0 0.035048 0.0389 0 0.94673 0.27202 0.075022 0.010327 4.5243 0.064438 7.7951e-005 0.82564 0.0055362 0.0062785 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.13403 0.91749 0.90217 0.0014005 0.98452 0.56824 0.0018867 0.42773 1.7941 1.7932 16.0074 144.9867 0.00018708 -85.6238 0.60095
1.705 0.98803 5.515e-005 3.8182 0.012027 2.2421e-005 0.0011545 0.18192 0.00065879 0.18257 0.16726 0 0.035045 0.0389 0 0.94682 0.27206 0.075037 0.010328 4.5249 0.064448 7.7965e-005 0.82563 0.0055367 0.0062791 0.0013927 0.98686 0.99165 3.0039e-006 1.2016e-005 0.13404 0.9177 0.90227 0.0014005 0.9846 0.56839 0.0018867 0.42774 1.7947 1.7938 16.0073 144.9867 0.00018692 -85.6241 0.60195
1.706 0.98803 5.5149e-005 3.8182 0.012027 2.2434e-005 0.0011545 0.18196 0.00065879 0.18262 0.1673 0 0.035043 0.0389 0 0.94691 0.2721 0.075051 0.01033 4.5255 0.064459 7.7979e-005 0.82562 0.0055373 0.0062797 0.0013926 0.98686 0.99165 3.0037e-006 1.2015e-005 0.13404 0.9179 0.90237 0.0014004 0.98469 0.56854 0.0018866 0.42775 1.7953 1.7944 16.0073 144.9867 0.00018676 -85.6245 0.60295
1.707 0.98803 5.5149e-005 3.8182 0.012027 2.2447e-005 0.0011545 0.182 0.00065879 0.18266 0.16734 0 0.03504 0.0389 0 0.947 0.27214 0.075065 0.010332 4.5261 0.06447 7.7993e-005 0.82561 0.0055378 0.0062802 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.13405 0.91811 0.90248 0.0014004 0.98477 0.56869 0.0018866 0.42777 1.7959 1.795 16.0073 144.9867 0.0001866 -85.6248 0.60395
1.708 0.98803 5.5149e-005 3.8182 0.012027 2.246e-005 0.0011545 0.18205 0.00065879 0.1827 0.16739 0 0.035038 0.0389 0 0.94709 0.27218 0.07508 0.010334 4.5267 0.06448 7.8007e-005 0.8256 0.0055384 0.0062808 0.0013925 0.98686 0.99165 3.0034e-006 1.2014e-005 0.13405 0.91831 0.90258 0.0014004 0.98485 0.56884 0.0018865 0.42778 1.7965 1.7956 16.0073 144.9868 0.00018644 -85.6251 0.60495
1.709 0.98803 5.5149e-005 3.8182 0.012027 2.2473e-005 0.0011545 0.18209 0.00065879 0.18274 0.16743 0 0.035035 0.0389 0 0.94718 0.27222 0.075094 0.010335 4.5273 0.064491 7.8021e-005 0.82559 0.0055389 0.0062813 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.13406 0.91852 0.90268 0.0014003 0.98493 0.56899 0.0018865 0.42779 1.7971 1.7962 16.0073 144.9868 0.00018628 -85.6254 0.60595
1.71 0.98803 5.5149e-005 3.8182 0.012027 2.2486e-005 0.0011545 0.18213 0.00065879 0.18279 0.16747 0 0.035033 0.0389 0 0.94727 0.27226 0.075109 0.010337 4.5279 0.064502 7.8035e-005 0.82558 0.0055394 0.0062819 0.0013924 0.98687 0.99165 3.0031e-006 1.2012e-005 0.13406 0.91872 0.90278 0.0014003 0.98501 0.56914 0.0018864 0.4278 1.7977 1.7968 16.0072 144.9868 0.00018612 -85.6257 0.60695
1.711 0.98803 5.5149e-005 3.8182 0.012027 2.25e-005 0.0011545 0.18218 0.00065879 0.18283 0.16751 0 0.03503 0.0389 0 0.94736 0.2723 0.075123 0.010339 4.5285 0.064512 7.8049e-005 0.82557 0.00554 0.0062825 0.0013923 0.98687 0.99165 3.0029e-006 1.2012e-005 0.13406 0.91892 0.90288 0.0014003 0.98509 0.56929 0.0018864 0.42782 1.7983 1.7974 16.0072 144.9868 0.00018596 -85.626 0.60795
1.712 0.98803 5.5149e-005 3.8182 0.012027 2.2513e-005 0.0011545 0.18222 0.00065879 0.18287 0.16755 0 0.035028 0.0389 0 0.94745 0.27234 0.075137 0.01034 4.5291 0.064523 7.8063e-005 0.82556 0.0055405 0.006283 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.13407 0.91912 0.90298 0.0014002 0.98516 0.56944 0.0018863 0.42783 1.7989 1.7979 16.0072 144.9868 0.0001858 -85.6263 0.60895
1.713 0.98803 5.5149e-005 3.8182 0.012027 2.2526e-005 0.0011545 0.18226 0.00065879 0.18292 0.16759 0 0.035025 0.0389 0 0.94754 0.27238 0.075152 0.010342 4.5297 0.064534 7.8077e-005 0.82554 0.0055411 0.0062836 0.0013921 0.98687 0.99165 3.0026e-006 1.201e-005 0.13407 0.91932 0.90308 0.0014002 0.98524 0.56959 0.0018863 0.42784 1.7995 1.7985 16.0072 144.9869 0.00018565 -85.6266 0.60995
1.714 0.98803 5.5149e-005 3.8182 0.012027 2.2539e-005 0.0011545 0.1823 0.00065879 0.18296 0.16763 0 0.035023 0.0389 0 0.94763 0.27242 0.075166 0.010344 4.5303 0.064544 7.8091e-005 0.82553 0.0055416 0.0062842 0.0013921 0.98687 0.99166 3.0024e-006 1.201e-005 0.13408 0.91953 0.90318 0.0014001 0.98532 0.56974 0.0018862 0.42786 1.8001 1.7991 16.0071 144.9869 0.00018549 -85.6269 0.61095
1.715 0.98803 5.5149e-005 3.8182 0.012027 2.2552e-005 0.0011545 0.18235 0.00065879 0.183 0.16767 0 0.035021 0.0389 0 0.94771 0.27246 0.075181 0.010346 4.5309 0.064555 7.8104e-005 0.82552 0.0055422 0.0062847 0.001392 0.98687 0.99166 3.0023e-006 1.2009e-005 0.13408 0.91973 0.90328 0.0014001 0.9854 0.56988 0.0018862 0.42787 1.8006 1.7997 16.0071 144.9869 0.00018534 -85.6272 0.61195
1.716 0.98803 5.5149e-005 3.8182 0.012027 2.2565e-005 0.0011545 0.18239 0.00065879 0.18304 0.16771 0 0.035018 0.0389 0 0.9478 0.2725 0.075195 0.010347 4.5315 0.064566 7.8118e-005 0.82551 0.0055427 0.0062853 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.13409 0.91992 0.90338 0.0014001 0.98547 0.57003 0.0018861 0.42788 1.8012 1.8003 16.0071 144.9869 0.00018518 -85.6275 0.61295
1.717 0.98803 5.5149e-005 3.8182 0.012027 2.2578e-005 0.0011545 0.18243 0.00065879 0.18309 0.16775 0 0.035016 0.0389 0 0.94789 0.27254 0.07521 0.010349 4.5321 0.064576 7.8132e-005 0.8255 0.0055433 0.0062859 0.0013919 0.98687 0.99166 3.002e-006 1.2008e-005 0.13409 0.92012 0.90347 0.0014 0.98555 0.57018 0.0018861 0.42789 1.8018 1.8009 16.0071 144.9869 0.00018503 -85.6278 0.61395
1.718 0.98803 5.5149e-005 3.8182 0.012027 2.2591e-005 0.0011545 0.18247 0.00065879 0.18313 0.16779 0 0.035013 0.0389 0 0.94798 0.27258 0.075224 0.010351 4.5328 0.064587 7.8146e-005 0.82549 0.0055438 0.0062864 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.1341 0.92032 0.90357 0.0014 0.98562 0.57033 0.001886 0.42791 1.8024 1.8015 16.0071 144.987 0.00018487 -85.6281 0.61495
1.719 0.98803 5.5149e-005 3.8182 0.012027 2.2604e-005 0.0011545 0.18252 0.00065879 0.18317 0.16783 0 0.035011 0.0389 0 0.94807 0.27262 0.075239 0.010352 4.5334 0.064598 7.816e-005 0.82548 0.0055444 0.006287 0.0013917 0.98687 0.99166 3.0017e-006 1.2007e-005 0.1341 0.92052 0.90367 0.0014 0.9857 0.57048 0.001886 0.42792 1.803 1.8021 16.007 144.987 0.00018472 -85.6284 0.61595
1.72 0.98803 5.5149e-005 3.8182 0.012027 2.2618e-005 0.0011545 0.18256 0.00065879 0.18321 0.16787 0 0.035008 0.0389 0 0.94816 0.27266 0.075253 0.010354 4.534 0.064609 7.8174e-005 0.82547 0.0055449 0.0062876 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.13411 0.92072 0.90377 0.0013999 0.98577 0.57063 0.0018859 0.42793 1.8036 1.8026 16.007 144.987 0.00018457 -85.6286 0.61695
1.721 0.98803 5.5148e-005 3.8182 0.012027 2.2631e-005 0.0011545 0.1826 0.00065879 0.18326 0.16791 0 0.035006 0.0389 0 0.94825 0.2727 0.075267 0.010356 4.5346 0.064619 7.8188e-005 0.82546 0.0055455 0.0062881 0.0013916 0.98687 0.99166 3.0014e-006 1.2005e-005 0.13411 0.92091 0.90386 0.0013999 0.98585 0.57078 0.0018859 0.42795 1.8041 1.8032 16.007 144.987 0.00018442 -85.6289 0.61795
1.722 0.98803 5.5148e-005 3.8182 0.012027 2.2644e-005 0.0011545 0.18264 0.00065879 0.1833 0.16795 0 0.035003 0.0389 0 0.94834 0.27274 0.075282 0.010358 4.5352 0.06463 7.8202e-005 0.82545 0.005546 0.0062887 0.0013915 0.98688 0.99166 3.0012e-006 1.2005e-005 0.13411 0.92111 0.90396 0.0013999 0.98592 0.57093 0.0018859 0.42796 1.8047 1.8038 16.007 144.987 0.00018426 -85.6292 0.61895
1.723 0.98803 5.5148e-005 3.8182 0.012027 2.2657e-005 0.0011545 0.18269 0.0006588 0.18334 0.16799 0 0.035001 0.0389 0 0.94843 0.27278 0.075296 0.010359 4.5358 0.064641 7.8216e-005 0.82544 0.0055466 0.0062892 0.0013915 0.98688 0.99166 3.0011e-006 1.2004e-005 0.13412 0.9213 0.90406 0.0013998 0.98599 0.57108 0.0018858 0.42797 1.8053 1.8044 16.0069 144.9871 0.00018411 -85.6295 0.61995
1.724 0.98803 5.5148e-005 3.8182 0.012027 2.267e-005 0.0011545 0.18273 0.0006588 0.18338 0.16803 0 0.034998 0.0389 0 0.94852 0.27282 0.075311 0.010361 4.5364 0.064651 7.823e-005 0.82543 0.0055471 0.0062898 0.0013914 0.98688 0.99166 3.0009e-006 1.2004e-005 0.13412 0.9215 0.90415 0.0013998 0.98607 0.57123 0.0018858 0.42798 1.8059 1.805 16.0069 144.9871 0.00018396 -85.6298 0.62095
1.725 0.98803 5.5148e-005 3.8182 0.012027 2.2683e-005 0.0011545 0.18277 0.0006588 0.18343 0.16807 0 0.034996 0.0389 0 0.94861 0.27286 0.075325 0.010363 4.537 0.064662 7.8244e-005 0.82542 0.0055477 0.0062904 0.0013913 0.98688 0.99166 3.0008e-006 1.2003e-005 0.13413 0.92169 0.90425 0.0013998 0.98614 0.57138 0.0018857 0.428 1.8064 1.8055 16.0069 144.9871 0.00018381 -85.6301 0.62195
1.726 0.98803 5.5148e-005 3.8182 0.012027 2.2696e-005 0.0011545 0.18281 0.0006588 0.18347 0.16811 0 0.034993 0.0389 0 0.9487 0.2729 0.07534 0.010364 4.5376 0.064673 7.8258e-005 0.82541 0.0055482 0.006291 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.13413 0.92188 0.90434 0.0013997 0.98621 0.57153 0.0018857 0.42801 1.807 1.8061 16.0069 144.9871 0.00018366 -85.6303 0.62295
1.727 0.98803 5.5148e-005 3.8182 0.012027 2.2709e-005 0.0011545 0.18286 0.0006588 0.18351 0.16815 0 0.034991 0.0389 0 0.94879 0.27294 0.075354 0.010366 4.5382 0.064683 7.8272e-005 0.82539 0.0055488 0.0062915 0.0013912 0.98688 0.99166 3.0005e-006 1.2002e-005 0.13414 0.92208 0.90444 0.0013997 0.98628 0.57168 0.0018856 0.42802 1.8076 1.8067 16.0069 144.9871 0.00018352 -85.6306 0.62395
1.728 0.98803 5.5148e-005 3.8182 0.012027 2.2722e-005 0.0011545 0.1829 0.0006588 0.18355 0.16819 0 0.034989 0.0389 0 0.94888 0.27298 0.075369 0.010368 4.5389 0.064694 7.8286e-005 0.82538 0.0055493 0.0062921 0.0013912 0.98688 0.99166 3.0003e-006 1.2001e-005 0.13414 0.92227 0.90453 0.0013997 0.98635 0.57183 0.0018856 0.42803 1.8081 1.8072 16.0068 144.9872 0.00018337 -85.6309 0.62495
1.729 0.98803 5.5148e-005 3.8182 0.012027 2.2736e-005 0.0011545 0.18294 0.0006588 0.18359 0.16823 0 0.034986 0.0389 0 0.94897 0.27302 0.075383 0.01037 4.5395 0.064705 7.83e-005 0.82537 0.0055499 0.0062927 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.13415 0.92246 0.90463 0.0013996 0.98642 0.57197 0.0018855 0.42805 1.8087 1.8078 16.0068 144.9872 0.00018322 -85.6311 0.62595
1.73 0.98803 5.5148e-005 3.8182 0.012027 2.2749e-005 0.0011545 0.18298 0.0006588 0.18364 0.16827 0 0.034984 0.0389 0 0.94906 0.27306 0.075398 0.010371 4.5401 0.064716 7.8314e-005 0.82536 0.0055504 0.0062932 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.13415 0.92265 0.90472 0.0013996 0.98649 0.57212 0.0018855 0.42806 1.8093 1.8084 16.0068 144.9872 0.00018307 -85.6314 0.62695
1.731 0.98803 5.5148e-005 3.8182 0.012027 2.2762e-005 0.0011545 0.18302 0.0006588 0.18368 0.16831 0 0.034981 0.0389 0 0.94915 0.2731 0.075412 0.010373 4.5407 0.064726 7.8328e-005 0.82535 0.005551 0.0062938 0.001391 0.98688 0.99166 2.9999e-006 1.1999e-005 0.13416 0.92284 0.90481 0.0013996 0.98656 0.57227 0.0018855 0.42807 1.8098 1.809 16.0068 144.9872 0.00018293 -85.6317 0.62795
1.732 0.98803 5.5148e-005 3.8182 0.012027 2.2775e-005 0.0011545 0.18307 0.0006588 0.18372 0.16834 0 0.034979 0.0389 0 0.94924 0.27314 0.075427 0.010375 4.5413 0.064737 7.8342e-005 0.82534 0.0055516 0.0062944 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.13416 0.92303 0.90491 0.0013995 0.98663 0.57242 0.0018854 0.42809 1.8104 1.8095 16.0067 144.9873 0.00018278 -85.6319 0.62895
1.733 0.98803 5.5148e-005 3.8182 0.012027 2.2788e-005 0.0011545 0.18311 0.0006588 0.18376 0.16838 0 0.034976 0.0389 0 0.94933 0.27318 0.075441 0.010376 4.5419 0.064748 7.8356e-005 0.82533 0.0055521 0.0062949 0.0013908 0.98688 0.99167 2.9996e-006 1.1998e-005 0.13416 0.92322 0.905 0.0013995 0.9867 0.57257 0.0018854 0.4281 1.811 1.8101 16.0067 144.9873 0.00018263 -85.6322 0.62995
1.734 0.98803 5.5148e-005 3.8182 0.012027 2.2801e-005 0.0011545 0.18315 0.0006588 0.1838 0.16842 0 0.034974 0.0389 0 0.94942 0.27322 0.075456 0.010378 4.5425 0.064758 7.837e-005 0.82532 0.0055527 0.0062955 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.13417 0.92341 0.90509 0.0013995 0.98677 0.57272 0.0018853 0.42811 1.8115 1.8106 16.0067 144.9873 0.00018249 -85.6325 0.63095
1.735 0.98803 5.5148e-005 3.8182 0.012027 2.2814e-005 0.0011545 0.18319 0.0006588 0.18385 0.16846 0 0.034971 0.0389 0 0.94951 0.27326 0.07547 0.01038 4.5432 0.064769 7.8384e-005 0.82531 0.0055532 0.0062961 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.13417 0.9236 0.90518 0.0013994 0.98684 0.57287 0.0018853 0.42812 1.8121 1.8112 16.0067 144.9873 0.00018234 -85.6327 0.63195
1.736 0.98803 5.5148e-005 3.8182 0.012027 2.2827e-005 0.0011545 0.18323 0.0006588 0.18389 0.1685 0 0.034969 0.0389 0 0.9496 0.2733 0.075485 0.010382 4.5438 0.06478 7.8398e-005 0.8253 0.0055538 0.0062966 0.0013907 0.98689 0.99167 2.9992e-006 1.1997e-005 0.13418 0.92378 0.90527 0.0013994 0.9869 0.57302 0.0018853 0.42814 1.8127 1.8118 16.0067 144.9873 0.0001822 -85.633 0.63295
1.737 0.98803 5.5147e-005 3.8182 0.012027 2.284e-005 0.0011545 0.18328 0.0006588 0.18393 0.16854 0 0.034967 0.0389 0 0.94969 0.27334 0.075499 0.010383 4.5444 0.064791 7.8412e-005 0.82529 0.0055543 0.0062972 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.13418 0.92397 0.90537 0.0013994 0.98697 0.57316 0.0018852 0.42815 1.8132 1.8123 16.0066 144.9874 0.00018206 -85.6332 0.63395
1.738 0.98803 5.5147e-005 3.8182 0.012027 2.2854e-005 0.0011545 0.18332 0.0006588 0.18397 0.16858 0 0.034964 0.0389 0 0.94978 0.27338 0.075514 0.010385 4.545 0.064801 7.8426e-005 0.82528 0.0055549 0.0062978 0.0013905 0.98689 0.99167 2.9989e-006 1.1996e-005 0.13419 0.92416 0.90546 0.0013993 0.98704 0.57331 0.0018852 0.42816 1.8138 1.8129 16.0066 144.9874 0.00018191 -85.6335 0.63495
1.739 0.98803 5.5147e-005 3.8182 0.012027 2.2867e-005 0.0011545 0.18336 0.0006588 0.18401 0.16862 0 0.034962 0.0389 0 0.94987 0.27342 0.075528 0.010387 4.5456 0.064812 7.844e-005 0.82527 0.0055554 0.0062983 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.13419 0.92434 0.90555 0.0013993 0.9871 0.57346 0.0018851 0.42817 1.8143 1.8134 16.0066 144.9874 0.00018177 -85.6337 0.63595
1.74 0.98803 5.5147e-005 3.8182 0.012027 2.288e-005 0.0011545 0.1834 0.0006588 0.18406 0.16866 0 0.034959 0.0389 0 0.94996 0.27346 0.075543 0.010389 4.5462 0.064823 7.8454e-005 0.82526 0.005556 0.0062989 0.0013904 0.98689 0.99167 2.9987e-006 1.1995e-005 0.1342 0.92453 0.90564 0.0013993 0.98717 0.57361 0.0018851 0.42819 1.8149 1.814 16.0066 144.9874 0.00018163 -85.634 0.63695
1.741 0.98803 5.5147e-005 3.8182 0.012027 2.2893e-005 0.0011545 0.18344 0.00065881 0.1841 0.1687 0 0.034957 0.0389 0 0.95005 0.2735 0.075557 0.01039 4.5469 0.064833 7.8468e-005 0.82524 0.0055565 0.0062995 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.1342 0.92471 0.90573 0.0013992 0.98723 0.57376 0.001885 0.4282 1.8154 1.8146 16.0065 144.9874 0.00018149 -85.6342 0.63795
1.742 0.98803 5.5147e-005 3.8182 0.012027 2.2906e-005 0.0011545 0.18348 0.00065881 0.18414 0.16874 0 0.034955 0.0389 0 0.95014 0.27354 0.075572 0.010392 4.5475 0.064844 7.8482e-005 0.82523 0.0055571 0.0063001 0.0013903 0.98689 0.99167 2.9984e-006 1.1994e-005 0.13421 0.92489 0.90582 0.0013992 0.9873 0.57391 0.001885 0.42821 1.816 1.8151 16.0065 144.9875 0.00018135 -85.6345 0.63895
1.743 0.98803 5.5147e-005 3.8182 0.012027 2.2919e-005 0.0011545 0.18353 0.00065881 0.18418 0.16878 0 0.034952 0.0389 0 0.95023 0.27359 0.075586 0.010394 4.5481 0.064855 7.8496e-005 0.82522 0.0055577 0.0063006 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.13421 0.92508 0.90591 0.0013992 0.98736 0.57405 0.001885 0.42822 1.8165 1.8157 16.0065 144.9875 0.00018121 -85.6347 0.63995
1.744 0.98803 5.5147e-005 3.8182 0.012027 2.2932e-005 0.0011545 0.18357 0.00065881 0.18422 0.16882 0 0.03495 0.0389 0 0.95032 0.27363 0.075601 0.010395 4.5487 0.064866 7.851e-005 0.82521 0.0055582 0.0063012 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.13421 0.92526 0.906 0.0013992 0.98742 0.5742 0.0018849 0.42824 1.8171 1.8162 16.0065 144.9875 0.00018106 -85.635 0.64095
1.745 0.98803 5.5147e-005 3.8182 0.012027 2.2945e-005 0.0011545 0.18361 0.00065881 0.18426 0.16886 0 0.034947 0.0389 0 0.95041 0.27367 0.075615 0.010397 4.5493 0.064876 7.8524e-005 0.8252 0.0055588 0.0063018 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.13422 0.92544 0.90609 0.0013991 0.98749 0.57435 0.0018849 0.42825 1.8176 1.8168 16.0064 144.9875 0.00018093 -85.6352 0.64195
1.746 0.98803 5.5147e-005 3.8182 0.012027 2.2958e-005 0.0011545 0.18365 0.00065881 0.18431 0.1689 0 0.034945 0.0389 0 0.9505 0.27371 0.07563 0.010399 4.55 0.064887 7.8538e-005 0.82519 0.0055593 0.0063024 0.0013901 0.98689 0.99167 2.9979e-006 1.1991e-005 0.13422 0.92562 0.90617 0.0013991 0.98755 0.5745 0.0018849 0.42826 1.8182 1.8173 16.0064 144.9875 0.00018079 -85.6355 0.64295
1.747 0.98804 5.5147e-005 3.8182 0.012027 2.2972e-005 0.0011545 0.18369 0.00065881 0.18435 0.16894 0 0.034942 0.0389 0 0.95059 0.27375 0.075644 0.010401 4.5506 0.064898 7.8552e-005 0.82518 0.0055599 0.0063029 0.00139 0.9869 0.99167 2.9978e-006 1.1991e-005 0.13423 0.9258 0.90626 0.0013991 0.98761 0.57465 0.0018848 0.42828 1.8187 1.8179 16.0064 144.9876 0.00018065 -85.6357 0.64395
1.748 0.98804 5.5147e-005 3.8182 0.012027 2.2985e-005 0.0011545 0.18373 0.00065881 0.18439 0.16897 0 0.03494 0.0389 0 0.95068 0.27379 0.075659 0.010402 4.5512 0.064909 7.8566e-005 0.82517 0.0055604 0.0063035 0.00139 0.9869 0.99167 2.9976e-006 1.199e-005 0.13423 0.92598 0.90635 0.001399 0.98768 0.57479 0.0018848 0.42829 1.8193 1.8184 16.0064 144.9876 0.00018051 -85.6359 0.64495
1.749 0.98804 5.5147e-005 3.8182 0.012026 2.2998e-005 0.0011545 0.18378 0.00065881 0.18443 0.16901 0 0.034938 0.0389 0 0.95077 0.27383 0.075673 0.010404 4.5518 0.064919 7.858e-005 0.82516 0.005561 0.0063041 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.13424 0.92616 0.90644 0.001399 0.98774 0.57494 0.0018847 0.4283 1.8198 1.819 16.0064 144.9876 0.00018037 -85.6362 0.64595
1.75 0.98804 5.5147e-005 3.8182 0.012026 2.3011e-005 0.0011545 0.18382 0.00065881 0.18447 0.16905 0 0.034935 0.0389 0 0.95086 0.27387 0.075688 0.010406 4.5524 0.06493 7.8594e-005 0.82515 0.0055616 0.0063046 0.0013899 0.9869 0.99167 2.9974e-006 1.1989e-005 0.13424 0.92634 0.90653 0.001399 0.9878 0.57509 0.0018847 0.42831 1.8203 1.8195 16.0063 144.9876 0.00018024 -85.6364 0.64695
1.751 0.98804 5.5147e-005 3.8182 0.012026 2.3024e-005 0.0011545 0.18386 0.00065881 0.18451 0.16909 0 0.034933 0.0389 0 0.95095 0.27391 0.075702 0.010407 4.5531 0.064941 7.8608e-005 0.82514 0.0055621 0.0063052 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.13425 0.92652 0.90661 0.001399 0.98786 0.57524 0.0018847 0.42833 1.8209 1.82 16.0063 144.9876 0.0001801 -85.6366 0.64795
1.752 0.98804 5.5146e-005 3.8182 0.012026 2.3037e-005 0.0011545 0.1839 0.00065881 0.18455 0.16913 0 0.03493 0.0389 0 0.95104 0.27395 0.075717 0.010409 4.5537 0.064952 7.8622e-005 0.82513 0.0055627 0.0063058 0.0013898 0.9869 0.99167 2.9971e-006 1.1988e-005 0.13425 0.9267 0.9067 0.0013989 0.98792 0.57539 0.0018846 0.42834 1.8214 1.8206 16.0063 144.9877 0.00017996 -85.6369 0.64895
1.753 0.98804 5.5146e-005 3.8182 0.012026 2.305e-005 0.0011545 0.18394 0.00065881 0.1846 0.16917 0 0.034928 0.0389 0 0.95113 0.27399 0.075731 0.010411 4.5543 0.064962 7.8636e-005 0.82512 0.0055632 0.0063064 0.0013897 0.9869 0.99167 2.997e-006 1.1988e-005 0.13426 0.92688 0.90679 0.0013989 0.98798 0.57553 0.0018846 0.42835 1.822 1.8211 16.0063 144.9877 0.00017983 -85.6371 0.64995
1.754 0.98804 5.5146e-005 3.8182 0.012026 2.3063e-005 0.0011545 0.18398 0.00065881 0.18464 0.16921 0 0.034926 0.0389 0 0.95122 0.27403 0.075746 0.010413 4.5549 0.064973 7.865e-005 0.82511 0.0055638 0.0063069 0.0013897 0.9869 0.99168 2.9969e-006 1.1987e-005 0.13426 0.92706 0.90687 0.0013989 0.98804 0.57568 0.0018846 0.42836 1.8225 1.8217 16.0062 144.9877 0.00017969 -85.6373 0.65095
1.755 0.98804 5.5146e-005 3.8182 0.012026 2.3076e-005 0.0011545 0.18402 0.00065881 0.18468 0.16925 0 0.034923 0.0389 0 0.95131 0.27407 0.07576 0.010414 4.5556 0.064984 7.8664e-005 0.82509 0.0055643 0.0063075 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.13427 0.92723 0.90696 0.0013988 0.9881 0.57583 0.0018845 0.42838 1.823 1.8222 16.0062 144.9877 0.00017956 -85.6376 0.65195
1.756 0.98804 5.5146e-005 3.8182 0.012026 2.309e-005 0.0011545 0.18407 0.00065881 0.18472 0.16929 0 0.034921 0.0389 0 0.9514 0.27411 0.075775 0.010416 4.5562 0.064995 7.8678e-005 0.82508 0.0055649 0.0063081 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.13427 0.92741 0.90704 0.0013988 0.98816 0.57598 0.0018845 0.42839 1.8236 1.8227 16.0062 144.9877 0.00017942 -85.6378 0.65295
1.757 0.98804 5.5146e-005 3.8182 0.012026 2.3103e-005 0.0011545 0.18411 0.00065881 0.18476 0.16932 0 0.034919 0.0389 0 0.95149 0.27415 0.075789 0.010418 4.5568 0.065005 7.8692e-005 0.82507 0.0055655 0.0063087 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.13427 0.92758 0.90713 0.0013988 0.98822 0.57612 0.0018844 0.4284 1.8241 1.8233 16.0062 144.9878 0.00017929 -85.638 0.65395
1.758 0.98804 5.5146e-005 3.8182 0.012026 2.3116e-005 0.0011545 0.18415 0.00065881 0.1848 0.16936 0 0.034916 0.0389 0 0.95158 0.27419 0.075804 0.01042 4.5574 0.065016 7.8706e-005 0.82506 0.005566 0.0063092 0.0013894 0.9869 0.99168 2.9964e-006 1.1986e-005 0.13428 0.92776 0.90721 0.0013988 0.98828 0.57627 0.0018844 0.42841 1.8246 1.8238 16.0061 144.9878 0.00017916 -85.6382 0.65495
1.759 0.98804 5.5146e-005 3.8182 0.012026 2.3129e-005 0.0011545 0.18419 0.00065881 0.18484 0.1694 0 0.034914 0.0389 0 0.95167 0.27423 0.075819 0.010421 4.5581 0.065027 7.872e-005 0.82505 0.0055666 0.0063098 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.13428 0.92793 0.9073 0.0013987 0.98833 0.57642 0.0018844 0.42843 1.8252 1.8243 16.0061 144.9878 0.00017902 -85.6385 0.65595
1.76 0.98804 5.5146e-005 3.8182 0.012026 2.3142e-005 0.0011545 0.18423 0.00065882 0.18488 0.16944 0 0.034911 0.0389 0 0.95176 0.27427 0.075833 0.010423 4.5587 0.065038 7.8734e-005 0.82504 0.0055671 0.0063104 0.0013893 0.9869 0.99168 2.9962e-006 1.1985e-005 0.13429 0.92811 0.90738 0.0013987 0.98839 0.57657 0.0018843 0.42844 1.8257 1.8249 16.0061 144.9878 0.00017889 -85.6387 0.65695
1.761 0.98804 5.5146e-005 3.8182 0.012026 2.3155e-005 0.0011545 0.18427 0.00065882 0.18493 0.16948 0 0.034909 0.0389 0 0.95185 0.27431 0.075848 0.010425 4.5593 0.065048 7.8748e-005 0.82503 0.0055677 0.006311 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.13429 0.92828 0.90747 0.0013987 0.98845 0.57671 0.0018843 0.42845 1.8262 1.8254 16.0061 144.9878 0.00017876 -85.6389 0.65795
1.762 0.98804 5.5146e-005 3.8182 0.012026 2.3168e-005 0.0011545 0.18431 0.00065882 0.18497 0.16952 0 0.034907 0.0389 0 0.95194 0.27435 0.075862 0.010426 4.5599 0.065059 7.8762e-005 0.82502 0.0055683 0.0063116 0.0013892 0.98691 0.99168 2.996e-006 1.1984e-005 0.1343 0.92845 0.90755 0.0013986 0.9885 0.57686 0.0018843 0.42847 1.8268 1.8259 16.006 144.9879 0.00017863 -85.6391 0.65895
1.763 0.98804 5.5146e-005 3.8182 0.012026 2.3181e-005 0.0011545 0.18435 0.00065882 0.18501 0.16956 0 0.034904 0.0389 0 0.95203 0.27439 0.075877 0.010428 4.5606 0.06507 7.8776e-005 0.82501 0.0055688 0.0063121 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.1343 0.92862 0.90763 0.0013986 0.98856 0.57701 0.0018842 0.42848 1.8273 1.8265 16.006 144.9879 0.0001785 -85.6393 0.65995
1.764 0.98804 5.5146e-005 3.8182 0.012026 2.3194e-005 0.0011545 0.18439 0.00065882 0.18505 0.1696 0 0.034902 0.0389 0 0.95212 0.27443 0.075891 0.01043 4.5612 0.065081 7.879e-005 0.825 0.0055694 0.0063127 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.13431 0.9288 0.90772 0.0013986 0.98862 0.57716 0.0018842 0.42849 1.8278 1.827 16.006 144.9879 0.00017837 -85.6395 0.66095
1.765 0.98804 5.5146e-005 3.8182 0.012026 2.3208e-005 0.0011545 0.18443 0.00065882 0.18509 0.16963 0 0.0349 0.0389 0 0.95221 0.27447 0.075906 0.010432 4.5618 0.065091 7.8804e-005 0.82499 0.0055699 0.0063133 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.13431 0.92897 0.9078 0.0013986 0.98867 0.5773 0.0018842 0.4285 1.8283 1.8275 16.006 144.9879 0.00017824 -85.6397 0.66195
1.766 0.98804 5.5146e-005 3.8182 0.012026 2.3221e-005 0.0011545 0.18448 0.00065882 0.18513 0.16967 0 0.034897 0.0389 0 0.9523 0.27451 0.075921 0.010433 4.5625 0.065102 7.8818e-005 0.82498 0.0055705 0.0063139 0.001389 0.98691 0.99168 2.9955e-006 1.1982e-005 0.13432 0.92914 0.90788 0.0013985 0.98873 0.57745 0.0018841 0.42852 1.8288 1.828 16.006 144.9879 0.00017811 -85.64 0.66295
1.767 0.98804 5.5146e-005 3.8182 0.012026 2.3234e-005 0.0011545 0.18452 0.00065882 0.18517 0.16971 0 0.034895 0.0389 0 0.95239 0.27455 0.075935 0.010435 4.5631 0.065113 7.8832e-005 0.82497 0.0055711 0.0063144 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.13432 0.92931 0.90796 0.0013985 0.98878 0.5776 0.0018841 0.42853 1.8294 1.8286 16.0059 144.988 0.00017798 -85.6402 0.66395
1.768 0.98804 5.5145e-005 3.8182 0.012026 2.3247e-005 0.0011545 0.18456 0.00065882 0.18521 0.16975 0 0.034892 0.0389 0 0.95248 0.2746 0.07595 0.010437 4.5637 0.065124 7.8846e-005 0.82496 0.0055716 0.006315 0.001389 0.98691 0.99168 2.9953e-006 1.1981e-005 0.13433 0.92948 0.90804 0.0013985 0.98884 0.57774 0.0018841 0.42854 1.8299 1.8291 16.0059 144.988 0.00017785 -85.6404 0.66495
1.769 0.98804 5.5145e-005 3.8182 0.012026 2.326e-005 0.0011545 0.1846 0.00065882 0.18525 0.16979 0 0.03489 0.0389 0 0.95257 0.27464 0.075964 0.010438 4.5643 0.065134 7.886e-005 0.82494 0.0055722 0.0063156 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.13433 0.92964 0.90813 0.0013985 0.98889 0.57789 0.001884 0.42855 1.8304 1.8296 16.0059 144.988 0.00017772 -85.6406 0.66595
1.77 0.98804 5.5145e-005 3.8182 0.012026 2.3273e-005 0.0011545 0.18464 0.00065882 0.18529 0.16983 0 0.034888 0.0389 0 0.95266 0.27468 0.075979 0.01044 4.565 0.065145 7.8875e-005 0.82493 0.0055728 0.0063162 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.13434 0.92981 0.90821 0.0013984 0.98895 0.57804 0.001884 0.42857 1.8309 1.8301 16.0059 144.988 0.00017759 -85.6408 0.66695
1.771 0.98804 5.5145e-005 3.8182 0.012026 2.3286e-005 0.0011545 0.18468 0.00065882 0.18533 0.16987 0 0.034885 0.0389 0 0.95275 0.27472 0.075993 0.010442 4.5656 0.065156 7.8889e-005 0.82492 0.0055733 0.0063168 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.13434 0.92998 0.90829 0.0013984 0.989 0.57818 0.001884 0.42858 1.8314 1.8306 16.0058 144.988 0.00017747 -85.641 0.66795
1.772 0.98804 5.5145e-005 3.8182 0.012026 2.3299e-005 0.0011545 0.18472 0.00065882 0.18537 0.1699 0 0.034883 0.0389 0 0.95284 0.27476 0.076008 0.010444 4.5662 0.065167 7.8903e-005 0.82491 0.0055739 0.0063173 0.0013888 0.98691 0.99168 2.9948e-006 1.1979e-005 0.13434 0.93015 0.90837 0.0013984 0.98905 0.57833 0.0018839 0.42859 1.832 1.8312 16.0058 144.9881 0.00017734 -85.6412 0.66895
1.773 0.98804 5.5145e-005 3.8182 0.012026 2.3312e-005 0.0011545 0.18476 0.00065882 0.18542 0.16994 0 0.034881 0.0389 0 0.95293 0.2748 0.076023 0.010445 4.5669 0.065177 7.8917e-005 0.8249 0.0055744 0.0063179 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.13435 0.93032 0.90845 0.0013984 0.9891 0.57848 0.0018839 0.4286 1.8325 1.8317 16.0058 144.9881 0.00017721 -85.6414 0.66995
1.774 0.98804 5.5145e-005 3.8182 0.012026 2.3326e-005 0.0011545 0.1848 0.00065882 0.18546 0.16998 0 0.034878 0.0389 0 0.95302 0.27484 0.076037 0.010447 4.5675 0.065188 7.8931e-005 0.82489 0.005575 0.0063185 0.0013887 0.98691 0.99168 2.9946e-006 1.1978e-005 0.13435 0.93048 0.90853 0.0013983 0.98916 0.57862 0.0018839 0.42862 1.833 1.8322 16.0058 144.9881 0.00017709 -85.6416 0.67095
1.775 0.98804 5.5145e-005 3.8182 0.012026 2.3339e-005 0.0011545 0.18484 0.00065882 0.1855 0.17002 0 0.034876 0.0389 0 0.95311 0.27488 0.076052 0.010449 4.5681 0.065199 7.8945e-005 0.82488 0.0055756 0.0063191 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.13436 0.93065 0.90861 0.0013983 0.98921 0.57877 0.0018838 0.42863 1.8335 1.8327 16.0057 144.9881 0.00017696 -85.6418 0.67195
1.776 0.98804 5.5145e-005 3.8182 0.012026 2.3352e-005 0.0011545 0.18488 0.00065882 0.18554 0.17006 0 0.034874 0.0389 0 0.9532 0.27492 0.076066 0.010451 4.5688 0.06521 7.8959e-005 0.82487 0.0055761 0.0063197 0.0013886 0.98691 0.99168 2.9944e-006 1.1978e-005 0.13436 0.93081 0.90869 0.0013983 0.98926 0.57892 0.0018838 0.42864 1.834 1.8332 16.0057 144.9881 0.00017684 -85.642 0.67295
1.777 0.98804 5.5145e-005 3.8182 0.012026 2.3365e-005 0.0011545 0.18492 0.00065882 0.18558 0.1701 0 0.034871 0.0389 0 0.95329 0.27496 0.076081 0.010452 4.5694 0.065221 7.8973e-005 0.82486 0.0055767 0.0063203 0.0013885 0.98691 0.99168 2.9943e-006 1.1977e-005 0.13437 0.93098 0.90877 0.0013983 0.98931 0.57906 0.0018838 0.42865 1.8345 1.8337 16.0057 144.9882 0.00017671 -85.6422 0.67395
1.778 0.98804 5.5145e-005 3.8182 0.012026 2.3378e-005 0.0011545 0.18496 0.00065882 0.18562 0.17013 0 0.034869 0.0389 0 0.95338 0.275 0.076096 0.010454 4.57 0.065231 7.8987e-005 0.82485 0.0055773 0.0063208 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.13437 0.93114 0.90885 0.0013982 0.98936 0.57921 0.0018837 0.42867 1.835 1.8342 16.0057 144.9882 0.00017659 -85.6424 0.67495
1.779 0.98804 5.5145e-005 3.8182 0.012026 2.3391e-005 0.0011545 0.185 0.00065882 0.18566 0.17017 0 0.034867 0.0389 0 0.95347 0.27504 0.07611 0.010456 4.5707 0.065242 7.9001e-005 0.82484 0.0055778 0.0063214 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.13438 0.93131 0.90893 0.0013982 0.98941 0.57936 0.0018837 0.42868 1.8355 1.8348 16.0056 144.9882 0.00017646 -85.6426 0.67595
1.78 0.98804 5.5145e-005 3.8182 0.012026 2.3404e-005 0.0011545 0.18505 0.00065883 0.1857 0.17021 0 0.034864 0.0389 0 0.95356 0.27508 0.076125 0.010458 4.5713 0.065253 7.9015e-005 0.82483 0.0055784 0.006322 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.13438 0.93147 0.90901 0.0013982 0.98946 0.5795 0.0018837 0.42869 1.836 1.8353 16.0056 144.9882 0.00017634 -85.6428 0.67695
1.781 0.98804 5.5145e-005 3.8182 0.012026 2.3417e-005 0.0011545 0.18509 0.00065883 0.18574 0.17025 0 0.034862 0.0389 0 0.95365 0.27512 0.076139 0.010459 4.5719 0.065264 7.9029e-005 0.82482 0.005579 0.0063226 0.0013884 0.98692 0.99169 2.9939e-006 1.1976e-005 0.13439 0.93163 0.90908 0.0013982 0.98951 0.57965 0.0018837 0.4287 1.8366 1.8358 16.0056 144.9882 0.00017622 -85.643 0.67795
1.782 0.98804 5.5145e-005 3.8182 0.012026 2.343e-005 0.0011545 0.18513 0.00065883 0.18578 0.17029 0 0.03486 0.0389 0 0.95374 0.27516 0.076154 0.010461 4.5726 0.065274 7.9043e-005 0.8248 0.0055795 0.0063232 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.13439 0.93179 0.90916 0.0013982 0.98956 0.5798 0.0018836 0.42872 1.8371 1.8363 16.0056 144.9883 0.00017609 -85.6431 0.67895
1.783 0.98804 5.5144e-005 3.8182 0.012026 2.3444e-005 0.0011545 0.18517 0.00065883 0.18582 0.17032 0 0.034857 0.0389 0 0.95383 0.2752 0.076169 0.010463 4.5732 0.065285 7.9057e-005 0.82479 0.0055801 0.0063237 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.1344 0.93195 0.90924 0.0013981 0.98961 0.57994 0.0018836 0.42873 1.8376 1.8368 16.0055 144.9883 0.00017597 -85.6433 0.67995
1.784 0.98804 5.5144e-005 3.8182 0.012026 2.3457e-005 0.0011545 0.18521 0.00065883 0.18586 0.17036 0 0.034855 0.0389 0 0.95393 0.27524 0.076183 0.010464 4.5739 0.065296 7.9072e-005 0.82478 0.0055807 0.0063243 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.1344 0.93212 0.90932 0.0013981 0.98966 0.58009 0.0018836 0.42874 1.8381 1.8373 16.0055 144.9883 0.00017585 -85.6435 0.68095
1.785 0.98804 5.5144e-005 3.8182 0.012026 2.347e-005 0.0011545 0.18525 0.00065883 0.1859 0.1704 0 0.034853 0.0389 0 0.95402 0.27529 0.076198 0.010466 4.5745 0.065307 7.9086e-005 0.82477 0.0055812 0.0063249 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.13441 0.93228 0.90939 0.0013981 0.98971 0.58023 0.0018835 0.42875 1.8386 1.8378 16.0055 144.9883 0.00017573 -85.6437 0.68195
1.786 0.98804 5.5144e-005 3.8182 0.012026 2.3483e-005 0.0011545 0.18529 0.00065883 0.18594 0.17044 0 0.03485 0.0389 0 0.95411 0.27533 0.076212 0.010468 4.5751 0.065318 7.91e-005 0.82476 0.0055818 0.0063255 0.0013881 0.98692 0.99169 2.9934e-006 1.1974e-005 0.13441 0.93244 0.90947 0.0013981 0.98976 0.58038 0.0018835 0.42877 1.8391 1.8383 16.0055 144.9883 0.00017561 -85.6439 0.68295
1.787 0.98804 5.5144e-005 3.8182 0.012026 2.3496e-005 0.0011545 0.18533 0.00065883 0.18598 0.17048 0 0.034848 0.0389 0 0.9542 0.27537 0.076227 0.01047 4.5758 0.065328 7.9114e-005 0.82475 0.0055824 0.0063261 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.13441 0.9326 0.90955 0.001398 0.98981 0.58053 0.0018835 0.42878 1.8396 1.8388 16.0054 144.9884 0.00017549 -85.6441 0.68395
1.788 0.98804 5.5144e-005 3.8182 0.012026 2.3509e-005 0.0011545 0.18537 0.00065883 0.18602 0.17051 0 0.034846 0.0389 0 0.95429 0.27541 0.076242 0.010471 4.5764 0.065339 7.9128e-005 0.82474 0.0055829 0.0063267 0.0013881 0.98692 0.99169 2.9932e-006 1.1973e-005 0.13442 0.93276 0.90962 0.001398 0.98986 0.58067 0.0018834 0.42879 1.8401 1.8393 16.0054 144.9884 0.00017537 -85.6443 0.68495
1.789 0.98804 5.5144e-005 3.8182 0.012026 2.3522e-005 0.0011545 0.18541 0.00065883 0.18606 0.17055 0 0.034843 0.0389 0 0.95438 0.27545 0.076256 0.010473 4.5771 0.06535 7.9142e-005 0.82473 0.0055835 0.0063272 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.13442 0.93291 0.9097 0.001398 0.9899 0.58082 0.0018834 0.4288 1.8406 1.8398 16.0054 144.9884 0.00017525 -85.6444 0.68595
1.79 0.98804 5.5144e-005 3.8182 0.012026 2.3535e-005 0.0011545 0.18545 0.00065883 0.1861 0.17059 0 0.034841 0.0389 0 0.95447 0.27549 0.076271 0.010475 4.5777 0.065361 7.9156e-005 0.82472 0.0055841 0.0063278 0.001388 0.98692 0.99169 2.993e-006 1.1972e-005 0.13443 0.93307 0.90978 0.001398 0.98995 0.58096 0.0018834 0.42882 1.8411 1.8403 16.0054 144.9884 0.00017513 -85.6446 0.68695
1.791 0.98804 5.5144e-005 3.8182 0.012026 2.3548e-005 0.0011545 0.18549 0.00065883 0.18614 0.17063 0 0.034839 0.0389 0 0.95456 0.27553 0.076286 0.010477 4.5783 0.065371 7.917e-005 0.82471 0.0055846 0.0063284 0.0013879 0.98692 0.99169 2.9929e-006 1.1972e-005 0.13443 0.93323 0.90985 0.001398 0.99 0.58111 0.0018834 0.42883 1.8416 1.8408 16.0053 144.9885 0.00017501 -85.6448 0.68795
1.792 0.98804 5.5144e-005 3.8182 0.012026 2.3562e-005 0.0011545 0.18553 0.00065883 0.18618 0.17066 0 0.034837 0.0389 0 0.95465 0.27557 0.0763 0.010478 4.579 0.065382 7.9184e-005 0.8247 0.0055852 0.006329 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.13444 0.93339 0.90993 0.0013979 0.99005 0.58126 0.0018833 0.42884 1.8421 1.8413 16.0053 144.9885 0.00017489 -85.645 0.68895
1.793 0.98804 5.5144e-005 3.8182 0.012026 2.3575e-005 0.0011545 0.18557 0.00065883 0.18622 0.1707 0 0.034834 0.0389 0 0.95474 0.27561 0.076315 0.01048 4.5796 0.065393 7.9198e-005 0.82469 0.0055858 0.0063296 0.0013878 0.98692 0.99169 2.9928e-006 1.1971e-005 0.13444 0.93354 0.91 0.0013979 0.99009 0.5814 0.0018833 0.42885 1.8425 1.8418 16.0053 144.9885 0.00017478 -85.6451 0.68995
1.794 0.98804 5.5144e-005 3.8182 0.012026 2.3588e-005 0.0011545 0.18561 0.00065883 0.18626 0.17074 0 0.034832 0.0389 0 0.95483 0.27565 0.076329 0.010482 4.5803 0.065404 7.9213e-005 0.82468 0.0055863 0.0063302 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.13445 0.9337 0.91008 0.0013979 0.99014 0.58155 0.0018833 0.42887 1.843 1.8423 16.0053 144.9885 0.00017466 -85.6453 0.69095
1.795 0.98804 5.5144e-005 3.8182 0.012026 2.3601e-005 0.0011545 0.18565 0.00065883 0.1863 0.17078 0 0.03483 0.0389 0 0.95492 0.27569 0.076344 0.010483 4.5809 0.065415 7.9227e-005 0.82466 0.0055869 0.0063308 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.13445 0.93386 0.91015 0.0013979 0.99018 0.58169 0.0018832 0.42888 1.8435 1.8428 16.0052 144.9885 0.00017454 -85.6455 0.69195
1.796 0.98804 5.5144e-005 3.8182 0.012026 2.3614e-005 0.0011545 0.18569 0.00065883 0.18634 0.17082 0 0.034827 0.0389 0 0.95501 0.27573 0.076359 0.010485 4.5815 0.065425 7.9241e-005 0.82465 0.0055875 0.0063313 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.13446 0.93401 0.91023 0.0013978 0.99023 0.58184 0.0018832 0.42889 1.844 1.8433 16.0052 144.9886 0.00017442 -85.6457 0.69295
1.797 0.98804 5.5144e-005 3.8182 0.012026 2.3627e-005 0.0011545 0.18573 0.00065883 0.18638 0.17085 0 0.034825 0.0389 0 0.9551 0.27577 0.076373 0.010487 4.5822 0.065436 7.9255e-005 0.82464 0.005588 0.0063319 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.13446 0.93417 0.9103 0.0013978 0.99027 0.58198 0.0018832 0.4289 1.8445 1.8437 16.0052 144.9886 0.00017431 -85.6458 0.69395
1.798 0.98804 5.5144e-005 3.8182 0.012026 2.364e-005 0.0011545 0.18577 0.00065883 0.18642 0.17089 0 0.034823 0.0389 0 0.95519 0.27581 0.076388 0.010489 4.5828 0.065447 7.9269e-005 0.82463 0.0055886 0.0063325 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.13447 0.93432 0.91037 0.0013978 0.99032 0.58213 0.0018832 0.42892 1.845 1.8442 16.0051 144.9886 0.00017419 -85.646 0.69495
1.799 0.98804 5.5143e-005 3.8182 0.012026 2.3653e-005 0.0011545 0.18581 0.00065884 0.18646 0.17093 0 0.03482 0.0389 0 0.95528 0.27585 0.076403 0.01049 4.5835 0.065458 7.9283e-005 0.82462 0.0055892 0.0063331 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.13447 0.93447 0.91045 0.0013978 0.99036 0.58227 0.0018831 0.42893 1.8455 1.8447 16.0051 144.9886 0.00017408 -85.6462 0.69595
1.8 0.98804 5.5143e-005 3.8182 0.012026 2.3666e-005 0.0011545 0.18585 0.00065884 0.1865 0.17097 0 0.034818 0.0389 0 0.95537 0.2759 0.076417 0.010492 4.5841 0.065469 7.9297e-005 0.82461 0.0055898 0.0063337 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.13448 0.93463 0.91052 0.0013978 0.99041 0.58242 0.0018831 0.42894 1.846 1.8452 16.0051 144.9886 0.00017396 -85.6463 0.69695
1.801 0.98804 5.5143e-005 3.8182 0.012026 2.368e-005 0.0011545 0.18589 0.00065884 0.18654 0.171 0 0.034816 0.0389 0 0.95547 0.27594 0.076432 0.010494 4.5848 0.065479 7.9311e-005 0.8246 0.0055903 0.0063343 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.13448 0.93478 0.91059 0.0013977 0.99045 0.58256 0.0018831 0.42895 1.8465 1.8457 16.0051 144.9887 0.00017385 -85.6465 0.69795
1.802 0.98804 5.5143e-005 3.8182 0.012026 2.3693e-005 0.0011545 0.18593 0.00065884 0.18658 0.17104 0 0.034814 0.0389 0 0.95556 0.27598 0.076447 0.010496 4.5854 0.06549 7.9326e-005 0.82459 0.0055909 0.0063349 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.13448 0.93493 0.91067 0.0013977 0.9905 0.58271 0.0018831 0.42897 1.8469 1.8462 16.005 144.9887 0.00017373 -85.6467 0.69895
1.803 0.98804 5.5143e-005 3.8182 0.012026 2.3706e-005 0.0011545 0.18597 0.00065884 0.18662 0.17108 0 0.034811 0.0389 0 0.95565 0.27602 0.076461 0.010497 4.5861 0.065501 7.934e-005 0.82458 0.0055915 0.0063355 0.0013875 0.98693 0.99169 2.9919e-006 1.1967e-005 0.13449 0.93508 0.91074 0.0013977 0.99054 0.58286 0.001883 0.42898 1.8474 1.8467 16.005 144.9887 0.00017362 -85.6468 0.69995
1.804 0.98804 5.5143e-005 3.8182 0.012026 2.3719e-005 0.0011545 0.18601 0.00065884 0.18666 0.17112 0 0.034809 0.0389 0 0.95574 0.27606 0.076476 0.010499 4.5867 0.065512 7.9354e-005 0.82457 0.005592 0.0063361 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.13449 0.93524 0.91081 0.0013977 0.99058 0.583 0.001883 0.42899 1.8479 1.8472 16.005 144.9887 0.00017351 -85.647 0.70095
1.805 0.98804 5.5143e-005 3.8182 0.012026 2.3732e-005 0.0011545 0.18605 0.00065884 0.1867 0.17115 0 0.034807 0.0389 0 0.95583 0.2761 0.076491 0.010501 4.5873 0.065523 7.9368e-005 0.82456 0.0055926 0.0063366 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.1345 0.93539 0.91088 0.0013977 0.99063 0.58315 0.001883 0.429 1.8484 1.8476 16.005 144.9887 0.00017339 -85.6472 0.70195
1.806 0.98804 5.5143e-005 3.8182 0.012026 2.3745e-005 0.0011545 0.18609 0.00065884 0.18674 0.17119 0 0.034805 0.0389 0 0.95592 0.27614 0.076505 0.010503 4.588 0.065534 7.9382e-005 0.82455 0.0055932 0.0063372 0.0013873 0.98693 0.99169 2.9916e-006 1.1966e-005 0.1345 0.93554 0.91095 0.0013976 0.99067 0.58329 0.001883 0.42902 1.8489 1.8481 16.0049 144.9888 0.00017328 -85.6473 0.70295
1.807 0.98804 5.5143e-005 3.8182 0.012026 2.3758e-005 0.0011546 0.18613 0.00065884 0.18678 0.17123 0 0.034802 0.0389 0 0.95601 0.27618 0.07652 0.010504 4.5886 0.065544 7.9396e-005 0.82454 0.0055938 0.0063378 0.0013873 0.98693 0.99169 2.9915e-006 1.1966e-005 0.13451 0.93569 0.91103 0.0013976 0.99071 0.58344 0.0018829 0.42903 1.8493 1.8486 16.0049 144.9888 0.00017317 -85.6475 0.70395
1.808 0.98804 5.5143e-005 3.8182 0.012026 2.3771e-005 0.0011546 0.18616 0.00065884 0.18682 0.17126 0 0.0348 0.0389 0 0.9561 0.27622 0.076535 0.010506 4.5893 0.065555 7.941e-005 0.82452 0.0055943 0.0063384 0.0013873 0.98693 0.9917 2.9914e-006 1.1966e-005 0.13451 0.93584 0.9111 0.0013976 0.99075 0.58358 0.0018829 0.42904 1.8498 1.8491 16.0049 144.9888 0.00017306 -85.6476 0.70495
1.809 0.98804 5.5143e-005 3.8182 0.012026 2.3784e-005 0.0011546 0.1862 0.00065884 0.18686 0.1713 0 0.034798 0.0389 0 0.95619 0.27626 0.076549 0.010508 4.5899 0.065566 7.9424e-005 0.82451 0.0055949 0.006339 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.13452 0.93599 0.91117 0.0013976 0.99079 0.58373 0.0018829 0.42905 1.8503 1.8496 16.0049 144.9888 0.00017294 -85.6478 0.70595
1.81 0.98804 5.5143e-005 3.8182 0.012026 2.3797e-005 0.0011546 0.18624 0.00065884 0.1869 0.17134 0 0.034795 0.0389 0 0.95628 0.2763 0.076564 0.010509 4.5906 0.065577 7.9439e-005 0.8245 0.0055955 0.0063396 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.13452 0.93613 0.91124 0.0013976 0.99084 0.58387 0.0018829 0.42907 1.8508 1.85 16.0048 144.9888 0.00017283 -85.648 0.70695
1.811 0.98804 5.5143e-005 3.8182 0.012026 2.3811e-005 0.0011546 0.18628 0.00065884 0.18694 0.17138 0 0.034793 0.0389 0 0.95637 0.27634 0.076579 0.010511 4.5912 0.065588 7.9453e-005 0.82449 0.005596 0.0063402 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.13453 0.93628 0.91131 0.0013975 0.99088 0.58402 0.0018828 0.42908 1.8512 1.8505 16.0048 144.9889 0.00017272 -85.6481 0.70795
1.812 0.98804 5.5143e-005 3.8182 0.012026 2.3824e-005 0.0011546 0.18632 0.00065884 0.18698 0.17141 0 0.034791 0.0389 0 0.95646 0.27638 0.076593 0.010513 4.5919 0.065598 7.9467e-005 0.82448 0.0055966 0.0063408 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.13453 0.93643 0.91138 0.0013975 0.99092 0.58416 0.0018828 0.42909 1.8517 1.851 16.0048 144.9889 0.00017261 -85.6483 0.70895
1.813 0.98804 5.5143e-005 3.8182 0.012026 2.3837e-005 0.0011546 0.18636 0.00065884 0.18702 0.17145 0 0.034789 0.0389 0 0.95656 0.27643 0.076608 0.010515 4.5925 0.065609 7.9481e-005 0.82447 0.0055972 0.0063414 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.13454 0.93658 0.91145 0.0013975 0.99096 0.5843 0.0018828 0.4291 1.8522 1.8515 16.0048 144.9889 0.0001725 -85.6484 0.70995
1.814 0.98804 5.5142e-005 3.8182 0.012026 2.385e-005 0.0011546 0.1864 0.00065884 0.18706 0.17149 0 0.034786 0.0389 0 0.95665 0.27647 0.076623 0.010516 4.5932 0.06562 7.9495e-005 0.82446 0.0055978 0.006342 0.0013871 0.98693 0.9917 2.9909e-006 1.1964e-005 0.13454 0.93672 0.91152 0.0013975 0.991 0.58445 0.0018828 0.42912 1.8527 1.8519 16.0047 144.9889 0.00017239 -85.6486 0.71095
1.815 0.98804 5.5142e-005 3.8182 0.012026 2.3863e-005 0.0011546 0.18644 0.00065884 0.1871 0.17152 0 0.034784 0.0389 0 0.95674 0.27651 0.076637 0.010518 4.5938 0.065631 7.9509e-005 0.82445 0.0055983 0.0063425 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.13455 0.93687 0.91159 0.0013975 0.99104 0.58459 0.0018827 0.42913 1.8531 1.8524 16.0047 144.9889 0.00017228 -85.6487 0.71195
1.816 0.98804 5.5142e-005 3.8182 0.012026 2.3876e-005 0.0011546 0.18648 0.00065884 0.18713 0.17156 0 0.034782 0.0389 0 0.95683 0.27655 0.076652 0.01052 4.5945 0.065642 7.9524e-005 0.82444 0.0055989 0.0063431 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.13455 0.93702 0.91166 0.0013975 0.99108 0.58474 0.0018827 0.42914 1.8536 1.8529 16.0047 144.989 0.00017217 -85.6489 0.71295
1.817 0.98804 5.5142e-005 3.8182 0.012026 2.3889e-005 0.0011546 0.18652 0.00065884 0.18717 0.1716 0 0.03478 0.0389 0 0.95692 0.27659 0.076667 0.010522 4.5951 0.065653 7.9538e-005 0.82443 0.0055995 0.0063437 0.0013869 0.98693 0.9917 2.9907e-006 1.1963e-005 0.13456 0.93716 0.91173 0.0013974 0.99112 0.58488 0.0018827 0.42915 1.8541 1.8533 16.0047 144.989 0.00017207 -85.649 0.71395
1.818 0.98804 5.5142e-005 3.8182 0.012026 2.3902e-005 0.0011546 0.18656 0.00065884 0.18721 0.17164 0 0.034777 0.0389 0 0.95701 0.27663 0.076681 0.010523 4.5958 0.065663 7.9552e-005 0.82442 0.0056001 0.0063443 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.13456 0.93731 0.9118 0.0013974 0.99116 0.58503 0.0018827 0.42917 1.8545 1.8538 16.0046 144.989 0.00017196 -85.6492 0.71495
1.819 0.98804 5.5142e-005 3.8182 0.012026 2.3915e-005 0.0011546 0.1866 0.00065884 0.18725 0.17167 0 0.034775 0.0389 0 0.9571 0.27667 0.076696 0.010525 4.5965 0.065674 7.9566e-005 0.82441 0.0056006 0.0063449 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.13457 0.93745 0.91186 0.0013974 0.9912 0.58517 0.0018826 0.42918 1.855 1.8543 16.0046 144.989 0.00017185 -85.6493 0.71595
1.82 0.98804 5.5142e-005 3.8182 0.012026 2.3929e-005 0.0011546 0.18664 0.00065885 0.18729 0.17171 0 0.034773 0.0389 0 0.95719 0.27671 0.076711 0.010527 4.5971 0.065685 7.958e-005 0.82439 0.0056012 0.0063455 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.13457 0.93759 0.91193 0.0013974 0.99124 0.58532 0.0018826 0.42919 1.8555 1.8548 16.0046 144.989 0.00017174 -85.6495 0.71695
1.821 0.98804 5.5142e-005 3.8182 0.012025 2.3942e-005 0.0011546 0.18668 0.00065885 0.18733 0.17175 0 0.034771 0.0389 0 0.95728 0.27675 0.076725 0.010529 4.5978 0.065696 7.9594e-005 0.82438 0.0056018 0.0063461 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.13457 0.93774 0.912 0.0013974 0.99127 0.58546 0.0018826 0.4292 1.8559 1.8552 16.0045 144.9891 0.00017164 -85.6496 0.71795
1.822 0.98804 5.5142e-005 3.8182 0.012025 2.3955e-005 0.0011546 0.18672 0.00065885 0.18737 0.17178 0 0.034768 0.0389 0 0.95737 0.27679 0.07674 0.01053 4.5984 0.065707 7.9608e-005 0.82437 0.0056024 0.0063467 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.13458 0.93788 0.91207 0.0013973 0.99131 0.5856 0.0018826 0.42922 1.8564 1.8557 16.0045 144.9891 0.00017153 -85.6497 0.71895
1.823 0.98804 5.5142e-005 3.8182 0.012025 2.3968e-005 0.0011546 0.18675 0.00065885 0.18741 0.17182 0 0.034766 0.0389 0 0.95746 0.27683 0.076755 0.010532 4.5991 0.065718 7.9623e-005 0.82436 0.0056029 0.0063473 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.13458 0.93802 0.91214 0.0013973 0.99135 0.58575 0.0018825 0.42923 1.8569 1.8561 16.0045 144.9891 0.00017142 -85.6499 0.71995
1.824 0.98804 5.5142e-005 3.8182 0.012025 2.3981e-005 0.0011546 0.18679 0.00065885 0.18745 0.17186 0 0.034764 0.0389 0 0.95756 0.27687 0.07677 0.010534 4.5997 0.065728 7.9637e-005 0.82435 0.0056035 0.0063479 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.13459 0.93817 0.9122 0.0013973 0.99139 0.58589 0.0018825 0.42924 1.8573 1.8566 16.0045 144.9891 0.00017132 -85.65 0.72095
1.825 0.98804 5.5142e-005 3.8182 0.012025 2.3994e-005 0.0011546 0.18683 0.00065885 0.18749 0.17189 0 0.034762 0.0389 0 0.95765 0.27692 0.076784 0.010535 4.6004 0.065739 7.9651e-005 0.82434 0.0056041 0.0063485 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.13459 0.93831 0.91227 0.0013973 0.99143 0.58604 0.0018825 0.42925 1.8578 1.8571 16.0044 144.9891 0.00017121 -85.6502 0.72195
1.826 0.98804 5.5142e-005 3.8182 0.012025 2.4007e-005 0.0011546 0.18687 0.00065885 0.18753 0.17193 0 0.034759 0.0389 0 0.95774 0.27696 0.076799 0.010537 4.601 0.06575 7.9665e-005 0.82433 0.0056047 0.0063491 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.1346 0.93845 0.91234 0.0013973 0.99146 0.58618 0.0018825 0.42926 1.8582 1.8575 16.0044 144.9892 0.00017111 -85.6503 0.72295
1.827 0.98804 5.5142e-005 3.8182 0.012025 2.402e-005 0.0011546 0.18691 0.00065885 0.18756 0.17197 0 0.034757 0.0389 0 0.95783 0.277 0.076814 0.010539 4.6017 0.065761 7.9679e-005 0.82432 0.0056052 0.0063497 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.1346 0.93859 0.9124 0.0013973 0.9915 0.58633 0.0018825 0.42928 1.8587 1.858 16.0044 144.9892 0.000171 -85.6505 0.72395
1.828 0.98804 5.5142e-005 3.8182 0.012025 2.4033e-005 0.0011546 0.18695 0.00065885 0.1876 0.172 0 0.034755 0.0389 0 0.95792 0.27704 0.076828 0.010541 4.6024 0.065772 7.9694e-005 0.82431 0.0056058 0.0063503 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.13461 0.93873 0.91247 0.0013972 0.99154 0.58647 0.0018824 0.42929 1.8592 1.8585 16.0044 144.9892 0.0001709 -85.6506 0.72495
1.829 0.98804 5.5142e-005 3.8182 0.012025 2.4047e-005 0.0011546 0.18699 0.00065885 0.18764 0.17204 0 0.034753 0.0389 0 0.95801 0.27708 0.076843 0.010542 4.603 0.065783 7.9708e-005 0.8243 0.0056064 0.0063509 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.13461 0.93887 0.91254 0.0013972 0.99157 0.58661 0.0018824 0.4293 1.8596 1.8589 16.0043 144.9892 0.00017079 -85.6507 0.72595
1.83 0.98804 5.5141e-005 3.8182 0.012025 2.406e-005 0.0011546 0.18703 0.00065885 0.18768 0.17208 0 0.034751 0.0389 0 0.9581 0.27712 0.076858 0.010544 4.6037 0.065793 7.9722e-005 0.82429 0.005607 0.0063515 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.13462 0.93901 0.9126 0.0013972 0.99161 0.58676 0.0018824 0.42931 1.8601 1.8594 16.0043 144.9892 0.00017069 -85.6509 0.72695
1.831 0.98804 5.5141e-005 3.8182 0.012025 2.4073e-005 0.0011546 0.18707 0.00065885 0.18772 0.17211 0 0.034748 0.0389 0 0.95819 0.27716 0.076873 0.010546 4.6043 0.065804 7.9736e-005 0.82428 0.0056075 0.006352 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.13462 0.93915 0.91267 0.0013972 0.99165 0.5869 0.0018824 0.42933 1.8605 1.8598 16.0043 144.9893 0.00017059 -85.651 0.72795
1.832 0.98804 5.5141e-005 3.8182 0.012025 2.4086e-005 0.0011546 0.1871 0.00065885 0.18776 0.17215 0 0.034746 0.0389 0 0.95828 0.2772 0.076887 0.010548 4.605 0.065815 7.975e-005 0.82426 0.0056081 0.0063526 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.13463 0.93929 0.91273 0.0013972 0.99168 0.58704 0.0018823 0.42934 1.861 1.8603 16.0042 144.9893 0.00017048 -85.6511 0.72895
1.833 0.98804 5.5141e-005 3.8182 0.012025 2.4099e-005 0.0011546 0.18714 0.00065885 0.1878 0.17219 0 0.034744 0.0389 0 0.95838 0.27724 0.076902 0.010549 4.6056 0.065826 7.9764e-005 0.82425 0.0056087 0.0063532 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.13463 0.93943 0.9128 0.0013972 0.99172 0.58719 0.0018823 0.42935 1.8614 1.8607 16.0042 144.9893 0.00017038 -85.6513 0.72995
1.834 0.98804 5.5141e-005 3.8182 0.012025 2.4112e-005 0.0011546 0.18718 0.00065885 0.18784 0.17222 0 0.034742 0.0389 0 0.95847 0.27728 0.076917 0.010551 4.6063 0.065837 7.9779e-005 0.82424 0.0056093 0.0063538 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.13464 0.93956 0.91286 0.0013971 0.99175 0.58733 0.0018823 0.42936 1.8619 1.8612 16.0042 144.9893 0.00017028 -85.6514 0.73095
1.835 0.98804 5.5141e-005 3.8182 0.012025 2.4125e-005 0.0011546 0.18722 0.00065885 0.18788 0.17226 0 0.034739 0.0389 0 0.95856 0.27732 0.076932 0.010553 4.607 0.065848 7.9793e-005 0.82423 0.0056099 0.0063544 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.13464 0.9397 0.91293 0.0013971 0.99179 0.58748 0.0018823 0.42938 1.8623 1.8617 16.0042 144.9893 0.00017018 -85.6515 0.73195
1.836 0.98804 5.5141e-005 3.8182 0.012025 2.4138e-005 0.0011546 0.18726 0.00065885 0.18791 0.1723 0 0.034737 0.0389 0 0.95865 0.27737 0.076946 0.010555 4.6076 0.065858 7.9807e-005 0.82422 0.0056104 0.006355 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.13465 0.93984 0.91299 0.0013971 0.99183 0.58762 0.0018823 0.42939 1.8628 1.8621 16.0041 144.9894 0.00017007 -85.6517 0.73295
1.837 0.98804 5.5141e-005 3.8182 0.012025 2.4151e-005 0.0011546 0.1873 0.00065885 0.18795 0.17233 0 0.034735 0.0389 0 0.95874 0.27741 0.076961 0.010556 4.6083 0.065869 7.9821e-005 0.82421 0.005611 0.0063556 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.13465 0.93998 0.91306 0.0013971 0.99186 0.58776 0.0018822 0.4294 1.8632 1.8626 16.0041 144.9894 0.00016997 -85.6518 0.73395
1.838 0.98804 5.5141e-005 3.8182 0.012025 2.4164e-005 0.0011546 0.18734 0.00065885 0.18799 0.17237 0 0.034733 0.0389 0 0.95883 0.27745 0.076976 0.010558 4.609 0.06588 7.9835e-005 0.8242 0.0056116 0.0063562 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.13466 0.94011 0.91312 0.0013971 0.99189 0.58791 0.0018822 0.42941 1.8637 1.863 16.0041 144.9894 0.00016987 -85.6519 0.73495
1.839 0.98804 5.5141e-005 3.8182 0.012025 2.4178e-005 0.0011546 0.18738 0.00065885 0.18803 0.17241 0 0.034731 0.0389 0 0.95892 0.27749 0.07699 0.01056 4.6096 0.065891 7.985e-005 0.82419 0.0056122 0.0063568 0.0013862 0.98694 0.9917 2.9891e-006 1.1956e-005 0.13466 0.94025 0.91319 0.0013971 0.99193 0.58805 0.0018822 0.42943 1.8641 1.8635 16.0041 144.9894 0.00016977 -85.6521 0.73595
1.84 0.98804 5.5141e-005 3.8182 0.012025 2.4191e-005 0.0011546 0.18741 0.00065885 0.18807 0.17244 0 0.034728 0.0389 0 0.95901 0.27753 0.077005 0.010562 4.6103 0.065902 7.9864e-005 0.82418 0.0056128 0.0063574 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.13467 0.94038 0.91325 0.0013971 0.99196 0.58819 0.0018822 0.42944 1.8646 1.8639 16.004 144.9895 0.00016967 -85.6522 0.73695
1.841 0.98804 5.5141e-005 3.8182 0.012025 2.4204e-005 0.0011546 0.18745 0.00065886 0.18811 0.17248 0 0.034726 0.0389 0 0.95911 0.27757 0.07702 0.010563 4.6109 0.065913 7.9878e-005 0.82417 0.0056133 0.006358 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.13467 0.94052 0.91331 0.001397 0.992 0.58834 0.0018822 0.42945 1.865 1.8644 16.004 144.9895 0.00016957 -85.6523 0.73795
1.842 0.98804 5.5141e-005 3.8182 0.012025 2.4217e-005 0.0011546 0.18749 0.00065886 0.18815 0.17251 0 0.034724 0.0389 0 0.9592 0.27761 0.077035 0.010565 4.6116 0.065924 7.9892e-005 0.82416 0.0056139 0.0063586 0.0013862 0.98694 0.9917 2.9889e-006 1.1955e-005 0.13467 0.94065 0.91338 0.001397 0.99203 0.58848 0.0018821 0.42946 1.8655 1.8648 16.004 144.9895 0.00016947 -85.6524 0.73895
1.843 0.98804 5.5141e-005 3.8182 0.012025 2.423e-005 0.0011546 0.18753 0.00065886 0.18818 0.17255 0 0.034722 0.0389 0 0.95929 0.27765 0.077049 0.010567 4.6123 0.065934 7.9906e-005 0.82415 0.0056145 0.0063592 0.0013861 0.98695 0.9917 2.9888e-006 1.1955e-005 0.13468 0.94079 0.91344 0.001397 0.99206 0.58862 0.0018821 0.42947 1.8659 1.8652 16.0039 144.9895 0.00016937 -85.6526 0.73995
1.844 0.98804 5.5141e-005 3.8182 0.012025 2.4243e-005 0.0011546 0.18757 0.00065886 0.18822 0.17259 0 0.03472 0.0389 0 0.95938 0.27769 0.077064 0.010569 4.6129 0.065945 7.9921e-005 0.82413 0.0056151 0.0063598 0.0013861 0.98695 0.9917 2.9888e-006 1.1955e-005 0.13468 0.94092 0.9135 0.001397 0.9921 0.58877 0.0018821 0.42949 1.8664 1.8657 16.0039 144.9895 0.00016927 -85.6527 0.74095
1.845 0.98804 5.514e-005 3.8182 0.012025 2.4256e-005 0.0011546 0.18761 0.00065886 0.18826 0.17262 0 0.034717 0.0389 0 0.95947 0.27773 0.077079 0.01057 4.6136 0.065956 7.9935e-005 0.82412 0.0056157 0.0063604 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.13469 0.94105 0.91357 0.001397 0.99213 0.58891 0.0018821 0.4295 1.8668 1.8661 16.0039 144.9896 0.00016918 -85.6528 0.74195
1.846 0.98804 5.514e-005 3.8182 0.012025 2.4269e-005 0.0011546 0.18764 0.00065886 0.1883 0.17266 0 0.034715 0.0389 0 0.95956 0.27778 0.077094 0.010572 4.6143 0.065967 7.9949e-005 0.82411 0.0056162 0.006361 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.13469 0.94119 0.91363 0.001397 0.99216 0.58905 0.0018821 0.42951 1.8673 1.8666 16.0039 144.9896 0.00016908 -85.6529 0.74295
1.847 0.98804 5.514e-005 3.8182 0.012025 2.4282e-005 0.0011546 0.18768 0.00065886 0.18834 0.1727 0 0.034713 0.0389 0 0.95965 0.27782 0.077108 0.010574 4.6149 0.065978 7.9963e-005 0.8241 0.0056168 0.0063616 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.1347 0.94132 0.91369 0.0013969 0.9922 0.58919 0.001882 0.42952 1.8677 1.867 16.0038 144.9896 0.00016898 -85.6531 0.74395
1.848 0.98804 5.514e-005 3.8182 0.012025 2.4296e-005 0.0011546 0.18772 0.00065886 0.18838 0.17273 0 0.034711 0.0389 0 0.95974 0.27786 0.077123 0.010575 4.6156 0.065989 7.9977e-005 0.82409 0.0056174 0.0063622 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.1347 0.94145 0.91375 0.0013969 0.99223 0.58934 0.001882 0.42954 1.8681 1.8675 16.0038 144.9896 0.00016888 -85.6532 0.74495
1.849 0.98804 5.514e-005 3.8182 0.012025 2.4309e-005 0.0011546 0.18776 0.00065886 0.18841 0.17277 0 0.034709 0.0389 0 0.95984 0.2779 0.077138 0.010577 4.6163 0.066 7.9992e-005 0.82408 0.005618 0.0063628 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.13471 0.94158 0.91381 0.0013969 0.99226 0.58948 0.001882 0.42955 1.8686 1.8679 16.0038 144.9896 0.00016879 -85.6533 0.74595
1.85 0.98804 5.514e-005 3.8182 0.012025 2.4322e-005 0.0011546 0.1878 0.00065886 0.18845 0.1728 0 0.034706 0.0389 0 0.95993 0.27794 0.077153 0.010579 4.6169 0.06601 8.0006e-005 0.82407 0.0056186 0.0063634 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.13471 0.94171 0.91388 0.0013969 0.99229 0.58962 0.001882 0.42956 1.869 1.8683 16.0038 144.9897 0.00016869 -85.6534 0.74695
1.851 0.98804 5.514e-005 3.8182 0.012025 2.4335e-005 0.0011546 0.18784 0.00065886 0.18849 0.17284 0 0.034704 0.0389 0 0.96002 0.27798 0.077168 0.010581 4.6176 0.066021 8.002e-005 0.82406 0.0056191 0.006364 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.13472 0.94184 0.91394 0.0013969 0.99232 0.58977 0.001882 0.42957 1.8695 1.8688 16.0037 144.9897 0.00016859 -85.6535 0.74795
1.852 0.98804 5.514e-005 3.8182 0.012025 2.4348e-005 0.0011546 0.18787 0.00065886 0.18853 0.17288 0 0.034702 0.0389 0 0.96011 0.27802 0.077182 0.010582 4.6183 0.066032 8.0034e-005 0.82405 0.0056197 0.0063646 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.13472 0.94197 0.914 0.0013969 0.99236 0.58991 0.0018819 0.42958 1.8699 1.8692 16.0037 144.9897 0.0001685 -85.6536 0.74895
1.853 0.98804 5.514e-005 3.8182 0.012025 2.4361e-005 0.0011546 0.18791 0.00065886 0.18857 0.17291 0 0.0347 0.0389 0 0.9602 0.27806 0.077197 0.010584 4.6189 0.066043 8.0049e-005 0.82404 0.0056203 0.0063652 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.13473 0.9421 0.91406 0.0013969 0.99239 0.59005 0.0018819 0.4296 1.8703 1.8697 16.0037 144.9897 0.0001684 -85.6538 0.74995
1.854 0.98804 5.514e-005 3.8182 0.012025 2.4374e-005 0.0011546 0.18795 0.00065886 0.1886 0.17295 0 0.034698 0.0389 0 0.96029 0.2781 0.077212 0.010586 4.6196 0.066054 8.0063e-005 0.82403 0.0056209 0.0063658 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.13473 0.94223 0.91412 0.0013968 0.99242 0.59019 0.0018819 0.42961 1.8708 1.8701 16.0036 144.9897 0.0001683 -85.6539 0.75095
1.855 0.98804 5.514e-005 3.8182 0.012025 2.4387e-005 0.0011546 0.18799 0.00065886 0.18864 0.17298 0 0.034696 0.0389 0 0.96038 0.27815 0.077227 0.010588 4.6203 0.066065 8.0077e-005 0.82402 0.0056215 0.0063664 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.13474 0.94236 0.91418 0.0013968 0.99245 0.59034 0.0018819 0.42962 1.8712 1.8705 16.0036 144.9898 0.00016821 -85.654 0.75195
1.856 0.98804 5.514e-005 3.8182 0.012025 2.44e-005 0.0011546 0.18803 0.00065886 0.18868 0.17302 0 0.034693 0.0389 0 0.96048 0.27819 0.077241 0.010589 4.6209 0.066076 8.0091e-005 0.824 0.0056221 0.006367 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.13474 0.94249 0.91424 0.0013968 0.99248 0.59048 0.0018819 0.42963 1.8716 1.871 16.0036 144.9898 0.00016811 -85.6541 0.75295
1.857 0.98804 5.514e-005 3.8182 0.012025 2.4414e-005 0.0011546 0.18806 0.00065886 0.18872 0.17306 0 0.034691 0.0389 0 0.96057 0.27823 0.077256 0.010591 4.6216 0.066086 8.0105e-005 0.82399 0.0056226 0.0063676 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.13475 0.94262 0.9143 0.0013968 0.99251 0.59062 0.0018819 0.42965 1.8721 1.8714 16.0036 144.9898 0.00016802 -85.6542 0.75395
1.858 0.98804 5.514e-005 3.8182 0.012025 2.4427e-005 0.0011546 0.1881 0.00065886 0.18876 0.17309 0 0.034689 0.0389 0 0.96066 0.27827 0.077271 0.010593 4.6223 0.066097 8.012e-005 0.82398 0.0056232 0.0063682 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.13475 0.94275 0.91436 0.0013968 0.99254 0.59076 0.0018818 0.42966 1.8725 1.8718 16.0035 144.9898 0.00016793 -85.6543 0.75495
1.859 0.98804 5.514e-005 3.8182 0.012025 2.444e-005 0.0011546 0.18814 0.00065886 0.18879 0.17313 0 0.034687 0.0389 0 0.96075 0.27831 0.077286 0.010595 4.623 0.066108 8.0134e-005 0.82397 0.0056238 0.0063688 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.13476 0.94287 0.91442 0.0013968 0.99257 0.59091 0.0018818 0.42967 1.8729 1.8723 16.0035 144.9898 0.00016783 -85.6544 0.75595
1.86 0.98804 5.514e-005 3.8182 0.012025 2.4453e-005 0.0011546 0.18818 0.00065886 0.18883 0.17316 0 0.034685 0.0389 0 0.96084 0.27835 0.077301 0.010596 4.6236 0.066119 8.0148e-005 0.82396 0.0056244 0.0063694 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.13476 0.943 0.91448 0.0013968 0.9926 0.59105 0.0018818 0.42968 1.8734 1.8727 16.0035 144.9899 0.00016774 -85.6546 0.75695
1.861 0.98804 5.5139e-005 3.8182 0.012025 2.4466e-005 0.0011546 0.18822 0.00065886 0.18887 0.1732 0 0.034683 0.0389 0 0.96093 0.27839 0.077315 0.010598 4.6243 0.06613 8.0162e-005 0.82395 0.005625 0.00637 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.13477 0.94313 0.91454 0.0013967 0.99263 0.59119 0.0018818 0.42969 1.8738 1.8731 16.0034 144.9899 0.00016764 -85.6547 0.75795
1.862 0.98804 5.5139e-005 3.8182 0.012025 2.4479e-005 0.0011546 0.18825 0.00065887 0.18891 0.17323 0 0.03468 0.0389 0 0.96103 0.27843 0.07733 0.0106 4.625 0.066141 8.0177e-005 0.82394 0.0056256 0.0063706 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.13477 0.94325 0.9146 0.0013967 0.99266 0.59133 0.0018818 0.42971 1.8742 1.8736 16.0034 144.9899 0.00016755 -85.6548 0.75895
1.863 0.98804 5.5139e-005 3.8182 0.012025 2.4492e-005 0.0011546 0.18829 0.00065887 0.18895 0.17327 0 0.034678 0.0389 0 0.96112 0.27847 0.077345 0.010602 4.6256 0.066152 8.0191e-005 0.82393 0.0056262 0.0063713 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.13478 0.94338 0.91466 0.0013967 0.99269 0.59148 0.0018817 0.42972 1.8746 1.874 16.0034 144.9899 0.00016746 -85.6549 0.75995
1.864 0.98804 5.5139e-005 3.8182 0.012025 2.4505e-005 0.0011546 0.18833 0.00065887 0.18898 0.17331 0 0.034676 0.0389 0 0.96121 0.27852 0.07736 0.010603 4.6263 0.066163 8.0205e-005 0.82392 0.0056267 0.0063719 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.13478 0.94351 0.91472 0.0013967 0.99272 0.59162 0.0018817 0.42973 1.8751 1.8744 16.0034 144.9899 0.00016737 -85.655 0.76095
1.865 0.98804 5.5139e-005 3.8182 0.012025 2.4518e-005 0.0011546 0.18837 0.00065887 0.18902 0.17334 0 0.034674 0.0389 0 0.9613 0.27856 0.077375 0.010605 4.627 0.066174 8.0219e-005 0.82391 0.0056273 0.0063725 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.13479 0.94363 0.91478 0.0013967 0.99275 0.59176 0.0018817 0.42974 1.8755 1.8748 16.0033 144.99 0.00016727 -85.6551 0.76195
1.866 0.98804 5.5139e-005 3.8182 0.012025 2.4531e-005 0.0011546 0.18841 0.00065887 0.18906 0.17338 0 0.034672 0.0389 0 0.96139 0.2786 0.077389 0.010607 4.6277 0.066184 8.0234e-005 0.8239 0.0056279 0.0063731 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.13479 0.94376 0.91483 0.0013967 0.99278 0.5919 0.0018817 0.42976 1.8759 1.8753 16.0033 144.99 0.00016718 -85.6552 0.76295
1.867 0.98804 5.5139e-005 3.8182 0.012025 2.4545e-005 0.0011546 0.18844 0.00065887 0.1891 0.17341 0 0.03467 0.0389 0 0.96148 0.27864 0.077404 0.010609 4.6283 0.066195 8.0248e-005 0.82388 0.0056285 0.0063737 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.1348 0.94388 0.91489 0.0013967 0.99281 0.59204 0.0018817 0.42977 1.8763 1.8757 16.0033 144.99 0.00016709 -85.6553 0.76395
1.868 0.98804 5.5139e-005 3.8182 0.012025 2.4558e-005 0.0011546 0.18848 0.00065887 0.18913 0.17345 0 0.034667 0.0389 0 0.96157 0.27868 0.077419 0.01061 4.629 0.066206 8.0262e-005 0.82387 0.0056291 0.0063743 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.1348 0.944 0.91495 0.0013967 0.99283 0.59219 0.0018817 0.42978 1.8768 1.8761 16.0032 144.99 0.000167 -85.6554 0.76495
1.869 0.98804 5.5139e-005 3.8182 0.012025 2.4571e-005 0.0011546 0.18852 0.00065887 0.18917 0.17348 0 0.034665 0.0389 0 0.96167 0.27872 0.077434 0.010612 4.6297 0.066217 8.0276e-005 0.82386 0.0056297 0.0063749 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.1348 0.94413 0.91501 0.0013966 0.99286 0.59233 0.0018816 0.42979 1.8772 1.8765 16.0032 144.99 0.00016691 -85.6555 0.76595
1.87 0.98804 5.5139e-005 3.8182 0.012025 2.4584e-005 0.0011546 0.18856 0.00065887 0.18921 0.17352 0 0.034663 0.0389 0 0.96176 0.27876 0.077449 0.010614 4.6304 0.066228 8.0291e-005 0.82385 0.0056303 0.0063755 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.13481 0.94425 0.91506 0.0013966 0.99289 0.59247 0.0018816 0.4298 1.8776 1.877 16.0032 144.9901 0.00016682 -85.6556 0.76695
1.871 0.98804 5.5139e-005 3.8182 0.012025 2.4597e-005 0.0011546 0.18859 0.00065887 0.18925 0.17355 0 0.034661 0.0389 0 0.96185 0.2788 0.077463 0.010616 4.631 0.066239 8.0305e-005 0.82384 0.0056308 0.0063761 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.13481 0.94437 0.91512 0.0013966 0.99292 0.59261 0.0018816 0.42982 1.878 1.8774 16.0032 144.9901 0.00016673 -85.6557 0.76795
1.872 0.98804 5.5139e-005 3.8182 0.012025 2.461e-005 0.0011546 0.18863 0.00065887 0.18929 0.17359 0 0.034659 0.0389 0 0.96194 0.27885 0.077478 0.010617 4.6317 0.06625 8.0319e-005 0.82383 0.0056314 0.0063767 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.13482 0.9445 0.91518 0.0013966 0.99295 0.59275 0.0018816 0.42983 1.8785 1.8778 16.0031 144.9901 0.00016664 -85.6558 0.76895
1.873 0.98804 5.5139e-005 3.8182 0.012025 2.4623e-005 0.0011546 0.18867 0.00065887 0.18932 0.17363 0 0.034657 0.0389 0 0.96203 0.27889 0.077493 0.010619 4.6324 0.066261 8.0333e-005 0.82382 0.005632 0.0063773 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.13482 0.94462 0.91524 0.0013966 0.99297 0.5929 0.0018816 0.42984 1.8789 1.8782 16.0031 144.9901 0.00016655 -85.6559 0.76995
1.874 0.98804 5.5139e-005 3.8182 0.012025 2.4636e-005 0.0011546 0.18871 0.00065887 0.18936 0.17366 0 0.034655 0.0389 0 0.96212 0.27893 0.077508 0.010621 4.6331 0.066271 8.0348e-005 0.82381 0.0056326 0.0063779 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.13483 0.94474 0.91529 0.0013966 0.993 0.59304 0.0018816 0.42985 1.8793 1.8786 16.0031 144.9901 0.00016646 -85.656 0.77095
1.875 0.98804 5.5139e-005 3.8182 0.012025 2.4649e-005 0.0011546 0.18874 0.00065887 0.1894 0.1737 0 0.034652 0.0389 0 0.96222 0.27897 0.077523 0.010623 4.6338 0.066282 8.0362e-005 0.8238 0.0056332 0.0063785 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.13483 0.94486 0.91535 0.0013966 0.99303 0.59318 0.0018815 0.42987 1.8797 1.8791 16.003 144.9902 0.00016637 -85.6561 0.77195
1.876 0.98804 5.5138e-005 3.8182 0.012025 2.4663e-005 0.0011546 0.18878 0.00065887 0.18944 0.17373 0 0.03465 0.0389 0 0.96231 0.27901 0.077537 0.010624 4.6344 0.066293 8.0376e-005 0.82379 0.0056338 0.0063791 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.13484 0.94498 0.91541 0.0013966 0.99305 0.59332 0.0018815 0.42988 1.8801 1.8795 16.003 144.9902 0.00016628 -85.6562 0.77295
1.877 0.98804 5.5138e-005 3.8182 0.012025 2.4676e-005 0.0011546 0.18882 0.00065887 0.18947 0.17377 0 0.034648 0.0389 0 0.9624 0.27905 0.077552 0.010626 4.6351 0.066304 8.039e-005 0.82378 0.0056344 0.0063797 0.0013853 0.98696 0.99171 2.9868e-006 1.1947e-005 0.13484 0.9451 0.91546 0.0013965 0.99308 0.59346 0.0018815 0.42989 1.8805 1.8799 16.003 144.9902 0.00016619 -85.6563 0.77395
1.878 0.98804 5.5138e-005 3.8182 0.012025 2.4689e-005 0.0011546 0.18886 0.00065887 0.18951 0.1738 0 0.034646 0.0389 0 0.96249 0.27909 0.077567 0.010628 4.6358 0.066315 8.0405e-005 0.82377 0.005635 0.0063803 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.13485 0.94522 0.91552 0.0013965 0.99311 0.5936 0.0018815 0.4299 1.881 1.8803 16.003 144.9902 0.00016611 -85.6564 0.77495
1.879 0.98804 5.5138e-005 3.8182 0.012025 2.4702e-005 0.0011546 0.18889 0.00065887 0.18955 0.17384 0 0.034644 0.0389 0 0.96258 0.27913 0.077582 0.01063 4.6365 0.066326 8.0419e-005 0.82375 0.0056355 0.006381 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.13485 0.94534 0.91557 0.0013965 0.99313 0.59375 0.0018815 0.42991 1.8814 1.8807 16.0029 144.9902 0.00016602 -85.6565 0.77595
1.88 0.98804 5.5138e-005 3.8182 0.012025 2.4715e-005 0.0011546 0.18893 0.00065887 0.18958 0.17387 0 0.034642 0.0389 0 0.96268 0.27918 0.077597 0.010631 4.6372 0.066337 8.0433e-005 0.82374 0.0056361 0.0063816 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.13486 0.94546 0.91563 0.0013965 0.99316 0.59389 0.0018815 0.42993 1.8818 1.8811 16.0029 144.9903 0.00016593 -85.6566 0.77695
1.881 0.98804 5.5138e-005 3.8182 0.012025 2.4728e-005 0.0011546 0.18897 0.00065887 0.18962 0.17391 0 0.03464 0.0389 0 0.96277 0.27922 0.077612 0.010633 4.6378 0.066348 8.0448e-005 0.82373 0.0056367 0.0063822 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.13486 0.94558 0.91569 0.0013965 0.99319 0.59403 0.0018815 0.42994 1.8822 1.8816 16.0029 144.9903 0.00016584 -85.6567 0.77795
1.882 0.98804 5.5138e-005 3.8182 0.012025 2.4741e-005 0.0011546 0.18901 0.00065887 0.18966 0.17394 0 0.034638 0.0389 0 0.96286 0.27926 0.077626 0.010635 4.6385 0.066359 8.0462e-005 0.82372 0.0056373 0.0063828 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.13487 0.9457 0.91574 0.0013965 0.99321 0.59417 0.0018814 0.42995 1.8826 1.882 16.0028 144.9903 0.00016576 -85.6568 0.77895
1.883 0.98804 5.5138e-005 3.8182 0.012025 2.4754e-005 0.0011546 0.18904 0.00065887 0.1897 0.17398 0 0.034635 0.0389 0 0.96295 0.2793 0.077641 0.010637 4.6392 0.06637 8.0476e-005 0.82371 0.0056379 0.0063834 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.13487 0.94582 0.9158 0.0013965 0.99324 0.59431 0.0018814 0.42996 1.883 1.8824 16.0028 144.9903 0.00016567 -85.6569 0.77995
1.884 0.98804 5.5138e-005 3.8182 0.012025 2.4767e-005 0.0011546 0.18908 0.00065888 0.18973 0.17401 0 0.034633 0.0389 0 0.96304 0.27934 0.077656 0.010638 4.6399 0.06638 8.049e-005 0.8237 0.0056385 0.006384 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.13488 0.94593 0.91585 0.0013965 0.99326 0.59445 0.0018814 0.42997 1.8834 1.8828 16.0028 144.9904 0.00016558 -85.657 0.78095
1.885 0.98804 5.5138e-005 3.8182 0.012025 2.478e-005 0.0011546 0.18912 0.00065888 0.18977 0.17405 0 0.034631 0.0389 0 0.96313 0.27938 0.077671 0.01064 4.6406 0.066391 8.0505e-005 0.82369 0.0056391 0.0063846 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.13488 0.94605 0.91591 0.0013964 0.99329 0.59459 0.0018814 0.42999 1.8838 1.8832 16.0028 144.9904 0.0001655 -85.6571 0.78195
1.886 0.98804 5.5138e-005 3.8182 0.012025 2.4794e-005 0.0011546 0.18915 0.00065888 0.18981 0.17408 0 0.034629 0.0389 0 0.96323 0.27942 0.077686 0.010642 4.6413 0.066402 8.0519e-005 0.82368 0.0056397 0.0063852 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.13489 0.94617 0.91596 0.0013964 0.99331 0.59473 0.0018814 0.43 1.8842 1.8836 16.0027 144.9904 0.00016541 -85.6572 0.78295
1.887 0.98804 5.5138e-005 3.8182 0.012025 2.4807e-005 0.0011546 0.18919 0.00065888 0.18985 0.17412 0 0.034627 0.0389 0 0.96332 0.27946 0.077701 0.010644 4.6419 0.066413 8.0533e-005 0.82367 0.0056403 0.0063858 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.13489 0.94629 0.91601 0.0013964 0.99334 0.59487 0.0018814 0.43001 1.8847 1.884 16.0027 144.9904 0.00016533 -85.6573 0.78395
1.888 0.98804 5.5138e-005 3.8182 0.012025 2.482e-005 0.0011546 0.18923 0.00065888 0.18988 0.17415 0 0.034625 0.0389 0 0.96341 0.27951 0.077715 0.010645 4.6426 0.066424 8.0548e-005 0.82366 0.0056409 0.0063864 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.1349 0.9464 0.91607 0.0013964 0.99337 0.59502 0.0018813 0.43002 1.8851 1.8844 16.0027 144.9904 0.00016524 -85.6574 0.78495
1.889 0.98804 5.5138e-005 3.8182 0.012025 2.4833e-005 0.0011546 0.18927 0.00065888 0.18992 0.17419 0 0.034623 0.0389 0 0.9635 0.27955 0.07773 0.010647 4.6433 0.066435 8.0562e-005 0.82365 0.0056414 0.006387 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.1349 0.94652 0.91612 0.0013964 0.99339 0.59516 0.0018813 0.43003 1.8855 1.8848 16.0026 144.9905 0.00016516 -85.6575 0.78595
1.89 0.98804 5.5138e-005 3.8182 0.012025 2.4846e-005 0.0011546 0.1893 0.00065888 0.18996 0.17422 0 0.034621 0.0389 0 0.96359 0.27959 0.077745 0.010649 4.644 0.066446 8.0576e-005 0.82363 0.005642 0.0063877 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.13491 0.94663 0.91618 0.0013964 0.99341 0.5953 0.0018813 0.43005 1.8859 1.8853 16.0026 144.9905 0.00016507 -85.6576 0.78695
1.891 0.98804 5.5138e-005 3.8182 0.012025 2.4859e-005 0.0011546 0.18934 0.00065888 0.18999 0.17426 0 0.034619 0.0389 0 0.96369 0.27963 0.07776 0.010651 4.6447 0.066457 8.059e-005 0.82362 0.0056426 0.0063883 0.001385 0.98696 0.99171 2.9861e-006 1.1944e-005 0.13491 0.94675 0.91623 0.0013964 0.99344 0.59544 0.0018813 0.43006 1.8863 1.8857 16.0026 144.9905 0.00016499 -85.6576 0.78795
1.892 0.98804 5.5137e-005 3.8182 0.012025 2.4872e-005 0.0011546 0.18938 0.00065888 0.19003 0.17429 0 0.034616 0.0389 0 0.96378 0.27967 0.077775 0.010652 4.6454 0.066468 8.0605e-005 0.82361 0.0056432 0.0063889 0.0013849 0.98696 0.99171 2.9861e-006 1.1944e-005 0.13492 0.94686 0.91628 0.0013964 0.99346 0.59558 0.0018813 0.43007 1.8867 1.8861 16.0026 144.9905 0.0001649 -85.6577 0.78895
1.893 0.98804 5.5137e-005 3.8182 0.012024 2.4885e-005 0.0011546 0.18941 0.00065888 0.19007 0.17433 0 0.034614 0.0389 0 0.96387 0.27971 0.07779 0.010654 4.646 0.066479 8.0619e-005 0.8236 0.0056438 0.0063895 0.0013849 0.98696 0.99171 2.986e-006 1.1944e-005 0.13492 0.94698 0.91634 0.0013964 0.99349 0.59572 0.0018813 0.43008 1.8871 1.8865 16.0025 144.9905 0.00016482 -85.6578 0.78995
1.894 0.98804 5.5137e-005 3.8182 0.012024 2.4898e-005 0.0011546 0.18945 0.00065888 0.1901 0.17436 0 0.034612 0.0389 0 0.96396 0.27975 0.077805 0.010656 4.6467 0.06649 8.0633e-005 0.82359 0.0056444 0.0063901 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.13493 0.94709 0.91639 0.0013964 0.99351 0.59586 0.0018813 0.4301 1.8875 1.8869 16.0025 144.9906 0.00016474 -85.6579 0.79095
1.895 0.98804 5.5137e-005 3.8182 0.012024 2.4912e-005 0.0011546 0.18949 0.00065888 0.19014 0.1744 0 0.03461 0.0389 0 0.96405 0.27979 0.07782 0.010657 4.6474 0.0665 8.0648e-005 0.82358 0.005645 0.0063907 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.13493 0.94721 0.91644 0.0013963 0.99354 0.596 0.0018812 0.43011 1.8879 1.8873 16.0025 144.9906 0.00016465 -85.658 0.79195
1.896 0.98804 5.5137e-005 3.8182 0.012024 2.4925e-005 0.0011546 0.18952 0.00065888 0.19018 0.17443 0 0.034608 0.0389 0 0.96414 0.27984 0.077834 0.010659 4.6481 0.066511 8.0662e-005 0.82357 0.0056456 0.0063913 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.13494 0.94732 0.91649 0.0013963 0.99356 0.59614 0.0018812 0.43012 1.8883 1.8877 16.0024 144.9906 0.00016457 -85.6581 0.79295
1.897 0.98804 5.5137e-005 3.8182 0.012024 2.4938e-005 0.0011546 0.18956 0.00065888 0.19021 0.17447 0 0.034606 0.0389 0 0.96424 0.27988 0.077849 0.010661 4.6488 0.066522 8.0676e-005 0.82356 0.0056462 0.0063919 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.13494 0.94743 0.91655 0.0013963 0.99358 0.59628 0.0018812 0.43013 1.8887 1.8881 16.0024 144.9906 0.00016449 -85.6582 0.79395
1.898 0.98804 5.5137e-005 3.8182 0.012024 2.4951e-005 0.0011546 0.1896 0.00065888 0.19025 0.1745 0 0.034604 0.0389 0 0.96433 0.27992 0.077864 0.010663 4.6495 0.066533 8.0691e-005 0.82355 0.0056468 0.0063926 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.13495 0.94755 0.9166 0.0013963 0.99361 0.59642 0.0018812 0.43014 1.8891 1.8885 16.0024 144.9906 0.0001644 -85.6583 0.79495
1.899 0.98804 5.5137e-005 3.8182 0.012024 2.4964e-005 0.0011546 0.18963 0.00065888 0.19029 0.17454 0 0.034602 0.0389 0 0.96442 0.27996 0.077879 0.010664 4.6502 0.066544 8.0705e-005 0.82354 0.0056474 0.0063932 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.13495 0.94766 0.91665 0.0013963 0.99363 0.59656 0.0018812 0.43016 1.8895 1.8889 16.0023 144.9907 0.00016432 -85.6583 0.79595
1.9 0.98804 5.5137e-005 3.8182 0.012024 2.4977e-005 0.0011546 0.18967 0.00065888 0.19033 0.17457 0 0.0346 0.0389 0 0.96451 0.28 0.077894 0.010666 4.6509 0.066555 8.0719e-005 0.82353 0.005648 0.0063938 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.13496 0.94777 0.9167 0.0013963 0.99365 0.5967 0.0018812 0.43017 1.8899 1.8893 16.0023 144.9907 0.00016424 -85.6584 0.79695
1.901 0.98804 5.5137e-005 3.8182 0.012024 2.499e-005 0.0011546 0.18971 0.00065888 0.19036 0.17461 0 0.034598 0.0389 0 0.9646 0.28004 0.077909 0.010668 4.6516 0.066566 8.0733e-005 0.82351 0.0056485 0.0063944 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.13496 0.94788 0.91676 0.0013963 0.99368 0.59684 0.0018812 0.43018 1.8903 1.8897 16.0023 144.9907 0.00016416 -85.6585 0.79795
1.902 0.98804 5.5137e-005 3.8182 0.012024 2.5003e-005 0.0011546 0.18974 0.00065888 0.1904 0.17464 0 0.034596 0.0389 0 0.9647 0.28008 0.077924 0.01067 4.6522 0.066577 8.0748e-005 0.8235 0.0056491 0.006395 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.13497 0.94799 0.91681 0.0013963 0.9937 0.59698 0.0018812 0.43019 1.8907 1.8901 16.0023 144.9907 0.00016408 -85.6586 0.79895
1.903 0.98804 5.5137e-005 3.8182 0.012024 2.5016e-005 0.0011546 0.18978 0.00065888 0.19044 0.17467 0 0.034594 0.0389 0 0.96479 0.28013 0.077938 0.010671 4.6529 0.066588 8.0762e-005 0.82349 0.0056497 0.0063956 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.13497 0.94811 0.91686 0.0013963 0.99372 0.59712 0.0018811 0.4302 1.8911 1.8905 16.0022 144.9907 0.000164 -85.6587 0.79995
1.904 0.98804 5.5137e-005 3.8182 0.012024 2.5029e-005 0.0011546 0.18982 0.00065888 0.19047 0.17471 0 0.034591 0.0389 0 0.96488 0.28017 0.077953 0.010673 4.6536 0.066599 8.0776e-005 0.82348 0.0056503 0.0063962 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.13498 0.94822 0.91691 0.0013962 0.99374 0.59727 0.0018811 0.43022 1.8915 1.8909 16.0022 144.9908 0.00016392 -85.6588 0.80095
1.905 0.98804 5.5137e-005 3.8182 0.012024 2.5043e-005 0.0011546 0.18985 0.00065888 0.19051 0.17474 0 0.034589 0.0389 0 0.96497 0.28021 0.077968 0.010675 4.6543 0.06661 8.0791e-005 0.82347 0.0056509 0.0063969 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.13498 0.94833 0.91696 0.0013962 0.99377 0.59741 0.0018811 0.43023 1.8919 1.8913 16.0022 144.9908 0.00016384 -85.6588 0.80195
1.906 0.98804 5.5137e-005 3.8182 0.012024 2.5056e-005 0.0011546 0.18989 0.00065888 0.19054 0.17478 0 0.034587 0.0389 0 0.96507 0.28025 0.077983 0.010677 4.655 0.066621 8.0805e-005 0.82346 0.0056515 0.0063975 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.13499 0.94844 0.91701 0.0013962 0.99379 0.59755 0.0018811 0.43024 1.8923 1.8917 16.0021 144.9908 0.00016376 -85.6589 0.80295
1.907 0.98804 5.5136e-005 3.8182 0.012024 2.5069e-005 0.0011546 0.18993 0.00065889 0.19058 0.17481 0 0.034585 0.0389 0 0.96516 0.28029 0.077998 0.010678 4.6557 0.066631 8.0819e-005 0.82345 0.0056521 0.0063981 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.13499 0.94855 0.91706 0.0013962 0.99381 0.59769 0.0018811 0.43025 1.8927 1.8921 16.0021 144.9908 0.00016368 -85.659 0.80395
1.908 0.98804 5.5136e-005 3.8182 0.012024 2.5082e-005 0.0011546 0.18996 0.00065889 0.19062 0.17485 0 0.034583 0.0389 0 0.96525 0.28033 0.078013 0.01068 4.6564 0.066642 8.0834e-005 0.82344 0.0056527 0.0063987 0.0013846 0.98696 0.99172 2.9854e-006 1.1941e-005 0.135 0.94866 0.91711 0.0013962 0.99383 0.59783 0.0018811 0.43026 1.893 1.8925 16.0021 144.9908 0.0001636 -85.6591 0.80495
1.909 0.98804 5.5136e-005 3.8182 0.012024 2.5095e-005 0.0011546 0.19 0.00065889 0.19065 0.17488 0 0.034581 0.0389 0 0.96534 0.28037 0.078028 0.010682 4.6571 0.066653 8.0848e-005 0.82343 0.0056533 0.0063993 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.135 0.94876 0.91716 0.0013962 0.99385 0.59797 0.0018811 0.43028 1.8934 1.8928 16.002 144.9909 0.00016352 -85.6592 0.80595
1.91 0.98804 5.5136e-005 3.8182 0.012024 2.5108e-005 0.0011546 0.19004 0.00065889 0.19069 0.17492 0 0.034579 0.0389 0 0.96543 0.28042 0.078043 0.010684 4.6578 0.066664 8.0862e-005 0.82342 0.0056539 0.0063999 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.135 0.94887 0.91721 0.0013962 0.99387 0.59811 0.0018811 0.43029 1.8938 1.8932 16.002 144.9909 0.00016344 -85.6592 0.80695
1.911 0.98804 5.5136e-005 3.8182 0.012024 2.5121e-005 0.0011546 0.19007 0.00065889 0.19073 0.17495 0 0.034577 0.0389 0 0.96553 0.28046 0.078058 0.010685 4.6585 0.066675 8.0877e-005 0.82341 0.0056545 0.0064005 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.13501 0.94898 0.91726 0.0013962 0.9939 0.59825 0.001881 0.4303 1.8942 1.8936 16.002 144.9909 0.00016336 -85.6593 0.80795
1.912 0.98804 5.5136e-005 3.8182 0.012024 2.5134e-005 0.0011546 0.19011 0.00065889 0.19076 0.17498 0 0.034575 0.0389 0 0.96562 0.2805 0.078073 0.010687 4.6592 0.066686 8.0891e-005 0.82339 0.0056551 0.0064012 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.13501 0.94909 0.91731 0.0013962 0.99392 0.59839 0.001881 0.43031 1.8946 1.894 16.002 144.9909 0.00016328 -85.6594 0.80895
1.913 0.98804 5.5136e-005 3.8182 0.012024 2.5147e-005 0.0011546 0.19015 0.00065889 0.1908 0.17502 0 0.034573 0.0389 0 0.96571 0.28054 0.078087 0.010689 4.6599 0.066697 8.0905e-005 0.82338 0.0056557 0.0064018 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.13502 0.9492 0.91736 0.0013962 0.99394 0.59852 0.001881 0.43032 1.895 1.8944 16.0019 144.9909 0.0001632 -85.6595 0.80995
1.914 0.98804 5.5136e-005 3.8182 0.012024 2.516e-005 0.0011546 0.19018 0.00065889 0.19084 0.17505 0 0.034571 0.0389 0 0.9658 0.28058 0.078102 0.010691 4.6606 0.066708 8.092e-005 0.82337 0.0056563 0.0064024 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.13502 0.9493 0.91741 0.0013962 0.99396 0.59866 0.001881 0.43034 1.8954 1.8948 16.0019 144.991 0.00016312 -85.6595 0.81095
1.915 0.98804 5.5136e-005 3.8182 0.012024 2.5174e-005 0.0011546 0.19022 0.00065889 0.19087 0.17509 0 0.034569 0.0389 0 0.96589 0.28062 0.078117 0.010692 4.6613 0.066719 8.0934e-005 0.82336 0.0056569 0.006403 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.13503 0.94941 0.91746 0.0013961 0.99398 0.5988 0.001881 0.43035 1.8958 1.8952 16.0019 144.991 0.00016305 -85.6596 0.81195
1.916 0.98804 5.5136e-005 3.8182 0.012024 2.5187e-005 0.0011546 0.19025 0.00065889 0.19091 0.17512 0 0.034567 0.0389 0 0.96599 0.28066 0.078132 0.010694 4.662 0.06673 8.0948e-005 0.82335 0.0056575 0.0064036 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.13503 0.94952 0.91751 0.0013961 0.994 0.59894 0.001881 0.43036 1.8962 1.8956 16.0018 144.991 0.00016297 -85.6597 0.81295
1.917 0.98804 5.5136e-005 3.8182 0.012024 2.52e-005 0.0011546 0.19029 0.00065889 0.19094 0.17516 0 0.034565 0.0389 0 0.96608 0.28071 0.078147 0.010696 4.6627 0.066741 8.0963e-005 0.82334 0.0056581 0.0064042 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.13504 0.94962 0.91756 0.0013961 0.99402 0.59908 0.001881 0.43037 1.8965 1.896 16.0018 144.991 0.00016289 -85.6598 0.81395
1.918 0.98804 5.5136e-005 3.8182 0.012024 2.5213e-005 0.0011546 0.19033 0.00065889 0.19098 0.17519 0 0.034563 0.0389 0 0.96617 0.28075 0.078162 0.010698 4.6634 0.066752 8.0977e-005 0.82333 0.0056587 0.0064049 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.13504 0.94973 0.91761 0.0013961 0.99404 0.59922 0.001881 0.43038 1.8969 1.8963 16.0018 144.991 0.00016281 -85.6598 0.81495
1.919 0.98804 5.5136e-005 3.8182 0.012024 2.5226e-005 0.0011546 0.19036 0.00065889 0.19102 0.17522 0 0.03456 0.0389 0 0.96626 0.28079 0.078177 0.0107 4.6641 0.066763 8.0991e-005 0.82332 0.0056593 0.0064055 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.13505 0.94984 0.91766 0.0013961 0.99406 0.59936 0.0018809 0.43039 1.8973 1.8967 16.0017 144.9911 0.00016274 -85.6599 0.81595
1.92 0.98804 5.5136e-005 3.8182 0.012024 2.5239e-005 0.0011546 0.1904 0.00065889 0.19105 0.17526 0 0.034558 0.0389 0 0.96636 0.28083 0.078192 0.010701 4.6648 0.066774 8.1006e-005 0.82331 0.0056599 0.0064061 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.13505 0.94994 0.91771 0.0013961 0.99408 0.5995 0.0018809 0.43041 1.8977 1.8971 16.0017 144.9911 0.00016266 -85.66 0.81695
1.921 0.98804 5.5136e-005 3.8182 0.012024 2.5252e-005 0.0011546 0.19044 0.00065889 0.19109 0.17529 0 0.034556 0.0389 0 0.96645 0.28087 0.078207 0.010703 4.6655 0.066784 8.102e-005 0.8233 0.0056605 0.0064067 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.13506 0.95005 0.91776 0.0013961 0.9941 0.59964 0.0018809 0.43042 1.8981 1.8975 16.0017 144.9911 0.00016259 -85.6601 0.81795
1.922 0.98804 5.5135e-005 3.8182 0.012024 2.5265e-005 0.0011546 0.19047 0.00065889 0.19113 0.17533 0 0.034554 0.0389 0 0.96654 0.28091 0.078222 0.010705 4.6662 0.066795 8.1034e-005 0.82329 0.0056611 0.0064073 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.13506 0.95015 0.9178 0.0013961 0.99412 0.59978 0.0018809 0.43043 1.8985 1.8979 16.0017 144.9911 0.00016251 -85.6601 0.81895
1.923 0.98804 5.5135e-005 3.8182 0.012024 2.5278e-005 0.0011546 0.19051 0.00065889 0.19116 0.17536 0 0.034552 0.0389 0 0.96663 0.28096 0.078237 0.010707 4.6669 0.066806 8.1049e-005 0.82327 0.0056617 0.006408 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.13507 0.95026 0.91785 0.0013961 0.99414 0.59992 0.0018809 0.43044 1.8988 1.8983 16.0016 144.9912 0.00016243 -85.6602 0.81995
1.924 0.98804 5.5135e-005 3.8182 0.012024 2.5292e-005 0.0011546 0.19054 0.00065889 0.1912 0.17539 0 0.03455 0.0389 0 0.96672 0.281 0.078251 0.010708 4.6676 0.066817 8.1063e-005 0.82326 0.0056623 0.0064086 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.13507 0.95036 0.9179 0.0013961 0.99416 0.60006 0.0018809 0.43045 1.8992 1.8986 16.0016 144.9912 0.00016236 -85.6603 0.82095
1.925 0.98804 5.5135e-005 3.8182 0.012024 2.5305e-005 0.0011546 0.19058 0.00065889 0.19123 0.17543 0 0.034548 0.0389 0 0.96682 0.28104 0.078266 0.01071 4.6683 0.066828 8.1077e-005 0.82325 0.0056629 0.0064092 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.13508 0.95046 0.91795 0.0013961 0.99418 0.6002 0.0018809 0.43047 1.8996 1.899 16.0016 144.9912 0.00016228 -85.6603 0.82195
1.926 0.98804 5.5135e-005 3.8182 0.012024 2.5318e-005 0.0011546 0.19062 0.00065889 0.19127 0.17546 0 0.034546 0.0389 0 0.96691 0.28108 0.078281 0.010712 4.669 0.066839 8.1092e-005 0.82324 0.0056635 0.0064098 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.13508 0.95057 0.918 0.001396 0.9942 0.60034 0.0018809 0.43048 1.9 1.8994 16.0015 144.9912 0.00016221 -85.6604 0.82295
1.927 0.98804 5.5135e-005 3.8182 0.012024 2.5331e-005 0.0011546 0.19065 0.00065889 0.19131 0.1755 0 0.034544 0.0389 0 0.967 0.28112 0.078296 0.010714 4.6697 0.06685 8.1106e-005 0.82323 0.0056641 0.0064104 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.13509 0.95067 0.91804 0.001396 0.99422 0.60048 0.0018809 0.43049 1.9004 1.8998 16.0015 144.9912 0.00016213 -85.6605 0.82395
1.928 0.98804 5.5135e-005 3.8182 0.012024 2.5344e-005 0.0011546 0.19069 0.00065889 0.19134 0.17553 0 0.034542 0.0389 0 0.96709 0.28116 0.078311 0.010715 4.6704 0.066861 8.112e-005 0.82322 0.0056647 0.0064111 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.13509 0.95077 0.91809 0.001396 0.99424 0.60062 0.0018808 0.4305 1.9007 1.9002 16.0015 144.9913 0.00016206 -85.6606 0.82495
1.929 0.98804 5.5135e-005 3.8182 0.012024 2.5357e-005 0.0011546 0.19072 0.00065889 0.19138 0.17556 0 0.03454 0.0389 0 0.96719 0.2812 0.078326 0.010717 4.6711 0.066872 8.1135e-005 0.82321 0.0056653 0.0064117 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.1351 0.95088 0.91814 0.001396 0.99426 0.60075 0.0018808 0.43051 1.9011 1.9005 16.0014 144.9913 0.00016198 -85.6606 0.82595
1.93 0.98804 5.5135e-005 3.8182 0.012024 2.537e-005 0.0011547 0.19076 0.0006589 0.19141 0.1756 0 0.034538 0.0389 0 0.96728 0.28125 0.078341 0.010719 4.6718 0.066883 8.1149e-005 0.8232 0.0056659 0.0064123 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.1351 0.95098 0.91818 0.001396 0.99428 0.60089 0.0018808 0.43053 1.9015 1.9009 16.0014 144.9913 0.00016191 -85.6607 0.82695
1.931 0.98804 5.5135e-005 3.8182 0.012024 2.5383e-005 0.0011547 0.19079 0.0006589 0.19145 0.17563 0 0.034536 0.0389 0 0.96737 0.28129 0.078356 0.010721 4.6725 0.066894 8.1163e-005 0.82319 0.0056665 0.0064129 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.13511 0.95108 0.91823 0.001396 0.9943 0.60103 0.0018808 0.43054 1.9019 1.9013 16.0014 144.9913 0.00016184 -85.6608 0.82795
1.932 0.98804 5.5135e-005 3.8182 0.012024 2.5396e-005 0.0011547 0.19083 0.0006589 0.19148 0.17566 0 0.034534 0.0389 0 0.96746 0.28133 0.078371 0.010722 4.6732 0.066905 8.1178e-005 0.82318 0.0056671 0.0064135 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.13511 0.95118 0.91828 0.001396 0.99432 0.60117 0.0018808 0.43055 1.9022 1.9017 16.0014 144.9913 0.00016176 -85.6608 0.82895
1.933 0.98804 5.5135e-005 3.8182 0.012024 2.5409e-005 0.0011547 0.19087 0.0006589 0.19152 0.1757 0 0.034532 0.0389 0 0.96756 0.28137 0.078386 0.010724 4.6739 0.066916 8.1192e-005 0.82317 0.0056677 0.0064142 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.13512 0.95128 0.91832 0.001396 0.99433 0.60131 0.0018808 0.43056 1.9026 1.9021 16.0013 144.9914 0.00016169 -85.6609 0.82995
1.934 0.98804 5.5135e-005 3.8182 0.012024 2.5423e-005 0.0011547 0.1909 0.0006589 0.19156 0.17573 0 0.03453 0.0389 0 0.96765 0.28141 0.078401 0.010726 4.6746 0.066927 8.1207e-005 0.82315 0.0056683 0.0064148 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.13512 0.95138 0.91837 0.001396 0.99435 0.60145 0.0018808 0.43057 1.903 1.9024 16.0013 144.9914 0.00016162 -85.661 0.83095
1.935 0.98804 5.5135e-005 3.8182 0.012024 2.5436e-005 0.0011547 0.19094 0.0006589 0.19159 0.17577 0 0.034528 0.0389 0 0.96774 0.28145 0.078416 0.010728 4.6753 0.066938 8.1221e-005 0.82314 0.0056689 0.0064154 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.13513 0.95148 0.91842 0.001396 0.99437 0.60159 0.0018808 0.43059 1.9034 1.9028 16.0013 144.9914 0.00016154 -85.661 0.83195
1.936 0.98804 5.5135e-005 3.8182 0.012024 2.5449e-005 0.0011547 0.19097 0.0006589 0.19163 0.1758 0 0.034526 0.0389 0 0.96783 0.2815 0.078431 0.010729 4.676 0.066949 8.1235e-005 0.82313 0.0056695 0.006416 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.13513 0.95158 0.91846 0.001396 0.99439 0.60173 0.0018808 0.4306 1.9037 1.9032 16.0012 144.9914 0.00016147 -85.6611 0.83295
1.937 0.98804 5.5135e-005 3.8182 0.012024 2.5462e-005 0.0011547 0.19101 0.0006589 0.19166 0.17583 0 0.034524 0.0389 0 0.96793 0.28154 0.078446 0.010731 4.6767 0.06696 8.125e-005 0.82312 0.0056701 0.0064167 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.13514 0.95168 0.91851 0.001396 0.99441 0.60186 0.0018807 0.43061 1.9041 1.9036 16.0012 144.9914 0.0001614 -85.6612 0.83395
1.938 0.98804 5.5134e-005 3.8182 0.012024 2.5475e-005 0.0011547 0.19104 0.0006589 0.1917 0.17587 0 0.034522 0.0389 0 0.96802 0.28158 0.078461 0.010733 4.6774 0.066971 8.1264e-005 0.82311 0.0056707 0.0064173 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.13514 0.95178 0.91856 0.0013959 0.99443 0.602 0.0018807 0.43062 1.9045 1.9039 16.0012 144.9915 0.00016133 -85.6612 0.83495
1.939 0.98804 5.5134e-005 3.8182 0.012024 2.5488e-005 0.0011547 0.19108 0.0006589 0.19173 0.1759 0 0.03452 0.0389 0 0.96811 0.28162 0.078476 0.010735 4.6781 0.066982 8.1278e-005 0.8231 0.0056713 0.0064179 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.13515 0.95188 0.9186 0.0013959 0.99444 0.60214 0.0018807 0.43063 1.9049 1.9043 16.0011 144.9915 0.00016126 -85.6613 0.83595
1.94 0.98804 5.5134e-005 3.8182 0.012024 2.5501e-005 0.0011547 0.19112 0.0006589 0.19177 0.17593 0 0.034518 0.0389 0 0.9682 0.28166 0.078491 0.010736 4.6788 0.066992 8.1293e-005 0.82309 0.0056719 0.0064185 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.13515 0.95198 0.91865 0.0013959 0.99446 0.60228 0.0018807 0.43064 1.9052 1.9047 16.0011 144.9915 0.00016118 -85.6613 0.83695
1.941 0.98804 5.5134e-005 3.8182 0.012024 2.5514e-005 0.0011547 0.19115 0.0006589 0.19181 0.17597 0 0.034516 0.0389 0 0.9683 0.2817 0.078505 0.010738 4.6795 0.067003 8.1307e-005 0.82308 0.0056725 0.0064191 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.13516 0.95208 0.91869 0.0013959 0.99448 0.60242 0.0018807 0.43066 1.9056 1.905 16.0011 144.9915 0.00016111 -85.6614 0.83795
1.942 0.98804 5.5134e-005 3.8182 0.012024 2.5527e-005 0.0011547 0.19119 0.0006589 0.19184 0.176 0 0.034514 0.0389 0 0.96839 0.28175 0.07852 0.01074 4.6802 0.067014 8.1322e-005 0.82307 0.0056731 0.0064198 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.13516 0.95218 0.91874 0.0013959 0.9945 0.60256 0.0018807 0.43067 1.906 1.9054 16.001 144.9915 0.00016104 -85.6615 0.83895
1.943 0.98804 5.5134e-005 3.8182 0.012024 2.554e-005 0.0011547 0.19122 0.0006589 0.19188 0.17603 0 0.034512 0.0389 0 0.96848 0.28179 0.078535 0.010742 4.681 0.067025 8.1336e-005 0.82306 0.0056737 0.0064204 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.13517 0.95228 0.91878 0.0013959 0.99451 0.6027 0.0018807 0.43068 1.9063 1.9058 16.001 144.9916 0.00016097 -85.6615 0.83995
1.944 0.98804 5.5134e-005 3.8182 0.012024 2.5554e-005 0.0011547 0.19126 0.0006589 0.19191 0.17607 0 0.03451 0.0389 0 0.96857 0.28183 0.07855 0.010743 4.6817 0.067036 8.135e-005 0.82305 0.0056743 0.006421 0.001384 0.98697 0.99172 2.9841e-006 1.1936e-005 0.13517 0.95237 0.91883 0.0013959 0.99453 0.60283 0.0018807 0.43069 1.9067 1.9061 16.001 144.9916 0.0001609 -85.6616 0.84095
1.945 0.98804 5.5134e-005 3.8182 0.012024 2.5567e-005 0.0011547 0.19129 0.0006589 0.19195 0.1761 0 0.034508 0.0389 0 0.96867 0.28187 0.078565 0.010745 4.6824 0.067047 8.1365e-005 0.82303 0.0056749 0.0064216 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.13518 0.95247 0.91887 0.0013959 0.99455 0.60297 0.0018807 0.4307 1.9071 1.9065 16.001 144.9916 0.00016083 -85.6617 0.84195
1.946 0.98804 5.5134e-005 3.8182 0.012024 2.558e-005 0.0011547 0.19133 0.0006589 0.19198 0.17613 0 0.034506 0.0389 0 0.96876 0.28191 0.07858 0.010747 4.6831 0.067058 8.1379e-005 0.82302 0.0056755 0.0064223 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.13518 0.95257 0.91892 0.0013959 0.99457 0.60311 0.0018807 0.43072 1.9074 1.9069 16.0009 144.9916 0.00016076 -85.6617 0.84295
1.947 0.98804 5.5134e-005 3.8182 0.012024 2.5593e-005 0.0011547 0.19136 0.0006589 0.19202 0.17617 0 0.034504 0.0389 0 0.96885 0.28195 0.078595 0.010749 4.6838 0.067069 8.1393e-005 0.82301 0.0056761 0.0064229 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.13519 0.95266 0.91896 0.0013959 0.99458 0.60325 0.0018806 0.43073 1.9078 1.9072 16.0009 144.9916 0.00016069 -85.6618 0.84395
1.948 0.98804 5.5134e-005 3.8182 0.012024 2.5606e-005 0.0011547 0.1914 0.0006589 0.19205 0.1762 0 0.034502 0.0389 0 0.96894 0.282 0.07861 0.01075 4.6845 0.06708 8.1408e-005 0.823 0.0056767 0.0064235 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.13519 0.95276 0.919 0.0013959 0.9946 0.60339 0.0018806 0.43074 1.9082 1.9076 16.0009 144.9917 0.00016062 -85.6618 0.84495
1.949 0.98804 5.5134e-005 3.8182 0.012024 2.5619e-005 0.0011547 0.19143 0.0006589 0.19209 0.17623 0 0.0345 0.0389 0 0.96904 0.28204 0.078625 0.010752 4.6852 0.067091 8.1422e-005 0.82299 0.0056773 0.0064241 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.1352 0.95286 0.91905 0.0013959 0.99462 0.60352 0.0018806 0.43075 1.9085 1.908 16.0008 144.9917 0.00016055 -85.6619 0.84595
1.95 0.98804 5.5134e-005 3.8182 0.012024 2.5632e-005 0.0011547 0.19147 0.0006589 0.19212 0.17627 0 0.034498 0.0389 0 0.96913 0.28208 0.07864 0.010754 4.6859 0.067102 8.1437e-005 0.82298 0.0056779 0.0064248 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.1352 0.95295 0.91909 0.0013959 0.99463 0.60366 0.0018806 0.43076 1.9089 1.9083 16.0008 144.9917 0.00016048 -85.662 0.84695
1.951 0.98804 5.5134e-005 3.8182 0.012024 2.5645e-005 0.0011547 0.19151 0.0006589 0.19216 0.1763 0 0.034496 0.0389 0 0.96922 0.28212 0.078655 0.010756 4.6866 0.067113 8.1451e-005 0.82297 0.0056785 0.0064254 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.13521 0.95305 0.91914 0.0013958 0.99465 0.6038 0.0018806 0.43077 1.9093 1.9087 16.0008 144.9917 0.00016041 -85.662 0.84795
1.952 0.98804 5.5134e-005 3.8182 0.012024 2.5658e-005 0.0011547 0.19154 0.0006589 0.19219 0.17633 0 0.034494 0.0389 0 0.96931 0.28216 0.07867 0.010757 4.6874 0.067124 8.1465e-005 0.82296 0.0056791 0.006426 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.13521 0.95314 0.91918 0.0013958 0.99467 0.60394 0.0018806 0.43079 1.9096 1.9091 16.0007 144.9917 0.00016034 -85.6621 0.84895
1.953 0.98804 5.5133e-005 3.8182 0.012024 2.5671e-005 0.0011547 0.19158 0.0006589 0.19223 0.17637 0 0.034492 0.0389 0 0.96941 0.2822 0.078685 0.010759 4.6881 0.067135 8.148e-005 0.82295 0.0056797 0.0064266 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.13522 0.95324 0.91922 0.0013958 0.99468 0.60408 0.0018806 0.4308 1.91 1.9094 16.0007 144.9918 0.00016027 -85.6621 0.84995
1.954 0.98804 5.5133e-005 3.8182 0.012024 2.5685e-005 0.0011547 0.19161 0.00065891 0.19227 0.1764 0 0.03449 0.0389 0 0.9695 0.28225 0.0787 0.010761 4.6888 0.067146 8.1494e-005 0.82294 0.0056803 0.0064273 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13522 0.95333 0.91927 0.0013958 0.9947 0.60421 0.0018806 0.43081 1.9103 1.9098 16.0007 144.9918 0.00016021 -85.6622 0.85095
1.955 0.98804 5.5133e-005 3.8182 0.012024 2.5698e-005 0.0011547 0.19165 0.00065891 0.1923 0.17643 0 0.034488 0.0389 0 0.96959 0.28229 0.078715 0.010763 4.6895 0.067157 8.1509e-005 0.82292 0.0056809 0.0064279 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13523 0.95343 0.91931 0.0013958 0.99471 0.60435 0.0018806 0.43082 1.9107 1.9102 16.0006 144.9918 0.00016014 -85.6622 0.85195
1.956 0.98804 5.5133e-005 3.8182 0.012024 2.5711e-005 0.0011547 0.19168 0.00065891 0.19234 0.17647 0 0.034486 0.0389 0 0.96968 0.28233 0.07873 0.010764 4.6902 0.067168 8.1523e-005 0.82291 0.0056815 0.0064285 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13523 0.95352 0.91935 0.0013958 0.99473 0.60449 0.0018806 0.43083 1.9111 1.9105 16.0006 144.9918 0.00016007 -85.6623 0.85295
1.957 0.98804 5.5133e-005 3.8182 0.012024 2.5724e-005 0.0011547 0.19172 0.00065891 0.19237 0.1765 0 0.034484 0.0389 0 0.96978 0.28237 0.078745 0.010766 4.6909 0.067179 8.1537e-005 0.8229 0.0056821 0.0064291 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.13524 0.95362 0.9194 0.0013958 0.99475 0.60463 0.0018806 0.43084 1.9114 1.9109 16.0006 144.9918 0.00016 -85.6624 0.85395
1.958 0.98804 5.5133e-005 3.8182 0.012024 2.5737e-005 0.0011547 0.19175 0.00065891 0.19241 0.17653 0 0.034482 0.0389 0 0.96987 0.28241 0.07876 0.010768 4.6916 0.06719 8.1552e-005 0.82289 0.0056827 0.0064298 0.0013839 0.98697 0.99172 2.9836e-006 1.1934e-005 0.13524 0.95371 0.91944 0.0013958 0.99476 0.60476 0.0018805 0.43086 1.9118 1.9112 16.0006 144.9919 0.00015994 -85.6624 0.85495
1.959 0.98804 5.5133e-005 3.8182 0.012024 2.575e-005 0.0011547 0.19179 0.00065891 0.19244 0.17657 0 0.03448 0.0389 0 0.96996 0.28245 0.078775 0.01077 4.6924 0.067201 8.1566e-005 0.82288 0.0056833 0.0064304 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.13525 0.9538 0.91948 0.0013958 0.99478 0.6049 0.0018805 0.43087 1.9121 1.9116 16.0005 144.9919 0.00015987 -85.6625 0.85595
1.96 0.98804 5.5133e-005 3.8182 0.012024 2.5763e-005 0.0011547 0.19182 0.00065891 0.19248 0.1766 0 0.034478 0.0389 0 0.97006 0.2825 0.07879 0.010771 4.6931 0.067212 8.1581e-005 0.82287 0.005684 0.006431 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.13525 0.9539 0.91952 0.0013958 0.99479 0.60504 0.0018805 0.43088 1.9125 1.912 16.0005 144.9919 0.0001598 -85.6625 0.85695
1.961 0.98804 5.5133e-005 3.8182 0.012024 2.5776e-005 0.0011547 0.19186 0.00065891 0.19251 0.17663 0 0.034476 0.0389 0 0.97015 0.28254 0.078805 0.010773 4.6938 0.067223 8.1595e-005 0.82286 0.0056846 0.0064317 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13526 0.95399 0.91957 0.0013958 0.99481 0.60518 0.0018805 0.43089 1.9129 1.9123 16.0005 144.9919 0.00015973 -85.6626 0.85795
1.962 0.98804 5.5133e-005 3.8182 0.012024 2.5789e-005 0.0011547 0.19189 0.00065891 0.19255 0.17667 0 0.034474 0.0389 0 0.97024 0.28258 0.07882 0.010775 4.6945 0.067234 8.1609e-005 0.82285 0.0056852 0.0064323 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13526 0.95408 0.91961 0.0013958 0.99482 0.60531 0.0018805 0.4309 1.9132 1.9127 16.0004 144.992 0.00015967 -85.6626 0.85895
1.963 0.98804 5.5133e-005 3.8182 0.012024 2.5803e-005 0.0011547 0.19193 0.00065891 0.19258 0.1767 0 0.034472 0.0389 0 0.97033 0.28262 0.078835 0.010777 4.6952 0.067245 8.1624e-005 0.82284 0.0056858 0.0064329 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13527 0.95417 0.91965 0.0013958 0.99484 0.60545 0.0018805 0.43092 1.9136 1.913 16.0004 144.992 0.0001596 -85.6627 0.85995
1.964 0.98804 5.5133e-005 3.8182 0.012024 2.5816e-005 0.0011547 0.19196 0.00065891 0.19262 0.17673 0 0.03447 0.0389 0 0.97043 0.28266 0.07885 0.010778 4.6959 0.067256 8.1638e-005 0.82283 0.0056864 0.0064335 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.13527 0.95426 0.91969 0.0013958 0.99486 0.60559 0.0018805 0.43093 1.9139 1.9134 16.0004 144.992 0.00015954 -85.6627 0.86095
1.965 0.98804 5.5133e-005 3.8182 0.012023 2.5829e-005 0.0011547 0.192 0.00065891 0.19265 0.17676 0 0.034468 0.0389 0 0.97052 0.28271 0.078865 0.01078 4.6967 0.067267 8.1653e-005 0.82281 0.005687 0.0064342 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.13528 0.95436 0.91974 0.0013958 0.99487 0.60573 0.0018805 0.43094 1.9143 1.9137 16.0003 144.992 0.00015947 -85.6628 0.86195
1.966 0.98804 5.5133e-005 3.8182 0.012023 2.5842e-005 0.0011547 0.19203 0.00065891 0.19268 0.1768 0 0.034466 0.0389 0 0.97061 0.28275 0.07888 0.010782 4.6974 0.067278 8.1667e-005 0.8228 0.0056876 0.0064348 0.0013838 0.98698 0.99172 2.9834e-006 1.1933e-005 0.13528 0.95445 0.91978 0.0013957 0.99489 0.60586 0.0018805 0.43095 1.9146 1.9141 16.0003 144.992 0.0001594 -85.6628 0.86295
1.967 0.98804 5.5133e-005 3.8182 0.012023 2.5855e-005 0.0011547 0.19207 0.00065891 0.19272 0.17683 0 0.034464 0.0389 0 0.9707 0.28279 0.078895 0.010784 4.6981 0.067289 8.1681e-005 0.82279 0.0056882 0.0064354 0.0013837 0.98698 0.99172 2.9834e-006 1.1933e-005 0.13529 0.95454 0.91982 0.0013957 0.9949 0.606 0.0018805 0.43096 1.915 1.9144 16.0003 144.9921 0.00015934 -85.6629 0.86395
1.968 0.98804 5.5133e-005 3.8182 0.012023 2.5868e-005 0.0011547 0.1921 0.00065891 0.19275 0.17686 0 0.034462 0.0389 0 0.9708 0.28283 0.07891 0.010786 4.6988 0.0673 8.1696e-005 0.82278 0.0056888 0.0064361 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.13529 0.95463 0.91986 0.0013957 0.99491 0.60614 0.0018805 0.43097 1.9153 1.9148 16.0002 144.9921 0.00015927 -85.6629 0.86495
1.969 0.98804 5.5132e-005 3.8182 0.012023 2.5881e-005 0.0011547 0.19213 0.00065891 0.19279 0.1769 0 0.03446 0.0389 0 0.97089 0.28287 0.078925 0.010787 4.6995 0.067311 8.171e-005 0.82277 0.0056894 0.0064367 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.1353 0.95472 0.9199 0.0013957 0.99493 0.60627 0.0018805 0.43099 1.9157 1.9152 16.0002 144.9921 0.00015921 -85.663 0.86595
1.97 0.98804 5.5132e-005 3.8182 0.012023 2.5894e-005 0.0011547 0.19217 0.00065891 0.19282 0.17693 0 0.034458 0.0389 0 0.97098 0.28291 0.07894 0.010789 4.7003 0.067322 8.1725e-005 0.82276 0.00569 0.0064373 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.1353 0.95481 0.91994 0.0013957 0.99494 0.60641 0.0018804 0.431 1.916 1.9155 16.0002 144.9921 0.00015914 -85.663 0.86695
1.971 0.98804 5.5132e-005 3.8182 0.012023 2.5907e-005 0.0011547 0.1922 0.00065891 0.19286 0.17696 0 0.034456 0.0389 0 0.97108 0.28296 0.078955 0.010791 4.701 0.067333 8.1739e-005 0.82275 0.0056906 0.006438 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.13531 0.9549 0.91998 0.0013957 0.99496 0.60655 0.0018804 0.43101 1.9164 1.9159 16.0001 144.9921 0.00015908 -85.6631 0.86795
1.972 0.98804 5.5132e-005 3.8182 0.012023 2.592e-005 0.0011547 0.19224 0.00065891 0.19289 0.17699 0 0.034454 0.0389 0 0.97117 0.283 0.07897 0.010793 4.7017 0.067344 8.1754e-005 0.82274 0.0056912 0.0064386 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13531 0.95499 0.92002 0.0013957 0.99497 0.60669 0.0018804 0.43102 1.9167 1.9162 16.0001 144.9922 0.00015901 -85.6631 0.86895
1.973 0.98804 5.5132e-005 3.8182 0.012023 2.5934e-005 0.0011547 0.19227 0.00065891 0.19293 0.17703 0 0.034453 0.0389 0 0.97126 0.28304 0.078985 0.010794 4.7024 0.067355 8.1768e-005 0.82273 0.0056919 0.0064392 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13532 0.95508 0.92006 0.0013957 0.99499 0.60682 0.0018804 0.43103 1.9171 1.9166 16.0001 144.9922 0.00015895 -85.6632 0.86995
1.974 0.98804 5.5132e-005 3.8182 0.012023 2.5947e-005 0.0011547 0.19231 0.00065891 0.19296 0.17706 0 0.034451 0.0389 0 0.97135 0.28308 0.079 0.010796 4.7032 0.067366 8.1782e-005 0.82272 0.0056925 0.0064398 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13532 0.95517 0.92011 0.0013957 0.995 0.60696 0.0018804 0.43104 1.9174 1.9169 16.0001 144.9922 0.00015889 -85.6632 0.87095
1.975 0.98804 5.5132e-005 3.8182 0.012023 2.596e-005 0.0011547 0.19234 0.00065891 0.193 0.17709 0 0.034449 0.0389 0 0.97145 0.28312 0.079015 0.010798 4.7039 0.067377 8.1797e-005 0.82271 0.0056931 0.0064405 0.0013836 0.98698 0.99173 2.9832e-006 1.1933e-005 0.13533 0.95526 0.92015 0.0013957 0.99502 0.6071 0.0018804 0.43106 1.9178 1.9173 16 144.9922 0.00015882 -85.6633 0.87195
1.976 0.98804 5.5132e-005 3.8182 0.012023 2.5973e-005 0.0011547 0.19238 0.00065891 0.19303 0.17712 0 0.034447 0.0389 0 0.97154 0.28317 0.07903 0.0108 4.7046 0.067388 8.1811e-005 0.82269 0.0056937 0.0064411 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.13533 0.95534 0.92019 0.0013957 0.99503 0.60723 0.0018804 0.43107 1.9181 1.9176 16 144.9922 0.00015876 -85.6633 0.87295
1.977 0.98804 5.5132e-005 3.8182 0.012023 2.5986e-005 0.0011547 0.19241 0.00065891 0.19307 0.17716 0 0.034445 0.0389 0 0.97163 0.28321 0.079045 0.010801 4.7053 0.067398 8.1826e-005 0.82268 0.0056943 0.0064417 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.13534 0.95543 0.92023 0.0013957 0.99504 0.60737 0.0018804 0.43108 1.9185 1.918 16 144.9923 0.0001587 -85.6634 0.87395
1.978 0.98804 5.5132e-005 3.8182 0.012023 2.5999e-005 0.0011547 0.19245 0.00065891 0.1931 0.17719 0 0.034443 0.0389 0 0.97173 0.28325 0.07906 0.010803 4.7061 0.067409 8.184e-005 0.82267 0.0056949 0.0064424 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.13534 0.95552 0.92027 0.0013957 0.99506 0.60751 0.0018804 0.43109 1.9188 1.9183 15.9999 144.9923 0.00015863 -85.6634 0.87495
1.979 0.98804 5.5132e-005 3.8182 0.012023 2.6012e-005 0.0011547 0.19248 0.00065892 0.19314 0.17722 0 0.034441 0.0389 0 0.97182 0.28329 0.079075 0.010805 4.7068 0.06742 8.1855e-005 0.82266 0.0056955 0.006443 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.13535 0.95561 0.92031 0.0013957 0.99507 0.60764 0.0018804 0.4311 1.9192 1.9187 15.9999 144.9923 0.00015857 -85.6635 0.87595
1.98 0.98804 5.5132e-005 3.8182 0.012023 2.6025e-005 0.0011547 0.19252 0.00065892 0.19317 0.17725 0 0.034439 0.0389 0 0.97191 0.28333 0.07909 0.010807 4.7075 0.067431 8.1869e-005 0.82265 0.0056961 0.0064436 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13535 0.95569 0.92035 0.0013957 0.99509 0.60778 0.0018804 0.43111 1.9195 1.919 15.9999 144.9923 0.00015851 -85.6635 0.87695
1.981 0.98804 5.5132e-005 3.8182 0.012023 2.6038e-005 0.0011547 0.19255 0.00065892 0.1932 0.17729 0 0.034437 0.0389 0 0.972 0.28337 0.079105 0.010808 4.7082 0.067442 8.1883e-005 0.82264 0.0056967 0.0064443 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13536 0.95578 0.92039 0.0013957 0.9951 0.60792 0.0018804 0.43113 1.9199 1.9193 15.9998 144.9923 0.00015844 -85.6636 0.87795
1.982 0.98804 5.5132e-005 3.8182 0.012023 2.6051e-005 0.0011547 0.19258 0.00065892 0.19324 0.17732 0 0.034435 0.0389 0 0.9721 0.28342 0.07912 0.01081 4.709 0.067453 8.1898e-005 0.82263 0.0056973 0.0064449 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13536 0.95587 0.92043 0.0013957 0.99511 0.60805 0.0018804 0.43114 1.9202 1.9197 15.9998 144.9924 0.00015838 -85.6636 0.87895
1.983 0.98804 5.5132e-005 3.8182 0.012023 2.6065e-005 0.0011547 0.19262 0.00065892 0.19327 0.17735 0 0.034433 0.0389 0 0.97219 0.28346 0.079136 0.010812 4.7097 0.067464 8.1912e-005 0.82262 0.005698 0.0064455 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.13537 0.95595 0.92047 0.0013956 0.99513 0.60819 0.0018803 0.43115 1.9205 1.92 15.9998 144.9924 0.00015832 -85.6637 0.87995
1.984 0.98804 5.5131e-005 3.8182 0.012023 2.6078e-005 0.0011547 0.19265 0.00065892 0.19331 0.17738 0 0.034431 0.0389 0 0.97228 0.2835 0.079151 0.010814 4.7104 0.067475 8.1927e-005 0.82261 0.0056986 0.0064462 0.0013836 0.98698 0.99173 2.9829e-006 1.1932e-005 0.13537 0.95604 0.9205 0.0013956 0.99514 0.60833 0.0018803 0.43116 1.9209 1.9204 15.9997 144.9924 0.00015826 -85.6637 0.88095
1.985 0.98804 5.5131e-005 3.8182 0.012023 2.6091e-005 0.0011547 0.19269 0.00065892 0.19334 0.17742 0 0.034429 0.0389 0 0.97238 0.28354 0.079166 0.010815 4.7111 0.067486 8.1941e-005 0.8226 0.0056992 0.0064468 0.0013835 0.98698 0.99173 2.9829e-006 1.1932e-005 0.13538 0.95613 0.92054 0.0013956 0.99515 0.60846 0.0018803 0.43117 1.9212 1.9207 15.9997 144.9924 0.0001582 -85.6638 0.88195
1.986 0.98804 5.5131e-005 3.8182 0.012023 2.6104e-005 0.0011547 0.19272 0.00065892 0.19338 0.17745 0 0.034427 0.0389 0 0.97247 0.28358 0.079181 0.010817 4.7119 0.067497 8.1956e-005 0.82258 0.0056998 0.0064474 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.13538 0.95621 0.92058 0.0013956 0.99517 0.6086 0.0018803 0.43118 1.9216 1.9211 15.9997 144.9924 0.00015814 -85.6638 0.88295
1.987 0.98804 5.5131e-005 3.8182 0.012023 2.6117e-005 0.0011547 0.19276 0.00065892 0.19341 0.17748 0 0.034425 0.0389 0 0.97256 0.28363 0.079196 0.010819 4.7126 0.067508 8.197e-005 0.82257 0.0057004 0.0064481 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.13539 0.9563 0.92062 0.0013956 0.99518 0.60873 0.0018803 0.4312 1.9219 1.9214 15.9996 144.9925 0.00015807 -85.6638 0.88395
1.988 0.98804 5.5131e-005 3.8182 0.012023 2.613e-005 0.0011547 0.19279 0.00065892 0.19344 0.17751 0 0.034423 0.0389 0 0.97266 0.28367 0.079211 0.010821 4.7133 0.067519 8.1985e-005 0.82256 0.005701 0.0064487 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13539 0.95638 0.92066 0.0013956 0.99519 0.60887 0.0018803 0.43121 1.9223 1.9217 15.9996 144.9925 0.00015801 -85.6639 0.88495
1.989 0.98804 5.5131e-005 3.8182 0.012023 2.6143e-005 0.0011547 0.19282 0.00065892 0.19348 0.17755 0 0.034422 0.0389 0 0.97275 0.28371 0.079226 0.010822 4.7141 0.06753 8.1999e-005 0.82255 0.0057016 0.0064493 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.1354 0.95647 0.9207 0.0013956 0.9952 0.60901 0.0018803 0.43122 1.9226 1.9221 15.9996 144.9925 0.00015795 -85.6639 0.88595
1.99 0.98804 5.5131e-005 3.8182 0.012023 2.6156e-005 0.0011547 0.19286 0.00065892 0.19351 0.17758 0 0.03442 0.0389 0 0.97284 0.28375 0.079241 0.010824 4.7148 0.067541 8.2013e-005 0.82254 0.0057022 0.00645 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.1354 0.95655 0.92074 0.0013956 0.99522 0.60914 0.0018803 0.43123 1.9229 1.9224 15.9995 144.9925 0.00015789 -85.664 0.88695
1.991 0.98804 5.5131e-005 3.8182 0.012023 2.6169e-005 0.0011547 0.19289 0.00065892 0.19355 0.17761 0 0.034418 0.0389 0 0.97293 0.28379 0.079256 0.010826 4.7155 0.067552 8.2028e-005 0.82253 0.0057029 0.0064506 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13541 0.95664 0.92078 0.0013956 0.99523 0.60928 0.0018803 0.43124 1.9233 1.9228 15.9995 144.9925 0.00015783 -85.664 0.88795
1.992 0.98804 5.5131e-005 3.8182 0.012023 2.6182e-005 0.0011547 0.19293 0.00065892 0.19358 0.17764 0 0.034416 0.0389 0 0.97303 0.28384 0.079271 0.010828 4.7162 0.067563 8.2042e-005 0.82252 0.0057035 0.0064512 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.13541 0.95672 0.92081 0.0013956 0.99524 0.60941 0.0018803 0.43125 1.9236 1.9231 15.9995 144.9926 0.00015777 -85.6641 0.88895
1.993 0.98804 5.5131e-005 3.8182 0.012023 2.6196e-005 0.0011547 0.19296 0.00065892 0.19361 0.17767 0 0.034414 0.0389 0 0.97312 0.28388 0.079286 0.01083 4.717 0.067574 8.2057e-005 0.82251 0.0057041 0.0064519 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13542 0.95681 0.92085 0.0013956 0.99526 0.60955 0.0018803 0.43126 1.924 1.9234 15.9994 144.9926 0.00015771 -85.6641 0.88995
1.994 0.98804 5.5131e-005 3.8182 0.012023 2.6209e-005 0.0011547 0.19299 0.00065892 0.19365 0.17771 0 0.034412 0.0389 0 0.97321 0.28392 0.079301 0.010831 4.7177 0.067585 8.2071e-005 0.8225 0.0057047 0.0064525 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13542 0.95689 0.92089 0.0013956 0.99527 0.60969 0.0018803 0.43128 1.9243 1.9238 15.9994 144.9926 0.00015765 -85.6641 0.89095
1.995 0.98804 5.5131e-005 3.8182 0.012023 2.6222e-005 0.0011547 0.19303 0.00065892 0.19368 0.17774 0 0.03441 0.0389 0 0.97331 0.28396 0.079316 0.010833 4.7184 0.067596 8.2086e-005 0.82249 0.0057053 0.0064532 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13543 0.95697 0.92093 0.0013956 0.99528 0.60982 0.0018803 0.43129 1.9246 1.9241 15.9994 144.9926 0.00015759 -85.6642 0.89195
1.996 0.98804 5.5131e-005 3.8182 0.012023 2.6235e-005 0.0011547 0.19306 0.00065892 0.19372 0.17777 0 0.034408 0.0389 0 0.9734 0.284 0.079331 0.010835 4.7192 0.067607 8.21e-005 0.82247 0.0057059 0.0064538 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.13543 0.95705 0.92097 0.0013956 0.99529 0.60996 0.0018803 0.4313 1.925 1.9245 15.9994 144.9926 0.00015753 -85.6642 0.89295
1.997 0.98804 5.5131e-005 3.8182 0.012023 2.6248e-005 0.0011547 0.1931 0.00065892 0.19375 0.1778 0 0.034406 0.0389 0 0.97349 0.28405 0.079346 0.010837 4.7199 0.067618 8.2115e-005 0.82246 0.0057065 0.0064544 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13544 0.95714 0.921 0.0013956 0.9953 0.61009 0.0018802 0.43131 1.9253 1.9248 15.9993 144.9927 0.00015747 -85.6643 0.89395
1.998 0.98804 5.5131e-005 3.8182 0.012023 2.6261e-005 0.0011547 0.19313 0.00065892 0.19378 0.17783 0 0.034404 0.0389 0 0.97359 0.28409 0.079361 0.010838 4.7206 0.067629 8.2129e-005 0.82245 0.0057071 0.0064551 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13544 0.95722 0.92104 0.0013956 0.99532 0.61023 0.0018802 0.43132 1.9256 1.9251 15.9993 144.9927 0.00015741 -85.6643 0.89495
1.999 0.98804 5.513e-005 3.8182 0.012023 2.6274e-005 0.0011547 0.19316 0.00065892 0.19382 0.17787 0 0.034402 0.0389 0 0.97368 0.28413 0.079376 0.01084 4.7214 0.06764 8.2144e-005 0.82244 0.0057078 0.0064557 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13545 0.9573 0.92108 0.0013956 0.99533 0.61036 0.0018802 0.43133 1.926 1.9255 15.9993 144.9927 0.00015735 -85.6644 0.89595
2 0.98804 5.513e-005 3.8182 0.012023 2.6287e-005 0.0011547 0.1932 0.00065892 0.19385 0.1779 0 0.034401 0.0389 0 0.97377 0.28417 0.079391 0.010842 4.7221 0.067651 8.2158e-005 0.82243 0.0057084 0.0064563 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13545 0.95738 0.92112 0.0013956 0.99534 0.6105 0.0018802 0.43135 1.9263 1.9258 15.9992 144.9927 0.0001573 -85.6644 0.89695
2.001 0.98804 5.513e-005 3.8182 0.012023 2.63e-005 0.0011547 0.19323 0.00065892 0.19389 0.17793 0 0.034399 0.0389 0 0.97387 0.28421 0.079407 0.010844 4.7228 0.067662 8.2173e-005 0.82242 0.005709 0.006457 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.13546 0.95747 0.92115 0.0013956 0.99535 0.61064 0.0018802 0.43136 1.9266 1.9261 15.9992 144.9928 0.00015724 -85.6644 0.89795
2.002 0.98804 5.513e-005 3.8182 0.012023 2.6313e-005 0.0011547 0.19327 0.00065892 0.19392 0.17796 0 0.034397 0.0389 0 0.97396 0.28426 0.079422 0.010845 4.7236 0.067673 8.2187e-005 0.82241 0.0057096 0.0064576 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.13546 0.95755 0.92119 0.0013955 0.99536 0.61077 0.0018802 0.43137 1.927 1.9265 15.9992 144.9928 0.00015718 -85.6645 0.89895
2.003 0.98804 5.513e-005 3.8182 0.012023 2.6327e-005 0.0011547 0.1933 0.00065892 0.19395 0.17799 0 0.034395 0.0389 0 0.97405 0.2843 0.079437 0.010847 4.7243 0.067684 8.2201e-005 0.8224 0.0057102 0.0064582 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.13547 0.95763 0.92123 0.0013955 0.99538 0.61091 0.0018802 0.43138 1.9273 1.9268 15.9991 144.9928 0.00015712 -85.6645 0.89995
2.004 0.98804 5.513e-005 3.8182 0.012023 2.634e-005 0.0011547 0.19333 0.00065893 0.19399 0.17803 0 0.034393 0.0389 0 0.97415 0.28434 0.079452 0.010849 4.7251 0.067695 8.2216e-005 0.82239 0.0057108 0.0064589 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.13547 0.95771 0.92126 0.0013955 0.99539 0.61104 0.0018802 0.43139 1.9276 1.9271 15.9991 144.9928 0.00015706 -85.6646 0.90095
2.005 0.98804 5.513e-005 3.8182 0.012023 2.6353e-005 0.0011547 0.19337 0.00065893 0.19402 0.17806 0 0.034391 0.0389 0 0.97424 0.28438 0.079467 0.010851 4.7258 0.067707 8.223e-005 0.82238 0.0057114 0.0064595 0.0013833 0.98698 0.99173 2.9825e-006 1.193e-005 0.13548 0.95779 0.9213 0.0013955 0.9954 0.61118 0.0018802 0.4314 1.928 1.9275 15.9991 144.9928 0.000157 -85.6646 0.90195
2.006 0.98804 5.513e-005 3.8182 0.012023 2.6366e-005 0.0011547 0.1934 0.00065893 0.19406 0.17809 0 0.034389 0.0389 0 0.97433 0.28442 0.079482 0.010852 4.7265 0.067718 8.2245e-005 0.82236 0.0057121 0.0064602 0.0013833 0.98698 0.99173 2.9825e-006 1.193e-005 0.13548 0.95787 0.92134 0.0013955 0.99541 0.61131 0.0018802 0.43141 1.9283 1.9278 15.999 144.9929 0.00015695 -85.6646 0.90295
2.007 0.98804 5.513e-005 3.8182 0.012023 2.6379e-005 0.0011547 0.19343 0.00065893 0.19409 0.17812 0 0.034387 0.0389 0 0.97442 0.28447 0.079497 0.010854 4.7273 0.067729 8.2259e-005 0.82235 0.0057127 0.0064608 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.13549 0.95795 0.92137 0.0013955 0.99542 0.61145 0.0018802 0.43143 1.9286 1.9281 15.999 144.9929 0.00015689 -85.6647 0.90395
2.008 0.98804 5.513e-005 3.8182 0.012023 2.6392e-005 0.0011547 0.19347 0.00065893 0.19412 0.17815 0 0.034385 0.0389 0 0.97452 0.28451 0.079512 0.010856 4.728 0.06774 8.2274e-005 0.82234 0.0057133 0.0064614 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.13549 0.95803 0.92141 0.0013955 0.99543 0.61158 0.0018802 0.43144 1.929 1.9285 15.999 144.9929 0.00015683 -85.6647 0.90495
2.009 0.98804 5.513e-005 3.8182 0.012023 2.6405e-005 0.0011547 0.1935 0.00065893 0.19416 0.17819 0 0.034383 0.0389 0 0.97461 0.28455 0.079527 0.010858 4.7287 0.067751 8.2288e-005 0.82233 0.0057139 0.0064621 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.1355 0.95811 0.92145 0.0013955 0.99545 0.61172 0.0018802 0.43145 1.9293 1.9288 15.9989 144.9929 0.00015678 -85.6647 0.90595
2.01 0.98804 5.513e-005 3.8182 0.012023 2.6418e-005 0.0011547 0.19354 0.00065893 0.19419 0.17822 0 0.034382 0.0389 0 0.9747 0.28459 0.079542 0.010859 4.7295 0.067762 8.2303e-005 0.82232 0.0057145 0.0064627 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.1355 0.95819 0.92148 0.0013955 0.99546 0.61185 0.0018802 0.43146 1.9296 1.9291 15.9989 144.9929 0.00015672 -85.6648 0.90695
2.011 0.98804 5.513e-005 3.8182 0.012023 2.6431e-005 0.0011547 0.19357 0.00065893 0.19422 0.17825 0 0.03438 0.0389 0 0.9748 0.28463 0.079557 0.010861 4.7302 0.067773 8.2317e-005 0.82231 0.0057151 0.0064634 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.13551 0.95827 0.92152 0.0013955 0.99547 0.61199 0.0018802 0.43147 1.9299 1.9295 15.9989 144.993 0.00015666 -85.6648 0.90795
2.012 0.98804 5.513e-005 3.8182 0.012023 2.6444e-005 0.0011547 0.1936 0.00065893 0.19426 0.17828 0 0.034378 0.0389 0 0.97489 0.28468 0.079572 0.010863 4.731 0.067784 8.2332e-005 0.8223 0.0057158 0.006464 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13551 0.95835 0.92155 0.0013955 0.99548 0.61212 0.0018802 0.43148 1.9303 1.9298 15.9988 144.993 0.00015661 -85.6649 0.90895
2.013 0.98804 5.513e-005 3.8182 0.012023 2.6458e-005 0.0011547 0.19364 0.00065893 0.19429 0.17831 0 0.034376 0.0389 0 0.97498 0.28472 0.079588 0.010865 4.7317 0.067795 8.2346e-005 0.82229 0.0057164 0.0064646 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13552 0.95843 0.92159 0.0013955 0.99549 0.61226 0.0018801 0.43149 1.9306 1.9301 15.9988 144.993 0.00015655 -85.6649 0.90995
2.014 0.98804 5.513e-005 3.8182 0.012023 2.6471e-005 0.0011547 0.19367 0.00065893 0.19432 0.17834 0 0.034374 0.0389 0 0.97508 0.28476 0.079603 0.010867 4.7324 0.067806 8.2361e-005 0.82228 0.005717 0.0064653 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13552 0.95851 0.92162 0.0013955 0.9955 0.61239 0.0018801 0.43151 1.9309 1.9304 15.9988 144.993 0.00015649 -85.6649 0.91095
2.015 0.98804 5.5129e-005 3.8182 0.012023 2.6484e-005 0.0011547 0.1937 0.00065893 0.19436 0.17838 0 0.034372 0.0389 0 0.97517 0.2848 0.079618 0.010868 4.7332 0.067817 8.2375e-005 0.82227 0.0057176 0.0064659 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13553 0.95858 0.92166 0.0013955 0.99551 0.61253 0.0018801 0.43152 1.9313 1.9308 15.9987 144.993 0.00015644 -85.665 0.91195
2.016 0.98804 5.5129e-005 3.8182 0.012023 2.6497e-005 0.0011547 0.19374 0.00065893 0.19439 0.17841 0 0.03437 0.0389 0 0.97526 0.28484 0.079633 0.01087 4.7339 0.067828 8.239e-005 0.82225 0.0057182 0.0064666 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.13554 0.95866 0.9217 0.0013955 0.99552 0.61266 0.0018801 0.43153 1.9316 1.9311 15.9987 144.9931 0.00015638 -85.665 0.91295
2.017 0.98804 5.5129e-005 3.8182 0.012023 2.651e-005 0.0011547 0.19377 0.00065893 0.19442 0.17844 0 0.034368 0.0389 0 0.97536 0.28489 0.079648 0.010872 4.7347 0.067839 8.2404e-005 0.82224 0.0057188 0.0064672 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13554 0.95874 0.92173 0.0013955 0.99553 0.6128 0.0018801 0.43154 1.9319 1.9314 15.9987 144.9931 0.00015633 -85.665 0.91395
2.018 0.98804 5.5129e-005 3.8182 0.012023 2.6523e-005 0.0011547 0.1938 0.00065893 0.19446 0.17847 0 0.034367 0.0389 0 0.97545 0.28493 0.079663 0.010874 4.7354 0.06785 8.2419e-005 0.82223 0.0057195 0.0064678 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13555 0.95882 0.92177 0.0013955 0.99554 0.61293 0.0018801 0.43155 1.9322 1.9317 15.9986 144.9931 0.00015627 -85.6651 0.91495
2.019 0.98804 5.5129e-005 3.8182 0.012023 2.6536e-005 0.0011547 0.19384 0.00065893 0.19449 0.1785 0 0.034365 0.0389 0 0.97554 0.28497 0.079678 0.010875 4.7361 0.067861 8.2433e-005 0.82222 0.0057201 0.0064685 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13555 0.95889 0.9218 0.0013955 0.99555 0.61307 0.0018801 0.43156 1.9326 1.9321 15.9986 144.9931 0.00015622 -85.6651 0.91595
2.02 0.98804 5.5129e-005 3.8182 0.012023 2.6549e-005 0.0011547 0.19387 0.00065893 0.19452 0.17853 0 0.034363 0.0389 0 0.97564 0.28501 0.079693 0.010877 4.7369 0.067872 8.2448e-005 0.82221 0.0057207 0.0064691 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13556 0.95897 0.92184 0.0013955 0.99557 0.6132 0.0018801 0.43158 1.9329 1.9324 15.9986 144.9931 0.00015616 -85.6651 0.91695
2.021 0.98804 5.5129e-005 3.8182 0.012023 2.6562e-005 0.0011547 0.1939 0.00065893 0.19456 0.17856 0 0.034361 0.0389 0 0.97573 0.28505 0.079708 0.010879 4.7376 0.067883 8.2462e-005 0.8222 0.0057213 0.0064698 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.13556 0.95905 0.92187 0.0013955 0.99558 0.61334 0.0018801 0.43159 1.9332 1.9327 15.9985 144.9932 0.00015611 -85.6652 0.91795
2.022 0.98804 5.5129e-005 3.8182 0.012023 2.6575e-005 0.0011547 0.19394 0.00065893 0.19459 0.1786 0 0.034359 0.0389 0 0.97582 0.2851 0.079724 0.010881 4.7384 0.067894 8.2477e-005 0.82219 0.0057219 0.0064704 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13557 0.95913 0.92191 0.0013955 0.99559 0.61347 0.0018801 0.4316 1.9335 1.933 15.9985 144.9932 0.00015605 -85.6652 0.91895
2.023 0.98804 5.5129e-005 3.8182 0.012023 2.6589e-005 0.0011547 0.19397 0.00065893 0.19462 0.17863 0 0.034357 0.0389 0 0.97592 0.28514 0.079739 0.010882 4.7391 0.067905 8.2491e-005 0.82218 0.0057226 0.006471 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13557 0.9592 0.92194 0.0013955 0.9956 0.61361 0.0018801 0.43161 1.9338 1.9334 15.9985 144.9932 0.000156 -85.6652 0.91995
2.024 0.98804 5.5129e-005 3.8182 0.012023 2.6602e-005 0.0011547 0.194 0.00065893 0.19466 0.17866 0 0.034355 0.0389 0 0.97601 0.28518 0.079754 0.010884 4.7399 0.067916 8.2506e-005 0.82217 0.0057232 0.0064717 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13558 0.95928 0.92197 0.0013955 0.99561 0.61374 0.0018801 0.43162 1.9342 1.9337 15.9984 144.9932 0.00015594 -85.6653 0.92095
2.025 0.98804 5.5129e-005 3.8182 0.012023 2.6615e-005 0.0011547 0.19404 0.00065893 0.19469 0.17869 0 0.034353 0.0389 0 0.9761 0.28522 0.079769 0.010886 4.7406 0.067927 8.252e-005 0.82216 0.0057238 0.0064723 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13558 0.95935 0.92201 0.0013954 0.99562 0.61388 0.0018801 0.43163 1.9345 1.934 15.9984 144.9932 0.00015589 -85.6653 0.92195
2.026 0.98804 5.5129e-005 3.8182 0.012023 2.6628e-005 0.0011547 0.19407 0.00065893 0.19472 0.17872 0 0.034352 0.0389 0 0.9762 0.28526 0.079784 0.010888 4.7414 0.067938 8.2535e-005 0.82214 0.0057244 0.006473 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13559 0.95943 0.92204 0.0013954 0.99563 0.61401 0.0018801 0.43164 1.9348 1.9343 15.9984 144.9933 0.00015583 -85.6653 0.92295
2.027 0.98804 5.5129e-005 3.8182 0.012023 2.6641e-005 0.0011547 0.1941 0.00065893 0.19476 0.17875 0 0.03435 0.0389 0 0.97629 0.28531 0.079799 0.010889 4.7421 0.067949 8.2549e-005 0.82213 0.005725 0.0064736 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.13559 0.9595 0.92208 0.0013954 0.99564 0.61414 0.0018801 0.43165 1.9351 1.9346 15.9983 144.9933 0.00015578 -85.6654 0.92395
2.028 0.98804 5.5129e-005 3.8182 0.012023 2.6654e-005 0.0011547 0.19414 0.00065893 0.19479 0.17878 0 0.034348 0.0389 0 0.97638 0.28535 0.079814 0.010891 4.7429 0.06796 8.2564e-005 0.82212 0.0057257 0.0064743 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.1356 0.95958 0.92211 0.0013954 0.99565 0.61428 0.0018801 0.43167 1.9354 1.935 15.9983 144.9933 0.00015573 -85.6654 0.92495
2.029 0.98804 5.5129e-005 3.8182 0.012023 2.6667e-005 0.0011547 0.19417 0.00065893 0.19482 0.17881 0 0.034346 0.0389 0 0.97648 0.28539 0.079829 0.010893 4.7436 0.067971 8.2578e-005 0.82211 0.0057263 0.0064749 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.1356 0.95965 0.92215 0.0013954 0.99566 0.61441 0.0018801 0.43168 1.9358 1.9353 15.9983 144.9933 0.00015567 -85.6654 0.92595
2.03 0.98804 5.5128e-005 3.8182 0.012023 2.668e-005 0.0011547 0.1942 0.00065894 0.19486 0.17885 0 0.034344 0.0389 0 0.97657 0.28543 0.079845 0.010895 4.7444 0.067982 8.2593e-005 0.8221 0.0057269 0.0064755 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.13561 0.95973 0.92218 0.0013954 0.99567 0.61455 0.0018801 0.43169 1.9361 1.9356 15.9982 144.9933 0.00015562 -85.6655 0.92695
2.031 0.98804 5.5128e-005 3.8182 0.012023 2.6693e-005 0.0011547 0.19423 0.00065894 0.19489 0.17888 0 0.034342 0.0389 0 0.97667 0.28548 0.07986 0.010897 4.7451 0.067993 8.2607e-005 0.82209 0.0057275 0.0064762 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.13561 0.9598 0.92221 0.0013954 0.99568 0.61468 0.0018801 0.4317 1.9364 1.9359 15.9982 144.9934 0.00015557 -85.6655 0.92795
2.032 0.98804 5.5128e-005 3.8182 0.012023 2.6706e-005 0.0011547 0.19427 0.00065894 0.19492 0.17891 0 0.03434 0.0389 0 0.97676 0.28552 0.079875 0.010898 4.7458 0.068004 8.2622e-005 0.82208 0.0057281 0.0064768 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.13562 0.95988 0.92225 0.0013954 0.99569 0.61481 0.00188 0.43171 1.9367 1.9362 15.9982 144.9934 0.00015551 -85.6655 0.92895
2.033 0.98804 5.5128e-005 3.8182 0.012023 2.672e-005 0.0011547 0.1943 0.00065894 0.19496 0.17894 0 0.034339 0.0389 0 0.97685 0.28556 0.07989 0.0109 4.7466 0.068015 8.2636e-005 0.82207 0.0057288 0.0064775 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.13562 0.95995 0.92228 0.0013954 0.9957 0.61495 0.00188 0.43172 1.937 1.9366 15.9982 144.9934 0.00015546 -85.6656 0.92995
2.034 0.98804 5.5128e-005 3.8182 0.012023 2.6733e-005 0.0011547 0.19433 0.00065894 0.19499 0.17897 0 0.034337 0.0389 0 0.97695 0.2856 0.079905 0.010902 4.7473 0.068026 8.2651e-005 0.82206 0.0057294 0.0064781 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.13563 0.96003 0.92231 0.0013954 0.99571 0.61508 0.00188 0.43173 1.9374 1.9369 15.9981 144.9934 0.00015541 -85.6656 0.93095
2.035 0.98804 5.5128e-005 3.8182 0.012023 2.6746e-005 0.0011547 0.19437 0.00065894 0.19502 0.179 0 0.034335 0.0389 0 0.97704 0.28564 0.07992 0.010904 4.7481 0.068037 8.2665e-005 0.82205 0.00573 0.0064788 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.13563 0.9601 0.92235 0.0013954 0.99572 0.61522 0.00188 0.43175 1.9377 1.9372 15.9981 144.9935 0.00015536 -85.6656 0.93195
2.036 0.98804 5.5128e-005 3.8182 0.012022 2.6759e-005 0.0011547 0.1944 0.00065894 0.19505 0.17903 0 0.034333 0.0389 0 0.97713 0.28569 0.079935 0.010905 4.7488 0.068048 8.268e-005 0.82203 0.0057306 0.0064794 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.13564 0.96017 0.92238 0.0013954 0.99572 0.61535 0.00188 0.43176 1.938 1.9375 15.9981 144.9935 0.00015531 -85.6656 0.93295
2.037 0.98804 5.5128e-005 3.8182 0.012022 2.6772e-005 0.0011547 0.19443 0.00065894 0.19509 0.17906 0 0.034331 0.0389 0 0.97723 0.28573 0.07995 0.010907 4.7496 0.068059 8.2694e-005 0.82202 0.0057312 0.0064801 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.13564 0.96025 0.92241 0.0013954 0.99573 0.61548 0.00188 0.43177 1.9383 1.9378 15.998 144.9935 0.00015525 -85.6657 0.93395
2.038 0.98804 5.5128e-005 3.8182 0.012022 2.6785e-005 0.0011547 0.19447 0.00065894 0.19512 0.17909 0 0.034329 0.0389 0 0.97732 0.28577 0.079966 0.010909 4.7504 0.06807 8.2709e-005 0.82201 0.0057319 0.0064807 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.13565 0.96032 0.92245 0.0013954 0.99574 0.61562 0.00188 0.43178 1.9386 1.9381 15.998 144.9935 0.0001552 -85.6657 0.93495
2.039 0.98804 5.5128e-005 3.8182 0.012022 2.6798e-005 0.0011547 0.1945 0.00065894 0.19515 0.17913 0 0.034328 0.0389 0 0.97741 0.28581 0.079981 0.010911 4.7511 0.068081 8.2723e-005 0.822 0.0057325 0.0064814 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.13565 0.96039 0.92248 0.0013954 0.99575 0.61575 0.00188 0.43179 1.9389 1.9385 15.998 144.9935 0.00015515 -85.6657 0.93595
2.04 0.98804 5.5128e-005 3.8182 0.012022 2.6811e-005 0.0011547 0.19453 0.00065894 0.19519 0.17916 0 0.034326 0.0389 0 0.97751 0.28585 0.079996 0.010912 4.7519 0.068092 8.2738e-005 0.82199 0.0057331 0.006482 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.13566 0.96046 0.92251 0.0013954 0.99576 0.61589 0.00188 0.4318 1.9392 1.9388 15.9979 144.9936 0.0001551 -85.6658 0.93695
2.041 0.98804 5.5128e-005 3.8182 0.012022 2.6824e-005 0.0011547 0.19456 0.00065894 0.19522 0.17919 0 0.034324 0.0389 0 0.9776 0.2859 0.080011 0.010914 4.7526 0.068103 8.2752e-005 0.82198 0.0057337 0.0064826 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13566 0.96053 0.92254 0.0013954 0.99577 0.61602 0.00188 0.43181 1.9396 1.9391 15.9979 144.9936 0.00015505 -85.6658 0.93795
2.042 0.98804 5.5128e-005 3.8182 0.012022 2.6837e-005 0.0011547 0.1946 0.00065894 0.19525 0.17922 0 0.034322 0.0389 0 0.97769 0.28594 0.080026 0.010916 4.7534 0.068114 8.2767e-005 0.82197 0.0057344 0.0064833 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13567 0.96061 0.92258 0.0013954 0.99578 0.61615 0.00188 0.43183 1.9399 1.9394 15.9979 144.9936 0.000155 -85.6658 0.93895
2.043 0.98804 5.5128e-005 3.8182 0.012022 2.685e-005 0.0011548 0.19463 0.00065894 0.19528 0.17925 0 0.03432 0.0389 0 0.97779 0.28598 0.080041 0.010918 4.7541 0.068125 8.2781e-005 0.82196 0.005735 0.0064839 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.13567 0.96068 0.92261 0.0013954 0.99579 0.61629 0.00188 0.43184 1.9402 1.9397 15.9978 144.9936 0.00015494 -85.6659 0.93995
2.044 0.98804 5.5128e-005 3.8182 0.012022 2.6864e-005 0.0011548 0.19466 0.00065894 0.19532 0.17928 0 0.034318 0.0389 0 0.97788 0.28602 0.080056 0.010919 4.7549 0.068137 8.2796e-005 0.82195 0.0057356 0.0064846 0.0013831 0.98699 0.99173 2.9818e-006 1.1927e-005 0.13568 0.96075 0.92264 0.0013954 0.9958 0.61642 0.00188 0.43185 1.9405 1.94 15.9978 144.9936 0.00015489 -85.6659 0.94095
2.045 0.98804 5.5127e-005 3.8182 0.012022 2.6877e-005 0.0011548 0.19469 0.00065894 0.19535 0.17931 0 0.034317 0.0389 0 0.97798 0.28607 0.080072 0.010921 4.7556 0.068148 8.281e-005 0.82194 0.0057362 0.0064852 0.001383 0.98699 0.99173 2.9818e-006 1.1927e-005 0.13568 0.96082 0.92267 0.0013954 0.99581 0.61655 0.00188 0.43186 1.9408 1.9403 15.9978 144.9937 0.00015484 -85.6659 0.94195
2.046 0.98804 5.5127e-005 3.8182 0.012022 2.689e-005 0.0011548 0.19473 0.00065894 0.19538 0.17934 0 0.034315 0.0389 0 0.97807 0.28611 0.080087 0.010923 4.7564 0.068159 8.2825e-005 0.82192 0.0057368 0.0064859 0.001383 0.98699 0.99173 2.9818e-006 1.1927e-005 0.13569 0.96089 0.9227 0.0013954 0.99582 0.61669 0.00188 0.43187 1.9411 1.9407 15.9977 144.9937 0.00015479 -85.6659 0.94295
2.047 0.98804 5.5127e-005 3.8182 0.012022 2.6903e-005 0.0011548 0.19476 0.00065894 0.19541 0.17937 0 0.034313 0.0389 0 0.97816 0.28615 0.080102 0.010925 4.7571 0.06817 8.2839e-005 0.82191 0.0057375 0.0064865 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13569 0.96096 0.92274 0.0013954 0.99582 0.61682 0.00188 0.43188 1.9414 1.941 15.9977 144.9937 0.00015474 -85.666 0.94395
2.048 0.98804 5.5127e-005 3.8182 0.012022 2.6916e-005 0.0011548 0.19479 0.00065894 0.19545 0.1794 0 0.034311 0.0389 0 0.97826 0.28619 0.080117 0.010927 4.7579 0.068181 8.2854e-005 0.8219 0.0057381 0.0064872 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.1357 0.96103 0.92277 0.0013954 0.99583 0.61695 0.00188 0.43189 1.9417 1.9413 15.9977 144.9937 0.00015469 -85.666 0.94495
2.049 0.98804 5.5127e-005 3.8182 0.012022 2.6929e-005 0.0011548 0.19483 0.00065894 0.19548 0.17943 0 0.034309 0.0389 0 0.97835 0.28624 0.080132 0.010928 4.7586 0.068192 8.2868e-005 0.82189 0.0057387 0.0064878 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.1357 0.9611 0.9228 0.0013954 0.99584 0.61709 0.00188 0.4319 1.942 1.9416 15.9976 144.9937 0.00015464 -85.666 0.94595
2.05 0.98804 5.5127e-005 3.8182 0.012022 2.6942e-005 0.0011548 0.19486 0.00065894 0.19551 0.17947 0 0.034307 0.0389 0 0.97844 0.28628 0.080147 0.01093 4.7594 0.068203 8.2883e-005 0.82188 0.0057393 0.0064885 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13571 0.96117 0.92283 0.0013954 0.99585 0.61722 0.00188 0.43192 1.9423 1.9419 15.9976 144.9938 0.00015459 -85.666 0.94695
2.051 0.98804 5.5127e-005 3.8182 0.012022 2.6955e-005 0.0011548 0.19489 0.00065894 0.19554 0.1795 0 0.034306 0.0389 0 0.97854 0.28632 0.080163 0.010932 4.7602 0.068214 8.2898e-005 0.82187 0.00574 0.0064891 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13571 0.96124 0.92286 0.0013954 0.99586 0.61735 0.00188 0.43193 1.9427 1.9422 15.9976 144.9938 0.00015454 -85.6661 0.94795
2.052 0.98804 5.5127e-005 3.8182 0.012022 2.6968e-005 0.0011548 0.19492 0.00065894 0.19558 0.17953 0 0.034304 0.0389 0 0.97863 0.28636 0.080178 0.010934 4.7609 0.068225 8.2912e-005 0.82186 0.0057406 0.0064898 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13572 0.96131 0.92289 0.0013954 0.99587 0.61749 0.00188 0.43194 1.943 1.9425 15.9975 144.9938 0.00015449 -85.6661 0.94895
2.053 0.98804 5.5127e-005 3.8182 0.012022 2.6981e-005 0.0011548 0.19496 0.00065894 0.19561 0.17956 0 0.034302 0.0389 0 0.97872 0.2864 0.080193 0.010935 4.7617 0.068236 8.2927e-005 0.82185 0.0057412 0.0064904 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.13572 0.96138 0.92293 0.0013953 0.99588 0.61762 0.00188 0.43195 1.9433 1.9428 15.9975 144.9938 0.00015444 -85.6661 0.94995
2.054 0.98804 5.5127e-005 3.8182 0.012022 2.6995e-005 0.0011548 0.19499 0.00065894 0.19564 0.17959 0 0.0343 0.0389 0 0.97882 0.28645 0.080208 0.010937 4.7624 0.068247 8.2941e-005 0.82184 0.0057418 0.0064911 0.001383 0.98699 0.99173 2.9817e-006 1.1926e-005 0.13573 0.96145 0.92296 0.0013953 0.99589 0.61775 0.0018799 0.43196 1.9436 1.9431 15.9975 144.9938 0.00015439 -85.6661 0.95095
2.055 0.98804 5.5127e-005 3.8182 0.012022 2.7008e-005 0.0011548 0.19502 0.00065894 0.19567 0.17962 0 0.034298 0.0389 0 0.97891 0.28649 0.080223 0.010939 4.7632 0.068258 8.2956e-005 0.82182 0.0057425 0.0064917 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13573 0.96152 0.92299 0.0013953 0.99589 0.61789 0.0018799 0.43197 1.9439 1.9434 15.9974 144.9939 0.00015435 -85.6662 0.95195
2.056 0.98804 5.5127e-005 3.8182 0.012022 2.7021e-005 0.0011548 0.19505 0.00065894 0.19571 0.17965 0 0.034297 0.0389 0 0.97901 0.28653 0.080238 0.010941 4.764 0.068269 8.297e-005 0.82181 0.0057431 0.0064924 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13574 0.96159 0.92302 0.0013953 0.9959 0.61802 0.0018799 0.43198 1.9442 1.9437 15.9974 144.9939 0.0001543 -85.6662 0.95295
2.057 0.98804 5.5127e-005 3.8182 0.012022 2.7034e-005 0.0011548 0.19508 0.00065895 0.19574 0.17968 0 0.034295 0.0389 0 0.9791 0.28657 0.080254 0.010942 4.7647 0.06828 8.2985e-005 0.8218 0.0057437 0.006493 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13574 0.96166 0.92305 0.0013953 0.99591 0.61815 0.0018799 0.43199 1.9445 1.944 15.9974 144.9939 0.00015425 -85.6662 0.95395
2.058 0.98804 5.5127e-005 3.8182 0.012022 2.7047e-005 0.0011548 0.19512 0.00065895 0.19577 0.17971 0 0.034293 0.0389 0 0.97919 0.28662 0.080269 0.010944 4.7655 0.068291 8.2999e-005 0.82179 0.0057443 0.0064937 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13575 0.96173 0.92308 0.0013953 0.99592 0.61828 0.0018799 0.43201 1.9448 1.9444 15.9973 144.9939 0.0001542 -85.6662 0.95495
2.059 0.98804 5.5127e-005 3.8182 0.012022 2.706e-005 0.0011548 0.19515 0.00065895 0.1958 0.17974 0 0.034291 0.0389 0 0.97929 0.28666 0.080284 0.010946 4.7662 0.068302 8.3014e-005 0.82178 0.005745 0.0064943 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13576 0.9618 0.92311 0.0013953 0.99593 0.61842 0.0018799 0.43202 1.9451 1.9447 15.9973 144.9939 0.00015415 -85.6663 0.95595
2.06 0.98804 5.5127e-005 3.8182 0.012022 2.7073e-005 0.0011548 0.19518 0.00065895 0.19584 0.17977 0 0.034289 0.0389 0 0.97938 0.2867 0.080299 0.010948 4.767 0.068313 8.3028e-005 0.82177 0.0057456 0.006495 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13576 0.96186 0.92314 0.0013953 0.99593 0.61855 0.0018799 0.43203 1.9454 1.945 15.9973 144.994 0.0001541 -85.6663 0.95695
2.061 0.98804 5.5126e-005 3.8182 0.012022 2.7086e-005 0.0011548 0.19521 0.00065895 0.19587 0.1798 0 0.034288 0.0389 0 0.97947 0.28674 0.080314 0.01095 4.7678 0.068324 8.3043e-005 0.82176 0.0057462 0.0064956 0.0013829 0.98699 0.99173 2.9816e-006 1.1926e-005 0.13577 0.96193 0.92317 0.0013953 0.99594 0.61868 0.0018799 0.43204 1.9457 1.9453 15.9972 144.994 0.00015405 -85.6663 0.95795
2.062 0.98804 5.5126e-005 3.8182 0.012022 2.7099e-005 0.0011548 0.19525 0.00065895 0.1959 0.17983 0 0.034286 0.0389 0 0.97957 0.28678 0.08033 0.010951 4.7685 0.068335 8.3058e-005 0.82175 0.0057468 0.0064963 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13577 0.962 0.9232 0.0013953 0.99595 0.61882 0.0018799 0.43205 1.946 1.9456 15.9972 144.994 0.00015401 -85.6663 0.95895
2.063 0.98804 5.5126e-005 3.8182 0.012022 2.7112e-005 0.0011548 0.19528 0.00065895 0.19593 0.17986 0 0.034284 0.0389 0 0.97966 0.28683 0.080345 0.010953 4.7693 0.068346 8.3072e-005 0.82174 0.0057475 0.0064969 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13578 0.96207 0.92323 0.0013953 0.99596 0.61895 0.0018799 0.43206 1.9463 1.9459 15.9972 144.994 0.00015396 -85.6664 0.95995
2.064 0.98804 5.5126e-005 3.8182 0.012022 2.7126e-005 0.0011548 0.19531 0.00065895 0.19597 0.17989 0 0.034282 0.0389 0 0.97976 0.28687 0.08036 0.010955 4.77 0.068357 8.3087e-005 0.82173 0.0057481 0.0064976 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13578 0.96213 0.92326 0.0013953 0.99597 0.61908 0.0018799 0.43207 1.9466 1.9462 15.9971 144.994 0.00015391 -85.6664 0.96095
2.065 0.98804 5.5126e-005 3.8182 0.012022 2.7139e-005 0.0011548 0.19534 0.00065895 0.196 0.17992 0 0.03428 0.0389 0 0.97985 0.28691 0.080375 0.010957 4.7708 0.068369 8.3101e-005 0.82171 0.0057487 0.0064982 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13579 0.9622 0.92329 0.0013953 0.99597 0.61921 0.0018799 0.43208 1.9469 1.9465 15.9971 144.9941 0.00015386 -85.6664 0.96195
2.066 0.98804 5.5126e-005 3.8182 0.012022 2.7152e-005 0.0011548 0.19537 0.00065895 0.19603 0.17995 0 0.034279 0.0389 0 0.97994 0.28695 0.08039 0.010958 4.7716 0.06838 8.3116e-005 0.8217 0.0057494 0.0064989 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13579 0.96227 0.92332 0.0013953 0.99598 0.61935 0.0018799 0.4321 1.9472 1.9468 15.9971 144.9941 0.00015382 -85.6664 0.96295
2.067 0.98804 5.5126e-005 3.8182 0.012022 2.7165e-005 0.0011548 0.19541 0.00065895 0.19606 0.17998 0 0.034277 0.0389 0 0.98004 0.287 0.080405 0.01096 4.7723 0.068391 8.313e-005 0.82169 0.00575 0.0064995 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.1358 0.96233 0.92335 0.0013953 0.99599 0.61948 0.0018799 0.43211 1.9475 1.9471 15.997 144.9941 0.00015377 -85.6665 0.96395
2.068 0.98804 5.5126e-005 3.8182 0.012022 2.7178e-005 0.0011548 0.19544 0.00065895 0.19609 0.18001 0 0.034275 0.0389 0 0.98013 0.28704 0.080421 0.010962 4.7731 0.068402 8.3145e-005 0.82168 0.0057506 0.0065002 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.1358 0.9624 0.92338 0.0013953 0.996 0.61961 0.0018799 0.43212 1.9478 1.9474 15.997 144.9941 0.00015372 -85.6665 0.96495
2.069 0.98804 5.5126e-005 3.8182 0.012022 2.7191e-005 0.0011548 0.19547 0.00065895 0.19613 0.18004 0 0.034273 0.0389 0 0.98022 0.28708 0.080436 0.010964 4.7739 0.068413 8.3159e-005 0.82167 0.0057512 0.0065008 0.0013829 0.98699 0.99173 2.9815e-006 1.1926e-005 0.13581 0.96247 0.92341 0.0013953 0.99601 0.61974 0.0018799 0.43213 1.9481 1.9477 15.997 144.9941 0.00015368 -85.6665 0.96595
2.07 0.98804 5.5126e-005 3.8182 0.012022 2.7204e-005 0.0011548 0.1955 0.00065895 0.19616 0.18007 0 0.034271 0.0389 0 0.98032 0.28712 0.080451 0.010965 4.7746 0.068424 8.3174e-005 0.82166 0.0057519 0.0065015 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13581 0.96253 0.92344 0.0013953 0.99601 0.61988 0.0018799 0.43214 1.9484 1.948 15.9969 144.9942 0.00015363 -85.6665 0.96695
2.071 0.98804 5.5126e-005 3.8182 0.012022 2.7217e-005 0.0011548 0.19554 0.00065895 0.19619 0.1801 0 0.03427 0.0389 0 0.98041 0.28717 0.080466 0.010967 4.7754 0.068435 8.3189e-005 0.82165 0.0057525 0.0065021 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13582 0.9626 0.92347 0.0013953 0.99602 0.62001 0.0018799 0.43215 1.9487 1.9483 15.9969 144.9942 0.00015358 -85.6666 0.96795
2.072 0.98804 5.5126e-005 3.8182 0.012022 2.723e-005 0.0011548 0.19557 0.00065895 0.19622 0.18014 0 0.034268 0.0389 0 0.98051 0.28721 0.080481 0.010969 4.7762 0.068446 8.3203e-005 0.82164 0.0057531 0.0065028 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13582 0.96266 0.9235 0.0013953 0.99603 0.62014 0.0018799 0.43216 1.949 1.9486 15.9969 144.9942 0.00015354 -85.6666 0.96895
2.073 0.98804 5.5126e-005 3.8182 0.012022 2.7243e-005 0.0011548 0.1956 0.00065895 0.19625 0.18017 0 0.034266 0.0389 0 0.9806 0.28725 0.080497 0.010971 4.7769 0.068457 8.3218e-005 0.82163 0.0057538 0.0065034 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13583 0.96273 0.92353 0.0013953 0.99604 0.62027 0.0018799 0.43217 1.9493 1.9489 15.9968 144.9942 0.00015349 -85.6666 0.96995
2.074 0.98804 5.5126e-005 3.8182 0.012022 2.7257e-005 0.0011548 0.19563 0.00065895 0.19629 0.1802 0 0.034264 0.0389 0 0.98069 0.28729 0.080512 0.010973 4.7777 0.068468 8.3232e-005 0.82162 0.0057544 0.0065041 0.0013829 0.98699 0.99173 2.9814e-006 1.1926e-005 0.13583 0.96279 0.92356 0.0013953 0.99604 0.6204 0.0018799 0.43218 1.9496 1.9492 15.9968 144.9943 0.00015344 -85.6666 0.97095
2.075 0.98804 5.5126e-005 3.8182 0.012022 2.727e-005 0.0011548 0.19566 0.00065895 0.19632 0.18023 0 0.034263 0.0389 0 0.98079 0.28734 0.080527 0.010974 4.7785 0.068479 8.3247e-005 0.8216 0.005755 0.0065047 0.0013829 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13584 0.96286 0.92359 0.0013953 0.99605 0.62054 0.0018799 0.4322 1.9499 1.9495 15.9968 144.9943 0.0001534 -85.6666 0.97195
2.076 0.98804 5.5125e-005 3.8182 0.012022 2.7283e-005 0.0011548 0.19569 0.00065895 0.19635 0.18026 0 0.034261 0.0389 0 0.98088 0.28738 0.080542 0.010976 4.7792 0.06849 8.3261e-005 0.82159 0.0057556 0.0065054 0.0013829 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13584 0.96292 0.92362 0.0013953 0.99606 0.62067 0.0018799 0.43221 1.9502 1.9498 15.9967 144.9943 0.00015335 -85.6667 0.97295
2.077 0.98804 5.5125e-005 3.8182 0.012022 2.7296e-005 0.0011548 0.19573 0.00065895 0.19638 0.18029 0 0.034259 0.0389 0 0.98098 0.28742 0.080557 0.010978 4.78 0.068501 8.3276e-005 0.82158 0.0057563 0.006506 0.0013829 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13585 0.96299 0.92365 0.0013953 0.99606 0.6208 0.0018799 0.43222 1.9505 1.9501 15.9967 144.9943 0.00015331 -85.6667 0.97395
2.078 0.98804 5.5125e-005 3.8182 0.012022 2.7309e-005 0.0011548 0.19576 0.00065895 0.19641 0.18032 0 0.034257 0.0389 0 0.98107 0.28746 0.080573 0.01098 4.7808 0.068512 8.329e-005 0.82157 0.0057569 0.0065067 0.0013829 0.98699 0.99173 2.9814e-006 1.1925e-005 0.13585 0.96305 0.92368 0.0013953 0.99607 0.62093 0.0018799 0.43223 1.9508 1.9504 15.9967 144.9943 0.00015326 -85.6667 0.97495
2.079 0.98804 5.5125e-005 3.8182 0.012022 2.7322e-005 0.0011548 0.19579 0.00065895 0.19644 0.18035 0 0.034255 0.0389 0 0.98116 0.28751 0.080588 0.010981 4.7815 0.068523 8.3305e-005 0.82156 0.0057575 0.0065074 0.0013829 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13586 0.96311 0.92371 0.0013953 0.99608 0.62106 0.0018799 0.43224 1.9511 1.9507 15.9966 144.9944 0.00015322 -85.6667 0.97595
2.08 0.98804 5.5125e-005 3.8182 0.012022 2.7335e-005 0.0011548 0.19582 0.00065895 0.19648 0.18038 0 0.034254 0.0389 0 0.98126 0.28755 0.080603 0.010983 4.7823 0.068534 8.332e-005 0.82155 0.0057582 0.006508 0.0013829 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13586 0.96318 0.92373 0.0013953 0.99609 0.6212 0.0018799 0.43225 1.9514 1.951 15.9966 144.9944 0.00015317 -85.6667 0.97695
2.081 0.98804 5.5125e-005 3.8182 0.012022 2.7348e-005 0.0011548 0.19585 0.00065895 0.19651 0.18041 0 0.034252 0.0389 0 0.98135 0.28759 0.080618 0.010985 4.7831 0.068546 8.3334e-005 0.82154 0.0057588 0.0065087 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13587 0.96324 0.92376 0.0013953 0.99609 0.62133 0.0018798 0.43226 1.9517 1.9513 15.9966 144.9944 0.00015313 -85.6668 0.97795
2.082 0.98804 5.5125e-005 3.8182 0.012022 2.7361e-005 0.0011548 0.19589 0.00065895 0.19654 0.18044 0 0.03425 0.0389 0 0.98145 0.28763 0.080634 0.010987 4.7839 0.068557 8.3349e-005 0.82153 0.0057594 0.0065093 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13587 0.96331 0.92379 0.0013953 0.9961 0.62146 0.0018798 0.43227 1.952 1.9516 15.9965 144.9944 0.00015308 -85.6668 0.97895
2.083 0.98804 5.5125e-005 3.8182 0.012022 2.7374e-005 0.0011548 0.19592 0.00065895 0.19657 0.18047 0 0.034248 0.0389 0 0.98154 0.28767 0.080649 0.010988 4.7846 0.068568 8.3363e-005 0.82152 0.00576 0.00651 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13588 0.96337 0.92382 0.0013953 0.99611 0.62159 0.0018798 0.43229 1.9523 1.9519 15.9965 144.9944 0.00015304 -85.6668 0.97995
2.084 0.98804 5.5125e-005 3.8182 0.012022 2.7387e-005 0.0011548 0.19595 0.00065896 0.1966 0.1805 0 0.034247 0.0389 0 0.98163 0.28772 0.080664 0.01099 4.7854 0.068579 8.3378e-005 0.8215 0.0057607 0.0065106 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13588 0.96343 0.92385 0.0013953 0.99611 0.62172 0.0018798 0.4323 1.9526 1.9521 15.9965 144.9945 0.00015299 -85.6668 0.98095
2.085 0.98804 5.5125e-005 3.8182 0.012022 2.7401e-005 0.0011548 0.19598 0.00065896 0.19663 0.18053 0 0.034245 0.0389 0 0.98173 0.28776 0.080679 0.010992 4.7862 0.06859 8.3392e-005 0.82149 0.0057613 0.0065113 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13589 0.96349 0.92388 0.0013953 0.99612 0.62185 0.0018798 0.43231 1.9529 1.9524 15.9964 144.9945 0.00015295 -85.6668 0.98195
2.086 0.98804 5.5125e-005 3.8182 0.012022 2.7414e-005 0.0011548 0.19601 0.00065896 0.19667 0.18056 0 0.034243 0.0389 0 0.98182 0.2878 0.080694 0.010994 4.7869 0.068601 8.3407e-005 0.82148 0.0057619 0.0065119 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13589 0.96356 0.9239 0.0013953 0.99613 0.62199 0.0018798 0.43232 1.9532 1.9527 15.9964 144.9945 0.0001529 -85.6669 0.98295
2.087 0.98804 5.5125e-005 3.8182 0.012022 2.7427e-005 0.0011548 0.19604 0.00065896 0.1967 0.18058 0 0.034241 0.0389 0 0.98192 0.28784 0.08071 0.010996 4.7877 0.068612 8.3422e-005 0.82147 0.0057626 0.0065126 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.1359 0.96362 0.92393 0.0013953 0.99613 0.62212 0.0018798 0.43233 1.9535 1.953 15.9963 144.9945 0.00015286 -85.6669 0.98395
2.088 0.98804 5.5125e-005 3.8182 0.012022 2.744e-005 0.0011548 0.19608 0.00065896 0.19673 0.18061 0 0.03424 0.0389 0 0.98201 0.28789 0.080725 0.010997 4.7885 0.068623 8.3436e-005 0.82146 0.0057632 0.0065132 0.0013828 0.98699 0.99173 2.9813e-006 1.1925e-005 0.13591 0.96368 0.92396 0.0013953 0.99614 0.62225 0.0018798 0.43234 1.9538 1.9533 15.9963 144.9945 0.00015281 -85.6669 0.98495
2.089 0.98804 5.5125e-005 3.8182 0.012022 2.7453e-005 0.0011548 0.19611 0.00065896 0.19676 0.18064 0 0.034238 0.0389 0 0.9821 0.28793 0.08074 0.010999 4.7893 0.068634 8.3451e-005 0.82145 0.0057638 0.0065139 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13591 0.96374 0.92399 0.0013953 0.99615 0.62238 0.0018798 0.43235 1.954 1.9536 15.9963 144.9946 0.00015277 -85.6669 0.98595
2.09 0.98804 5.5125e-005 3.8182 0.012022 2.7466e-005 0.0011548 0.19614 0.00065896 0.19679 0.18067 0 0.034236 0.0389 0 0.9822 0.28797 0.080755 0.011001 4.79 0.068645 8.3465e-005 0.82144 0.0057645 0.0065146 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13592 0.96381 0.92402 0.0013952 0.99615 0.62251 0.0018798 0.43236 1.9543 1.9539 15.9962 144.9946 0.00015273 -85.6669 0.98695
2.091 0.98804 5.5124e-005 3.8182 0.012022 2.7479e-005 0.0011548 0.19617 0.00065896 0.19682 0.1807 0 0.034234 0.0389 0 0.98229 0.28801 0.080771 0.011003 4.7908 0.068656 8.348e-005 0.82143 0.0057651 0.0065152 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13592 0.96387 0.92404 0.0013952 0.99616 0.62264 0.0018798 0.43237 1.9546 1.9542 15.9962 144.9946 0.00015268 -85.667 0.98795
2.092 0.98804 5.5124e-005 3.8182 0.012022 2.7492e-005 0.0011548 0.1962 0.00065896 0.19686 0.18073 0 0.034233 0.0389 0 0.98239 0.28806 0.080786 0.011004 4.7916 0.068667 8.3495e-005 0.82142 0.0057657 0.0065159 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13593 0.96393 0.92407 0.0013952 0.99617 0.62277 0.0018798 0.43239 1.9549 1.9545 15.9962 144.9946 0.00015264 -85.667 0.98895
2.093 0.98804 5.5124e-005 3.8182 0.012022 2.7505e-005 0.0011548 0.19623 0.00065896 0.19689 0.18076 0 0.034231 0.0389 0 0.98248 0.2881 0.080801 0.011006 4.7924 0.068678 8.3509e-005 0.82141 0.0057664 0.0065165 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13593 0.96399 0.9241 0.0013952 0.99617 0.62291 0.0018798 0.4324 1.9552 1.9548 15.9961 144.9946 0.0001526 -85.667 0.98995
2.094 0.98804 5.5124e-005 3.8182 0.012022 2.7518e-005 0.0011548 0.19626 0.00065896 0.19692 0.18079 0 0.034229 0.0389 0 0.98257 0.28814 0.080816 0.011008 4.7931 0.068689 8.3524e-005 0.82139 0.005767 0.0065172 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13594 0.96405 0.92413 0.0013952 0.99618 0.62304 0.0018798 0.43241 1.9555 1.9551 15.9961 144.9947 0.00015255 -85.667 0.99095
2.095 0.98804 5.5124e-005 3.8182 0.012022 2.7532e-005 0.0011548 0.1963 0.00065896 0.19695 0.18082 0 0.034227 0.0389 0 0.98267 0.28818 0.080832 0.01101 4.7939 0.0687 8.3538e-005 0.82138 0.0057676 0.0065178 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13594 0.96411 0.92415 0.0013952 0.99619 0.62317 0.0018798 0.43242 1.9558 1.9554 15.9961 144.9947 0.00015251 -85.667 0.99195
2.096 0.98804 5.5124e-005 3.8182 0.012022 2.7545e-005 0.0011548 0.19633 0.00065896 0.19698 0.18085 0 0.034226 0.0389 0 0.98276 0.28823 0.080847 0.011012 4.7947 0.068712 8.3553e-005 0.82137 0.0057683 0.0065185 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13595 0.96417 0.92418 0.0013952 0.99619 0.6233 0.0018798 0.43243 1.9561 1.9556 15.996 144.9947 0.00015247 -85.667 0.99295
2.097 0.98804 5.5124e-005 3.8182 0.012022 2.7558e-005 0.0011548 0.19636 0.00065896 0.19701 0.18088 0 0.034224 0.0389 0 0.98286 0.28827 0.080862 0.011013 4.7955 0.068723 8.3567e-005 0.82136 0.0057689 0.0065192 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13595 0.96423 0.92421 0.0013952 0.9962 0.62343 0.0018798 0.43244 1.9564 1.9559 15.996 144.9947 0.00015242 -85.6671 0.99395
2.098 0.98804 5.5124e-005 3.8182 0.012022 2.7571e-005 0.0011548 0.19639 0.00065896 0.19704 0.18091 0 0.034222 0.0389 0 0.98295 0.28831 0.080877 0.011015 4.7963 0.068734 8.3582e-005 0.82135 0.0057695 0.0065198 0.0013828 0.98699 0.99173 2.9812e-006 1.1925e-005 0.13596 0.96429 0.92424 0.0013952 0.99621 0.62356 0.0018798 0.43245 1.9566 1.9562 15.996 144.9947 0.00015238 -85.6671 0.99495
2.099 0.98804 5.5124e-005 3.8182 0.012022 2.7584e-005 0.0011548 0.19642 0.00065896 0.19708 0.18094 0 0.03422 0.0389 0 0.98304 0.28835 0.080892 0.011017 4.797 0.068745 8.3597e-005 0.82134 0.0057702 0.0065205 0.0013828 0.98699 0.99173 2.9811e-006 1.1924e-005 0.13596 0.96435 0.92426 0.0013952 0.99621 0.62369 0.0018798 0.43246 1.9569 1.9565 15.9959 144.9948 0.00015234 -85.6671 0.99595
2.1 0.98804 5.5124e-005 3.8182 0.012022 2.7597e-005 0.0011548 0.19645 0.00065896 0.19711 0.18097 0 0.034219 0.0389 0 0.98314 0.2884 0.080908 0.011019 4.7978 0.068756 8.3611e-005 0.82133 0.0057708 0.0065211 0.0013828 0.98699 0.99173 2.9812e-006 1.1924e-005 0.13597 0.96441 0.92429 0.0013952 0.99622 0.62382 0.0018798 0.43247 1.9572 1.9568 15.9959 144.9948 0.0001523 -85.6642 0.99695
2.101 0.98804 5.5124e-005 3.8182 0.012022 2.761e-005 0.0011548 0.19648 0.00065896 0.19714 0.181 0 0.034217 0.0389 0 0.98323 0.28844 0.080923 0.01102 4.7986 0.068767 8.3626e-005 0.82132 0.0057714 0.0065218 0.0064727 0.98324 0.991 1.4517e-005 5.3332e-005 0.13597 0.96442 0.92432 0.0027731 0.99621 0.62394 0.0023953 0.43243 1.9575 1.9571 15.9959 144.9948 0.00015226 -76.1614 0.99795
2.102 0.98804 5.5124e-005 3.8182 0.012022 2.7623e-005 0.0011548 0.19651 0.00065896 0.19717 0.18103 0 0.034215 0.0389 0 0.98333 0.28848 0.080938 0.011022 4.7994 0.068778 8.364e-005 0.82131 0.0057721 0.0065225 0.026218 0.97172 0.98767 6.5967e-005 0.00022946 0.13598 0.96421 0.92434 0.0053004 0.99616 0.62403 0.003336 0.43231 1.9578 1.9574 15.9958 144.9947 0.00015225 -67.1475 0.99895
2.103 0.98804 5.5124e-005 3.8182 0.012022 2.7636e-005 0.0011548 0.19655 0.00065896 0.1972 0.18106 0 0.034213 0.0389 0 0.98342 0.28852 0.080953 0.011024 4.8001 0.068789 8.3655e-005 0.82129 0.0057727 0.0065231 0.094864 0.94723 0.97733 0.00028436 0.00091302 0.13598 0.96345 0.92437 0.0092472 0.99589 0.62412 0.0044248 0.43215 1.9581 1.9577 15.9957 144.9947 0.00015226 -58.0161 0.99995
2.104 0.98804 5.5124e-005 3.8182 0.012022 2.7649e-005 0.0011548 0.19658 0.00065896 0.19723 0.18109 0 0.034212 0.0389 0 0.98352 0.28857 0.080969 0.011026 4.8009 0.0688 8.367e-005 0.82128 0.0057733 0.0065238 0.4879 0.85636 0.93875 0.0021782 0.0054736 0.13599 0.96143 0.92439 0.015752 0.99179 0.62413 0.0056237 0.43196 1.9584 1.9579 15.9965 144.9947 0.0001523 -37.2253 0.15622
2.105 0.98804 5.5124e-005 3.8182 0.012022 2.7662e-005 0.0011548 0.19661 0.00065896 0.19726 0.18112 0 0.03421 0.0389 0 0.98361 0.28861 0.080984 0.011027 4.8017 0.068811 8.3684e-005 0.82127 0.005774 0.0065244 0.99959 0.0021784 0.71215 0.93681 0.99582 0.13599 0.92788 0.92144 0.33227 0.96436 0.61042 0.044026 0.43175 1.9166 0.96054 16.0004 144.9944 0.00023298 23.9777 0.0019535
2.106 0.98804 5.5124e-005 3.8182 0.012022 2.7676e-005 0.0011548 0.19664 0.00065896 0.19729 0.18115 0 0.034208 0.0389 0 0.9837 0.28865 0.080999 0.011029 4.8025 0.068822 8.3699e-005 0.82126 0.0057746 0.0065251 0.99929 1.4442e-006 0.52836 0.99636 0.99924 0.136 0.8878 0.90357 0.59961 0.9372 0.59341 0.094467 0.43154 1.7331 0.58754 16 144.9931 0.00034163 18.0845 0.0029535
2.107 0.98804 5.5123e-005 3.8182 0.012022 2.7689e-005 0.0011548 0.19667 0.00065896 0.19732 0.18118 0 0.034206 0.0389 0 0.9838 0.28869 0.081015 0.011031 4.8033 0.068833 8.3713e-005 0.82125 0.0057752 0.0065257 0.99865 5.9553e-010 0.3925 0.9931 0.99797 0.136 0.85064 0.88049 0.71157 0.91081 0.57728 0.13104 0.43134 1.5574 0.56034 15.9996 144.9914 0.00040945 12.1529 0.0039535
2.108 0.98804 5.5123e-005 3.8182 0.012021 2.7702e-005 0.0011548 0.1967 0.00065896 0.19736 0.18121 0 0.034205 0.0389 0 0.98389 0.28874 0.08103 0.011033 4.8041 0.068844 8.3728e-005 0.82124 0.0057759 0.0065264 0.99791 -8.6359e-011 0.29206 0.98653 0.99592 0.13601 0.81704 0.85502 0.75852 0.88516 0.56231 0.15879 0.43113 1.4106 0.59654 15.9993 144.9898 0.00045965 8.1973 0.0049535
2.109 0.98804 5.5123e-005 3.8182 0.012021 2.7715e-005 0.0011548 0.19673 0.00065896 0.19739 0.18124 0 0.034203 0.0389 0 0.98399 0.28878 0.081045 0.011035 4.8048 0.068856 8.3743e-005 0.82123 0.0057765 0.0065271 0.9972 7.5257e-011 0.21769 0.97827 0.99341 0.13601 0.78668 0.82854 0.77654 0.86025 0.54855 0.18142 0.43093 1.2937 0.65289 15.999 144.9881 0.00049789 5.5539 0.0059535
2.11 0.98804 5.5123e-005 3.8182 0.012021 2.7728e-005 0.0011548 0.19676 0.00065896 0.19742 0.18126 0 0.034201 0.0389 0 0.98408 0.28882 0.08106 0.011036 4.8056 0.068867 8.3757e-005 0.82122 0.0057771 0.0065277 0.99651 1.3531e-011 0.1625 0.96889 0.99057 0.13602 0.75904 0.80194 0.77997 0.83604 0.53588 0.20068 0.43072 1.2038 0.71406 15.9987 144.9866 0.00052692 3.5536 0.0069535
2.111 0.98804 5.5123e-005 3.8182 0.012021 2.7741e-005 0.0011548 0.19679 0.00065896 0.19745 0.18129 0 0.0342 0.0389 0 0.98418 0.28886 0.081076 0.011038 4.8064 0.068878 8.3772e-005 0.82121 0.0057778 0.0065284 0.99578 9.8485e-011 0.12148 0.95837 0.98734 0.13603 0.73376 0.77587 0.77515 0.81251 0.52424 0.21741 0.43052 1.1369 0.77225 15.9984 144.9851 0.00054882 1.8517 0.0079535
2.112 0.98804 5.5123e-005 3.8182 0.012021 2.7754e-005 0.0011548 0.19683 0.00065896 0.19748 0.18132 0 0.034198 0.0389 0 0.98427 0.28891 0.081091 0.01104 4.8072 0.068889 8.3786e-005 0.82119 0.0057784 0.0065291 0.99498 4.9308e-011 0.090953 0.94643 0.98356 0.13603 0.71059 0.75077 0.76516 0.78966 0.51358 0.23205 0.43031 1.0885 0.82331 15.9981 144.9837 0.00056532 0.27796 0.0089535
2.113 0.98804 5.5123e-005 3.8182 0.012021 2.7767e-005 0.0011548 0.19686 0.00065897 0.19751 0.18135 0 0.034196 0.0389 0 0.98436 0.28895 0.081106 0.011042 4.808 0.0689 8.3801e-005 0.82118 0.005779 0.0065297 0.99405 3.6151e-011 0.068216 0.93257 0.979 0.13604 0.68939 0.72699 0.75157 0.76746 0.50387 0.24487 0.43011 1.0546 0.8655 15.9978 144.9824 0.00057784 -1.2648 0.0099535
2.114 0.98804 5.5123e-005 3.8182 0.012021 2.778e-005 0.0011548 0.19689 0.00065897 0.19754 0.18138 0 0.034194 0.0389 0 0.98446 0.28899 0.081121 0.011043 4.8088 0.068911 8.3816e-005 0.82117 0.0057797 0.0065304 0.99291 -1.5658e-010 0.051264 0.9161 0.97333 0.13604 0.67008 0.70476 0.73516 0.7459 0.49513 0.25602 0.4299 1.0317 0.89881 15.9976 144.9812 0.00058748 -2.8465 0.010953
2.115 0.98804 5.5123e-005 3.8182 0.012021 2.7793e-005 0.0011548 0.19692 0.00065897 0.19757 0.18141 0 0.034193 0.0389 0 0.98455 0.28904 0.081137 0.011045 4.8095 0.068922 8.383e-005 0.82116 0.0057803 0.006531 0.99146 1.6827e-011 0.038617 0.8961 0.96606 0.13605 0.6526 0.68429 0.71624 0.72495 0.48736 0.2656 0.4297 1.0167 0.92423 15.9973 144.98 0.00059501 -4.5324 0.011953
2.116 0.98804 5.5123e-005 3.8182 0.012021 2.7807e-005 0.0011548 0.19695 0.00065897 0.1976 0.18144 0 0.034191 0.0389 0 0.98465 0.28908 0.081152 0.011047 4.8103 0.068933 8.3845e-005 0.82115 0.0057809 0.0065317 0.9895 1.9148e-010 0.029178 0.87121 0.9565 0.13605 0.63695 0.66579 0.69481 0.70462 0.48059 0.27364 0.4295 1.0074 0.94322 15.9971 144.979 0.00060096 -6.3975 0.012953
2.117 0.98804 5.5123e-005 3.8182 0.012021 2.782e-005 0.0011548 0.19698 0.00065897 0.19763 0.18147 0 0.034189 0.0389 0 0.98474 0.28912 0.081167 0.011049 4.8111 0.068944 8.386e-005 0.82114 0.0057816 0.0065324 0.98667 3.2637e-010 0.022134 0.83949 0.94336 0.13606 0.62317 0.64946 0.67064 0.68489 0.47487 0.28016 0.42929 1.0019 0.95725 15.9968 144.978 0.00060566 -8.5402 0.013953
2.118 0.98804 5.5123e-005 3.8182 0.012021 2.7833e-005 0.0011548 0.19701 0.00065897 0.19766 0.1815 0 0.034188 0.0389 0 0.98484 0.28916 0.081182 0.011051 4.8119 0.068955 8.3874e-005 0.82113 0.0057822 0.006533 0.98229 -8.4587e-011 0.016886 0.79795 0.92476 0.13606 0.61133 0.63552 0.64333 0.66576 0.47023 0.28515 0.42909 0.99918 0.96764 15.9966 144.9771 0.00060928 -11.0969 0.014953
2.119 0.98804 5.5123e-005 3.8182 0.012021 2.7846e-005 0.0011548 0.19704 0.00065897 0.1977 0.18153 0 0.034186 0.0389 0 0.98493 0.28921 0.081198 0.011052 4.8127 0.068966 8.3889e-005 0.82112 0.0057829 0.0065337 0.97483 5.7113e-011 0.012992 0.74212 0.89733 0.13607 0.60151 0.6242 0.61241 0.64725 0.46669 0.28857 0.42888 0.99823 0.97544 15.9964 144.9763 0.00061186 -14.2551 0.015953
2.12 0.98804 5.5123e-005 3.8182 0.012021 2.7859e-005 0.0011548 0.19707 0.00065897 0.19773 0.18156 0 0.034184 0.0389 0 0.98502 0.28925 0.081213 0.011054 4.8135 0.068978 8.3903e-005 0.82111 0.0057835 0.0065343 0.96075 -2.6464e-011 0.010132 0.66548 0.85543 0.13607 0.59378 0.61572 0.57754 0.62943 0.46421 0.29042 0.42868 0.99846 0.9815 15.9962 144.9756 0.00061336 -18.2453 0.016953
2.121 0.98804 5.5123e-005 3.8182 0.012021 2.7872e-005 0.0011548 0.1971 0.00065897 0.19776 0.18159 0 0.034182 0.0389 0 0.98512 0.28929 0.081228 0.011056 4.8143 0.068989 8.3918e-005 0.8211 0.0057841 0.006535 0.93163 1.0102e-011 0.0080766 0.5599 0.78998 0.13608 0.58804 0.61007 0.53873 0.61249 0.46265 0.2908 0.42848 0.9995 0.98657 15.996 144.9751 0.00061367 -23.2489 0.017953
2.122 0.98804 5.5122e-005 3.8182 0.012021 2.7885e-005 0.0011548 0.19713 0.00065897 0.19779 0.18161 0 0.034181 0.0389 0 0.98521 0.28933 0.081244 0.011058 4.8151 0.069 8.3933e-005 0.82108 0.0057848 0.0065357 0.86989 3.42e-012 0.0066626 0.4206 0.68896 0.13608 0.58398 0.60688 0.49597 0.59696 0.46178 0.28992 0.42827 1.0011 0.99079 15.9959 144.9746 0.00061293 -29.1348 0.018953
2.123 0.98804 5.5122e-005 3.8182 0.012021 2.7898e-005 0.0011548 0.19716 0.00065897 0.19782 0.18164 0 0.034179 0.0389 0 0.98531 0.28938 0.081259 0.011059 4.8158 0.069011 8.3947e-005 0.82107 0.0057854 0.0065363 0.7555 4.7756e-013 0.0057426 0.26115 0.5455 0.13609 0.5811 0.60524 0.44773 0.58412 0.46135 0.28793 0.42807 1.003 0.99429 15.9957 144.9742 0.0006115 -35.1909 0.019953
2.124 0.98804 5.5122e-005 3.8182 0.012021 2.7911e-005 0.0011548 0.19719 0.00065897 0.19785 0.18167 0 0.034177 0.0389 0 0.9854 0.28942 0.081274 0.011061 4.8166 0.069022 8.3962e-005 0.82106 0.005786 0.006537 0.59916 4.0976e-005 0.0051701 0.12319 0.37518 0.13609 0.57897 0.60429 0.39094 0.57581 0.46118 0.28471 0.42787 1.0051 0.99734 15.9956 144.9739 0.00060979 -40.5544 0.020953
2.125 0.98804 5.5122e-005 3.8182 0.012021 2.7924e-005 0.0011548 0.19723 0.00065897 0.19788 0.1817 0 0.034176 0.0389 0 0.9855 0.28946 0.081289 0.011063 4.8174 0.069033 8.3976e-005 0.82105 0.0057867 0.0065377 0.44496 0.00056688 0.0050027 0.042027 0.21696 0.1361 0.57737 0.60389 0.32472 0.57238 0.46115 0.27994 0.42767 1.0074 1.0001 15.9956 144.9737 0.00060801 -44.9429 0.021953
2.126 0.98804 5.5122e-005 3.8182 0.012021 2.7937e-005 0.0011548 0.19726 0.00065897 0.19791 0.18173 0 0.034174 0.0389 0 0.98559 0.2895 0.081305 0.011065 4.8182 0.069044 8.3991e-005 0.82104 0.0057873 0.0065383 0.32443 0.0014858 0.0052281 0.010841 0.10416 0.1361 0.57619 0.6043 0.25316 0.57204 0.46119 0.27333 0.42748 1.0097 1.0028 15.9955 144.9735 0.00060618 -48.4479 0.022953
2.127 0.98804 5.5122e-005 3.8182 0.012021 2.7951e-005 0.0011548 0.19729 0.00065897 0.19794 0.18176 0 0.034172 0.0389 0 0.98568 0.28955 0.08132 0.011066 4.819 0.069055 8.4006e-005 0.82103 0.005788 0.006539 0.24137 0.0029394 0.005844 0.0028101 0.04224 0.13611 0.57535 0.60551 0.18421 0.57296 0.46127 0.26473 0.42729 1.012 1.0053 15.9955 144.9734 0.00060432 -51.2191 0.023953
2.128 0.98804 5.5122e-005 3.8182 0.012021 2.7964e-005 0.0011548 0.19732 0.00065897 0.19797 0.18179 0 0.034171 0.0389 0 0.98578 0.28959 0.081335 0.011068 4.8198 0.069066 8.402e-005 0.82102 0.0057886 0.0065397 0.18629 0.0050224 0.0068386 0.0011675 0.015508 0.13611 0.5748 0.6072 0.12568 0.57427 0.46138 0.25424 0.4271 1.0144 1.0078 15.9954 144.9733 0.00060244 -53.4168 0.024953
2.129 0.98804 5.5122e-005 3.8182 0.012021 2.7977e-005 0.0011548 0.19735 0.00065897 0.198 0.18182 0 0.034169 0.0389 0 0.98587 0.28963 0.081351 0.01107 4.8206 0.069077 8.4035e-005 0.82101 0.0057892 0.0065403 0.14902 0.0077924 0.0081946 0.00074042 0.0060142 0.13612 0.57448 0.60909 0.081676 0.57567 0.46149 0.24211 0.42691 1.0167 1.0103 15.9954 144.9732 0.00060055 -55.1992 0.025953
2.13 0.98804 5.5122e-005 3.8182 0.012021 2.799e-005 0.0011548 0.19738 0.00065897 0.19803 0.18185 0 0.034167 0.0389 0 0.98597 0.28967 0.081366 0.011072 4.8214 0.069088 8.405e-005 0.821 0.0057899 0.006541 0.1225 0.01129 0.0098968 0.000545 0.0029772 0.13612 0.57434 0.61104 0.051951 0.57704 0.46161 0.22864 0.42673 1.0191 1.0127 15.9954 144.9732 0.00059865 -56.7026 0.026953
2.131 0.98804 5.5122e-005 3.8182 0.012021 2.8003e-005 0.0011548 0.19741 0.00065897 0.19806 0.18187 0 0.034165 0.0389 0 0.98606 0.28972 0.081381 0.011074 4.8222 0.0691 8.4064e-005 0.82098 0.0057905 0.0065416 0.10252 0.015562 0.01194 0.00042289 0.0019322 0.13613 0.57435 0.61299 0.033591 0.57836 0.46174 0.21412 0.42655 1.0215 1.0151 15.9954 144.9731 0.00059673 -58.03 0.027953
2.132 0.98804 5.5122e-005 3.8182 0.012021 2.8016e-005 0.0011548 0.19744 0.00065897 0.19809 0.1819 0 0.034164 0.0389 0 0.98616 0.28976 0.081397 0.011075 4.823 0.069111 8.4079e-005 0.82097 0.0057912 0.0065423 0.086703 0.020676 0.014328 0.00033732 0.0014522 0.13614 0.5745 0.61493 0.022997 0.57963 0.46186 0.19882 0.42638 1.0239 1.0175 15.9954 144.9731 0.00059481 -59.2503 0.028953
2.133 0.98804 5.5122e-005 3.8182 0.012021 2.8029e-005 0.0011548 0.19747 0.00065897 0.19812 0.18193 0 0.034162 0.0389 0 0.98625 0.2898 0.081412 0.011077 4.8238 0.069122 8.4094e-005 0.82096 0.0057918 0.006543 0.073759 0.026724 0.017079 0.00027275 0.0011527 0.13614 0.57476 0.61686 0.017106 0.58085 0.46199 0.18295 0.42621 1.0263 1.0199 15.9954 144.9731 0.00059289 -60.4049 0.029953
2.134 0.98804 5.5122e-005 3.8182 0.012021 2.8042e-005 0.0011548 0.1975 0.00065897 0.19815 0.18196 0 0.03416 0.0389 0 0.98635 0.28985 0.081427 0.011079 4.8246 0.069133 8.4108e-005 0.82095 0.0057924 0.0065436 0.062954 0.033824 0.020216 0.00022287 0.00093328 0.13615 0.57513 0.61877 0.013793 0.58202 0.46212 0.16676 0.42604 1.0287 1.0223 15.9954 144.9731 0.00059097 -61.5166 0.030953
2.135 0.98804 5.5122e-005 3.8182 0.012021 2.8055e-005 0.0011548 0.19753 0.00065897 0.19818 0.18199 0 0.034159 0.0389 0 0.98644 0.28989 0.081442 0.011081 4.8253 0.069144 8.4123e-005 0.82094 0.0057931 0.0065443 0.053846 0.042113 0.02377 0.00018327 0.00076299 0.13615 0.57559 0.62067 0.011785 0.58314 0.46225 0.15045 0.42587 1.031 1.0247 15.9954 144.973 0.00058904 -62.597 0.031953
2.136 0.98804 5.5122e-005 3.8182 0.012021 2.8068e-005 0.0011548 0.19756 0.00065897 0.19821 0.18202 0 0.034157 0.0389 0 0.98653 0.28993 0.081458 0.011082 4.8261 0.069155 8.4137e-005 0.82093 0.0057937 0.006545 0.046133 0.051743 0.027773 0.00015149 0.0006279 0.13616 0.57614 0.62255 0.010412 0.58423 0.46239 0.13425 0.42571 1.0334 1.0271 15.9954 144.973 0.0005871 -63.6514 0.032953
2.137 0.98804 5.5121e-005 3.8182 0.012021 2.8081e-005 0.0011548 0.19759 0.00065897 0.19825 0.18205 0 0.034155 0.0389 0 0.98663 0.28997 0.081473 0.011084 4.8269 0.069166 8.4152e-005 0.82092 0.0057943 0.0065456 0.039588 0.062879 0.032266 0.00012583 0.00051952 0.13616 0.57677 0.62441 0.0093556 0.58529 0.46252 0.1184 0.42555 1.0358 1.0295 15.9954 144.973 0.00058517 -64.6822 0.033953
2.138 0.98804 5.5121e-005 3.8182 0.012021 2.8095e-005 0.0011548 0.19762 0.00065897 0.19828 0.18207 0 0.034154 0.0389 0 0.98672 0.29002 0.081488 0.011086 4.8277 0.069177 8.4167e-005 0.82091 0.005795 0.0065463 0.034032 0.075692 0.037291 0.00010496 0.00043196 0.13617 0.57747 0.62625 0.0084772 0.58632 0.46265 0.10313 0.4254 1.0381 1.0319 15.9955 144.9729 0.00058323 -65.6905 0.034953
2.139 0.98804 5.5121e-005 3.8182 0.012021 2.8108e-005 0.0011548 0.19765 0.00065897 0.19831 0.1821 0 0.034152 0.0389 0 0.98682 0.29006 0.081504 0.011088 4.8285 0.069188 8.4181e-005 0.8209 0.0057956 0.006547 0.029312 0.090356 0.042893 8.7934e-005 0.00036085 0.13617 0.57823 0.62808 0.007718 0.58733 0.46278 0.088657 0.42525 1.0405 1.0343 15.9955 144.9729 0.0005813 -66.6764 0.035953
2.14 0.98804 5.5121e-005 3.8182 0.012021 2.8121e-005 0.0011548 0.19768 0.00065897 0.19834 0.18213 0 0.03415 0.0389 0 0.98691 0.2901 0.081519 0.01109 4.8293 0.069199 8.4196e-005 0.82088 0.0057963 0.0065476 0.025301 0.10704 0.049125 7.3981e-005 0.00030282 0.13618 0.57905 0.6299 0.0070508 0.58833 0.46292 0.075179 0.4251 1.0429 1.0367 15.9955 144.9729 0.00057936 -67.6398 0.036953
2.141 0.98804 5.5121e-005 3.8182 0.012021 2.8134e-005 0.0011548 0.19771 0.00065897 0.19837 0.18216 0 0.034149 0.0389 0 0.98701 0.29014 0.081534 0.011091 4.8301 0.06921 8.4211e-005 0.82087 0.0057969 0.0065483 0.021892 0.12592 0.056044 6.2514e-005 0.00025531 0.13618 0.57991 0.63169 0.0064607 0.58932 0.46305 0.062862 0.42496 1.0452 1.0391 15.9956 144.9729 0.00057742 -68.5801 0.037953
2.142 0.98804 5.5121e-005 3.8182 0.012021 2.8147e-005 0.0011548 0.19774 0.00065897 0.1984 0.18219 0 0.034147 0.0389 0 0.9871 0.29019 0.08155 0.011093 4.8309 0.069222 8.4225e-005 0.82086 0.0057975 0.006549 0.018993 0.14712 0.063712 5.3057e-005 0.00021625 0.13619 0.58082 0.63347 0.0059364 0.59031 0.46319 0.051829 0.42483 1.0476 1.0415 15.9956 144.9728 0.00057548 -69.4964 0.038953
2.143 0.98804 5.5121e-005 3.8182 0.012021 2.816e-005 0.0011548 0.19777 0.00065898 0.19843 0.18222 0 0.034145 0.0389 0 0.9872 0.29023 0.081565 0.011095 4.8317 0.069233 8.424e-005 0.82085 0.0057982 0.0065496 0.016527 0.17076 0.072199 4.5239e-005 0.00018405 0.13619 0.58177 0.63524 0.0054697 0.5913 0.46333 0.042151 0.4247 1.05 1.0438 15.9957 144.9728 0.00057354 -70.3879 0.039953
2.144 0.98804 5.5121e-005 3.8182 0.012021 2.8173e-005 0.0011548 0.1978 0.00065898 0.19846 0.18225 0 0.034144 0.0389 0 0.98729 0.29027 0.08158 0.011097 4.8325 0.069244 8.4255e-005 0.82084 0.0057988 0.0065503 0.01443 0.19692 0.081582 3.8758e-005 0.00015742 0.1362 0.58274 0.63698 0.0050538 0.5923 0.46346 0.033847 0.42458 1.0523 1.0462 15.9957 144.9728 0.0005716 -71.253 0.040953
2.145 0.98804 5.5121e-005 3.8182 0.012021 2.8186e-005 0.0011548 0.19783 0.00065898 0.19849 0.18227 0 0.034142 0.0389 0 0.98739 0.29032 0.081596 0.011098 4.8333 0.069255 8.4269e-005 0.82083 0.0057995 0.006551 0.012644 0.22563 0.09194 3.3374e-005 0.00013535 0.1362 0.58375 0.63871 0.0046828 0.59332 0.4636 0.026883 0.42446 1.0547 1.0486 15.9958 144.9727 0.00056966 -72.0905 0.041953
2.146 0.98804 5.5121e-005 3.8182 0.012021 2.8199e-005 0.0011548 0.19786 0.00065898 0.19852 0.1823 0 0.03414 0.0389 0 0.98748 0.29036 0.081611 0.0111 4.8341 0.069266 8.4284e-005 0.82082 0.0058001 0.0065516 0.011124 0.25683 0.10336 2.889e-005 0.00011701 0.13621 0.58479 0.64043 0.0043516 0.59435 0.46374 0.021181 0.42435 1.057 1.0509 15.9958 144.9727 0.00056773 -72.8987 0.042953
2.147 0.98804 5.5121e-005 3.8182 0.012021 2.8212e-005 0.0011549 0.19789 0.00065898 0.19855 0.18233 0 0.034139 0.0389 0 0.98757 0.2904 0.081626 0.011102 4.8349 0.069277 8.4298e-005 0.82081 0.0058008 0.0065523 0.0098298 0.29042 0.11591 2.5148e-005 0.00010173 0.13621 0.58584 0.64213 0.004056 0.5954 0.46388 0.016621 0.42424 1.0594 1.0533 15.9959 144.9727 0.00056579 -73.6761 0.043953
2.148 0.98804 5.5121e-005 3.8182 0.012021 2.8226e-005 0.0011549 0.19792 0.00065898 0.19858 0.18236 0 0.034137 0.0389 0 0.98767 0.29044 0.081642 0.011104 4.8357 0.069288 8.4313e-005 0.8208 0.0058014 0.006553 0.0087265 0.32621 0.12967 2.2019e-005 8.8973e-005 0.13622 0.58692 0.64382 0.0037922 0.59648 0.46402 0.01306 0.42414 1.0617 1.0557 15.996 144.9727 0.00056386 -74.4212 0.044953
2.149 0.98804 5.5121e-005 3.8182 0.012021 2.8239e-005 0.0011549 0.19795 0.00065898 0.19861 0.18239 0 0.034135 0.0389 0 0.98776 0.29049 0.081657 0.011106 4.8365 0.069299 8.4328e-005 0.82079 0.005802 0.0065536 0.0077855 0.36391 0.14469 1.9396e-005 7.8294e-005 0.13622 0.58801 0.64549 0.0035568 0.59759 0.46417 0.010342 0.42405 1.064 1.058 15.996 144.9726 0.00056193 -75.1327 0.045953
2.15 0.98804 5.5121e-005 3.8182 0.012021 2.8252e-005 0.0011549 0.19798 0.00065898 0.19864 0.18242 0 0.034134 0.0389 0 0.98786 0.29053 0.081672 0.011107 4.8373 0.06931 8.4342e-005 0.82077 0.0058027 0.0065543 0.0069825 0.40318 0.16101 1.7192e-005 6.9334e-005 0.13623 0.58911 0.64714 0.0033469 0.59873 0.46431 0.0083095 0.42396 1.0664 1.0604 15.9961 144.9726 0.00056 -75.8092 0.046953
2.151 0.98804 5.5121e-005 3.8182 0.012021 2.8265e-005 0.0011549 0.19801 0.00065898 0.19867 0.18245 0 0.034132 0.0389 0 0.98795 0.29057 0.081687 0.011109 4.8381 0.069322 8.4357e-005 0.82076 0.0058033 0.006555 0.0062962 0.44357 0.17863 1.5337e-005 6.1802e-005 0.13624 0.59022 0.64878 0.0031599 0.59991 0.46446 0.0068178 0.42387 1.0687 1.0627 15.9962 144.9726 0.00055808 -76.4501 0.047953
2.152 0.98804 5.512e-005 3.8182 0.012021 2.8278e-005 0.0011549 0.19804 0.00065898 0.1987 0.18247 0 0.03413 0.0389 0 0.98805 0.29061 0.081703 0.011111 4.8389 0.069333 8.4372e-005 0.82075 0.005804 0.0065556 0.0057095 0.48462 0.19751 1.3771e-005 5.5449e-005 0.13624 0.59135 0.65041 0.0029932 0.60112 0.46461 0.0057376 0.4238 1.071 1.0651 15.9962 144.9726 0.00055616 -77.0546 0.048953
2.153 0.98804 5.512e-005 3.8182 0.012021 2.8291e-005 0.0011549 0.19807 0.00065898 0.19873 0.1825 0 0.034129 0.0389 0 0.98814 0.29066 0.081718 0.011113 4.8397 0.069344 8.4386e-005 0.82074 0.0058046 0.0065563 0.0052069 0.52579 0.21759 1.2446e-005 5.008e-005 0.13625 0.59248 0.65202 0.0028449 0.60238 0.46476 0.0049611 0.42372 1.0734 1.0674 15.9963 144.9725 0.00055424 -77.6225 0.049953
2.154 0.98804 5.512e-005 3.8182 0.012021 2.8304e-005 0.0011549 0.1981 0.00065898 0.19876 0.18253 0 0.034127 0.0389 0 0.98824 0.2907 0.081733 0.011114 4.8405 0.069355 8.4401e-005 0.82073 0.0058053 0.006557 0.0047758 0.56657 0.23877 1.1323e-005 4.5531e-005 0.13625 0.59361 0.65362 0.0027129 0.60367 0.46491 0.0044026 0.42366 1.0757 1.0698 15.9964 144.9725 0.00055233 -78.1539 0.050953
2.155 0.98804 5.512e-005 3.8182 0.012021 2.8317e-005 0.0011549 0.19813 0.00065898 0.19879 0.18256 0 0.034125 0.0389 0 0.98833 0.29074 0.081749 0.011116 4.8413 0.069366 8.4416e-005 0.82072 0.0058059 0.0065577 0.0044055 0.60643 0.26091 1.0366e-005 4.1663e-005 0.13626 0.59476 0.6552 0.0025955 0.605 0.46506 0.0039971 0.42359 1.078 1.0721 15.9965 144.9725 0.00055043 -78.6493 0.051953
2.156 0.98804 5.512e-005 3.8182 0.012021 2.833e-005 0.0011549 0.19816 0.00065898 0.19882 0.18259 0 0.034124 0.0389 0 0.98843 0.29079 0.081764 0.011118 4.8421 0.069377 8.443e-005 0.82071 0.0058065 0.0065583 0.0040866 0.64489 0.28387 9.5514e-006 3.8367e-005 0.13626 0.5959 0.65677 0.0024911 0.60638 0.46521 0.0036973 0.42354 1.0803 1.0745 15.9966 144.9725 0.00054853 -79.1095 0.052953
2.157 0.98804 5.512e-005 3.8182 0.012021 2.8343e-005 0.0011549 0.19819 0.00065898 0.19885 0.18261 0 0.034122 0.0389 0 0.98852 0.29083 0.081779 0.01112 4.8429 0.069388 8.4445e-005 0.8207 0.0058072 0.006559 0.0038115 0.68154 0.30748 8.8542e-006 3.5551e-005 0.13627 0.59705 0.65833 0.0023984 0.60779 0.46537 0.00347 0.42348 1.0827 1.0768 15.9967 144.9725 0.00054663 -79.5355 0.053953
2.158 0.98804 5.512e-005 3.8182 0.012021 2.8356e-005 0.0011549 0.19822 0.00065898 0.19888 0.18264 0 0.03412 0.0389 0 0.98862 0.29087 0.081795 0.011122 4.8437 0.069399 8.446e-005 0.82069 0.0058078 0.0065597 0.0035741 0.71603 0.33156 8.2557e-006 3.3136e-005 0.13627 0.59821 0.65987 0.0023159 0.60924 0.46553 0.0032923 0.42343 1.085 1.0791 15.9967 144.9724 0.00054475 -79.9285 0.054953
2.159 0.98804 5.512e-005 3.8182 0.012021 2.837e-005 0.0011549 0.19825 0.00065898 0.19891 0.18267 0 0.034119 0.0389 0 0.98871 0.29091 0.08181 0.011123 4.8445 0.06941 8.4474e-005 0.82067 0.0058085 0.0065603 0.0033682 0.74811 0.35595 7.7415e-006 3.1059e-005 0.13628 0.59936 0.6614 0.0022425 0.61074 0.46568 0.0031494 0.42339 1.0873 1.0815 15.9968 144.9724 0.00054287 -80.2902 0.055953
2.16 0.98804 5.512e-005 3.8182 0.012021 2.8383e-005 0.0011549 0.19828 0.00065898 0.19894 0.1827 0 0.034117 0.0389 0 0.9888 0.29096 0.081826 0.011125 4.8453 0.069421 8.4489e-005 0.82066 0.0058091 0.006561 0.0031894 0.7776 0.38048 7.2979e-006 2.927e-005 0.13628 0.60051 0.66292 0.0021773 0.61226 0.46584 0.0030313 0.42335 1.0896 1.0838 15.9969 144.9724 0.000541 -80.622 0.056953
2.161 0.98804 5.512e-005 3.8182 0.012021 2.8396e-005 0.0011549 0.19831 0.00065898 0.19897 0.18273 0 0.034115 0.0389 0 0.9889 0.291 0.081841 0.011127 4.8462 0.069433 8.4504e-005 0.82065 0.0058098 0.0065617 0.003034 0.80441 0.40499 6.9141e-006 2.7722e-005 0.13629 0.60167 0.66442 0.0021193 0.61383 0.466 0.0029317 0.42331 1.0919 1.0861 15.997 144.9724 0.00053913 -80.9258 0.057953
2.162 0.98804 5.512e-005 3.8182 0.012021 2.8409e-005 0.0011549 0.19834 0.00065898 0.199 0.18276 0 0.034114 0.0389 0 0.98899 0.29104 0.081856 0.011129 4.847 0.069444 8.4518e-005 0.82064 0.0058104 0.0065623 0.0028985 0.82853 0.42935 6.5808e-006 2.638e-005 0.13629 0.60282 0.66591 0.0020677 0.61542 0.46617 0.0028463 0.42327 1.0942 1.0884 15.9971 144.9724 0.00053727 -81.2033 0.058953
2.163 0.98804 5.512e-005 3.8182 0.012021 2.8422e-005 0.0011549 0.19837 0.00065898 0.19903 0.18278 0 0.034112 0.0389 0 0.98909 0.29109 0.081872 0.01113 4.8478 0.069455 8.4533e-005 0.82063 0.005811 0.006563 0.0027801 0.85004 0.45343 6.2912e-006 2.5214e-005 0.1363 0.60397 0.66739 0.0020218 0.61705 0.46633 0.0027723 0.42324 1.0965 1.0907 15.9972 144.9724 0.00053542 -81.4564 0.059953
2.164 0.98804 5.512e-005 3.8182 0.012021 2.8435e-005 0.0011549 0.1984 0.00065898 0.19906 0.18281 0 0.034111 0.0389 0 0.98918 0.29113 0.081887 0.011132 4.8486 0.069466 8.4548e-005 0.82062 0.0058117 0.0065637 0.0026766 0.86903 0.47712 6.0393e-006 2.4197e-005 0.1363 0.60513 0.66886 0.0019808 0.6187 0.46649 0.0027077 0.42321 1.0988 1.093 15.9973 144.9724 0.00053358 -81.6868 0.060953
2.165 0.98804 5.512e-005 3.8182 0.012021 2.8448e-005 0.0011549 0.19843 0.00065898 0.19908 0.18284 0 0.034109 0.0389 0 0.98928 0.29117 0.081902 0.011134 4.8494 0.069477 8.4562e-005 0.82061 0.0058123 0.0065644 0.002586 0.88566 0.50033 5.8187e-006 2.3308e-005 0.13631 0.60628 0.67031 0.0019443 0.62038 0.46666 0.002651 0.42318 1.1011 1.0953 15.9974 144.9724 0.00053175 -81.8962 0.061953
2.166 0.98804 5.512e-005 3.8182 0.012021 2.8461e-005 0.0011549 0.19846 0.00065898 0.19911 0.18287 0 0.034107 0.0389 0 0.98937 0.29121 0.081918 0.011136 4.8502 0.069488 8.4577e-005 0.8206 0.005813 0.006565 0.0025058 0.90012 0.52298 5.6247e-006 2.2529e-005 0.13631 0.60743 0.67175 0.0019118 0.62208 0.46682 0.002601 0.42316 1.1033 1.0977 15.9975 144.9724 0.00052992 -82.0865 0.062953
2.167 0.98804 5.512e-005 3.8182 0.012021 2.8474e-005 0.0011549 0.19849 0.00065898 0.19914 0.1829 0 0.034106 0.0389 0 0.98947 0.29126 0.081933 0.011138 4.851 0.069499 8.4592e-005 0.82059 0.0058136 0.0065657 0.0024354 0.91259 0.54501 5.4546e-006 2.1845e-005 0.13632 0.60858 0.67318 0.0018828 0.62381 0.46699 0.0025567 0.42313 1.1056 1.1 15.9976 144.9724 0.00052811 -82.2592 0.063953
2.168 0.98804 5.5119e-005 3.8182 0.012021 2.8487e-005 0.0011549 0.19852 0.00065898 0.19917 0.18292 0 0.034104 0.0389 0 0.98956 0.2913 0.081948 0.011139 4.8518 0.06951 8.4606e-005 0.82057 0.0058143 0.0065664 0.0023731 0.9233 0.56637 5.305e-006 2.1243e-005 0.13633 0.60972 0.6746 0.0018568 0.62555 0.46716 0.0025174 0.42311 1.1079 1.1023 15.9977 144.9724 0.0005263 -82.4158 0.064953
2.169 0.98804 5.5119e-005 3.8182 0.012021 2.85e-005 0.0011549 0.19855 0.00065898 0.1992 0.18295 0 0.034102 0.0389 0 0.98966 0.29134 0.081964 0.011141 4.8526 0.069521 8.4621e-005 0.82056 0.0058149 0.006567 0.002318 0.93242 0.58703 5.1727e-006 2.0711e-005 0.13633 0.61087 0.676 0.0018336 0.62731 0.46732 0.0024826 0.42309 1.1102 1.1045 15.9977 144.9724 0.0005245 -82.5578 0.065953
2.17 0.98804 5.5119e-005 3.8182 0.012021 2.8514e-005 0.0011549 0.19858 0.00065898 0.19923 0.18298 0 0.034101 0.0389 0 0.98975 0.29139 0.081979 0.011143 4.8534 0.069533 8.4636e-005 0.82055 0.0058156 0.0065677 0.0022692 0.94017 0.60696 5.0557e-006 2.024e-005 0.13634 0.61201 0.6774 0.0018128 0.62908 0.46749 0.0024515 0.42307 1.1124 1.1068 15.9978 144.9724 0.00052271 -82.6865 0.066953
2.171 0.98804 5.5119e-005 3.8182 0.012021 2.8527e-005 0.0011549 0.19861 0.00065898 0.19926 0.18301 0 0.034099 0.0389 0 0.98985 0.29143 0.081994 0.011145 4.8542 0.069544 8.465e-005 0.82054 0.0058162 0.0065684 0.0022257 0.94672 0.62613 4.9519e-006 1.9823e-005 0.13634 0.61315 0.67878 0.0017942 0.63086 0.46766 0.0024238 0.42305 1.1147 1.1091 15.9979 144.9724 0.00052093 -82.8033 0.067953
2.172 0.98804 5.5119e-005 3.8182 0.012021 2.854e-005 0.0011549 0.19864 0.00065898 0.19929 0.18303 0 0.034097 0.0389 0 0.98994 0.29147 0.08201 0.011146 4.855 0.069555 8.4665e-005 0.82053 0.0058168 0.0065691 0.0021871 0.95223 0.64456 4.8596e-006 1.9452e-005 0.13635 0.61429 0.68015 0.0017775 0.63266 0.46783 0.0023991 0.42304 1.117 1.1114 15.998 144.9724 0.00051916 -82.9092 0.068953
2.173 0.98804 5.5119e-005 3.8182 0.012021 2.8553e-005 0.0011549 0.19867 0.00065899 0.19932 0.18306 0 0.034096 0.0389 0 0.99004 0.29151 0.082025 0.011148 4.8559 0.069566 8.468e-005 0.82052 0.0058175 0.0065697 0.0021525 0.95685 0.66223 4.7774e-006 1.9121e-005 0.13635 0.61542 0.68152 0.0017624 0.63446 0.468 0.0023769 0.42302 1.1192 1.1137 15.9981 144.9724 0.0005174 -83.0053 0.069953
2.174 0.98804 5.5119e-005 3.8182 0.012021 2.8566e-005 0.0011549 0.1987 0.00065899 0.19935 0.18309 0 0.034094 0.0389 0 0.99013 0.29156 0.08204 0.01115 4.8567 0.069577 8.4694e-005 0.82051 0.0058181 0.0065704 0.0021216 0.96072 0.67914 4.7038e-006 1.8826e-005 0.13636 0.61655 0.68287 0.0017489 0.63627 0.46817 0.0023571 0.42301 1.1215 1.116 15.9982 144.9724 0.00051565 -83.0926 0.070953
2.175 0.98804 5.5119e-005 3.8182 0.012021 2.8579e-005 0.0011549 0.19873 0.00065899 0.19938 0.18312 0 0.034093 0.0389 0 0.99023 0.2916 0.082056 0.011152 4.8575 0.069588 8.4709e-005 0.8205 0.0058188 0.0065711 0.0020939 0.96396 0.69531 4.6379e-006 1.8561e-005 0.13636 0.61768 0.6842 0.0017366 0.63808 0.46834 0.0023392 0.423 1.1237 1.1182 15.9983 144.9724 0.0005139 -83.172 0.071953
2.176 0.98804 5.5119e-005 3.8182 0.012021 2.8592e-005 0.0011549 0.19876 0.00065899 0.19941 0.18315 0 0.034091 0.0389 0 0.99032 0.29164 0.082071 0.011154 4.8583 0.069599 8.4724e-005 0.82049 0.0058194 0.0065718 0.0020689 0.96665 0.71075 4.5788e-006 1.8324e-005 0.13637 0.61881 0.68553 0.0017256 0.6399 0.46851 0.0023231 0.42298 1.126 1.1205 15.9984 144.9724 0.00051217 -83.2442 0.072953
2.177 0.98804 5.5119e-005 3.8182 0.012021 2.8605e-005 0.0011549 0.19878 0.00065899 0.19944 0.18317 0 0.034089 0.0389 0 0.99042 0.29169 0.082087 0.011155 4.8591 0.06961 8.4738e-005 0.82047 0.0058201 0.0065724 0.0020465 0.96891 0.72548 4.5255e-006 1.811e-005 0.13637 0.61993 0.68685 0.0017155 0.64173 0.46869 0.0023086 0.42297 1.1282 1.1228 15.9985 144.9724 0.00051044 -83.3101 0.073953
2.178 0.98804 5.5119e-005 3.8182 0.012021 2.8618e-005 0.0011549 0.19881 0.00065899 0.19947 0.1832 0 0.034088 0.0389 0 0.99051 0.29173 0.082102 0.011157 4.8599 0.069622 8.4753e-005 0.82046 0.0058207 0.0065731 0.0020261 0.97078 0.73952 4.4774e-006 1.7916e-005 0.13638 0.62105 0.68816 0.0017064 0.64355 0.46886 0.0022955 0.42296 1.1305 1.125 15.9986 144.9724 0.00050873 -83.3703 0.074953
2.179 0.98804 5.5119e-005 3.8182 0.01202 2.8631e-005 0.0011549 0.19884 0.00065899 0.1995 0.18323 0 0.034086 0.0389 0 0.99061 0.29177 0.082117 0.011159 4.8607 0.069633 8.4768e-005 0.82045 0.0058214 0.0065738 0.0020077 0.97235 0.75288 4.4339e-006 1.7742e-005 0.13638 0.62217 0.68946 0.0016982 0.64538 0.46903 0.0022836 0.42295 1.1327 1.1273 15.9987 144.9724 0.00050702 -83.4253 0.075953
2.18 0.98804 5.5119e-005 3.8182 0.01202 2.8644e-005 0.0011549 0.19887 0.00065899 0.19953 0.18326 0 0.034084 0.0389 0 0.9907 0.29181 0.082133 0.011161 4.8615 0.069644 8.4782e-005 0.82044 0.005822 0.0065745 0.0019911 0.97365 0.76558 4.3943e-006 1.7583e-005 0.13639 0.62328 0.69074 0.0016906 0.6472 0.4692 0.0022728 0.42294 1.135 1.1295 15.9988 144.9724 0.00050532 -83.4758 0.076953
2.181 0.98804 5.5119e-005 3.8182 0.01202 2.8658e-005 0.0011549 0.1989 0.00065899 0.19956 0.18328 0 0.034083 0.0389 0 0.99079 0.29186 0.082148 0.011162 4.8624 0.069655 8.4797e-005 0.82043 0.0058227 0.0065751 0.0019758 0.97474 0.77766 4.3584e-006 1.7439e-005 0.13639 0.62439 0.69202 0.0016837 0.64903 0.46937 0.002263 0.42293 1.1372 1.1318 15.9989 144.9724 0.00050364 -83.5221 0.077953
2.182 0.98804 5.5119e-005 3.8182 0.01202 2.8671e-005 0.0011549 0.19893 0.00065899 0.19959 0.18331 0 0.034081 0.0389 0 0.99089 0.2919 0.082163 0.011164 4.8632 0.069666 8.4812e-005 0.82042 0.0058233 0.0065758 0.0019618 0.97566 0.78914 4.3255e-006 1.7307e-005 0.1364 0.6255 0.69329 0.0016774 0.65085 0.46955 0.002254 0.42292 1.1394 1.134 15.9989 144.9724 0.00050196 -83.5648 0.078953
2.183 0.98804 5.5118e-005 3.8182 0.01202 2.8684e-005 0.0011549 0.19896 0.00065899 0.19961 0.18334 0 0.03408 0.0389 0 0.99098 0.29194 0.082179 0.011166 4.864 0.069677 8.4826e-005 0.82041 0.005824 0.0065765 0.001949 0.97642 0.80003 4.2953e-006 1.7185e-005 0.13641 0.6266 0.69454 0.0016716 0.65267 0.46972 0.0022458 0.42292 1.1416 1.1363 15.999 144.9724 0.00050029 -83.6042 0.079953
2.184 0.98804 5.5118e-005 3.8182 0.01202 2.8697e-005 0.0011549 0.19899 0.00065899 0.19964 0.18337 0 0.034078 0.0389 0 0.99108 0.29199 0.082194 0.011168 4.8648 0.069688 8.4841e-005 0.8204 0.0058246 0.0065771 0.0019373 0.97707 0.81037 4.2676e-006 1.7074e-005 0.13641 0.6277 0.69579 0.0016662 0.65449 0.46989 0.0022382 0.42291 1.1439 1.1385 15.9991 144.9724 0.00049863 -83.6407 0.080953
2.185 0.98804 5.5118e-005 3.8182 0.01202 2.871e-005 0.0011549 0.19902 0.00065899 0.19967 0.1834 0 0.034076 0.0389 0 0.99117 0.29203 0.08221 0.01117 4.8656 0.069699 8.4856e-005 0.82039 0.0058253 0.0065778 0.0019264 0.97762 0.82017 4.2421e-006 1.6972e-005 0.13642 0.6288 0.69703 0.0016613 0.6563 0.47006 0.0022312 0.4229 1.1461 1.1407 15.9992 144.9724 0.00049697 -83.6746 0.081953
2.186 0.98804 5.5118e-005 3.8182 0.01202 2.8723e-005 0.0011549 0.19905 0.00065899 0.1997 0.18342 0 0.034075 0.0389 0 0.99127 0.29207 0.082225 0.011171 4.8664 0.06971 8.4871e-005 0.82037 0.0058259 0.0065785 0.0019164 0.97808 0.82946 4.2184e-006 1.6877e-005 0.13642 0.6299 0.69825 0.0016566 0.65811 0.47024 0.0022248 0.4229 1.1483 1.143 15.9993 144.9724 0.00049533 -83.7061 0.082953
2.187 0.98804 5.5118e-005 3.8182 0.01202 2.8736e-005 0.0011549 0.19908 0.00065899 0.19973 0.18345 0 0.034073 0.0389 0 0.99136 0.29211 0.08224 0.011173 4.8673 0.069722 8.4885e-005 0.82036 0.0058266 0.0065792 0.0019071 0.97848 0.83826 4.1965e-006 1.6789e-005 0.13643 0.63099 0.69947 0.0016524 0.65992 0.47041 0.0022188 0.42289 1.1505 1.1452 15.9994 144.9724 0.0004937 -83.7355 0.083953
2.188 0.98804 5.5118e-005 3.8182 0.01202 2.8749e-005 0.0011549 0.19911 0.00065899 0.19976 0.18348 0 0.034072 0.0389 0 0.99146 0.29216 0.082256 0.011175 4.8681 0.069733 8.49e-005 0.82035 0.0058272 0.0065799 0.0018983 0.97882 0.8466 4.176e-006 1.6707e-005 0.13643 0.63208 0.70068 0.0016484 0.66172 0.47058 0.0022132 0.42288 1.1527 1.1474 15.9995 144.9724 0.00049207 -83.763 0.084953
2.189 0.98804 5.5118e-005 3.8182 0.01202 2.8762e-005 0.0011549 0.19914 0.00065899 0.19979 0.18351 0 0.03407 0.0389 0 0.99155 0.2922 0.082271 0.011177 4.8689 0.069744 8.4915e-005 0.82034 0.0058279 0.0065805 0.0018902 0.97911 0.8545 4.1569e-006 1.663e-005 0.13644 0.63316 0.70188 0.0016446 0.66352 0.47076 0.002208 0.42288 1.1549 1.1497 15.9996 144.9724 0.00049046 -83.7889 0.085953
2.19 0.98804 5.5118e-005 3.8182 0.01202 2.8775e-005 0.0011549 0.19916 0.00065899 0.19982 0.18353 0 0.034068 0.0389 0 0.99165 0.29224 0.082286 0.011178 4.8697 0.069755 8.4929e-005 0.82033 0.0058285 0.0065812 0.0018826 0.97937 0.86197 4.139e-006 1.6558e-005 0.13644 0.63425 0.70307 0.0016411 0.66532 0.47093 0.0022032 0.42287 1.1571 1.1519 15.9997 144.9724 0.00048885 -83.8133 0.086953
2.191 0.98804 5.5118e-005 3.8182 0.01202 2.8788e-005 0.0011549 0.19919 0.00065899 0.19985 0.18356 0 0.034067 0.0389 0 0.99174 0.29229 0.082302 0.01118 4.8705 0.069766 8.4944e-005 0.82032 0.0058291 0.0065819 0.0018754 0.97959 0.86905 4.1221e-006 1.6491e-005 0.13645 0.63533 0.70425 0.0016378 0.6671 0.4711 0.0021986 0.42287 1.1593 1.1541 15.9997 144.9724 0.00048725 -83.8363 0.087953
2.192 0.98804 5.5118e-005 3.8182 0.01202 2.8802e-005 0.0011549 0.19922 0.00065899 0.19988 0.18359 0 0.034065 0.0389 0 0.99184 0.29233 0.082317 0.011182 4.8714 0.069777 8.4959e-005 0.82031 0.0058298 0.0065826 0.0018686 0.97978 0.87574 4.1061e-006 1.6427e-005 0.13645 0.6364 0.70543 0.0016346 0.66888 0.47128 0.0021943 0.42286 1.1615 1.1563 15.9998 144.9725 0.00048566 -83.8582 0.088953
2.193 0.98804 5.5118e-005 3.8182 0.01202 2.8815e-005 0.0011549 0.19925 0.00065899 0.19991 0.18361 0 0.034064 0.0389 0 0.99193 0.29237 0.082333 0.011184 4.8722 0.069788 8.4973e-005 0.8203 0.0058304 0.0065832 0.0018622 0.97996 0.88207 4.0911e-006 1.6366e-005 0.13646 0.63747 0.70659 0.0016316 0.67066 0.47145 0.0021902 0.42286 1.1637 1.1585 15.9999 144.9725 0.00048408 -83.879 0.089953
2.194 0.98804 5.5118e-005 3.8182 0.01202 2.8828e-005 0.0011549 0.19928 0.00065899 0.19993 0.18364 0 0.034062 0.0389 0 0.99203 0.29242 0.082348 0.011186 4.873 0.069799 8.4988e-005 0.82029 0.0058311 0.0065839 0.0018561 0.98011 0.88806 4.0767e-006 1.6309e-005 0.13646 0.63854 0.70775 0.0016288 0.67243 0.47163 0.0021863 0.42285 1.1659 1.1607 16 144.9725 0.00048251 -83.8988 0.090953
2.195 0.98804 5.5118e-005 3.8182 0.01202 2.8841e-005 0.0011549 0.19931 0.00065899 0.19996 0.18367 0 0.03406 0.0389 0 0.99212 0.29246 0.082363 0.011187 4.8738 0.069811 8.5003e-005 0.82027 0.0058317 0.0065846 0.0018502 0.98026 0.89372 4.063e-006 1.6254e-005 0.13647 0.63961 0.70889 0.0016261 0.67419 0.4718 0.0021827 0.42285 1.168 1.1629 16.0001 144.9725 0.00048094 -83.9177 0.091953
2.196 0.98804 5.5118e-005 3.8182 0.01202 2.8854e-005 0.0011549 0.19934 0.00065899 0.19999 0.1837 0 0.034059 0.0389 0 0.99222 0.2925 0.082379 0.011189 4.8746 0.069822 8.5017e-005 0.82026 0.0058324 0.0065853 0.0018447 0.98038 0.89908 4.05e-006 1.6202e-005 0.13647 0.64067 0.71003 0.0016235 0.67595 0.47197 0.0021792 0.42284 1.1702 1.1651 16.0002 144.9725 0.00047939 -83.9358 0.092953
2.197 0.98804 5.5118e-005 3.8182 0.01202 2.8867e-005 0.0011549 0.19937 0.00065899 0.20002 0.18372 0 0.034057 0.0389 0 0.99231 0.29254 0.082394 0.011191 4.8755 0.069833 8.5032e-005 0.82025 0.005833 0.0065859 0.0018393 0.9805 0.90413 4.0375e-006 1.6152e-005 0.13648 0.64173 0.71116 0.001621 0.6777 0.47215 0.0021758 0.42284 1.1724 1.1673 16.0002 144.9725 0.00047784 -83.9533 0.093953
2.198 0.98804 5.5117e-005 3.8182 0.01202 2.888e-005 0.0011549 0.1994 0.00065899 0.20005 0.18375 0 0.034056 0.0389 0 0.99241 0.29259 0.08241 0.011193 4.8763 0.069844 8.5047e-005 0.82024 0.0058337 0.0065866 0.0018342 0.98061 0.90892 4.0255e-006 1.6104e-005 0.13649 0.64279 0.71228 0.0016186 0.67945 0.47232 0.0021726 0.42284 1.1745 1.1695 16.0003 144.9725 0.0004763 -83.9701 0.094953
2.199 0.98804 5.5117e-005 3.8182 0.01202 2.8893e-005 0.0011549 0.19942 0.00065899 0.20008 0.18378 0 0.034054 0.0389 0 0.9925 0.29263 0.082425 0.011194 4.8771 0.069855 8.5062e-005 0.82023 0.0058343 0.0065873 0.0018292 0.98071 0.91344 4.014e-006 1.6057e-005 0.13649 0.64384 0.71339 0.0016163 0.68119 0.47249 0.0021695 0.42283 1.1767 1.1716 16.0004 144.9725 0.00047477 -83.9864 0.095953
2.2 0.98804 5.5117e-005 3.8182 0.01202 2.8906e-005 0.0011549 0.19945 0.00065899 0.20011 0.18381 0 0.034052 0.0389 0 0.9926 0.29267 0.08244 0.011196 4.8779 0.069866 8.5076e-005 0.82022 0.005835 0.006588 0.0018245 0.9808 0.9177 4.0028e-006 1.6013e-005 0.1365 0.6449 0.7145 0.0016141 0.68292 0.47267 0.0021665 0.42283 1.1789 1.1738 16.0005 144.9725 0.00047325 -84.0021 0.096953
2.201 0.98804 5.5117e-005 3.8182 0.01202 2.8919e-005 0.0011549 0.19948 0.00065899 0.20014 0.18383 0 0.034051 0.0389 0 0.99269 0.29272 0.082456 0.011198 4.8787 0.069877 8.5091e-005 0.82021 0.0058356 0.0065886 0.0018199 0.98089 0.92174 3.992e-006 1.5969e-005 0.1365 0.64594 0.7156 0.0016119 0.68464 0.47284 0.0021636 0.42283 1.181 1.176 16.0006 144.9725 0.00047174 -84.0174 0.097953
2.202 0.98804 5.5117e-005 3.8182 0.01202 2.8932e-005 0.0011549 0.19951 0.00065899 0.20017 0.18386 0 0.034049 0.0389 0 0.99279 0.29276 0.082471 0.0112 4.8796 0.069888 8.5106e-005 0.8202 0.0058363 0.0065893 0.0018154 0.98097 0.92555 3.9815e-006 1.5927e-005 0.13651 0.64699 0.71669 0.0016098 0.68636 0.47302 0.0021608 0.42282 1.1832 1.1782 16.0006 144.9725 0.00047023 -84.0322 0.098953
2.203 0.98804 5.5117e-005 3.8182 0.01202 2.8946e-005 0.0011549 0.19954 0.00065899 0.20019 0.18389 0 0.034048 0.0389 0 0.99288 0.2928 0.082487 0.011202 4.8804 0.0699 8.512e-005 0.82019 0.0058369 0.00659 0.001811 0.98104 0.92915 3.9713e-006 1.5887e-005 0.13651 0.64803 0.71777 0.0016078 0.68807 0.47319 0.0021581 0.42282 1.1853 1.1803 16.0007 144.9725 0.00046874 -84.0467 0.099953
2.204 0.98804 5.5117e-005 3.8182 0.01202 2.8959e-005 0.0011549 0.19957 0.00065899 0.20022 0.18391 0 0.034046 0.0389 0 0.99298 0.29285 0.082502 0.011203 4.8812 0.069911 8.5135e-005 0.82017 0.0058376 0.0065907 0.0018068 0.98112 0.93255 3.9614e-006 1.5847e-005 0.13652 0.64907 0.71884 0.0016058 0.68977 0.47336 0.0021555 0.42282 1.1875 1.1825 16.0008 144.9725 0.00046725 -84.0608 0.10095
2.205 0.98804 5.5117e-005 3.8182 0.01202 2.8972e-005 0.0011549 0.1996 0.000659 0.20025 0.18394 0 0.034044 0.0389 0 0.99307 0.29289 0.082517 0.011205 4.882 0.069922 8.515e-005 0.82016 0.0058382 0.0065914 0.0018027 0.98119 0.93575 3.9518e-006 1.5808e-005 0.13652 0.6501 0.7199 0.0016039 0.69147 0.47354 0.0021529 0.42281 1.1896 1.1846 16.0009 144.9726 0.00046577 -84.0745 0.10195
2.206 0.98804 5.5117e-005 3.8182 0.01202 2.8985e-005 0.0011549 0.19963 0.000659 0.20028 0.18397 0 0.034043 0.0389 0 0.99317 0.29293 0.082533 0.011207 4.8829 0.069933 8.5164e-005 0.82015 0.0058389 0.006592 0.0017986 0.98125 0.93879 3.9424e-006 1.5771e-005 0.13653 0.65113 0.72096 0.001602 0.69316 0.47371 0.0021504 0.42281 1.1917 1.1868 16.001 144.9726 0.0004643 -84.088 0.10295
2.207 0.98804 5.5117e-005 3.8182 0.01202 2.8998e-005 0.0011549 0.19965 0.000659 0.20031 0.184 0 0.034041 0.0389 0 0.99326 0.29297 0.082548 0.011209 4.8837 0.069944 8.5179e-005 0.82014 0.0058396 0.0065927 0.0017947 0.98131 0.94165 3.9332e-006 1.5734e-005 0.13653 0.65216 0.72201 0.0016001 0.69484 0.47389 0.0021479 0.42281 1.1939 1.1889 16.001 144.9726 0.00046283 -84.1012 0.10395
2.208 0.98804 5.5117e-005 3.8182 0.01202 2.9011e-005 0.0011549 0.19968 0.000659 0.20034 0.18402 0 0.03404 0.0389 0 0.99336 0.29302 0.082564 0.01121 4.8845 0.069955 8.5194e-005 0.82013 0.0058402 0.0065934 0.0017908 0.98138 0.94435 3.9242e-006 1.5698e-005 0.13654 0.65319 0.72305 0.0015983 0.69652 0.47406 0.0021455 0.42281 1.196 1.1911 16.0011 144.9726 0.00046138 -84.1141 0.10495
2.209 0.98804 5.5117e-005 3.8182 0.01202 2.9024e-005 0.0011549 0.19971 0.000659 0.20037 0.18405 0 0.034038 0.0389 0 0.99345 0.29306 0.082579 0.011212 4.8853 0.069966 8.5209e-005 0.82012 0.0058409 0.0065941 0.0017871 0.98144 0.9469 3.9153e-006 1.5662e-005 0.13654 0.65421 0.72409 0.0015965 0.69819 0.47424 0.0021432 0.42281 1.1981 1.1932 16.0012 144.9726 0.00045993 -84.1268 0.10595
2.21 0.98804 5.5117e-005 3.8182 0.01202 2.9037e-005 0.0011549 0.19974 0.000659 0.2004 0.18408 0 0.034037 0.0389 0 0.99355 0.2931 0.082595 0.011214 4.8862 0.069977 8.5223e-005 0.82011 0.0058415 0.0065948 0.0017834 0.98149 0.94931 3.9067e-006 1.5628e-005 0.13655 0.65523 0.72512 0.0015948 0.69985 0.47441 0.0021409 0.4228 1.2003 1.1954 16.0013 144.9726 0.00045849 -84.1393 0.10695
2.211 0.98804 5.5117e-005 3.8182 0.01202 2.905e-005 0.0011549 0.19977 0.000659 0.20042 0.1841 0 0.034035 0.0389 0 0.99364 0.29315 0.08261 0.011216 4.887 0.069989 8.5238e-005 0.8201 0.0058422 0.0065954 0.0017797 0.98155 0.95158 3.8982e-006 1.5594e-005 0.13655 0.65624 0.72614 0.0015931 0.7015 0.47458 0.0021386 0.4228 1.2024 1.1975 16.0014 144.9726 0.00045705 -84.1516 0.10795
2.212 0.98804 5.5117e-005 3.8182 0.01202 2.9063e-005 0.0011549 0.1998 0.000659 0.20045 0.18413 0 0.034033 0.0389 0 0.99374 0.29319 0.082625 0.011218 4.8878 0.07 8.5253e-005 0.82009 0.0058428 0.0065961 0.0017762 0.9816 0.95373 3.8899e-006 1.556e-005 0.13656 0.65726 0.72715 0.0015914 0.70315 0.47476 0.0021364 0.4228 1.2045 1.1996 16.0014 144.9726 0.00045563 -84.1637 0.10895
2.213 0.98804 5.5116e-005 3.8182 0.01202 2.9076e-005 0.0011549 0.19983 0.000659 0.20048 0.18416 0 0.034032 0.0389 0 0.99384 0.29323 0.082641 0.011219 4.8887 0.070011 8.5267e-005 0.82007 0.0058435 0.0065968 0.0017726 0.98166 0.95575 3.8817e-006 1.5528e-005 0.13657 0.65827 0.72816 0.0015897 0.70479 0.47493 0.0021342 0.4228 1.2066 1.2018 16.0015 144.9726 0.00045421 -84.1756 0.10995
2.214 0.98804 5.5116e-005 3.8182 0.01202 2.909e-005 0.0011549 0.19985 0.000659 0.20051 0.18419 0 0.03403 0.0389 0 0.99393 0.29328 0.082656 0.011221 4.8895 0.070022 8.5282e-005 0.82006 0.0058441 0.0065975 0.0017692 0.98171 0.95766 3.8736e-006 1.5495e-005 0.13657 0.65927 0.72916 0.0015881 0.70642 0.47511 0.0021321 0.4228 1.2087 1.2039 16.0016 144.9726 0.0004528 -84.1874 0.11095
2.215 0.98804 5.5116e-005 3.8182 0.01202 2.9103e-005 0.0011549 0.19988 0.000659 0.20054 0.18421 0 0.034029 0.0389 0 0.99403 0.29332 0.082672 0.011223 4.8903 0.070033 8.5297e-005 0.82005 0.0058448 0.0065982 0.0017658 0.98176 0.95946 3.8656e-006 1.5463e-005 0.13658 0.66028 0.73015 0.0015865 0.70805 0.47528 0.00213 0.4228 1.2108 1.206 16.0017 144.9726 0.0004514 -84.199 0.11195
2.216 0.98804 5.5116e-005 3.8182 0.01202 2.9116e-005 0.0011549 0.19991 0.000659 0.20057 0.18424 0 0.034027 0.0389 0 0.99412 0.29336 0.082687 0.011225 4.8911 0.070044 8.5312e-005 0.82004 0.0058454 0.0065988 0.0017624 0.98181 0.96117 3.8578e-006 1.5432e-005 0.13658 0.66128 0.73113 0.0015849 0.70966 0.47545 0.0021279 0.4228 1.2129 1.2081 16.0017 144.9727 0.00045 -84.2104 0.11295
2.217 0.98804 5.5116e-005 3.8182 0.01202 2.9129e-005 0.0011549 0.19994 0.000659 0.20059 0.18427 0 0.034026 0.0389 0 0.99422 0.29341 0.082702 0.011226 4.892 0.070055 8.5326e-005 0.82003 0.0058461 0.0065995 0.0017591 0.98186 0.96277 3.8501e-006 1.5401e-005 0.13659 0.66228 0.73211 0.0015833 0.71127 0.47563 0.0021258 0.42279 1.215 1.2102 16.0018 144.9727 0.00044861 -84.2218 0.11395
2.218 0.98804 5.5116e-005 3.8182 0.01202 2.9142e-005 0.0011549 0.19997 0.000659 0.20062 0.18429 0 0.034024 0.0389 0 0.99431 0.29345 0.082718 0.011228 4.8928 0.070067 8.5341e-005 0.82002 0.0058467 0.0066002 0.0017558 0.98191 0.96429 3.8425e-006 1.5371e-005 0.13659 0.66327 0.73308 0.0015818 0.71288 0.4758 0.0021238 0.42279 1.2171 1.2123 16.0019 144.9727 0.00044723 -84.2329 0.11495
2.219 0.98804 5.5116e-005 3.8182 0.01202 2.9155e-005 0.0011549 0.2 0.000659 0.20065 0.18432 0 0.034022 0.0389 0 0.99441 0.29349 0.082733 0.01123 4.8936 0.070078 8.5356e-005 0.82001 0.0058474 0.0066009 0.0017526 0.98196 0.96572 3.835e-006 1.5341e-005 0.1366 0.66426 0.73405 0.0015802 0.71447 0.47598 0.0021218 0.42279 1.2192 1.2144 16.0019 144.9727 0.00044586 -84.244 0.11595
2.22 0.98804 5.5116e-005 3.8182 0.01202 2.9168e-005 0.0011549 0.20003 0.000659 0.20068 0.18435 0 0.034021 0.0389 0 0.9945 0.29353 0.082749 0.011232 4.8945 0.070089 8.537e-005 0.82 0.005848 0.0066016 0.0017494 0.982 0.96707 3.8276e-006 1.5311e-005 0.1366 0.66525 0.73501 0.0015787 0.71606 0.47615 0.0021198 0.42279 1.2212 1.2165 16.002 144.9727 0.0004445 -84.2549 0.11695
2.221 0.98804 5.5116e-005 3.8182 0.01202 2.9181e-005 0.0011549 0.20005 0.000659 0.20071 0.18437 0 0.034019 0.0389 0 0.9946 0.29358 0.082764 0.011234 4.8953 0.0701 8.5385e-005 0.81999 0.0058487 0.0066022 0.0017463 0.98205 0.96834 3.8202e-006 1.5282e-005 0.13661 0.66624 0.73596 0.0015773 0.71765 0.47633 0.0021178 0.42279 1.2233 1.2186 16.0021 144.9727 0.00044314 -84.2657 0.11795
2.222 0.98804 5.5116e-005 3.8182 0.01202 2.9194e-005 0.0011549 0.20008 0.000659 0.20074 0.1844 0 0.034018 0.0389 0 0.99469 0.29362 0.08278 0.011235 4.8961 0.070111 8.54e-005 0.81997 0.0058493 0.0066029 0.0017432 0.98209 0.96954 3.813e-006 1.5253e-005 0.13661 0.66722 0.7369 0.0015758 0.71922 0.4765 0.0021159 0.42279 1.2254 1.2207 16.0022 144.9727 0.00044179 -84.2764 0.11895
2.223 0.98804 5.5116e-005 3.8182 0.01202 2.9207e-005 0.0011549 0.20011 0.000659 0.20076 0.18443 0 0.034016 0.0389 0 0.99479 0.29366 0.082795 0.011237 4.897 0.070122 8.5415e-005 0.81996 0.00585 0.0066036 0.0017401 0.98214 0.97068 3.8059e-006 1.5224e-005 0.13662 0.6682 0.73784 0.0015743 0.72079 0.47667 0.002114 0.42279 1.2274 1.2228 16.0022 144.9727 0.00044044 -84.287 0.11995
2.224 0.98804 5.5116e-005 3.8182 0.01202 2.922e-005 0.0011549 0.20014 0.000659 0.20079 0.18445 0 0.034015 0.0389 0 0.99488 0.29371 0.08281 0.011239 4.8978 0.070133 8.5429e-005 0.81995 0.0058506 0.0066043 0.0017371 0.98218 0.97175 3.7988e-006 1.5196e-005 0.13662 0.66918 0.73877 0.0015729 0.72235 0.47685 0.0021121 0.42279 1.2295 1.2249 16.0023 144.9727 0.00043911 -84.2975 0.12095
2.225 0.98804 5.5116e-005 3.8182 0.01202 2.9234e-005 0.0011549 0.20017 0.000659 0.20082 0.18448 0 0.034013 0.0389 0 0.99498 0.29375 0.082826 0.011241 4.8986 0.070145 8.5444e-005 0.81994 0.0058513 0.006605 0.0017341 0.98222 0.97276 3.7918e-006 1.5168e-005 0.13663 0.67015 0.7397 0.0015714 0.7239 0.47702 0.0021102 0.42279 1.2316 1.2269 16.0024 144.9727 0.00043778 -84.3079 0.12195
2.226 0.98804 5.5116e-005 3.8182 0.01202 2.9247e-005 0.0011549 0.2002 0.000659 0.20085 0.18451 0 0.034012 0.0389 0 0.99507 0.29379 0.082841 0.011242 4.8995 0.070156 8.5459e-005 0.81993 0.005852 0.0066057 0.0017311 0.98227 0.97371 3.7849e-006 1.5141e-005 0.13664 0.67112 0.74062 0.00157 0.72545 0.4772 0.0021084 0.42279 1.2336 1.229 16.0024 144.9728 0.00043646 -84.3182 0.12295
2.227 0.98804 5.5116e-005 3.8182 0.01202 2.926e-005 0.0011549 0.20022 0.000659 0.20088 0.18453 0 0.03401 0.0389 0 0.99517 0.29384 0.082857 0.011244 4.9003 0.070167 8.5473e-005 0.81992 0.0058526 0.0066063 0.0017282 0.98231 0.97461 3.7781e-006 1.5113e-005 0.13664 0.67209 0.74153 0.0015686 0.72699 0.47737 0.0021065 0.42279 1.2357 1.2311 16.0025 144.9728 0.00043514 -84.3284 0.12395
2.228 0.98804 5.5115e-005 3.8182 0.01202 2.9273e-005 0.0011549 0.20025 0.000659 0.20091 0.18456 0 0.034008 0.0389 0 0.99526 0.29388 0.082872 0.011246 4.9011 0.070178 8.5488e-005 0.81991 0.0058533 0.006607 0.0017253 0.98235 0.97546 3.7714e-006 1.5086e-005 0.13665 0.67305 0.74244 0.0015672 0.72852 0.47754 0.0021047 0.42279 1.2377 1.2331 16.0026 144.9728 0.00043383 -84.3385 0.12495
2.229 0.98804 5.5115e-005 3.8182 0.01202 2.9286e-005 0.0011549 0.20028 0.000659 0.20093 0.18459 0 0.034007 0.0389 0 0.99536 0.29392 0.082888 0.011248 4.902 0.070189 8.5503e-005 0.8199 0.0058539 0.0066077 0.0017224 0.98239 0.97626 3.7647e-006 1.506e-005 0.13665 0.67402 0.74334 0.0015659 0.73005 0.47772 0.0021029 0.42279 1.2398 1.2352 16.0026 144.9728 0.00043253 -84.3485 0.12595
2.23 0.98804 5.5115e-005 3.8182 0.01202 2.9299e-005 0.0011549 0.20031 0.000659 0.20096 0.18461 0 0.034005 0.0389 0 0.99545 0.29397 0.082903 0.01125 4.9028 0.0702 8.5518e-005 0.81989 0.0058546 0.0066084 0.0017196 0.98243 0.97701 3.7581e-006 1.5033e-005 0.13666 0.67497 0.74424 0.0015645 0.73156 0.47789 0.0021012 0.42279 1.2418 1.2373 16.0027 144.9728 0.00043124 -84.3584 0.12695
2.231 0.98804 5.5115e-005 3.8182 0.01202 2.9312e-005 0.0011549 0.20034 0.000659 0.20099 0.18464 0 0.034004 0.0389 0 0.99555 0.29401 0.082919 0.011251 4.9037 0.070211 8.5532e-005 0.81987 0.0058552 0.0066091 0.0017168 0.98247 0.97772 3.7515e-006 1.5007e-005 0.13666 0.67593 0.74513 0.0015632 0.73308 0.47807 0.0020994 0.4228 1.2438 1.2393 16.0028 144.9728 0.00042995 -84.3682 0.12795
2.232 0.98804 5.5115e-005 3.8182 0.01202 2.9325e-005 0.0011549 0.20036 0.000659 0.20102 0.18467 0 0.034002 0.0389 0 0.99564 0.29405 0.082934 0.011253 4.9045 0.070222 8.5547e-005 0.81986 0.0058559 0.0066098 0.001714 0.98251 0.9784 3.7451e-006 1.4981e-005 0.13667 0.67688 0.74601 0.0015618 0.73458 0.47824 0.0020977 0.4228 1.2459 1.2414 16.0028 144.9728 0.00042867 -84.378 0.12895
2.233 0.98804 5.5115e-005 3.8182 0.01202 2.9338e-005 0.0011549 0.20039 0.000659 0.20105 0.18469 0 0.034001 0.0389 0 0.99574 0.2941 0.082949 0.011255 4.9053 0.070234 8.5562e-005 0.81985 0.0058565 0.0066104 0.0017113 0.98255 0.97903 3.7387e-006 1.4955e-005 0.13667 0.67783 0.74689 0.0015605 0.73608 0.47842 0.0020959 0.4228 1.2479 1.2434 16.0029 144.9728 0.00042739 -84.3876 0.12995
2.234 0.98804 5.5115e-005 3.8182 0.01202 2.9351e-005 0.0011549 0.20042 0.000659 0.20107 0.18472 0 0.033999 0.0389 0 0.99583 0.29414 0.082965 0.011257 4.9062 0.070245 8.5577e-005 0.81984 0.0058572 0.0066111 0.0017085 0.98259 0.97963 3.7324e-006 1.493e-005 0.13668 0.67878 0.74776 0.0015592 0.73757 0.47859 0.0020942 0.4228 1.2499 1.2454 16.003 144.9728 0.00042613 -84.3972 0.13095
2.235 0.98804 5.5115e-005 3.8182 0.01202 2.9364e-005 0.0011549 0.20045 0.000659 0.2011 0.18475 0 0.033998 0.0389 0 0.99593 0.29418 0.08298 0.011259 4.907 0.070256 8.5591e-005 0.81983 0.0058579 0.0066118 0.0017058 0.98263 0.9802 3.7261e-006 1.4905e-005 0.13668 0.67973 0.74863 0.0015579 0.73905 0.47876 0.0020925 0.4228 1.2519 1.2475 16.003 144.9729 0.00042486 -84.4067 0.13195
2.236 0.98804 5.5115e-005 3.8182 0.01202 2.9378e-005 0.0011549 0.20048 0.000659 0.20113 0.18477 0 0.033996 0.0389 0 0.99603 0.29422 0.082996 0.01126 4.9078 0.070267 8.5606e-005 0.81982 0.0058585 0.0066125 0.0017031 0.98267 0.98073 3.7199e-006 1.488e-005 0.13669 0.68067 0.74949 0.0015566 0.74052 0.47894 0.0020908 0.4228 1.254 1.2495 16.0031 144.9729 0.00042361 -84.4161 0.13295
2.237 0.98804 5.5115e-005 3.8182 0.01202 2.9391e-005 0.0011549 0.2005 0.000659 0.20116 0.1848 0 0.033995 0.0389 0 0.99612 0.29427 0.083011 0.011262 4.9087 0.070278 8.5621e-005 0.81981 0.0058592 0.0066132 0.0017005 0.9827 0.98123 3.7138e-006 1.4856e-005 0.13669 0.68161 0.75035 0.0015554 0.74199 0.47911 0.0020892 0.4228 1.256 1.2515 16.0032 144.9729 0.00042236 -84.4254 0.13395
2.238 0.98804 5.5115e-005 3.8182 0.01202 2.9404e-005 0.0011549 0.20053 0.00065901 0.20119 0.18483 0 0.033993 0.0389 0 0.99622 0.29431 0.083027 0.011264 4.9095 0.070289 8.5636e-005 0.8198 0.0058598 0.0066139 0.0016979 0.98274 0.98171 3.7077e-006 1.4831e-005 0.1367 0.68254 0.75119 0.0015541 0.74345 0.47929 0.0020875 0.4228 1.258 1.2535 16.0032 144.9729 0.00042112 -84.4347 0.13495
2.239 0.98804 5.5115e-005 3.8182 0.01202 2.9417e-005 0.0011549 0.20056 0.00065901 0.20121 0.18485 0 0.033992 0.0389 0 0.99631 0.29435 0.083042 0.011266 4.9104 0.0703 8.565e-005 0.81979 0.0058605 0.0066145 0.0016953 0.98278 0.98216 3.7017e-006 1.4807e-005 0.13671 0.68347 0.75204 0.0015529 0.74491 0.47946 0.0020859 0.42281 1.26 1.2556 16.0033 144.9729 0.00041989 -84.4439 0.13595
2.24 0.98804 5.5115e-005 3.8182 0.01202 2.943e-005 0.0011549 0.20059 0.00065901 0.20124 0.18488 0 0.03399 0.0389 0 0.99641 0.2944 0.083058 0.011267 4.9112 0.070312 8.5665e-005 0.81977 0.0058611 0.0066152 0.0016928 0.98281 0.98258 3.6957e-006 1.4783e-005 0.13671 0.6844 0.75288 0.0015516 0.74635 0.47963 0.0020843 0.42281 1.262 1.2576 16.0034 144.9729 0.00041866 -84.453 0.13695
2.241 0.98804 5.5115e-005 3.8182 0.01202 2.9443e-005 0.0011549 0.20062 0.00065901 0.20127 0.1849 0 0.033988 0.0389 0 0.9965 0.29444 0.083073 0.011269 4.912 0.070323 8.568e-005 0.81976 0.0058618 0.0066159 0.0016902 0.98285 0.98298 3.6898e-006 1.476e-005 0.13672 0.68533 0.75371 0.0015504 0.7478 0.47981 0.0020827 0.42281 1.264 1.2596 16.0034 144.9729 0.00041744 -84.462 0.13795
2.242 0.98804 5.5115e-005 3.8182 0.01202 2.9456e-005 0.0011549 0.20064 0.00065901 0.2013 0.18493 0 0.033987 0.0389 0 0.9966 0.29448 0.083089 0.011271 4.9129 0.070334 8.5694e-005 0.81975 0.0058624 0.0066166 0.0016877 0.98288 0.98336 3.6839e-006 1.4736e-005 0.13672 0.68626 0.75454 0.0015492 0.74923 0.47998 0.0020811 0.42281 1.2659 1.2616 16.0035 144.9729 0.00041622 -84.471 0.13895
2.243 0.98804 5.5115e-005 3.8182 0.01202 2.9469e-005 0.0011549 0.20067 0.00065901 0.20133 0.18496 0 0.033985 0.0389 0 0.99669 0.29453 0.083104 0.011273 4.9137 0.070345 8.5709e-005 0.81974 0.0058631 0.0066173 0.0016852 0.98292 0.98372 3.6781e-006 1.4713e-005 0.13673 0.68718 0.75536 0.001548 0.75066 0.48016 0.0020795 0.42281 1.2679 1.2636 16.0035 144.9729 0.00041501 -84.4799 0.13995
2.244 0.98804 5.5114e-005 3.8182 0.01202 2.9482e-005 0.0011549 0.2007 0.00065901 0.20135 0.18498 0 0.033984 0.0389 0 0.99679 0.29457 0.083119 0.011275 4.9146 0.070356 8.5724e-005 0.81973 0.0058638 0.006618 0.0016828 0.98295 0.98406 3.6724e-006 1.469e-005 0.13673 0.6881 0.75618 0.0015468 0.75208 0.48033 0.002078 0.42282 1.2699 1.2656 16.0036 144.973 0.00041381 -84.4887 0.14095
2.245 0.98804 5.5114e-005 3.8182 0.01202 2.9495e-005 0.001155 0.20073 0.00065901 0.20138 0.18501 0 0.033982 0.0389 0 0.99688 0.29461 0.083135 0.011276 4.9154 0.070367 8.5739e-005 0.81972 0.0058644 0.0066187 0.0016803 0.98299 0.98438 3.6667e-006 1.4668e-005 0.13674 0.68901 0.75699 0.0015456 0.75349 0.48051 0.0020764 0.42282 1.2719 1.2676 16.0037 144.973 0.00041262 -84.4974 0.14195
2.246 0.98804 5.5114e-005 3.8182 0.01202 2.9508e-005 0.001155 0.20076 0.00065901 0.20141 0.18504 0 0.033981 0.0389 0 0.99698 0.29466 0.08315 0.011278 4.9162 0.070378 8.5753e-005 0.81971 0.0058651 0.0066193 0.0016779 0.98302 0.98468 3.6611e-006 1.4645e-005 0.13674 0.68993 0.7578 0.0015444 0.75489 0.48068 0.0020749 0.42282 1.2739 1.2696 16.0037 144.973 0.00041142 -84.5061 0.14295
2.247 0.98804 5.5114e-005 3.8182 0.01202 2.9522e-005 0.001155 0.20078 0.00065901 0.20144 0.18506 0 0.033979 0.0389 0 0.99707 0.2947 0.083166 0.01128 4.9171 0.07039 8.5768e-005 0.8197 0.0058657 0.00662 0.0016755 0.98306 0.98496 3.6555e-006 1.4623e-005 0.13675 0.69084 0.7586 0.0015432 0.75629 0.48085 0.0020734 0.42282 1.2758 1.2715 16.0038 144.973 0.00041024 -84.5147 0.14395
2.248 0.98804 5.5114e-005 3.8182 0.01202 2.9535e-005 0.001155 0.20081 0.00065901 0.20146 0.18509 0 0.033978 0.0389 0 0.99717 0.29474 0.083181 0.011282 4.9179 0.070401 8.5783e-005 0.81969 0.0058664 0.0066207 0.0016731 0.98309 0.98523 3.65e-006 1.4601e-005 0.13675 0.69174 0.7594 0.0015421 0.75769 0.48103 0.0020718 0.42282 1.2778 1.2735 16.0038 144.973 0.00040906 -84.5232 0.14495
2.249 0.98804 5.5114e-005 3.8182 0.012019 2.9548e-005 0.001155 0.20084 0.00065901 0.20149 0.18511 0 0.033976 0.0389 0 0.99726 0.29479 0.083197 0.011283 4.9188 0.070412 8.5798e-005 0.81967 0.005867 0.0066214 0.0016707 0.98312 0.98548 3.6446e-006 1.4579e-005 0.13676 0.69265 0.76019 0.0015409 0.75907 0.4812 0.0020704 0.42283 1.2798 1.2755 16.0039 144.973 0.00040789 -84.5317 0.14595
2.25 0.98804 5.5114e-005 3.8182 0.012019 2.9561e-005 0.001155 0.20087 0.00065901 0.20152 0.18514 0 0.033975 0.0389 0 0.99736 0.29483 0.083212 0.011285 4.9196 0.070423 8.5812e-005 0.81966 0.0058677 0.0066221 0.0016684 0.98316 0.98572 3.6392e-006 1.4557e-005 0.13676 0.69355 0.76098 0.0015398 0.76045 0.48138 0.0020689 0.42283 1.2817 1.2775 16.004 144.973 0.00040673 -84.5401 0.14695
2.251 0.98804 5.5114e-005 3.8182 0.012019 2.9574e-005 0.001155 0.20089 0.00065901 0.20155 0.18517 0 0.033973 0.0389 0 0.99746 0.29487 0.083228 0.011287 4.9205 0.070434 8.5827e-005 0.81965 0.0058684 0.0066228 0.001666 0.98319 0.98595 3.6338e-006 1.4536e-005 0.13677 0.69445 0.76176 0.0015387 0.76182 0.48155 0.0020674 0.42283 1.2837 1.2794 16.004 144.973 0.00040557 -84.5484 0.14795
2.252 0.98804 5.5114e-005 3.8182 0.012019 2.9587e-005 0.001155 0.20092 0.00065901 0.20158 0.18519 0 0.033972 0.0389 0 0.99755 0.29492 0.083243 0.011289 4.9213 0.070445 8.5842e-005 0.81964 0.005869 0.0066235 0.0016638 0.98322 0.98617 3.6285e-006 1.4515e-005 0.13678 0.69535 0.76254 0.0015376 0.76319 0.48172 0.002066 0.42284 1.2856 1.2814 16.0041 144.973 0.00040441 -84.5567 0.14895
2.253 0.98804 5.5114e-005 3.8182 0.012019 2.96e-005 0.001155 0.20095 0.00065901 0.2016 0.18522 0 0.03397 0.0389 0 0.99765 0.29496 0.083259 0.011291 4.9222 0.070456 8.5857e-005 0.81963 0.0058697 0.0066241 0.0016615 0.98325 0.98637 3.6232e-006 1.4493e-005 0.13678 0.69624 0.76331 0.0015365 0.76454 0.4819 0.0020645 0.42284 1.2876 1.2834 16.0041 144.9731 0.00040327 -84.5649 0.14995
2.254 0.98804 5.5114e-005 3.8182 0.012019 2.9613e-005 0.001155 0.20098 0.00065901 0.20163 0.18525 0 0.033969 0.0389 0 0.99774 0.295 0.083274 0.011292 4.923 0.070468 8.5871e-005 0.81962 0.0058703 0.0066248 0.0016593 0.98328 0.98656 3.618e-006 1.4473e-005 0.13679 0.69713 0.76408 0.0015354 0.7659 0.48207 0.0020631 0.42284 1.2895 1.2853 16.0042 144.9731 0.00040212 -84.573 0.15095
2.255 0.98804 5.5114e-005 3.8182 0.012019 2.9626e-005 0.001155 0.201 0.00065901 0.20166 0.18527 0 0.033967 0.0389 0 0.99784 0.29505 0.08329 0.011294 4.9239 0.070479 8.5886e-005 0.81961 0.005871 0.0066255 0.0016571 0.98331 0.98674 3.6128e-006 1.4452e-005 0.13679 0.69802 0.76484 0.0015344 0.76724 0.48225 0.0020617 0.42284 1.2914 1.2873 16.0043 144.9731 0.00040099 -84.5811 0.15195
2.256 0.98804 5.5114e-005 3.8182 0.012019 2.9639e-005 0.001155 0.20103 0.00065901 0.20169 0.1853 0 0.033966 0.0389 0 0.99793 0.29509 0.083305 0.011296 4.9247 0.07049 8.5901e-005 0.8196 0.0058717 0.0066262 0.0016549 0.98334 0.98691 3.6077e-006 1.4431e-005 0.1368 0.69891 0.7656 0.0015333 0.76858 0.48242 0.0020603 0.42285 1.2934 1.2892 16.0043 144.9731 0.00039986 -84.5891 0.15295
2.257 0.98804 5.5114e-005 3.8182 0.012019 2.9652e-005 0.001155 0.20106 0.00065901 0.20171 0.18532 0 0.033964 0.0389 0 0.99803 0.29513 0.083321 0.011298 4.9256 0.070501 8.5916e-005 0.81958 0.0058723 0.0066269 0.0016527 0.98338 0.98708 3.6026e-006 1.4411e-005 0.1368 0.69979 0.76635 0.0015322 0.76991 0.48259 0.0020589 0.42285 1.2953 1.2911 16.0044 144.9731 0.00039873 -84.5971 0.15395
2.258 0.98804 5.5114e-005 3.8182 0.012019 2.9666e-005 0.001155 0.20109 0.00065901 0.20174 0.18535 0 0.033963 0.0389 0 0.99812 0.29518 0.083336 0.0113 4.9264 0.070512 8.593e-005 0.81957 0.005873 0.0066276 0.0016506 0.98341 0.98723 3.5976e-006 1.4391e-005 0.13681 0.70067 0.7671 0.0015311 0.77123 0.48277 0.0020575 0.42286 1.2972 1.2931 16.0044 144.9731 0.00039762 -84.605 0.15495
2.259 0.98804 5.5113e-005 3.8182 0.012019 2.9679e-005 0.001155 0.20111 0.00065901 0.20177 0.18538 0 0.033961 0.0389 0 0.99822 0.29522 0.083352 0.011301 4.9272 0.070523 8.5945e-005 0.81956 0.0058736 0.0066283 0.0016484 0.98343 0.98738 3.5926e-006 1.4371e-005 0.13681 0.70155 0.76784 0.0015301 0.77255 0.48294 0.0020561 0.42286 1.2991 1.295 16.0045 144.9731 0.0003965 -84.6128 0.15595
2.26 0.98804 5.5113e-005 3.8182 0.012019 2.9692e-005 0.001155 0.20114 0.00065901 0.2018 0.1854 0 0.03396 0.0389 0 0.99831 0.29526 0.083367 0.011303 4.9281 0.070535 8.596e-005 0.81955 0.0058743 0.006629 0.0016463 0.98346 0.98752 3.5877e-006 1.4351e-005 0.13682 0.70242 0.76858 0.001529 0.77386 0.48312 0.0020548 0.42286 1.301 1.2969 16.0045 144.9731 0.0003954 -84.6205 0.15695
2.261 0.98804 5.5113e-005 3.8182 0.012019 2.9705e-005 0.001155 0.20117 0.00065901 0.20182 0.18543 0 0.033958 0.0389 0 0.99841 0.29531 0.083383 0.011305 4.9289 0.070546 8.5975e-005 0.81954 0.005875 0.0066297 0.0016442 0.98349 0.98765 3.5828e-006 1.4332e-005 0.13682 0.70329 0.76932 0.001528 0.77517 0.48329 0.0020534 0.42287 1.3029 1.2989 16.0046 144.9732 0.00039429 -84.6282 0.15795
2.262 0.98804 5.5113e-005 3.8182 0.012019 2.9718e-005 0.001155 0.2012 0.00065901 0.20185 0.18545 0 0.033957 0.0389 0 0.99851 0.29535 0.083398 0.011307 4.9298 0.070557 8.5989e-005 0.81953 0.0058756 0.0066303 0.0016421 0.98352 0.98777 3.578e-006 1.4312e-005 0.13683 0.70416 0.77005 0.0015269 0.77647 0.48346 0.0020521 0.42287 1.3048 1.3008 16.0046 144.9732 0.0003932 -84.6359 0.15895
2.263 0.98804 5.5113e-005 3.8182 0.012019 2.9731e-005 0.001155 0.20122 0.00065901 0.20188 0.18548 0 0.033955 0.0389 0 0.9986 0.29539 0.083414 0.011308 4.9306 0.070568 8.6004e-005 0.81952 0.0058763 0.006631 0.0016399 0.98355 0.98789 3.5732e-006 1.4293e-005 0.13683 0.70503 0.77078 0.0015259 0.77776 0.48364 0.0020508 0.42287 1.3067 1.3027 16.0047 144.9732 0.00039211 -84.6435 0.15995
2.264 0.98804 5.5113e-005 3.8182 0.012019 2.9744e-005 0.001155 0.20125 0.00065901 0.20191 0.1855 0 0.033954 0.0389 0 0.9987 0.29544 0.083429 0.01131 4.9315 0.070579 8.6019e-005 0.81951 0.0058769 0.0066317 0.0016379 0.98358 0.988 3.5684e-006 1.4274e-005 0.13684 0.70589 0.7715 0.0015249 0.77904 0.48381 0.0020494 0.42288 1.3086 1.3046 16.0047 144.9732 0.00039103 -84.651 0.16095
2.265 0.98804 5.5113e-005 3.8182 0.012019 2.9757e-005 0.001155 0.20128 0.00065901 0.20193 0.18553 0 0.033952 0.0389 0 0.99879 0.29548 0.083444 0.011312 4.9323 0.07059 8.6034e-005 0.8195 0.0058776 0.0066324 0.0016358 0.98361 0.98811 3.5637e-006 1.4255e-005 0.13685 0.70675 0.77222 0.0015239 0.78032 0.48399 0.0020481 0.42288 1.3105 1.3065 16.0048 144.9732 0.00038995 -84.6584 0.16195
2.266 0.98804 5.5113e-005 3.8182 0.012019 2.977e-005 0.001155 0.20131 0.00065901 0.20196 0.18556 0 0.033951 0.0389 0 0.99889 0.29552 0.08346 0.011314 4.9332 0.070601 8.6048e-005 0.81948 0.0058783 0.0066331 0.0016338 0.98364 0.98821 3.5591e-006 1.4237e-005 0.13685 0.70761 0.77293 0.0015229 0.78159 0.48416 0.0020468 0.42289 1.3124 1.3084 16.0048 144.9732 0.00038887 -84.6658 0.16295
2.267 0.98804 5.5113e-005 3.8182 0.012019 2.9783e-005 0.001155 0.20133 0.00065901 0.20199 0.18558 0 0.033949 0.0389 0 0.99898 0.29557 0.083475 0.011316 4.9341 0.070613 8.6063e-005 0.81947 0.0058789 0.0066338 0.0016318 0.98366 0.98831 3.5545e-006 1.4218e-005 0.13686 0.70847 0.77364 0.001522 0.78286 0.48433 0.0020456 0.42289 1.3143 1.3103 16.0049 144.9732 0.0003878 -84.6732 0.16395
2.268 0.98804 5.5113e-005 3.8182 0.012019 2.9796e-005 0.001155 0.20136 0.00065901 0.20202 0.18561 0 0.033948 0.0389 0 0.99908 0.29561 0.083491 0.011317 4.9349 0.070624 8.6078e-005 0.81946 0.0058796 0.0066345 0.0016298 0.98369 0.9884 3.5499e-006 1.42e-005 0.13686 0.70932 0.77434 0.0015211 0.78412 0.48451 0.0020443 0.42289 1.3162 1.3122 16.005 144.9732 0.00038674 -84.6805 0.16495
2.269 0.98804 5.5113e-005 3.8182 0.012019 2.9809e-005 0.001155 0.20139 0.00065901 0.20204 0.18563 0 0.033946 0.0389 0 0.99917 0.29565 0.083506 0.011319 4.9358 0.070635 8.6093e-005 0.81945 0.0058802 0.0066352 0.0016279 0.98372 0.98848 3.5454e-006 1.4182e-005 0.13687 0.71017 0.77505 0.0015201 0.78537 0.48468 0.002043 0.4229 1.3181 1.3141 16.005 144.9733 0.00038569 -84.6877 0.16595
2.27 0.98804 5.5113e-005 3.8182 0.012019 2.9823e-005 0.001155 0.20142 0.00065901 0.20207 0.18566 0 0.033945 0.0389 0 0.99927 0.29569 0.083522 0.011321 4.9366 0.070646 8.6107e-005 0.81944 0.0058809 0.0066359 0.001626 0.98374 0.98857 3.5408e-006 1.4164e-005 0.13687 0.71102 0.77574 0.0015192 0.78662 0.48485 0.0020418 0.4229 1.3199 1.316 16.0051 144.9733 0.00038463 -84.6949 0.16695
2.271 0.98804 5.5113e-005 3.8182 0.012019 2.9836e-005 0.001155 0.20144 0.00065901 0.2021 0.18569 0 0.033943 0.0389 0 0.99937 0.29574 0.083537 0.011323 4.9375 0.070657 8.6122e-005 0.81943 0.0058816 0.0066365 0.0016241 0.98377 0.98864 3.5364e-006 1.4146e-005 0.13688 0.71187 0.77643 0.0015183 0.78786 0.48503 0.0020406 0.42291 1.3218 1.3179 16.0051 144.9733 0.00038359 -84.702 0.16795
2.272 0.98804 5.5113e-005 3.8182 0.012019 2.9849e-005 0.001155 0.20147 0.00065902 0.20212 0.18571 0 0.033942 0.0389 0 0.99946 0.29578 0.083553 0.011324 4.9383 0.070668 8.6137e-005 0.81942 0.0058822 0.0066372 0.0016222 0.9838 0.98872 3.5319e-006 1.4128e-005 0.13688 0.71271 0.77712 0.0015173 0.78909 0.4852 0.0020393 0.42291 1.3237 1.3197 16.0052 144.9733 0.00038255 -84.7091 0.16895
2.273 0.98804 5.5113e-005 3.8182 0.012019 2.9862e-005 0.001155 0.2015 0.00065902 0.20215 0.18574 0 0.03394 0.0389 0 0.99956 0.29582 0.083568 0.011326 4.9392 0.070679 8.6152e-005 0.81941 0.0058829 0.0066379 0.0016204 0.98382 0.98879 3.5275e-006 1.4111e-005 0.13689 0.71355 0.77781 0.0015164 0.79032 0.48538 0.0020381 0.42292 1.3255 1.3216 16.0052 144.9733 0.00038151 -84.7161 0.16995
2.274 0.98804 5.5112e-005 3.8182 0.012019 2.9875e-005 0.001155 0.20152 0.00065902 0.20218 0.18576 0 0.033939 0.0389 0 0.99965 0.29587 0.083584 0.011328 4.94 0.070691 8.6167e-005 0.8194 0.0058835 0.0066386 0.0016185 0.98385 0.98886 3.5232e-006 1.4093e-005 0.13689 0.71439 0.77849 0.0015154 0.79154 0.48555 0.0020369 0.42292 1.3274 1.3235 16.0053 144.9733 0.00038048 -84.723 0.17095
2.275 0.98804 5.5112e-005 3.8182 0.012019 2.9888e-005 0.001155 0.20155 0.00065902 0.20221 0.18579 0 0.033937 0.0389 0 0.99975 0.29591 0.083599 0.01133 4.9409 0.070702 8.6181e-005 0.81938 0.0058842 0.0066393 0.0016167 0.98388 0.98892 3.5189e-006 1.4076e-005 0.1369 0.71523 0.77916 0.0015145 0.79275 0.48572 0.0020357 0.42293 1.3292 1.3253 16.0053 144.9733 0.00037945 -84.7299 0.17195
2.276 0.98804 5.5112e-005 3.8182 0.012019 2.9901e-005 0.001155 0.20158 0.00065902 0.20223 0.18581 0 0.033936 0.0389 0 0.99984 0.29595 0.083615 0.011332 4.9417 0.070713 8.6196e-005 0.81937 0.0058849 0.00664 0.0016149 0.9839 0.98898 3.5146e-006 1.4059e-005 0.13691 0.71606 0.77984 0.0015136 0.79396 0.4859 0.0020345 0.42293 1.3311 1.3272 16.0054 144.9733 0.00037843 -84.7368 0.17295
2.277 0.98804 5.5112e-005 3.8182 0.012019 2.9914e-005 0.001155 0.20161 0.00065902 0.20226 0.18584 0 0.033934 0.0389 0 0.99994 0.296 0.08363 0.011333 4.9426 0.070724 8.6211e-005 0.81936 0.0058855 0.0066407 0.001613 0.98393 0.98904 3.5104e-006 1.4042e-005 0.13691 0.71689 0.78051 0.0015126 0.79516 0.48607 0.0020333 0.42294 1.3329 1.3291 16.0054 144.9734 0.00037742 -84.7436 0.17395
2.278 0.98804 5.5112e-005 3.8182 0.012019 2.9927e-005 0.001155 0.20163 0.00065902 0.20229 0.18587 0 0.033933 0.0389 0 1 0.29604 0.083646 0.011335 4.9435 0.070735 8.6226e-005 0.81935 0.0058862 0.0066414 0.0016111 0.98395 0.9891 3.5062e-006 1.4025e-005 0.13692 0.71772 0.78117 0.0015117 0.79636 0.48624 0.0020322 0.42294 1.3347 1.3309 16.0055 144.9734 0.00037641 -84.7503 0.17495
2.279 0.98804 5.5112e-005 3.8182 0.012019 2.994e-005 0.001155 0.20166 0.00065902 0.20231 0.18589 0 0.033931 0.0389 0 1.0001 0.29608 0.083661 0.011337 4.9443 0.070746 8.624e-005 0.81934 0.0058869 0.0066421 0.0016092 0.98398 0.98915 3.5021e-006 1.4009e-005 0.13692 0.71854 0.78183 0.0015107 0.79755 0.48642 0.002031 0.42295 1.3366 1.3327 16.0055 144.9734 0.00037541 -84.757 0.17595
2.28 0.98804 5.5112e-005 3.8182 0.012019 2.9953e-005 0.001155 0.20169 0.00065902 0.20234 0.18592 0 0.03393 0.0389 0 1.0002 0.29613 0.083677 0.011339 4.9452 0.070758 8.6255e-005 0.81933 0.0058875 0.0066428 0.0016074 0.984 0.9892 3.498e-006 1.3992e-005 0.13693 0.71936 0.78249 0.0015098 0.79873 0.48659 0.0020299 0.42295 1.3384 1.3346 16.0055 144.9734 0.00037441 -84.7637 0.17695
2.281 0.98804 5.5112e-005 3.8182 0.012019 2.9967e-005 0.001155 0.20171 0.00065902 0.20237 0.18594 0 0.033928 0.0389 0 1.0003 0.29617 0.083693 0.011341 4.946 0.070769 8.627e-005 0.81932 0.0058882 0.0066435 0.0016056 0.98402 0.98925 3.4939e-006 1.3976e-005 0.13693 0.72018 0.78314 0.001509 0.79991 0.48676 0.0020287 0.42296 1.3402 1.3364 16.0056 144.9734 0.00037341 -84.7702 0.17795
2.282 0.98804 5.5112e-005 3.8182 0.012019 2.998e-005 0.001155 0.20174 0.00065902 0.20239 0.18597 0 0.033927 0.0389 0 1.0004 0.29622 0.083708 0.011342 4.9469 0.07078 8.6285e-005 0.81931 0.0058888 0.0066442 0.0016038 0.98405 0.9893 3.4899e-006 1.396e-005 0.13694 0.721 0.78379 0.0015082 0.80108 0.48694 0.0020276 0.42296 1.342 1.3383 16.0056 144.9734 0.00037242 -84.7768 0.17895
2.283 0.98804 5.5112e-005 3.8182 0.012019 2.9993e-005 0.001155 0.20177 0.00065902 0.20242 0.18599 0 0.033925 0.0389 0 1.0005 0.29626 0.083724 0.011344 4.9477 0.070791 8.6299e-005 0.8193 0.0058895 0.0066448 0.001602 0.98407 0.98934 3.4859e-006 1.3944e-005 0.13694 0.72182 0.78444 0.0015074 0.80224 0.48711 0.0020265 0.42297 1.3439 1.3401 16.0057 144.9734 0.00037144 -84.7833 0.17995
2.284 0.98804 5.5112e-005 3.8182 0.012019 3.0006e-005 0.001155 0.20179 0.00065902 0.20245 0.18602 0 0.033924 0.0389 0 1.0006 0.2963 0.083739 0.011346 4.9486 0.070802 8.6314e-005 0.81928 0.0058902 0.0066455 0.0016003 0.9841 0.98939 3.482e-006 1.3928e-005 0.13695 0.72263 0.78508 0.0015065 0.8034 0.48729 0.0020254 0.42297 1.3457 1.3419 16.0057 144.9735 0.00037046 -84.7897 0.18095
2.285 0.98804 5.5112e-005 3.8182 0.012019 3.0019e-005 0.001155 0.20182 0.00065902 0.20248 0.18604 0 0.033922 0.0389 0 1.0007 0.29635 0.083755 0.011348 4.9495 0.070813 8.6329e-005 0.81927 0.0058908 0.0066462 0.0015986 0.98412 0.98943 3.478e-006 1.3912e-005 0.13695 0.72344 0.78572 0.0015057 0.80455 0.48746 0.0020243 0.42298 1.3475 1.3437 16.0058 144.9735 0.00036948 -84.7961 0.18195
2.286 0.98804 5.5112e-005 3.8182 0.012019 3.0032e-005 0.001155 0.20185 0.00065902 0.2025 0.18607 0 0.033921 0.0389 0 1.0008 0.29639 0.08377 0.011349 4.9503 0.070824 8.6344e-005 0.81926 0.0058915 0.0066469 0.001597 0.98414 0.98947 3.4741e-006 1.3897e-005 0.13696 0.72425 0.78635 0.0015049 0.8057 0.48763 0.0020232 0.42298 1.3493 1.3456 16.0058 144.9735 0.00036851 -84.8024 0.18295
2.287 0.98804 5.5112e-005 3.8182 0.012019 3.0045e-005 0.001155 0.20187 0.00065902 0.20253 0.18609 0 0.033919 0.0389 0 1.0009 0.29643 0.083786 0.011351 4.9512 0.070836 8.6359e-005 0.81925 0.0058922 0.0066476 0.0015954 0.98416 0.9895 3.4702e-006 1.3881e-005 0.13697 0.72505 0.78698 0.0015042 0.80684 0.48781 0.0020221 0.42299 1.3511 1.3474 16.0059 144.9735 0.00036755 -84.8087 0.18395
2.288 0.98804 5.5112e-005 3.8182 0.012019 3.0058e-005 0.001155 0.2019 0.00065902 0.20256 0.18612 0 0.033918 0.0389 0 1.001 0.29648 0.083801 0.011353 4.952 0.070847 8.6373e-005 0.81924 0.0058928 0.0066483 0.0015938 0.98419 0.98954 3.4664e-006 1.3866e-005 0.13697 0.72586 0.78761 0.0015034 0.80797 0.48798 0.002021 0.423 1.3529 1.3492 16.0059 144.9735 0.00036659 -84.815 0.18495
2.289 0.98804 5.5111e-005 3.8182 0.012019 3.0071e-005 0.001155 0.20193 0.00065902 0.20258 0.18615 0 0.033917 0.0389 0 1.0011 0.29652 0.083817 0.011355 4.9529 0.070858 8.6388e-005 0.81923 0.0058935 0.006649 0.0015922 0.98421 0.98958 3.4626e-006 1.3851e-005 0.13698 0.72666 0.78824 0.0015026 0.8091 0.48815 0.00202 0.423 1.3547 1.351 16.006 144.9735 0.00036563 -84.8212 0.18595
2.29 0.98804 5.5111e-005 3.8182 0.012019 3.0084e-005 0.001155 0.20196 0.00065902 0.20261 0.18617 0 0.033915 0.0389 0 1.0012 0.29656 0.083832 0.011357 4.9538 0.070869 8.6403e-005 0.81922 0.0058941 0.0066497 0.0015907 0.98423 0.98961 3.4588e-006 1.3836e-005 0.13698 0.72745 0.78886 0.0015018 0.81022 0.48833 0.0020189 0.42301 1.3564 1.3528 16.006 144.9735 0.00036468 -84.8273 0.18695
2.291 0.98804 5.5111e-005 3.8182 0.012019 3.0097e-005 0.001155 0.20198 0.00065902 0.20264 0.1862 0 0.033914 0.0389 0 1.0013 0.29661 0.083848 0.011358 4.9546 0.07088 8.6418e-005 0.81921 0.0058948 0.0066504 0.0015891 0.98425 0.98964 3.455e-006 1.3821e-005 0.13699 0.72825 0.78947 0.0015009 0.81134 0.4885 0.0020179 0.42301 1.3582 1.3546 16.006 144.9736 0.00036373 -84.8334 0.18795
2.292 0.98804 5.5111e-005 3.8182 0.012019 3.011e-005 0.001155 0.20201 0.00065902 0.20266 0.18622 0 0.033912 0.0389 0 1.0014 0.29665 0.083863 0.01136 4.9555 0.070891 8.6432e-005 0.81919 0.0058955 0.0066511 0.0015875 0.98428 0.98967 3.4513e-006 1.3806e-005 0.13699 0.72904 0.79009 0.0015001 0.81245 0.48867 0.0020168 0.42302 1.36 1.3564 16.0061 144.9736 0.00036279 -84.8395 0.18895
2.293 0.98804 5.5111e-005 3.8182 0.012019 3.0124e-005 0.001155 0.20204 0.00065902 0.20269 0.18625 0 0.033911 0.0389 0 1.0015 0.29669 0.083879 0.011362 4.9564 0.070903 8.6447e-005 0.81918 0.0058961 0.0066518 0.0015859 0.9843 0.9897 3.4477e-006 1.3791e-005 0.137 0.72983 0.7907 0.0014992 0.81355 0.48885 0.0020158 0.42303 1.3618 1.3581 16.0061 144.9736 0.00036186 -84.8455 0.18995
2.294 0.98804 5.5111e-005 3.8182 0.012019 3.0137e-005 0.001155 0.20206 0.00065902 0.20272 0.18627 0 0.033909 0.0389 0 1.0016 0.29674 0.083894 0.011364 4.9572 0.070914 8.6462e-005 0.81917 0.0058968 0.0066525 0.0015843 0.98432 0.98973 3.444e-006 1.3777e-005 0.137 0.73062 0.79131 0.0014984 0.81465 0.48902 0.0020148 0.42303 1.3635 1.3599 16.0062 144.9736 0.00036092 -84.8514 0.19095
2.295 0.98804 5.5111e-005 3.8182 0.012019 3.015e-005 0.001155 0.20209 0.00065902 0.20274 0.1863 0 0.033908 0.0389 0 1.0017 0.29678 0.08391 0.011366 4.9581 0.070925 8.6477e-005 0.81916 0.0058975 0.0066532 0.0015827 0.98434 0.98976 3.4404e-006 1.3762e-005 0.13701 0.73141 0.79191 0.0014976 0.81574 0.48919 0.0020138 0.42304 1.3653 1.3617 16.0062 144.9736 0.00036 -84.8573 0.19195
2.296 0.98804 5.5111e-005 3.8182 0.012019 3.0163e-005 0.001155 0.20212 0.00065902 0.20277 0.18632 0 0.033906 0.0389 0 1.0018 0.29682 0.083925 0.011367 4.959 0.070936 8.6492e-005 0.81915 0.0058981 0.0066539 0.0015811 0.98436 0.98979 3.4369e-006 1.3748e-005 0.13701 0.73219 0.79251 0.0014968 0.81683 0.48937 0.0020128 0.42304 1.3671 1.3635 16.0063 144.9736 0.00035907 -84.8632 0.19295
2.297 0.98804 5.5111e-005 3.8182 0.012019 3.0176e-005 0.001155 0.20214 0.00065902 0.2028 0.18635 0 0.033905 0.0389 0 1.0019 0.29687 0.083941 0.011369 4.9598 0.070947 8.6506e-005 0.81914 0.0058988 0.0066546 0.0015795 0.98438 0.98981 3.4334e-006 1.3734e-005 0.13702 0.73297 0.79311 0.001496 0.81791 0.48954 0.0020118 0.42305 1.3688 1.3652 16.0063 144.9736 0.00035816 -84.869 0.19395
2.298 0.98804 5.5111e-005 3.8182 0.012019 3.0189e-005 0.001155 0.20217 0.00065902 0.20282 0.18637 0 0.033903 0.0389 0 1.0019 0.29691 0.083956 0.011371 4.9607 0.070958 8.6521e-005 0.81913 0.0058995 0.0066552 0.0015779 0.9844 0.98984 3.4299e-006 1.372e-005 0.13703 0.73375 0.7937 0.0014952 0.81899 0.48971 0.0020108 0.42306 1.3706 1.367 16.0063 144.9737 0.00035724 -84.8748 0.19495
2.299 0.98804 5.5111e-005 3.8182 0.012019 3.0202e-005 0.001155 0.2022 0.00065902 0.20285 0.1864 0 0.033902 0.0389 0 1.002 0.29695 0.083972 0.011373 4.9615 0.07097 8.6536e-005 0.81912 0.0059001 0.0066559 0.0015763 0.98442 0.98986 3.4264e-006 1.3706e-005 0.13703 0.73452 0.79429 0.0014945 0.82005 0.48989 0.0020098 0.42306 1.3723 1.3688 16.0064 144.9737 0.00035633 -84.8806 0.19595
2.3 0.98804 5.5111e-005 3.8182 0.012019 3.0215e-005 0.001155 0.20222 0.00065902 0.20288 0.18642 0 0.0339 0.0389 0 1.0021 0.297 0.083987 0.011374 4.9624 0.070981 8.6551e-005 0.81911 0.0059008 0.0066566 0.0015748 0.98444 0.98989 3.423e-006 1.3692e-005 0.13704 0.7353 0.79488 0.0014938 0.82112 0.49006 0.0020088 0.42307 1.3741 1.3705 16.0064 144.9737 0.00035543 -84.8863 0.19695
2.301 0.98804 5.5111e-005 3.8182 0.012019 3.0228e-005 0.001155 0.20225 0.00065902 0.2029 0.18645 0 0.033899 0.0389 0 1.0022 0.29704 0.084003 0.011376 4.9633 0.070992 8.6565e-005 0.81909 0.0059015 0.0066573 0.0015733 0.98446 0.98991 3.4195e-006 1.3678e-005 0.13704 0.73607 0.79546 0.0014931 0.82218 0.49023 0.0020078 0.42308 1.3758 1.3723 16.0065 144.9737 0.00035453 -84.8919 0.19795
2.302 0.98804 5.5111e-005 3.8182 0.012019 3.0241e-005 0.001155 0.20228 0.00065902 0.20293 0.18647 0 0.033898 0.0389 0 1.0023 0.29708 0.084019 0.011378 4.9642 0.071003 8.658e-005 0.81908 0.0059021 0.006658 0.0015719 0.98448 0.98993 3.4161e-006 1.3665e-005 0.13705 0.73684 0.79604 0.0014924 0.82323 0.4904 0.0020069 0.42308 1.3775 1.374 16.0065 144.9737 0.00035363 -84.8975 0.19895
2.303 0.98804 5.5111e-005 3.8182 0.012019 3.0254e-005 0.001155 0.2023 0.00065902 0.20296 0.1865 0 0.033896 0.0389 0 1.0024 0.29713 0.084034 0.01138 4.965 0.071014 8.6595e-005 0.81907 0.0059028 0.0066587 0.0015705 0.9845 0.98996 3.4128e-006 1.3651e-005 0.13705 0.7376 0.79662 0.0014918 0.82427 0.49058 0.0020059 0.42309 1.3793 1.3758 16.0065 144.9737 0.00035274 -84.9031 0.19995
2.304 0.98804 5.511e-005 3.8182 0.012019 3.0268e-005 0.001155 0.20233 0.00065902 0.20298 0.18652 0 0.033895 0.0389 0 1.0025 0.29717 0.08405 0.011382 4.9659 0.071025 8.661e-005 0.81906 0.0059035 0.0066594 0.0015691 0.98452 0.98998 3.4094e-006 1.3638e-005 0.13706 0.73837 0.79719 0.0014911 0.82531 0.49075 0.002005 0.4231 1.381 1.3775 16.0066 144.9737 0.00035185 -84.9086 0.20095
2.305 0.98804 5.511e-005 3.8182 0.012019 3.0281e-005 0.001155 0.20236 0.00065902 0.20301 0.18655 0 0.033893 0.0389 0 1.0026 0.29721 0.084065 0.011383 4.9668 0.071037 8.6625e-005 0.81905 0.0059041 0.0066601 0.0015677 0.98454 0.99 3.4061e-006 1.3625e-005 0.13706 0.73913 0.79777 0.0014904 0.82635 0.49092 0.0020041 0.4231 1.3827 1.3792 16.0066 144.9738 0.00035097 -84.9141 0.20195
2.306 0.98804 5.511e-005 3.8182 0.012019 3.0294e-005 0.001155 0.20238 0.00065902 0.20304 0.18657 0 0.033892 0.0389 0 1.0027 0.29726 0.084081 0.011385 4.9676 0.071048 8.6639e-005 0.81904 0.0059048 0.0066608 0.0015664 0.98456 0.99002 3.4028e-006 1.3612e-005 0.13707 0.73989 0.79833 0.0014897 0.82738 0.4911 0.0020031 0.42311 1.3844 1.381 16.0067 144.9738 0.00035009 -84.9195 0.20295
2.307 0.98804 5.511e-005 3.8182 0.012019 3.0307e-005 0.001155 0.20241 0.00065903 0.20306 0.1866 0 0.03389 0.0389 0 1.0028 0.2973 0.084096 0.011387 4.9685 0.071059 8.6654e-005 0.81903 0.0059054 0.0066615 0.001565 0.98458 0.99004 3.3995e-006 1.3599e-005 0.13707 0.74065 0.7989 0.001489 0.8284 0.49127 0.0020022 0.42312 1.3862 1.3827 16.0067 144.9738 0.00034922 -84.9249 0.20395
2.308 0.98804 5.511e-005 3.8182 0.012019 3.032e-005 0.001155 0.20243 0.00065903 0.20309 0.18662 0 0.033889 0.0389 0 1.0029 0.29734 0.084112 0.011389 4.9694 0.07107 8.6669e-005 0.81902 0.0059061 0.0066622 0.0015637 0.9846 0.99005 3.3963e-006 1.3586e-005 0.13708 0.7414 0.79946 0.0014883 0.82942 0.49144 0.0020013 0.42313 1.3879 1.3844 16.0067 144.9738 0.00034835 -84.9303 0.20495
2.309 0.98804 5.511e-005 3.8182 0.012019 3.0333e-005 0.001155 0.20246 0.00065903 0.20312 0.18665 0 0.033887 0.0389 0 1.003 0.29739 0.084127 0.01139 4.9702 0.071081 8.6684e-005 0.81901 0.0059068 0.0066629 0.0015624 0.98462 0.99007 3.3931e-006 1.3573e-005 0.13709 0.74215 0.80002 0.0014876 0.83043 0.49162 0.0020004 0.42313 1.3896 1.3861 16.0068 144.9738 0.00034748 -84.9356 0.20595
2.31 0.98804 5.511e-005 3.8182 0.012019 3.0346e-005 0.001155 0.20249 0.00065903 0.20314 0.18667 0 0.033886 0.0389 0 1.0031 0.29743 0.084143 0.011392 4.9711 0.071092 8.6699e-005 0.81899 0.0059074 0.0066636 0.001561 0.98464 0.99009 3.39e-006 1.356e-005 0.13709 0.7429 0.80058 0.0014868 0.83144 0.49179 0.0019995 0.42314 1.3913 1.3879 16.0068 144.9738 0.00034662 -84.9409 0.20695
2.311 0.98804 5.511e-005 3.8182 0.012019 3.0359e-005 0.001155 0.20251 0.00065903 0.20317 0.1867 0 0.033885 0.0389 0 1.0032 0.29747 0.084158 0.011394 4.972 0.071103 8.6713e-005 0.81898 0.0059081 0.0066643 0.0015596 0.98466 0.99011 3.3868e-006 1.3548e-005 0.1371 0.74365 0.80113 0.0014861 0.83244 0.49196 0.0019986 0.42315 1.393 1.3896 16.0069 144.9738 0.00034577 -84.9461 0.20795
2.312 0.98804 5.511e-005 3.8182 0.012019 3.0372e-005 0.001155 0.20254 0.00065903 0.20319 0.18672 0 0.033883 0.0389 0 1.0033 0.29752 0.084174 0.011396 4.9728 0.071115 8.6728e-005 0.81897 0.0059088 0.006665 0.0015582 0.98467 0.99013 3.3837e-006 1.3535e-005 0.1371 0.7444 0.80168 0.0014853 0.83343 0.49213 0.0019977 0.42315 1.3947 1.3913 16.0069 144.9739 0.00034491 -84.9513 0.20895
2.313 0.98804 5.511e-005 3.8182 0.012019 3.0385e-005 0.001155 0.20257 0.00065903 0.20322 0.18675 0 0.033882 0.0389 0 1.0034 0.29756 0.08419 0.011398 4.9737 0.071126 8.6743e-005 0.81896 0.0059094 0.0066657 0.0015567 0.98469 0.99014 3.3807e-006 1.3523e-005 0.13711 0.74514 0.80223 0.0014846 0.83442 0.49231 0.0019968 0.42316 1.3964 1.393 16.0069 144.9739 0.00034407 -84.9565 0.20995
2.314 0.98804 5.511e-005 3.8182 0.012019 3.0398e-005 0.001155 0.20259 0.00065903 0.20325 0.18677 0 0.03388 0.0389 0 1.0035 0.2976 0.084205 0.011399 4.9746 0.071137 8.6758e-005 0.81895 0.0059101 0.0066664 0.0015554 0.98471 0.99016 3.3776e-006 1.3511e-005 0.13711 0.74588 0.80277 0.0014839 0.83541 0.49248 0.001996 0.42317 1.398 1.3947 16.007 144.9739 0.00034322 -84.9616 0.21095
2.315 0.98804 5.511e-005 3.8182 0.012019 3.0411e-005 0.001155 0.20262 0.00065903 0.20327 0.1868 0 0.033879 0.0389 0 1.0036 0.29765 0.084221 0.011401 4.9755 0.071148 8.6773e-005 0.81894 0.0059108 0.0066671 0.001554 0.98473 0.99017 3.3746e-006 1.3499e-005 0.13712 0.74662 0.80331 0.0014832 0.83639 0.49265 0.0019951 0.42318 1.3997 1.3964 16.007 144.9739 0.00034238 -84.9667 0.21195
2.316 0.98804 5.511e-005 3.8182 0.012019 3.0425e-005 0.001155 0.20264 0.00065903 0.2033 0.18682 0 0.033877 0.0389 0 1.0037 0.29769 0.084236 0.011403 4.9763 0.071159 8.6787e-005 0.81893 0.0059114 0.0066678 0.0015527 0.98475 0.99019 3.3716e-006 1.3486e-005 0.13712 0.74736 0.80385 0.0014825 0.83736 0.49282 0.0019943 0.42318 1.4014 1.398 16.007 144.9739 0.00034154 -84.9717 0.21295
2.317 0.98804 5.511e-005 3.8182 0.012019 3.0438e-005 0.001155 0.20267 0.00065903 0.20333 0.18685 0 0.033876 0.0389 0 1.0038 0.29774 0.084252 0.011405 4.9772 0.07117 8.6802e-005 0.81892 0.0059121 0.0066685 0.0015513 0.98476 0.99021 3.3686e-006 1.3475e-005 0.13713 0.74809 0.80439 0.0014819 0.83833 0.493 0.0019934 0.42319 1.4031 1.3997 16.0071 144.9739 0.00034071 -84.9767 0.21395
2.318 0.98804 5.511e-005 3.8182 0.012019 3.0451e-005 0.001155 0.2027 0.00065903 0.20335 0.18687 0 0.033875 0.0389 0 1.0039 0.29778 0.084267 0.011407 4.9781 0.071182 8.6817e-005 0.81891 0.0059128 0.0066692 0.00155 0.98478 0.99022 3.3656e-006 1.3463e-005 0.13713 0.74882 0.80492 0.0014813 0.83929 0.49317 0.0019926 0.4232 1.4047 1.4014 16.0071 144.9739 0.00033988 -84.9817 0.21495
2.319 0.98804 5.5109e-005 3.8182 0.012019 3.0464e-005 0.001155 0.20272 0.00065903 0.20338 0.1869 0 0.033873 0.0389 0 1.004 0.29782 0.084283 0.011408 4.979 0.071193 8.6832e-005 0.81889 0.0059135 0.0066699 0.0015488 0.9848 0.99023 3.3627e-006 1.3451e-005 0.13714 0.74955 0.80545 0.0014807 0.84025 0.49334 0.0019917 0.42321 1.4064 1.4031 16.0071 144.974 0.00033906 -84.9866 0.21595
2.32 0.98804 5.5109e-005 3.8182 0.012018 3.0477e-005 0.001155 0.20275 0.00065903 0.2034 0.18692 0 0.033872 0.0389 0 1.0041 0.29787 0.084298 0.01141 4.9798 0.071204 8.6847e-005 0.81888 0.0059141 0.0066706 0.0015475 0.98481 0.99025 3.3598e-006 1.3439e-005 0.13715 0.75028 0.80598 0.0014801 0.8412 0.49351 0.0019909 0.42321 1.4081 1.4048 16.0072 144.974 0.00033824 -84.9915 0.21695
2.321 0.98804 5.5109e-005 3.8182 0.012018 3.049e-005 0.001155 0.20278 0.00065903 0.20343 0.18695 0 0.03387 0.0389 0 1.0042 0.29791 0.084314 0.011412 4.9807 0.071215 8.6861e-005 0.81887 0.0059148 0.0066713 0.0015463 0.98483 0.99026 3.3569e-006 1.3428e-005 0.13715 0.751 0.8065 0.0014796 0.84215 0.49369 0.0019901 0.42322 1.4097 1.4064 16.0072 144.974 0.00033742 -84.9963 0.21795
2.322 0.98804 5.5109e-005 3.8182 0.012018 3.0503e-005 0.001155 0.2028 0.00065903 0.20346 0.18697 0 0.033869 0.0389 0 1.0042 0.29795 0.08433 0.011414 4.9816 0.071226 8.6876e-005 0.81886 0.0059155 0.006672 0.0015451 0.98485 0.99028 3.354e-006 1.3416e-005 0.13716 0.75173 0.80702 0.001479 0.84309 0.49386 0.0019893 0.42323 1.4114 1.4081 16.0072 144.974 0.00033661 -85.0012 0.21895
2.323 0.98804 5.5109e-005 3.8182 0.012018 3.0516e-005 0.001155 0.20283 0.00065903 0.20348 0.187 0 0.033867 0.0389 0 1.0043 0.298 0.084345 0.011415 4.9825 0.071237 8.6891e-005 0.81885 0.0059161 0.0066727 0.0015439 0.98487 0.99029 3.3512e-006 1.3405e-005 0.13716 0.75245 0.80754 0.0014784 0.84403 0.49403 0.0019885 0.42324 1.413 1.4097 16.0073 144.974 0.0003358 -85.0059 0.21995
2.324 0.98804 5.5109e-005 3.8182 0.012018 3.0529e-005 0.001155 0.20285 0.00065903 0.20351 0.18702 0 0.033866 0.0389 0 1.0044 0.29804 0.084361 0.011417 4.9833 0.071249 8.6906e-005 0.81884 0.0059168 0.0066734 0.0015428 0.98488 0.9903 3.3484e-006 1.3394e-005 0.13717 0.75317 0.80806 0.0014778 0.84496 0.4942 0.0019877 0.42325 1.4147 1.4114 16.0073 144.974 0.000335 -85.0107 0.22095
2.325 0.98804 5.5109e-005 3.8182 0.012018 3.0542e-005 0.001155 0.20288 0.00065903 0.20353 0.18704 0 0.033865 0.0389 0 1.0045 0.29808 0.084376 0.011419 4.9842 0.07126 8.6921e-005 0.81883 0.0059175 0.0066741 0.0015416 0.9849 0.99032 3.3456e-006 1.3382e-005 0.13717 0.75388 0.80857 0.0014772 0.84589 0.49438 0.0019869 0.42325 1.4163 1.413 16.0073 144.9741 0.0003342 -85.0154 0.22195
2.326 0.98804 5.5109e-005 3.8182 0.012018 3.0555e-005 0.001155 0.20291 0.00065903 0.20356 0.18707 0 0.033863 0.0389 0 1.0046 0.29813 0.084392 0.011421 4.9851 0.071271 8.6935e-005 0.81882 0.0059181 0.0066748 0.0015404 0.98491 0.99033 3.3428e-006 1.3371e-005 0.13718 0.7546 0.80908 0.0014766 0.84681 0.49455 0.0019861 0.42326 1.4179 1.4147 16.0074 144.9741 0.0003334 -85.0201 0.22295
2.327 0.98804 5.5109e-005 3.8182 0.012018 3.0569e-005 0.001155 0.20293 0.00065903 0.20359 0.18709 0 0.033862 0.0389 0 1.0047 0.29817 0.084407 0.011423 4.986 0.071282 8.695e-005 0.8188 0.0059188 0.0066755 0.0015392 0.98493 0.99034 3.34e-006 1.336e-005 0.13718 0.75531 0.80959 0.001476 0.84772 0.49472 0.0019853 0.42327 1.4196 1.4163 16.0074 144.9741 0.00033261 -85.0247 0.22395
2.328 0.98804 5.5109e-005 3.8182 0.012018 3.0582e-005 0.001155 0.20296 0.00065903 0.20361 0.18712 0 0.03386 0.0389 0 1.0048 0.29821 0.084423 0.011424 4.9869 0.071293 8.6965e-005 0.81879 0.0059195 0.0066762 0.001538 0.98495 0.99036 3.3373e-006 1.335e-005 0.13719 0.75602 0.8101 0.0014754 0.84863 0.49489 0.0019845 0.42328 1.4212 1.418 16.0074 144.9741 0.00033182 -85.0293 0.22495
2.329 0.98804 5.5109e-005 3.8182 0.012018 3.0595e-005 0.001155 0.20298 0.00065903 0.20364 0.18714 0 0.033859 0.0389 0 1.0049 0.29826 0.084439 0.011426 4.9877 0.071304 8.698e-005 0.81878 0.0059201 0.0066769 0.0015368 0.98496 0.99037 3.3346e-006 1.3339e-005 0.1372 0.75672 0.8106 0.0014747 0.84954 0.49507 0.0019837 0.42329 1.4228 1.4196 16.0075 144.9741 0.00033104 -85.0339 0.22595
2.33 0.98804 5.5109e-005 3.8182 0.012018 3.0608e-005 0.001155 0.20301 0.00065903 0.20366 0.18717 0 0.033857 0.0389 0 1.005 0.2983 0.084454 0.011428 4.9886 0.071316 8.6995e-005 0.81877 0.0059208 0.0066776 0.0015357 0.98498 0.99038 3.332e-006 1.3328e-005 0.1372 0.75743 0.8111 0.0014741 0.85044 0.49524 0.001983 0.42329 1.4244 1.4212 16.0075 144.9741 0.00033025 -85.0384 0.22695
2.331 0.98804 5.5109e-005 3.8182 0.012018 3.0621e-005 0.001155 0.20304 0.00065903 0.20369 0.18719 0 0.033856 0.0389 0 1.0051 0.29834 0.08447 0.01143 4.9895 0.071327 8.7009e-005 0.81876 0.0059215 0.0066783 0.0015345 0.98499 0.99039 3.3293e-006 1.3317e-005 0.13721 0.75813 0.8116 0.0014735 0.85134 0.49541 0.0019822 0.4233 1.426 1.4229 16.0075 144.9742 0.00032948 -85.0429 0.22795
2.332 0.98804 5.5109e-005 3.8182 0.012018 3.0634e-005 0.001155 0.20306 0.00065903 0.20372 0.18722 0 0.033855 0.0389 0 1.0052 0.29839 0.084485 0.011432 4.9904 0.071338 8.7024e-005 0.81875 0.0059221 0.006679 0.0015333 0.98501 0.9904 3.3267e-006 1.3307e-005 0.13721 0.75883 0.8121 0.0014729 0.85223 0.49558 0.0019815 0.42331 1.4276 1.4245 16.0076 144.9742 0.0003287 -85.0474 0.22895
2.333 0.98804 5.5109e-005 3.8182 0.012018 3.0647e-005 0.001155 0.20309 0.00065903 0.20374 0.18724 0 0.033853 0.0389 0 1.0053 0.29843 0.084501 0.011433 4.9913 0.071349 8.7039e-005 0.81874 0.0059228 0.0066797 0.0015321 0.98502 0.99041 3.3241e-006 1.3297e-005 0.13722 0.75953 0.81259 0.0014723 0.85311 0.49576 0.0019807 0.42332 1.4293 1.4261 16.0076 144.9742 0.00032793 -85.0518 0.22995
2.334 0.98804 5.5109e-005 3.8182 0.012018 3.066e-005 0.001155 0.20311 0.00065903 0.20377 0.18727 0 0.033852 0.0389 0 1.0054 0.29848 0.084516 0.011435 4.9921 0.07136 8.7054e-005 0.81873 0.0059235 0.0066804 0.001531 0.98504 0.99043 3.3215e-006 1.3286e-005 0.13722 0.76023 0.81308 0.0014717 0.85399 0.49593 0.00198 0.42333 1.4309 1.4277 16.0076 144.9742 0.00032717 -85.0562 0.23095
2.335 0.98804 5.5108e-005 3.8182 0.012018 3.0673e-005 0.001155 0.20314 0.00065903 0.20379 0.18729 0 0.03385 0.0389 0 1.0055 0.29852 0.084532 0.011437 4.993 0.071371 8.7069e-005 0.81872 0.0059242 0.0066811 0.0015299 0.98505 0.99044 3.3189e-006 1.3276e-005 0.13723 0.76092 0.81357 0.0014712 0.85487 0.4961 0.0019792 0.42334 1.4325 1.4293 16.0077 144.9742 0.0003264 -85.0606 0.23195
2.336 0.98804 5.5108e-005 3.8182 0.012018 3.0686e-005 0.001155 0.20317 0.00065903 0.20382 0.18731 0 0.033849 0.0389 0 1.0056 0.29856 0.084548 0.011439 4.9939 0.071383 8.7083e-005 0.8187 0.0059248 0.0066818 0.0015287 0.98507 0.99045 3.3164e-006 1.3266e-005 0.13723 0.76162 0.81405 0.0014706 0.85574 0.49627 0.0019785 0.42334 1.434 1.4309 16.0077 144.9742 0.00032564 -85.0649 0.23295
2.337 0.98804 5.5108e-005 3.8182 0.012018 3.0699e-005 0.0011551 0.20319 0.00065903 0.20385 0.18734 0 0.033848 0.0389 0 1.0057 0.29861 0.084563 0.01144 4.9948 0.071394 8.7098e-005 0.81869 0.0059255 0.0066825 0.0015277 0.98508 0.99046 3.3139e-006 1.3256e-005 0.13724 0.76231 0.81454 0.0014701 0.8566 0.49644 0.0019778 0.42335 1.4356 1.4325 16.0077 144.9742 0.00032489 -85.0692 0.23395
2.338 0.98804 5.5108e-005 3.8182 0.012018 3.0712e-005 0.0011551 0.20322 0.00065903 0.20387 0.18736 0 0.033846 0.0389 0 1.0058 0.29865 0.084579 0.011442 4.9957 0.071405 8.7113e-005 0.81868 0.0059262 0.0066832 0.0015266 0.9851 0.99047 3.3113e-006 1.3246e-005 0.13724 0.76299 0.81502 0.0014696 0.85746 0.49662 0.0019771 0.42336 1.4372 1.4341 16.0077 144.9743 0.00032414 -85.0735 0.23495
2.339 0.98804 5.5108e-005 3.8182 0.012018 3.0726e-005 0.0011551 0.20324 0.00065903 0.2039 0.18739 0 0.033845 0.0389 0 1.0059 0.29869 0.084594 0.011444 4.9965 0.071416 8.7128e-005 0.81867 0.0059268 0.0066839 0.0015255 0.98511 0.99048 3.3089e-006 1.3236e-005 0.13725 0.76368 0.81549 0.001469 0.85832 0.49679 0.0019764 0.42337 1.4388 1.4357 16.0078 144.9743 0.00032339 -85.0778 0.23595
2.34 0.98804 5.5108e-005 3.8182 0.012018 3.0739e-005 0.0011551 0.20327 0.00065903 0.20392 0.18741 0 0.033843 0.0389 0 1.006 0.29874 0.08461 0.011446 4.9974 0.071427 8.7143e-005 0.81866 0.0059275 0.0066846 0.0015245 0.98513 0.99049 3.3064e-006 1.3226e-005 0.13726 0.76436 0.81597 0.0014685 0.85917 0.49696 0.0019756 0.42338 1.4404 1.4373 16.0078 144.9743 0.00032264 -85.082 0.23695
2.341 0.98804 5.5108e-005 3.8182 0.012018 3.0752e-005 0.0011551 0.20329 0.00065903 0.20395 0.18744 0 0.033842 0.0389 0 1.0061 0.29878 0.084626 0.011448 4.9983 0.071438 8.7157e-005 0.81865 0.0059282 0.0066853 0.0015234 0.98514 0.9905 3.304e-006 1.3216e-005 0.13726 0.76504 0.81644 0.001468 0.86002 0.49713 0.0019749 0.42339 1.442 1.4389 16.0078 144.9743 0.0003219 -85.0861 0.23795
2.342 0.98804 5.5108e-005 3.8182 0.012018 3.0765e-005 0.0011551 0.20332 0.00065903 0.20397 0.18746 0 0.033841 0.0389 0 1.0062 0.29882 0.084641 0.011449 4.9992 0.07145 8.7172e-005 0.81864 0.0059288 0.006686 0.0015224 0.98515 0.99051 3.3015e-006 1.3206e-005 0.13727 0.76572 0.81691 0.0014675 0.86086 0.4973 0.0019742 0.4234 1.4435 1.4405 16.0079 144.9743 0.00032116 -85.0903 0.23895
2.343 0.98804 5.5108e-005 3.8182 0.012018 3.0778e-005 0.0011551 0.20335 0.00065903 0.204 0.18748 0 0.033839 0.0389 0 1.0063 0.29887 0.084657 0.011451 5.0001 0.071461 8.7187e-005 0.81863 0.0059295 0.0066867 0.0015213 0.98517 0.99052 3.2991e-006 1.3197e-005 0.13727 0.7664 0.81738 0.001467 0.86169 0.49747 0.0019736 0.4234 1.4451 1.4421 16.0079 144.9743 0.00032043 -85.0944 0.23995
2.344 0.98804 5.5108e-005 3.8182 0.012018 3.0791e-005 0.0011551 0.20337 0.00065904 0.20403 0.18751 0 0.033838 0.0389 0 1.0064 0.29891 0.084672 0.011453 5.001 0.071472 8.7202e-005 0.81862 0.0059302 0.0066874 0.0015203 0.98518 0.99053 3.2967e-006 1.3187e-005 0.13728 0.76708 0.81785 0.0014664 0.86253 0.49765 0.0019729 0.42341 1.4467 1.4436 16.0079 144.9744 0.0003197 -85.0985 0.24095
2.345 0.98804 5.5108e-005 3.8182 0.012018 3.0804e-005 0.0011551 0.2034 0.00065904 0.20405 0.18753 0 0.033836 0.0389 0 1.0065 0.29896 0.084688 0.011455 5.0019 0.071483 8.7217e-005 0.8186 0.0059309 0.0066881 0.0015193 0.9852 0.99054 3.2944e-006 1.3178e-005 0.13728 0.76775 0.81831 0.0014659 0.86335 0.49782 0.0019722 0.42342 1.4482 1.4452 16.0079 144.9744 0.00031897 -85.1025 0.24195
2.346 0.98804 5.5108e-005 3.8182 0.012018 3.0817e-005 0.0011551 0.20342 0.00065904 0.20408 0.18756 0 0.033835 0.0389 0 1.0066 0.299 0.084703 0.011457 5.0027 0.071494 8.7232e-005 0.81859 0.0059315 0.0066888 0.0015183 0.98521 0.99055 3.292e-006 1.3168e-005 0.13729 0.76842 0.81878 0.0014654 0.86418 0.49799 0.0019715 0.42343 1.4498 1.4468 16.008 144.9744 0.00031825 -85.1066 0.24295
2.347 0.98804 5.5108e-005 3.8182 0.012018 3.083e-005 0.0011551 0.20345 0.00065904 0.2041 0.18758 0 0.033834 0.0389 0 1.0067 0.29904 0.084719 0.011458 5.0036 0.071505 8.7246e-005 0.81858 0.0059322 0.0066895 0.0015173 0.98522 0.99056 3.2897e-006 1.3159e-005 0.13729 0.76909 0.81923 0.0014649 0.86499 0.49816 0.0019708 0.42344 1.4513 1.4483 16.008 144.9744 0.00031753 -85.1106 0.24395
2.348 0.98804 5.5108e-005 3.8182 0.012018 3.0843e-005 0.0011551 0.20347 0.00065904 0.20413 0.18761 0 0.033832 0.0389 0 1.0067 0.29909 0.084735 0.01146 5.0045 0.071517 8.7261e-005 0.81857 0.0059329 0.0066902 0.0015163 0.98524 0.99057 3.2874e-006 1.315e-005 0.1373 0.76976 0.81969 0.0014644 0.86581 0.49833 0.0019702 0.42345 1.4529 1.4499 16.008 144.9744 0.00031681 -85.1145 0.24495
2.349 0.98804 5.5108e-005 3.8182 0.012018 3.0856e-005 0.0011551 0.2035 0.00065904 0.20415 0.18763 0 0.033831 0.0389 0 1.0068 0.29913 0.08475 0.011462 5.0054 0.071528 8.7276e-005 0.81856 0.0059335 0.0066909 0.0015153 0.98525 0.99058 3.2851e-006 1.3141e-005 0.13731 0.77042 0.82015 0.0014639 0.86661 0.4985 0.0019695 0.42346 1.4544 1.4514 16.0081 144.9744 0.0003161 -85.1185 0.24595
2.35 0.98804 5.5107e-005 3.8182 0.012018 3.0869e-005 0.0011551 0.20353 0.00065904 0.20418 0.18765 0 0.033829 0.0389 0 1.0069 0.29917 0.084766 0.011464 5.0063 0.071539 8.7291e-005 0.81855 0.0059342 0.0066916 0.0015143 0.98526 0.99059 3.2828e-006 1.3132e-005 0.13731 0.77109 0.8206 0.0014633 0.86742 0.49868 0.0019689 0.42347 1.4559 1.453 16.0081 144.9745 0.00031539 -85.1224 0.24695
2.351 0.98804 5.5107e-005 3.8182 0.012018 3.0883e-005 0.0011551 0.20355 0.00065904 0.20421 0.18768 0 0.033828 0.0389 0 1.007 0.29922 0.084781 0.011465 5.0072 0.07155 8.7306e-005 0.81854 0.0059349 0.0066923 0.0015133 0.98528 0.9906 3.2806e-006 1.3123e-005 0.13732 0.77175 0.82105 0.0014628 0.86822 0.49885 0.0019682 0.42348 1.4575 1.4545 16.0081 144.9745 0.00031468 -85.1262 0.24795
2.352 0.98804 5.5107e-005 3.8182 0.012018 3.0896e-005 0.0011551 0.20358 0.00065904 0.20423 0.1877 0 0.033827 0.0389 0 1.0071 0.29926 0.084797 0.011467 5.0081 0.071561 8.732e-005 0.81853 0.0059356 0.006693 0.0015123 0.98529 0.99061 3.2784e-006 1.3114e-005 0.13732 0.77241 0.8215 0.0014623 0.86901 0.49902 0.0019676 0.42348 1.459 1.4561 16.0081 144.9745 0.00031398 -85.1301 0.24895
2.353 0.98804 5.5107e-005 3.8182 0.012018 3.0909e-005 0.0011551 0.2036 0.00065904 0.20426 0.18773 0 0.033825 0.0389 0 1.0072 0.2993 0.084813 0.011469 5.009 0.071573 8.7335e-005 0.81851 0.0059362 0.0066937 0.0015114 0.9853 0.99062 3.2761e-006 1.3105e-005 0.13733 0.77306 0.82194 0.0014619 0.8698 0.49919 0.0019669 0.42349 1.4605 1.4576 16.0082 144.9745 0.00031328 -85.1339 0.24995
2.354 0.98804 5.5107e-005 3.8182 0.012018 3.0922e-005 0.0011551 0.20363 0.00065904 0.20428 0.18775 0 0.033824 0.0389 0 1.0073 0.29935 0.084828 0.011471 5.0098 0.071584 8.735e-005 0.8185 0.0059369 0.0066944 0.0015104 0.98532 0.99063 3.2739e-006 1.3096e-005 0.13733 0.77372 0.82239 0.0014614 0.87059 0.49936 0.0019663 0.4235 1.462 1.4591 16.0082 144.9745 0.00031258 -85.1377 0.25095
2.355 0.98804 5.5107e-005 3.8182 0.012018 3.0935e-005 0.0011551 0.20365 0.00065904 0.20431 0.18777 0 0.033822 0.0389 0 1.0074 0.29939 0.084844 0.011473 5.0107 0.071595 8.7365e-005 0.81849 0.0059376 0.0066951 0.0015095 0.98533 0.99063 3.2718e-006 1.3087e-005 0.13734 0.77437 0.82283 0.0014609 0.87137 0.49953 0.0019657 0.42351 1.4636 1.4607 16.0082 144.9745 0.00031189 -85.1415 0.25195
2.356 0.98804 5.5107e-005 3.8182 0.012018 3.0948e-005 0.0011551 0.20368 0.00065904 0.20433 0.1878 0 0.033821 0.0389 0 1.0075 0.29944 0.084859 0.011474 5.0116 0.071606 8.738e-005 0.81848 0.0059383 0.0066958 0.0015085 0.98534 0.99064 3.2696e-006 1.3079e-005 0.13734 0.77502 0.82327 0.0014604 0.87214 0.4997 0.001965 0.42352 1.4651 1.4622 16.0082 144.9746 0.0003112 -85.1452 0.25295
2.357 0.98804 5.5107e-005 3.8182 0.012018 3.0961e-005 0.0011551 0.2037 0.00065904 0.20436 0.18782 0 0.03382 0.0389 0 1.0076 0.29948 0.084875 0.011476 5.0125 0.071617 8.7395e-005 0.81847 0.0059389 0.0066965 0.0015076 0.98535 0.99065 3.2675e-006 1.307e-005 0.13735 0.77567 0.82371 0.0014599 0.87291 0.49988 0.0019644 0.42353 1.4666 1.4637 16.0083 144.9746 0.00031051 -85.1489 0.25395
2.358 0.98804 5.5107e-005 3.8182 0.012018 3.0974e-005 0.0011551 0.20373 0.00065904 0.20438 0.18785 0 0.033818 0.0389 0 1.0077 0.29952 0.084891 0.011478 5.0134 0.071628 8.7409e-005 0.81846 0.0059396 0.0066972 0.0015067 0.98537 0.99066 3.2653e-006 1.3061e-005 0.13735 0.77632 0.82414 0.0014595 0.87368 0.50005 0.0019638 0.42354 1.4681 1.4652 16.0083 144.9746 0.00030983 -85.1526 0.25495
2.359 0.98804 5.5107e-005 3.8182 0.012018 3.0987e-005 0.0011551 0.20375 0.00065904 0.20441 0.18787 0 0.033817 0.0389 0 1.0078 0.29957 0.084906 0.01148 5.0143 0.07164 8.7424e-005 0.81845 0.0059403 0.0066979 0.0015057 0.98538 0.99067 3.2632e-006 1.3053e-005 0.13736 0.77696 0.82457 0.001459 0.87444 0.50022 0.0019632 0.42355 1.4696 1.4667 16.0083 144.9746 0.00030914 -85.1562 0.25595
2.36 0.98804 5.5107e-005 3.8182 0.012018 3.1e-005 0.0011551 0.20378 0.00065904 0.20443 0.18789 0 0.033816 0.0389 0 1.0079 0.29961 0.084922 0.011482 5.0152 0.071651 8.7439e-005 0.81844 0.0059409 0.0066986 0.0015048 0.98539 0.99068 3.2611e-006 1.3045e-005 0.13737 0.7776 0.825 0.0014585 0.8752 0.50039 0.0019626 0.42356 1.4711 1.4682 16.0083 144.9746 0.00030847 -85.1599 0.25695
2.361 0.98804 5.5107e-005 3.8182 0.012018 3.1013e-005 0.0011551 0.2038 0.00065904 0.20446 0.18792 0 0.033814 0.0389 0 1.008 0.29965 0.084937 0.011483 5.0161 0.071662 8.7454e-005 0.81843 0.0059416 0.0066993 0.0015039 0.9854 0.99069 3.259e-006 1.3036e-005 0.13737 0.77824 0.82543 0.0014581 0.87596 0.50056 0.001962 0.42357 1.4726 1.4697 16.0084 144.9746 0.00030779 -85.1635 0.25795
2.362 0.98804 5.5107e-005 3.8182 0.012018 3.1026e-005 0.0011551 0.20383 0.00065904 0.20448 0.18794 0 0.033813 0.0389 0 1.0081 0.2997 0.084953 0.011485 5.017 0.071673 8.7469e-005 0.81841 0.0059423 0.0067 0.001503 0.98541 0.99069 3.257e-006 1.3028e-005 0.13738 0.77888 0.82586 0.0014576 0.87671 0.50073 0.0019614 0.42358 1.4741 1.4712 16.0084 144.9747 0.00030712 -85.167 0.25895
2.363 0.98804 5.5107e-005 3.8182 0.012018 3.104e-005 0.0011551 0.20386 0.00065904 0.20451 0.18797 0 0.033811 0.0389 0 1.0082 0.29974 0.084969 0.011487 5.0179 0.071684 8.7483e-005 0.8184 0.005943 0.0067007 0.0015022 0.98543 0.9907 3.2549e-006 1.302e-005 0.13738 0.77952 0.82628 0.0014572 0.87745 0.5009 0.0019608 0.42359 1.4756 1.4727 16.0084 144.9747 0.00030645 -85.1706 0.25995
2.364 0.98804 5.5107e-005 3.8182 0.012018 3.1053e-005 0.0011551 0.20388 0.00065904 0.20453 0.18799 0 0.03381 0.0389 0 1.0083 0.29978 0.084984 0.011489 5.0188 0.071695 8.7498e-005 0.81839 0.0059436 0.0067014 0.0015013 0.98544 0.99071 3.2529e-006 1.3012e-005 0.13739 0.78016 0.82671 0.0014567 0.87819 0.50107 0.0019602 0.4236 1.477 1.4742 16.0084 144.9747 0.00030579 -85.1741 0.26095
2.365 0.98804 5.5106e-005 3.8182 0.012018 3.1066e-005 0.0011551 0.20391 0.00065904 0.20456 0.18801 0 0.033809 0.0389 0 1.0084 0.29983 0.085 0.01149 5.0197 0.071707 8.7513e-005 0.81838 0.0059443 0.0067021 0.0015004 0.98545 0.99072 3.2509e-006 1.3004e-005 0.13739 0.78079 0.82713 0.0014563 0.87893 0.50125 0.0019596 0.42361 1.4785 1.4757 16.0084 144.9747 0.00030513 -85.1776 0.26195
2.366 0.98804 5.5106e-005 3.8182 0.012018 3.1079e-005 0.0011551 0.20393 0.00065904 0.20459 0.18804 0 0.033807 0.0389 0 1.0085 0.29987 0.085016 0.011492 5.0206 0.071718 8.7528e-005 0.81837 0.005945 0.0067029 0.0014995 0.98546 0.99073 3.2489e-006 1.2996e-005 0.1374 0.78142 0.82755 0.0014558 0.87966 0.50142 0.0019591 0.42362 1.48 1.4772 16.0085 144.9747 0.00030447 -85.1811 0.26295
2.367 0.98804 5.5106e-005 3.8182 0.012018 3.1092e-005 0.0011551 0.20396 0.00065904 0.20461 0.18806 0 0.033806 0.0389 0 1.0086 0.29992 0.085031 0.011494 5.0215 0.071729 8.7543e-005 0.81836 0.0059457 0.0067036 0.0014987 0.98547 0.99073 3.2469e-006 1.2988e-005 0.1374 0.78205 0.82796 0.0014554 0.88039 0.50159 0.0019585 0.42363 1.4815 1.4787 16.0085 144.9747 0.00030381 -85.1845 0.26395
2.368 0.98804 5.5106e-005 3.8182 0.012018 3.1105e-005 0.0011551 0.20398 0.00065904 0.20464 0.18809 0 0.033805 0.0389 0 1.0087 0.29996 0.085047 0.011496 5.0223 0.07174 8.7558e-005 0.81835 0.0059463 0.0067043 0.0014978 0.98548 0.99074 3.245e-006 1.298e-005 0.13741 0.78267 0.82838 0.001455 0.88111 0.50176 0.0019579 0.42364 1.4829 1.4802 16.0085 144.9748 0.00030316 -85.1879 0.26495
2.369 0.98804 5.5106e-005 3.8182 0.012018 3.1118e-005 0.0011551 0.20401 0.00065904 0.20466 0.18811 0 0.033803 0.0389 0 1.0088 0.3 0.085062 0.011498 5.0232 0.071751 8.7572e-005 0.81834 0.005947 0.006705 0.0014969 0.98549 0.99075 3.243e-006 1.2972e-005 0.13742 0.7833 0.82879 0.0014545 0.88183 0.50193 0.0019574 0.42365 1.4844 1.4816 16.0085 144.9748 0.00030251 -85.1913 0.26595
2.37 0.98804 5.5106e-005 3.8182 0.012018 3.1131e-005 0.0011551 0.20403 0.00065904 0.20469 0.18813 0 0.033802 0.0389 0 1.0089 0.30005 0.085078 0.011499 5.0241 0.071762 8.7587e-005 0.81833 0.0059477 0.0067057 0.0014961 0.98551 0.99076 3.2411e-006 1.2964e-005 0.13742 0.78392 0.8292 0.0014541 0.88255 0.5021 0.0019568 0.42366 1.4859 1.4831 16.0086 144.9748 0.00030186 -85.1947 0.26695
2.371 0.98804 5.5106e-005 3.8182 0.012018 3.1144e-005 0.0011551 0.20406 0.00065904 0.20471 0.18816 0 0.0338 0.0389 0 1.009 0.30009 0.085094 0.011501 5.025 0.071774 8.7602e-005 0.81831 0.0059484 0.0067064 0.0014953 0.98552 0.99076 3.2392e-006 1.2957e-005 0.13743 0.78454 0.82961 0.0014537 0.88326 0.50227 0.0019562 0.42367 1.4873 1.4846 16.0086 144.9748 0.00030122 -85.198 0.26795
2.372 0.98804 5.5106e-005 3.8182 0.012018 3.1157e-005 0.0011551 0.20408 0.00065904 0.20474 0.18818 0 0.033799 0.0389 0 1.0091 0.30013 0.085109 0.011503 5.0259 0.071785 8.7617e-005 0.8183 0.005949 0.0067071 0.0014944 0.98553 0.99077 3.2373e-006 1.2949e-005 0.13743 0.78516 0.83001 0.0014532 0.88396 0.50244 0.0019557 0.42368 1.4888 1.486 16.0086 144.9748 0.00030058 -85.2014 0.26895
2.373 0.98804 5.5106e-005 3.8182 0.012018 3.117e-005 0.0011551 0.20411 0.00065904 0.20476 0.1882 0 0.033798 0.0389 0 1.0092 0.30018 0.085125 0.011505 5.0268 0.071796 8.7632e-005 0.81829 0.0059497 0.0067078 0.0014936 0.98554 0.99078 3.2354e-006 1.2942e-005 0.13744 0.78578 0.83042 0.0014528 0.88467 0.50261 0.0019551 0.42369 1.4902 1.4875 16.0086 144.9748 0.00029994 -85.2047 0.26995
2.374 0.98804 5.5106e-005 3.8182 0.012018 3.1183e-005 0.0011551 0.20413 0.00065904 0.20479 0.18823 0 0.033796 0.0389 0 1.0092 0.30022 0.08514 0.011507 5.0277 0.071807 8.7647e-005 0.81828 0.0059504 0.0067085 0.0014928 0.98555 0.99079 3.2335e-006 1.2934e-005 0.13744 0.7864 0.83082 0.0014524 0.88537 0.50278 0.0019546 0.4237 1.4917 1.4889 16.0086 144.9749 0.00029931 -85.2079 0.27095
2.375 0.98804 5.5106e-005 3.8182 0.012018 3.1197e-005 0.0011551 0.20416 0.00065904 0.20481 0.18825 0 0.033795 0.0389 0 1.0093 0.30027 0.085156 0.011508 5.0286 0.071818 8.7661e-005 0.81827 0.0059511 0.0067092 0.001492 0.98556 0.99079 3.2317e-006 1.2927e-005 0.13745 0.78701 0.83122 0.001452 0.88606 0.50295 0.0019541 0.42371 1.4931 1.4904 16.0087 144.9749 0.00029868 -85.2112 0.27195
2.376 0.98804 5.5106e-005 3.8182 0.012018 3.121e-005 0.0011551 0.20418 0.00065904 0.20484 0.18828 0 0.033794 0.0389 0 1.0094 0.30031 0.085172 0.01151 5.0295 0.07183 8.7676e-005 0.81826 0.0059517 0.0067099 0.0014912 0.98557 0.9908 3.2298e-006 1.2919e-005 0.13745 0.78762 0.83162 0.0014516 0.88675 0.50312 0.0019535 0.42372 1.4945 1.4918 16.0087 144.9749 0.00029805 -85.2144 0.27295
2.377 0.98804 5.5106e-005 3.8182 0.012018 3.1223e-005 0.0011551 0.20421 0.00065904 0.20486 0.1883 0 0.033792 0.0389 0 1.0095 0.30035 0.085187 0.011512 5.0304 0.071841 8.7691e-005 0.81825 0.0059524 0.0067106 0.0014904 0.98558 0.99081 3.228e-006 1.2912e-005 0.13746 0.78823 0.83202 0.0014512 0.88744 0.50329 0.001953 0.42373 1.496 1.4933 16.0087 144.9749 0.00029742 -85.2176 0.27395
2.378 0.98804 5.5106e-005 3.8182 0.012018 3.1236e-005 0.0011551 0.20423 0.00065904 0.20489 0.18832 0 0.033791 0.0389 0 1.0096 0.3004 0.085203 0.011514 5.0313 0.071852 8.7706e-005 0.81824 0.0059531 0.0067113 0.0014896 0.98559 0.99081 3.2262e-006 1.2905e-005 0.13747 0.78884 0.83241 0.0014508 0.88812 0.50346 0.0019525 0.42374 1.4974 1.4947 16.0087 144.9749 0.0002968 -85.2208 0.27495
2.379 0.98804 5.5106e-005 3.8182 0.012018 3.1249e-005 0.0011551 0.20426 0.00065904 0.20491 0.18835 0 0.03379 0.0389 0 1.0097 0.30044 0.085219 0.011516 5.0322 0.071863 8.7721e-005 0.81822 0.0059538 0.006712 0.0014888 0.9856 0.99082 3.2244e-006 1.2898e-005 0.13747 0.78945 0.83281 0.0014504 0.8888 0.50363 0.0019519 0.42375 1.4988 1.4961 16.0087 144.9749 0.00029618 -85.2239 0.27595
2.38 0.98804 5.5105e-005 3.8182 0.012018 3.1262e-005 0.0011551 0.20428 0.00065904 0.20494 0.18837 0 0.033788 0.0389 0 1.0098 0.30048 0.085234 0.011517 5.0331 0.071874 8.7736e-005 0.81821 0.0059544 0.0067127 0.0014881 0.98561 0.99083 3.2226e-006 1.289e-005 0.13748 0.79005 0.8332 0.00145 0.88947 0.50381 0.0019514 0.42376 1.5002 1.4976 16.0088 144.975 0.00029556 -85.227 0.27695
2.381 0.98804 5.5105e-005 3.8182 0.012018 3.1275e-005 0.0011551 0.20431 0.00065904 0.20496 0.18839 0 0.033787 0.0389 0 1.0099 0.30053 0.08525 0.011519 5.034 0.071885 8.775e-005 0.8182 0.0059551 0.0067135 0.0014873 0.98562 0.99084 3.2208e-006 1.2883e-005 0.13748 0.79065 0.83359 0.0014496 0.89014 0.50398 0.0019509 0.42377 1.5017 1.499 16.0088 144.975 0.00029495 -85.2302 0.27795
2.382 0.98804 5.5105e-005 3.8182 0.012018 3.1288e-005 0.0011551 0.20433 0.00065905 0.20499 0.18842 0 0.033786 0.0389 0 1.01 0.30057 0.085266 0.011521 5.0349 0.071897 8.7765e-005 0.81819 0.0059558 0.0067142 0.0014866 0.98563 0.99084 3.219e-006 1.2876e-005 0.13749 0.79125 0.83398 0.0014492 0.89081 0.50415 0.0019504 0.42378 1.5031 1.5004 16.0088 144.975 0.00029434 -85.2332 0.27895
2.383 0.98804 5.5105e-005 3.8182 0.012018 3.1301e-005 0.0011551 0.20436 0.00065905 0.20501 0.18844 0 0.033784 0.0389 0 1.0101 0.30062 0.085281 0.011523 5.0358 0.071908 8.778e-005 0.81818 0.0059565 0.0067149 0.0014858 0.98564 0.99085 3.2173e-006 1.2869e-005 0.13749 0.79185 0.83436 0.0014488 0.89147 0.50432 0.0019499 0.42379 1.5045 1.5018 16.0088 144.975 0.00029373 -85.2363 0.27995
2.384 0.98804 5.5105e-005 3.8182 0.012018 3.1314e-005 0.0011551 0.20438 0.00065905 0.20504 0.18846 0 0.033783 0.0389 0 1.0102 0.30066 0.085297 0.011524 5.0367 0.071919 8.7795e-005 0.81817 0.0059571 0.0067156 0.0014851 0.98565 0.99086 3.2156e-006 1.2862e-005 0.1375 0.79245 0.83475 0.0014484 0.89213 0.50449 0.0019494 0.4238 1.5059 1.5033 16.0088 144.975 0.00029312 -85.2393 0.28095
2.385 0.98804 5.5105e-005 3.8182 0.012018 3.1327e-005 0.0011551 0.20441 0.00065905 0.20506 0.18849 0 0.033782 0.0389 0 1.0103 0.3007 0.085312 0.011526 5.0376 0.07193 8.781e-005 0.81816 0.0059578 0.0067163 0.0014843 0.98566 0.99086 3.2139e-006 1.2856e-005 0.1375 0.79304 0.83513 0.0014481 0.89279 0.50466 0.0019489 0.42381 1.5073 1.5047 16.0089 144.975 0.00029252 -85.2424 0.28195
2.386 0.98804 5.5105e-005 3.8182 0.012018 3.134e-005 0.0011551 0.20443 0.00065905 0.20509 0.18851 0 0.03378 0.0389 0 1.0104 0.30075 0.085328 0.011528 5.0385 0.071941 8.7825e-005 0.81815 0.0059585 0.006717 0.0014836 0.98567 0.99087 3.2121e-006 1.2849e-005 0.13751 0.79364 0.83551 0.0014477 0.89344 0.50483 0.0019484 0.42382 1.5087 1.5061 16.0089 144.9751 0.00029192 -85.2453 0.28295
2.387 0.98804 5.5105e-005 3.8182 0.012018 3.1354e-005 0.0011551 0.20446 0.00065905 0.20511 0.18853 0 0.033779 0.0389 0 1.0105 0.30079 0.085344 0.01153 5.0394 0.071952 8.784e-005 0.81814 0.0059592 0.0067177 0.0014828 0.98568 0.99088 3.2105e-006 1.2842e-005 0.13752 0.79423 0.83589 0.0014473 0.89408 0.505 0.0019479 0.42383 1.5101 1.5075 16.0089 144.9751 0.00029132 -85.2483 0.28395
2.388 0.98804 5.5105e-005 3.8182 0.012018 3.1367e-005 0.0011551 0.20448 0.00065905 0.20513 0.18856 0 0.033777 0.0389 0 1.0106 0.30083 0.085359 0.011532 5.0404 0.071964 8.7854e-005 0.81812 0.0059598 0.0067184 0.0014821 0.98569 0.99088 3.2088e-006 1.2835e-005 0.13752 0.79482 0.83626 0.0014469 0.89473 0.50517 0.0019474 0.42384 1.5115 1.5089 16.0089 144.9751 0.00029073 -85.2513 0.28495
2.389 0.98804 5.5105e-005 3.8182 0.012018 3.138e-005 0.0011551 0.20451 0.00065905 0.20516 0.18858 0 0.033776 0.0389 0 1.0107 0.30088 0.085375 0.011533 5.0413 0.071975 8.7869e-005 0.81811 0.0059605 0.0067191 0.0014814 0.9857 0.99089 3.2071e-006 1.2829e-005 0.13753 0.7954 0.83664 0.0014466 0.89537 0.50534 0.0019469 0.42385 1.5129 1.5103 16.0089 144.9751 0.00029013 -85.2542 0.28595
2.39 0.98804 5.5105e-005 3.8182 0.012017 3.1393e-005 0.0011551 0.20453 0.00065905 0.20518 0.1886 0 0.033775 0.0389 0 1.0108 0.30092 0.085391 0.011535 5.0422 0.071986 8.7884e-005 0.8181 0.0059612 0.0067198 0.0014806 0.98571 0.99089 3.2055e-006 1.2822e-005 0.13753 0.79599 0.83701 0.0014462 0.896 0.50551 0.0019464 0.42386 1.5142 1.5117 16.0089 144.9751 0.00028954 -85.2571 0.28695
2.391 0.98804 5.5105e-005 3.8182 0.012017 3.1406e-005 0.0011551 0.20455 0.00065905 0.20521 0.18863 0 0.033773 0.0389 0 1.0109 0.30097 0.085406 0.011537 5.0431 0.071997 8.7899e-005 0.81809 0.0059619 0.0067205 0.0014799 0.98572 0.9909 3.2038e-006 1.2815e-005 0.13754 0.79657 0.83738 0.0014458 0.89663 0.50568 0.001946 0.42387 1.5156 1.5131 16.009 144.9751 0.00028896 -85.26 0.28795
2.392 0.98804 5.5105e-005 3.8182 0.012017 3.1419e-005 0.0011551 0.20458 0.00065905 0.20523 0.18865 0 0.033772 0.0389 0 1.011 0.30101 0.085422 0.011539 5.044 0.072008 8.7914e-005 0.81808 0.0059626 0.0067212 0.0014792 0.98573 0.99091 3.2022e-006 1.2809e-005 0.13754 0.79716 0.83775 0.0014455 0.89726 0.50585 0.0019455 0.42388 1.517 1.5144 16.009 144.9752 0.00028837 -85.2629 0.28895
2.393 0.98804 5.5105e-005 3.8182 0.012017 3.1432e-005 0.0011551 0.2046 0.00065905 0.20526 0.18867 0 0.033771 0.0389 0 1.0111 0.30105 0.085438 0.011541 5.0449 0.07202 8.7929e-005 0.81807 0.0059632 0.006722 0.0014785 0.98574 0.99091 3.2006e-006 1.2803e-005 0.13755 0.79774 0.83812 0.0014451 0.89789 0.50602 0.001945 0.42389 1.5184 1.5158 16.009 144.9752 0.00028779 -85.2657 0.28995
2.394 0.98804 5.5105e-005 3.8182 0.012017 3.1445e-005 0.0011551 0.20463 0.00065905 0.20528 0.1887 0 0.033769 0.0389 0 1.0112 0.3011 0.085453 0.011542 5.0458 0.072031 8.7943e-005 0.81806 0.0059639 0.0067227 0.0014778 0.98575 0.99092 3.199e-006 1.2796e-005 0.13755 0.79831 0.83849 0.0014447 0.89851 0.50619 0.0019446 0.4239 1.5197 1.5172 16.009 144.9752 0.00028721 -85.2685 0.29095
2.395 0.98804 5.5104e-005 3.8182 0.012017 3.1458e-005 0.0011551 0.20465 0.00065905 0.20531 0.18872 0 0.033768 0.0389 0 1.0113 0.30114 0.085469 0.011544 5.0467 0.072042 8.7958e-005 0.81805 0.0059646 0.0067234 0.0014771 0.98576 0.99093 3.1974e-006 1.279e-005 0.13756 0.79889 0.83885 0.0014444 0.89912 0.50636 0.0019441 0.42391 1.5211 1.5186 16.009 144.9752 0.00028664 -85.2713 0.29195
2.396 0.98804 5.5104e-005 3.8182 0.012017 3.1471e-005 0.0011551 0.20468 0.00065905 0.20533 0.18874 0 0.033767 0.0389 0 1.0114 0.30119 0.085484 0.011546 5.0476 0.072053 8.7973e-005 0.81803 0.0059653 0.0067241 0.0014764 0.98577 0.99093 3.1958e-006 1.2783e-005 0.13757 0.79947 0.83922 0.001444 0.89974 0.50653 0.0019436 0.42392 1.5225 1.5199 16.009 144.9752 0.00028606 -85.2741 0.29295
2.397 0.98804 5.5104e-005 3.8182 0.012017 3.1484e-005 0.0011551 0.2047 0.00065905 0.20536 0.18877 0 0.033765 0.0389 0 1.0115 0.30123 0.0855 0.011548 5.0485 0.072064 8.7988e-005 0.81802 0.0059659 0.0067248 0.0014758 0.98578 0.99094 3.1943e-006 1.2777e-005 0.13757 0.80004 0.83958 0.0014437 0.90035 0.5067 0.0019432 0.42393 1.5238 1.5213 16.0091 144.9752 0.00028549 -85.2769 0.29395
2.398 0.98804 5.5104e-005 3.8182 0.012017 3.1497e-005 0.0011551 0.20473 0.00065905 0.20538 0.18879 0 0.033764 0.0389 0 1.0116 0.30127 0.085516 0.011549 5.0494 0.072075 8.8003e-005 0.81801 0.0059666 0.0067255 0.0014751 0.98578 0.99094 3.1927e-006 1.2771e-005 0.13758 0.80061 0.83994 0.0014433 0.90095 0.50687 0.0019427 0.42394 1.5252 1.5227 16.0091 144.9753 0.00028492 -85.2796 0.29495
2.399 0.98804 5.5104e-005 3.8182 0.012017 3.1511e-005 0.0011551 0.20475 0.00065905 0.20541 0.18881 0 0.033763 0.0389 0 1.0117 0.30132 0.085531 0.011551 5.0503 0.072087 8.8018e-005 0.818 0.0059673 0.0067262 0.0014745 0.98579 0.99095 3.1912e-006 1.2765e-005 0.13758 0.80118 0.8403 0.001443 0.90155 0.50703 0.0019423 0.42395 1.5265 1.524 16.0091 144.9753 0.00028436 -85.2823 0.29595
2.4 0.98804 5.5104e-005 3.8182 0.012017 3.1524e-005 0.0011551 0.20478 0.00065905 0.20543 0.18884 0 0.033761 0.0389 0 1.0118 0.30136 0.085547 0.011553 5.0512 0.072098 8.8032e-005 0.81799 0.005968 0.0067269 0.0014738 0.9858 0.99096 3.1897e-006 1.2759e-005 0.13759 0.80175 0.84065 0.0014427 0.90215 0.5072 0.0019418 0.42396 1.5279 1.5254 16.0091 144.9753 0.00028379 -85.285 0.29695
2.401 0.98804 5.5104e-005 3.8182 0.012017 3.1537e-005 0.0011551 0.2048 0.00065905 0.20546 0.18886 0 0.03376 0.0389 0 1.0118 0.3014 0.085563 0.011555 5.0521 0.072109 8.8047e-005 0.81798 0.0059686 0.0067276 0.0014731 0.98581 0.99096 3.1881e-006 1.2753e-005 0.13759 0.80231 0.84101 0.0014423 0.90275 0.50737 0.0019414 0.42398 1.5292 1.5267 16.0091 144.9753 0.00028323 -85.2877 0.29795
2.402 0.98804 5.5104e-005 3.8182 0.012017 3.155e-005 0.0011551 0.20483 0.00065905 0.20548 0.18888 0 0.033759 0.0389 0 1.0119 0.30145 0.085578 0.011557 5.0531 0.07212 8.8062e-005 0.81797 0.0059693 0.0067283 0.0014725 0.98582 0.99097 3.1866e-006 1.2747e-005 0.1376 0.80288 0.84136 0.001442 0.90334 0.50754 0.0019409 0.42399 1.5306 1.5281 16.0091 144.9753 0.00028268 -85.2904 0.29895
2.403 0.98804 5.5104e-005 3.8182 0.012017 3.1563e-005 0.0011551 0.20485 0.00065905 0.2055 0.18891 0 0.033757 0.0389 0 1.012 0.30149 0.085594 0.011558 5.054 0.072131 8.8077e-005 0.81796 0.00597 0.0067291 0.0014718 0.98583 0.99097 3.1852e-006 1.2741e-005 0.1376 0.80344 0.84171 0.0014417 0.90393 0.50771 0.0019405 0.424 1.5319 1.5294 16.0091 144.9754 0.00028212 -85.293 0.29995
2.404 0.98804 5.5104e-005 3.8182 0.012017 3.1576e-005 0.0011551 0.20487 0.00065905 0.20553 0.18893 0 0.033756 0.0389 0 1.0121 0.30154 0.08561 0.01156 5.0549 0.072142 8.8092e-005 0.81795 0.0059707 0.0067298 0.0014712 0.98584 0.99098 3.1837e-006 1.2735e-005 0.13761 0.804 0.84206 0.0014413 0.90451 0.50788 0.0019401 0.42401 1.5332 1.5308 16.0092 144.9754 0.00028157 -85.2957 0.30095
2.405 0.98804 5.5104e-005 3.8182 0.012017 3.1589e-005 0.0011551 0.2049 0.00065905 0.20555 0.18895 0 0.033755 0.0389 0 1.0122 0.30158 0.085625 0.011562 5.0558 0.072154 8.8107e-005 0.81793 0.0059714 0.0067305 0.0014705 0.98585 0.99098 3.1822e-006 1.2729e-005 0.13762 0.80456 0.84241 0.001441 0.90509 0.50805 0.0019396 0.42402 1.5346 1.5321 16.0092 144.9754 0.00028102 -85.2983 0.30195
2.406 0.98804 5.5104e-005 3.8182 0.012017 3.1602e-005 0.0011551 0.20492 0.00065905 0.20558 0.18898 0 0.033753 0.0389 0 1.0123 0.30162 0.085641 0.011564 5.0567 0.072165 8.8122e-005 0.81792 0.005972 0.0067312 0.0014699 0.98585 0.99099 3.1808e-006 1.2723e-005 0.13762 0.80512 0.84276 0.0014407 0.90567 0.50822 0.0019392 0.42403 1.5359 1.5334 16.0092 144.9754 0.00028047 -85.3009 0.30295
2.407 0.98804 5.5104e-005 3.8182 0.012017 3.1615e-005 0.0011551 0.20495 0.00065905 0.2056 0.189 0 0.033752 0.0389 0 1.0124 0.30167 0.085657 0.011566 5.0576 0.072176 8.8136e-005 0.81791 0.0059727 0.0067319 0.0014692 0.98586 0.991 3.1793e-006 1.2717e-005 0.13763 0.80567 0.8431 0.0014403 0.90624 0.50839 0.0019388 0.42404 1.5372 1.5348 16.0092 144.9754 0.00027992 -85.3034 0.30395
2.408 0.98804 5.5104e-005 3.8182 0.012017 3.1628e-005 0.0011551 0.20497 0.00065905 0.20563 0.18902 0 0.033751 0.0389 0 1.0125 0.30171 0.085672 0.011567 5.0585 0.072187 8.8151e-005 0.8179 0.0059734 0.0067326 0.0014686 0.98587 0.991 3.1779e-006 1.2712e-005 0.13763 0.80623 0.84345 0.00144 0.90681 0.50856 0.0019384 0.42405 1.5385 1.5361 16.0092 144.9754 0.00027938 -85.306 0.30495
2.409 0.98804 5.5104e-005 3.8182 0.012017 3.1641e-005 0.0011551 0.205 0.00065905 0.20565 0.18905 0 0.03375 0.0389 0 1.0126 0.30175 0.085688 0.011569 5.0594 0.072198 8.8166e-005 0.81789 0.0059741 0.0067333 0.001468 0.98588 0.99101 3.1765e-006 1.2706e-005 0.13764 0.80678 0.84379 0.0014397 0.90738 0.50873 0.001938 0.42406 1.5398 1.5374 16.0092 144.9755 0.00027884 -85.3085 0.30595
2.41 0.98804 5.5103e-005 3.8182 0.012017 3.1654e-005 0.0011551 0.20502 0.00065905 0.20567 0.18907 0 0.033748 0.0389 0 1.0127 0.3018 0.085704 0.011571 5.0604 0.07221 8.8181e-005 0.81788 0.0059748 0.006734 0.0014673 0.98589 0.99101 3.175e-006 1.27e-005 0.13764 0.80733 0.84413 0.0014394 0.90795 0.5089 0.0019375 0.42407 1.5411 1.5387 16.0092 144.9755 0.0002783 -85.311 0.30695
2.411 0.98804 5.5103e-005 3.8182 0.012017 3.1668e-005 0.0011551 0.20504 0.00065905 0.2057 0.18909 0 0.033747 0.0389 0 1.0128 0.30184 0.085719 0.011573 5.0613 0.072221 8.8196e-005 0.81787 0.0059754 0.0067347 0.0014667 0.98589 0.99102 3.1736e-006 1.2695e-005 0.13765 0.80788 0.84447 0.001439 0.90851 0.50907 0.0019371 0.42408 1.5425 1.5401 16.0093 144.9755 0.00027776 -85.3135 0.30795
2.412 0.98804 5.5103e-005 3.8182 0.012017 3.1681e-005 0.0011551 0.20507 0.00065905 0.20572 0.18911 0 0.033746 0.0389 0 1.0129 0.30189 0.085735 0.011574 5.0622 0.072232 8.8211e-005 0.81786 0.0059761 0.0067355 0.0014661 0.9859 0.99102 3.1723e-006 1.2689e-005 0.13765 0.80843 0.84481 0.0014387 0.90906 0.50924 0.0019367 0.42409 1.5438 1.5414 16.0093 144.9755 0.00027723 -85.316 0.30895
2.413 0.98804 5.5103e-005 3.8182 0.012017 3.1694e-005 0.0011551 0.20509 0.00065905 0.20575 0.18914 0 0.033744 0.0389 0 1.013 0.30193 0.085751 0.011576 5.0631 0.072243 8.8226e-005 0.81785 0.0059768 0.0067362 0.0014655 0.98591 0.99103 3.1709e-006 1.2684e-005 0.13766 0.80897 0.84514 0.0014384 0.90962 0.5094 0.0019363 0.42411 1.5451 1.5427 16.0093 144.9755 0.0002767 -85.3185 0.30995
2.414 0.98804 5.5103e-005 3.8182 0.012017 3.1707e-005 0.0011551 0.20512 0.00065905 0.20577 0.18916 0 0.033743 0.0389 0 1.0131 0.30197 0.085766 0.011578 5.064 0.072254 8.824e-005 0.81783 0.0059775 0.0067369 0.001465 0.98592 0.99103 3.1695e-006 1.2678e-005 0.13767 0.80952 0.84548 0.0014381 0.91017 0.50957 0.0019359 0.42412 1.5464 1.544 16.0093 144.9755 0.00027617 -85.3209 0.31095
2.415 0.98804 5.5103e-005 3.8182 0.012017 3.172e-005 0.0011551 0.20514 0.00065905 0.2058 0.18918 0 0.033742 0.0389 0 1.0132 0.30202 0.085782 0.01158 5.0649 0.072265 8.8255e-005 0.81782 0.0059782 0.0067376 0.0014644 0.98593 0.99104 3.1681e-006 1.2673e-005 0.13767 0.81006 0.84581 0.0014378 0.91071 0.50974 0.0019355 0.42413 1.5476 1.5453 16.0093 144.9756 0.00027564 -85.3233 0.31195
2.416 0.98804 5.5103e-005 3.8182 0.012017 3.1733e-005 0.0011551 0.20517 0.00065905 0.20582 0.18921 0 0.03374 0.0389 0 1.0133 0.30206 0.085798 0.011582 5.0659 0.072277 8.827e-005 0.81781 0.0059788 0.0067383 0.0014638 0.98593 0.99104 3.1668e-006 1.2667e-005 0.13768 0.8106 0.84614 0.0014375 0.91126 0.50991 0.0019351 0.42414 1.5489 1.5466 16.0093 144.9756 0.00027512 -85.3257 0.31295
2.417 0.98804 5.5103e-005 3.8182 0.012017 3.1746e-005 0.0011551 0.20519 0.00065905 0.20584 0.18923 0 0.033739 0.0389 0 1.0134 0.30211 0.085813 0.011583 5.0668 0.072288 8.8285e-005 0.8178 0.0059795 0.006739 0.0014633 0.98594 0.99105 3.1654e-006 1.2662e-005 0.13768 0.81114 0.84647 0.0014372 0.9118 0.51008 0.0019347 0.42415 1.5502 1.5479 16.0093 144.9756 0.0002746 -85.3281 0.31395
2.418 0.98804 5.5103e-005 3.8182 0.012017 3.1759e-005 0.0011551 0.20521 0.00065905 0.20587 0.18925 0 0.033738 0.0389 0 1.0135 0.30215 0.085829 0.011585 5.0677 0.072299 8.83e-005 0.81779 0.0059802 0.0067397 0.0014627 0.98595 0.99105 3.1641e-006 1.2656e-005 0.13769 0.81167 0.8468 0.0014369 0.91234 0.51025 0.0019343 0.42416 1.5515 1.5492 16.0093 144.9756 0.00027408 -85.3305 0.31495
2.419 0.98804 5.5103e-005 3.8182 0.012017 3.1772e-005 0.0011551 0.20524 0.00065905 0.20589 0.18927 0 0.033736 0.0389 0 1.0136 0.30219 0.085845 0.011587 5.0686 0.07231 8.8315e-005 0.81778 0.0059809 0.0067404 0.0014621 0.98596 0.99106 3.1628e-006 1.2651e-005 0.13769 0.81221 0.84713 0.0014367 0.91287 0.51042 0.0019339 0.42417 1.5528 1.5505 16.0093 144.9756 0.00027356 -85.3329 0.31595
2.42 0.98804 5.5103e-005 3.8182 0.012017 3.1785e-005 0.0011551 0.20526 0.00065905 0.20592 0.1893 0 0.033735 0.0389 0 1.0137 0.30224 0.08586 0.011589 5.0695 0.072321 8.833e-005 0.81777 0.0059816 0.0067412 0.0014616 0.98596 0.99106 3.1615e-006 1.2646e-005 0.1377 0.81274 0.84746 0.0014364 0.9134 0.51059 0.0019336 0.42418 1.5541 1.5517 16.0094 144.9757 0.00027305 -85.3352 0.31695
2.421 0.98804 5.5103e-005 3.8182 0.012017 3.1798e-005 0.0011551 0.20529 0.00065905 0.20594 0.18932 0 0.033734 0.0389 0 1.0138 0.30228 0.085876 0.011591 5.0704 0.072333 8.8344e-005 0.81776 0.0059822 0.0067419 0.001461 0.98597 0.99107 3.1602e-006 1.2641e-005 0.1377 0.81327 0.84778 0.0014361 0.91393 0.51076 0.0019332 0.42419 1.5553 1.553 16.0094 144.9757 0.00027253 -85.3375 0.31795
2.422 0.98804 5.5103e-005 3.8182 0.012017 3.1811e-005 0.0011551 0.20531 0.00065906 0.20597 0.18934 0 0.033732 0.0389 0 1.0139 0.30233 0.085892 0.011592 5.0714 0.072344 8.8359e-005 0.81774 0.0059829 0.0067426 0.0014604 0.98598 0.99107 3.1589e-006 1.2636e-005 0.13771 0.8138 0.8481 0.0014358 0.91445 0.51092 0.0019328 0.42421 1.5566 1.5543 16.0094 144.9757 0.00027202 -85.3398 0.31895
2.423 0.98804 5.5103e-005 3.8182 0.012017 3.1825e-005 0.0011551 0.20533 0.00065906 0.20599 0.18937 0 0.033731 0.0389 0 1.014 0.30237 0.085907 0.011594 5.0723 0.072355 8.8374e-005 0.81773 0.0059836 0.0067433 0.0014598 0.98599 0.99108 3.1576e-006 1.2631e-005 0.13772 0.81433 0.84842 0.0014355 0.91497 0.51109 0.0019324 0.42422 1.5579 1.5556 16.0094 144.9757 0.00027152 -85.3421 0.31995
2.424 0.98804 5.5103e-005 3.8182 0.012017 3.1838e-005 0.0011552 0.20536 0.00065906 0.20601 0.18939 0 0.03373 0.0389 0 1.0141 0.30241 0.085923 0.011596 5.0732 0.072366 8.8389e-005 0.81772 0.0059843 0.006744 0.0014592 0.98599 0.99108 3.1564e-006 1.2625e-005 0.13772 0.81486 0.84874 0.0014352 0.91549 0.51126 0.0019321 0.42423 1.5591 1.5568 16.0094 144.9757 0.00027101 -85.3444 0.32095
2.425 0.98804 5.5102e-005 3.8182 0.012017 3.1851e-005 0.0011552 0.20538 0.00065906 0.20604 0.18941 0 0.033729 0.0389 0 1.0142 0.30246 0.085939 0.011598 5.0741 0.072377 8.8404e-005 0.81771 0.005985 0.0067447 0.0014587 0.986 0.99109 3.1551e-006 1.262e-005 0.13773 0.81539 0.84906 0.0014349 0.91601 0.51143 0.0019317 0.42424 1.5604 1.5581 16.0094 144.9757 0.00027051 -85.3466 0.32195
2.426 0.98804 5.5102e-005 3.8182 0.012017 3.1864e-005 0.0011552 0.20541 0.00065906 0.20606 0.18943 0 0.033727 0.0389 0 1.0143 0.3025 0.085954 0.011599 5.075 0.072388 8.8419e-005 0.8177 0.0059856 0.0067454 0.0014581 0.98601 0.99109 3.1539e-006 1.2615e-005 0.13773 0.81591 0.84938 0.0014346 0.91652 0.5116 0.0019313 0.42425 1.5616 1.5594 16.0094 144.9758 0.00027001 -85.3489 0.32295
2.427 0.98804 5.5102e-005 3.8182 0.012017 3.1877e-005 0.0011552 0.20543 0.00065906 0.20609 0.18946 0 0.033726 0.0389 0 1.0144 0.30255 0.08597 0.011601 5.076 0.0724 8.8434e-005 0.81769 0.0059863 0.0067462 0.0014575 0.98602 0.9911 3.1526e-006 1.261e-005 0.13774 0.81643 0.8497 0.0014343 0.91703 0.51177 0.0019309 0.42426 1.5629 1.5606 16.0094 144.9758 0.00026951 -85.3511 0.32395
2.428 0.98804 5.5102e-005 3.8182 0.012017 3.189e-005 0.0011552 0.20545 0.00065906 0.20611 0.18948 0 0.033725 0.0389 0 1.0145 0.30259 0.085986 0.011603 5.0769 0.072411 8.8448e-005 0.81768 0.005987 0.0067469 0.001457 0.98602 0.9911 3.1514e-006 1.2606e-005 0.13774 0.81695 0.85001 0.001434 0.91753 0.51193 0.0019306 0.42427 1.5641 1.5619 16.0094 144.9758 0.00026901 -85.3533 0.32495
2.429 0.98804 5.5102e-005 3.8182 0.012017 3.1903e-005 0.0011552 0.20548 0.00065906 0.20613 0.1895 0 0.033723 0.0389 0 1.0146 0.30263 0.086001 0.011605 5.0778 0.072422 8.8463e-005 0.81767 0.0059877 0.0067476 0.0014565 0.98603 0.99111 3.1502e-006 1.2601e-005 0.13775 0.81747 0.85032 0.0014338 0.91803 0.5121 0.0019302 0.42428 1.5654 1.5631 16.0094 144.9758 0.00026852 -85.3555 0.32595
2.43 0.98804 5.5102e-005 3.8182 0.012017 3.1916e-005 0.0011552 0.2055 0.00065906 0.20616 0.18952 0 0.033722 0.0389 0 1.0146 0.30268 0.086017 0.011607 5.0787 0.072433 8.8478e-005 0.81766 0.0059884 0.0067483 0.0014559 0.98604 0.99111 3.1489e-006 1.2596e-005 0.13775 0.81799 0.85063 0.0014335 0.91853 0.51227 0.0019299 0.4243 1.5666 1.5644 16.0095 144.9758 0.00026802 -85.3577 0.32695
2.431 0.98804 5.5102e-005 3.8182 0.012017 3.1929e-005 0.0011552 0.20553 0.00065906 0.20618 0.18955 0 0.033721 0.0389 0 1.0147 0.30272 0.086033 0.011608 5.0796 0.072444 8.8493e-005 0.81764 0.0059891 0.006749 0.0014554 0.98604 0.99112 3.1477e-006 1.2591e-005 0.13776 0.81851 0.85094 0.0014332 0.91903 0.51244 0.0019295 0.42431 1.5679 1.5656 16.0095 144.9759 0.00026753 -85.3598 0.32795
2.432 0.98804 5.5102e-005 3.8182 0.012017 3.1942e-005 0.0011552 0.20555 0.00065906 0.20621 0.18957 0 0.033719 0.0389 0 1.0148 0.30276 0.086049 0.01161 5.0806 0.072456 8.8508e-005 0.81763 0.0059897 0.0067497 0.0014549 0.98605 0.99112 3.1465e-006 1.2586e-005 0.13777 0.81902 0.85125 0.001433 0.91952 0.51261 0.0019292 0.42432 1.5691 1.5669 16.0095 144.9759 0.00026705 -85.362 0.32895
2.433 0.98804 5.5102e-005 3.8182 0.012017 3.1955e-005 0.0011552 0.20557 0.00065906 0.20623 0.18959 0 0.033718 0.0389 0 1.0149 0.30281 0.086064 0.011612 5.0815 0.072467 8.8523e-005 0.81762 0.0059904 0.0067504 0.0014544 0.98606 0.99112 3.1454e-006 1.2581e-005 0.13777 0.81953 0.85156 0.0014327 0.92001 0.51278 0.0019288 0.42433 1.5703 1.5681 16.0095 144.9759 0.00026656 -85.3641 0.32995
2.434 0.98804 5.5102e-005 3.8182 0.012017 3.1968e-005 0.0011552 0.2056 0.00065906 0.20625 0.18962 0 0.033717 0.0389 0 1.015 0.30285 0.08608 0.011614 5.0824 0.072478 8.8538e-005 0.81761 0.0059911 0.0067512 0.0014539 0.98606 0.99113 3.1442e-006 1.2577e-005 0.13778 0.82004 0.85187 0.0014324 0.9205 0.51294 0.0019285 0.42434 1.5716 1.5694 16.0095 144.9759 0.00026608 -85.3662 0.33095
2.435 0.98804 5.5102e-005 3.8182 0.012017 3.1981e-005 0.0011552 0.20562 0.00065906 0.20628 0.18964 0 0.033716 0.0389 0 1.0151 0.3029 0.086096 0.011616 5.0833 0.072489 8.8553e-005 0.8176 0.0059918 0.0067519 0.0014535 0.98607 0.99113 3.143e-006 1.2572e-005 0.13778 0.82055 0.85217 0.0014322 0.92098 0.51311 0.0019281 0.42435 1.5728 1.5706 16.0095 144.9759 0.00026559 -85.3683 0.33195
2.436 0.98804 5.5102e-005 3.8182 0.012017 3.1995e-005 0.0011552 0.20565 0.00065906 0.2063 0.18966 0 0.033714 0.0389 0 1.0152 0.30294 0.086111 0.011617 5.0843 0.0725 8.8567e-005 0.81759 0.0059925 0.0067526 0.001453 0.98608 0.99114 3.1418e-006 1.2567e-005 0.13779 0.82106 0.85248 0.0014319 0.92147 0.51328 0.0019278 0.42436 1.574 1.5718 16.0095 144.9759 0.00026511 -85.3704 0.33295
2.437 0.98804 5.5102e-005 3.8182 0.012017 3.2008e-005 0.0011552 0.20567 0.00065906 0.20632 0.18968 0 0.033713 0.0389 0 1.0153 0.30298 0.086127 0.011619 5.0852 0.072511 8.8582e-005 0.81758 0.0059931 0.0067533 0.0014525 0.98608 0.99114 3.1407e-006 1.2563e-005 0.13779 0.82157 0.85278 0.0014317 0.92194 0.51345 0.0019274 0.42438 1.5752 1.5731 16.0095 144.976 0.00026464 -85.3725 0.33395
2.438 0.98804 5.5102e-005 3.8182 0.012017 3.2021e-005 0.0011552 0.20569 0.00065906 0.20635 0.18971 0 0.033712 0.0389 0 1.0154 0.30303 0.086143 0.011621 5.0861 0.072523 8.8597e-005 0.81757 0.0059938 0.006754 0.001452 0.98609 0.99115 3.1396e-006 1.2558e-005 0.1378 0.82207 0.85308 0.0014314 0.92242 0.51362 0.0019271 0.42439 1.5765 1.5743 16.0095 144.976 0.00026416 -85.3745 0.33495
2.439 0.98804 5.5102e-005 3.8182 0.012017 3.2034e-005 0.0011552 0.20572 0.00065906 0.20637 0.18973 0 0.03371 0.0389 0 1.0155 0.30307 0.086158 0.011623 5.087 0.072534 8.8612e-005 0.81755 0.0059945 0.0067547 0.0014515 0.9861 0.99115 3.1384e-006 1.2554e-005 0.1378 0.82257 0.85338 0.0014312 0.92289 0.51378 0.0019268 0.4244 1.5777 1.5755 16.0095 144.976 0.00026369 -85.3766 0.33595
2.44 0.98804 5.5101e-005 3.8182 0.012017 3.2047e-005 0.0011552 0.20574 0.00065906 0.2064 0.18975 0 0.033709 0.0389 0 1.0156 0.30312 0.086174 0.011625 5.088 0.072545 8.8627e-005 0.81754 0.0059952 0.0067554 0.001451 0.9861 0.99116 3.1373e-006 1.2549e-005 0.13781 0.82308 0.85368 0.0014309 0.92336 0.51395 0.0019264 0.42441 1.5789 1.5767 16.0095 144.976 0.00026322 -85.3786 0.33695
2.441 0.98804 5.5101e-005 3.8182 0.012017 3.206e-005 0.0011552 0.20576 0.00065906 0.20642 0.18977 0 0.033708 0.0389 0 1.0157 0.30316 0.08619 0.011626 5.0889 0.072556 8.8642e-005 0.81753 0.0059959 0.0067562 0.0014505 0.98611 0.99116 3.1362e-006 1.2545e-005 0.13782 0.82358 0.85397 0.0014307 0.92383 0.51412 0.0019261 0.42442 1.5801 1.5779 16.0095 144.976 0.00026275 -85.3806 0.33795
2.442 0.98804 5.5101e-005 3.8182 0.012017 3.2073e-005 0.0011552 0.20579 0.00065906 0.20644 0.1898 0 0.033707 0.0389 0 1.0158 0.3032 0.086205 0.011628 5.0898 0.072567 8.8657e-005 0.81752 0.0059966 0.0067569 0.00145 0.98612 0.99116 3.1351e-006 1.254e-005 0.13782 0.82407 0.85427 0.0014304 0.92429 0.51429 0.0019258 0.42443 1.5813 1.5791 16.0096 144.9761 0.00026228 -85.3826 0.33895
2.443 0.98804 5.5101e-005 3.8182 0.012017 3.2086e-005 0.0011552 0.20581 0.00065906 0.20647 0.18982 0 0.033705 0.0389 0 1.0159 0.30325 0.086221 0.01163 5.0908 0.072578 8.8671e-005 0.81751 0.0059972 0.0067576 0.0014495 0.98612 0.99117 3.134e-006 1.2536e-005 0.13783 0.82457 0.85456 0.0014302 0.92475 0.51445 0.0019255 0.42445 1.5825 1.5803 16.0096 144.9761 0.00026182 -85.3846 0.33995
2.444 0.98804 5.5101e-005 3.8182 0.012017 3.2099e-005 0.0011552 0.20584 0.00065906 0.20649 0.18984 0 0.033704 0.0389 0 1.016 0.30329 0.086237 0.011632 5.0917 0.07259 8.8686e-005 0.8175 0.0059979 0.0067583 0.001449 0.98613 0.99117 3.1329e-006 1.2532e-005 0.13783 0.82507 0.85486 0.0014299 0.92521 0.51462 0.0019251 0.42446 1.5837 1.5815 16.0096 144.9761 0.00026135 -85.3866 0.34095
2.445 0.98804 5.5101e-005 3.8182 0.012017 3.2112e-005 0.0011552 0.20586 0.00065906 0.20651 0.18986 0 0.033703 0.0389 0 1.0161 0.30334 0.086253 0.011633 5.0926 0.072601 8.8701e-005 0.81749 0.0059986 0.006759 0.0014485 0.98613 0.99118 3.1318e-006 1.2527e-005 0.13784 0.82556 0.85515 0.0014297 0.92567 0.51479 0.0019248 0.42447 1.5849 1.5827 16.0096 144.9761 0.00026089 -85.3885 0.34195
2.446 0.98804 5.5101e-005 3.8182 0.012017 3.2125e-005 0.0011552 0.20588 0.00065906 0.20654 0.18988 0 0.033701 0.0389 0 1.0162 0.30338 0.086268 0.011635 5.0935 0.072612 8.8716e-005 0.81748 0.0059993 0.0067597 0.001448 0.98614 0.99118 3.1307e-006 1.2523e-005 0.13784 0.82605 0.85544 0.0014294 0.92612 0.51496 0.0019245 0.42448 1.5861 1.5839 16.0096 144.9761 0.00026043 -85.3905 0.34295
2.447 0.98804 5.5101e-005 3.8182 0.012017 3.2138e-005 0.0011552 0.20591 0.00065906 0.20656 0.18991 0 0.0337 0.0389 0 1.0163 0.30342 0.086284 0.011637 5.0945 0.072623 8.8731e-005 0.81747 0.006 0.0067605 0.0014476 0.98615 0.99118 3.1297e-006 1.2519e-005 0.13785 0.82654 0.85573 0.0014292 0.92657 0.51512 0.0019242 0.42449 1.5872 1.5851 16.0096 144.9761 0.00025998 -85.3924 0.34395
2.448 0.98804 5.5101e-005 3.8182 0.012017 3.2152e-005 0.0011552 0.20593 0.00065906 0.20658 0.18993 0 0.033699 0.0389 0 1.0164 0.30347 0.0863 0.011639 5.0954 0.072634 8.8746e-005 0.81745 0.0060007 0.0067612 0.0014471 0.98615 0.99119 3.1286e-006 1.2514e-005 0.13786 0.82703 0.85602 0.0014289 0.92702 0.51529 0.0019239 0.4245 1.5884 1.5863 16.0096 144.9762 0.00025952 -85.3943 0.34495
2.449 0.98804 5.5101e-005 3.8182 0.012017 3.2165e-005 0.0011552 0.20595 0.00065906 0.20661 0.18995 0 0.033698 0.0389 0 1.0165 0.30351 0.086315 0.011641 5.0963 0.072646 8.8761e-005 0.81744 0.0060013 0.0067619 0.0014467 0.98616 0.99119 3.1275e-006 1.251e-005 0.13786 0.82752 0.8563 0.0014287 0.92746 0.51546 0.0019236 0.42452 1.5896 1.5875 16.0096 144.9762 0.00025907 -85.3962 0.34595
2.45 0.98804 5.5101e-005 3.8182 0.012017 3.2178e-005 0.0011552 0.20598 0.00065906 0.20663 0.18997 0 0.033696 0.0389 0 1.0166 0.30356 0.086331 0.011642 5.0973 0.072657 8.8776e-005 0.81743 0.006002 0.0067626 0.0014462 0.98616 0.9912 3.1265e-006 1.2506e-005 0.13787 0.82801 0.85659 0.0014284 0.9279 0.51563 0.0019233 0.42453 1.5908 1.5887 16.0096 144.9762 0.00025862 -85.3981 0.34695
2.451 0.98804 5.5101e-005 3.8182 0.012017 3.2191e-005 0.0011552 0.206 0.00065906 0.20666 0.19 0 0.033695 0.0389 0 1.0167 0.3036 0.086347 0.011644 5.0982 0.072668 8.879e-005 0.81742 0.0060027 0.0067633 0.0014458 0.98617 0.9912 3.1255e-006 1.2502e-005 0.13787 0.82849 0.85687 0.0014282 0.92834 0.51579 0.0019229 0.42454 1.592 1.5899 16.0096 144.9762 0.00025817 -85.4 0.34795
2.452 0.98804 5.5101e-005 3.8182 0.012017 3.2204e-005 0.0011552 0.20602 0.00065906 0.20668 0.19002 0 0.033694 0.0389 0 1.0168 0.30364 0.086362 0.011646 5.0991 0.072679 8.8805e-005 0.81741 0.0060034 0.006764 0.0014453 0.98618 0.9912 3.1244e-006 1.2498e-005 0.13788 0.82897 0.85716 0.001428 0.92878 0.51596 0.0019226 0.42455 1.5931 1.591 16.0096 144.9762 0.00025772 -85.4018 0.34895
2.453 0.98804 5.5101e-005 3.8182 0.012017 3.2217e-005 0.0011552 0.20605 0.00065906 0.2067 0.19004 0 0.033693 0.0389 0 1.0169 0.30369 0.086378 0.011648 5.1001 0.07269 8.882e-005 0.8174 0.0060041 0.0067648 0.0014449 0.98618 0.99121 3.1234e-006 1.2494e-005 0.13788 0.82946 0.85744 0.0014278 0.92921 0.51613 0.0019223 0.42456 1.5943 1.5922 16.0096 144.9763 0.00025728 -85.4037 0.34995
2.454 0.98804 5.5101e-005 3.8182 0.012017 3.223e-005 0.0011552 0.20607 0.00065906 0.20673 0.19006 0 0.033691 0.0389 0 1.017 0.30373 0.086394 0.01165 5.101 0.072701 8.8835e-005 0.81739 0.0060048 0.0067655 0.0014445 0.98619 0.99121 3.1224e-006 1.249e-005 0.13789 0.82994 0.85772 0.0014276 0.92964 0.51629 0.001922 0.42457 1.5955 1.5934 16.0096 144.9763 0.00025683 -85.4055 0.35095
2.455 0.98804 5.51e-005 3.8182 0.012017 3.2243e-005 0.0011552 0.2061 0.00065906 0.20675 0.19009 0 0.03369 0.0389 0 1.0171 0.30378 0.08641 0.011651 5.1019 0.072713 8.885e-005 0.81738 0.0060054 0.0067662 0.001444 0.98619 0.99121 3.1214e-006 1.2486e-005 0.13789 0.83041 0.858 0.0014273 0.93007 0.51646 0.0019217 0.42459 1.5966 1.5946 16.0096 144.9763 0.00025639 -85.4073 0.35195
2.456 0.98804 5.51e-005 3.8182 0.012017 3.2256e-005 0.0011552 0.20612 0.00065906 0.20677 0.19011 0 0.033689 0.0389 0 1.0172 0.30382 0.086425 0.011653 5.1029 0.072724 8.8865e-005 0.81737 0.0060061 0.0067669 0.0014436 0.9862 0.99122 3.1204e-006 1.2482e-005 0.1379 0.83089 0.85828 0.0014271 0.9305 0.51663 0.0019215 0.4246 1.5978 1.5957 16.0096 144.9763 0.00025595 -85.4091 0.35295
2.457 0.98804 5.51e-005 3.8182 0.012017 3.2269e-005 0.0011552 0.20614 0.00065906 0.2068 0.19013 0 0.033688 0.0389 0 1.0173 0.30386 0.086441 0.011655 5.1038 0.072735 8.888e-005 0.81735 0.0060068 0.0067676 0.0014432 0.98621 0.99122 3.1194e-006 1.2478e-005 0.13791 0.83137 0.85855 0.0014269 0.93092 0.5168 0.0019212 0.42461 1.5989 1.5969 16.0096 144.9763 0.00025551 -85.4109 0.35395
2.458 0.98804 5.51e-005 3.8182 0.012017 3.2282e-005 0.0011552 0.20617 0.00065906 0.20682 0.19015 0 0.033686 0.0389 0 1.0174 0.30391 0.086457 0.011657 5.1047 0.072746 8.8895e-005 0.81734 0.0060075 0.0067684 0.0014427 0.98621 0.99123 3.1184e-006 1.2474e-005 0.13791 0.83184 0.85883 0.0014267 0.93134 0.51696 0.0019209 0.42462 1.6001 1.598 16.0096 144.9763 0.00025508 -85.4127 0.35495
2.459 0.98804 5.51e-005 3.8182 0.012017 3.2295e-005 0.0011552 0.20619 0.00065906 0.20684 0.19017 0 0.033685 0.0389 0 1.0175 0.30395 0.086472 0.011658 5.1057 0.072757 8.8909e-005 0.81733 0.0060082 0.0067691 0.0014423 0.98622 0.99123 3.1175e-006 1.247e-005 0.13792 0.83232 0.8591 0.0014264 0.93176 0.51713 0.0019206 0.42463 1.6012 1.5992 16.0096 144.9764 0.00025464 -85.4145 0.35595
2.46 0.98804 5.51e-005 3.8182 0.012016 3.2308e-005 0.0011552 0.20621 0.00065906 0.20687 0.1902 0 0.033684 0.0389 0 1.0176 0.304 0.086488 0.01166 5.1066 0.072769 8.8924e-005 0.81732 0.0060089 0.0067698 0.0014419 0.98622 0.99123 3.1165e-006 1.2466e-005 0.13792 0.83279 0.85938 0.0014262 0.93218 0.5173 0.0019203 0.42465 1.6024 1.6004 16.0097 144.9764 0.00025421 -85.4162 0.35695
2.461 0.98804 5.51e-005 3.8182 0.012016 3.2322e-005 0.0011552 0.20624 0.00065906 0.20689 0.19022 0 0.033682 0.0389 0 1.0176 0.30404 0.086504 0.011662 5.1075 0.07278 8.8939e-005 0.81731 0.0060096 0.0067705 0.0014415 0.98623 0.99124 3.1155e-006 1.2462e-005 0.13793 0.83326 0.85965 0.001426 0.93259 0.51746 0.00192 0.42466 1.6035 1.6015 16.0097 144.9764 0.00025378 -85.418 0.35795
2.462 0.98805 5.51e-005 3.8182 0.012016 3.2335e-005 0.0011552 0.20626 0.00065906 0.20691 0.19024 0 0.033681 0.0389 0 1.0177 0.30408 0.08652 0.011664 5.1085 0.072791 8.8954e-005 0.8173 0.0060102 0.0067712 0.0014411 0.98623 0.99124 3.1146e-006 1.2458e-005 0.13793 0.83372 0.85992 0.0014258 0.933 0.51763 0.0019197 0.42467 1.6047 1.6026 16.0097 144.9764 0.00025335 -85.4197 0.35895
2.463 0.98805 5.51e-005 3.8182 0.012016 3.2348e-005 0.0011552 0.20628 0.00065907 0.20694 0.19026 0 0.03368 0.0389 0 1.0178 0.30413 0.086535 0.011666 5.1094 0.072802 8.8969e-005 0.81729 0.0060109 0.0067719 0.0014406 0.98624 0.99124 3.1136e-006 1.2454e-005 0.13794 0.83419 0.86019 0.0014256 0.93341 0.5178 0.0019194 0.42468 1.6058 1.6038 16.0097 144.9764 0.00025293 -85.4214 0.35995
2.464 0.98805 5.51e-005 3.8182 0.012016 3.2361e-005 0.0011552 0.20631 0.00065907 0.20696 0.19028 0 0.033679 0.0389 0 1.0179 0.30417 0.086551 0.011667 5.1103 0.072813 8.8984e-005 0.81728 0.0060116 0.0067727 0.0014402 0.98624 0.99125 3.1127e-006 1.2451e-005 0.13794 0.83466 0.86046 0.0014253 0.93381 0.51796 0.0019192 0.42469 1.6069 1.6049 16.0097 144.9765 0.0002525 -85.4231 0.36095
2.465 0.98805 5.51e-005 3.8182 0.012016 3.2374e-005 0.0011552 0.20633 0.00065907 0.20698 0.19031 0 0.033677 0.0389 0 1.018 0.30422 0.086567 0.011669 5.1113 0.072825 8.8999e-005 0.81726 0.0060123 0.0067734 0.0014398 0.98625 0.99125 3.1117e-006 1.2447e-005 0.13795 0.83512 0.86073 0.0014251 0.93421 0.51813 0.0019189 0.4247 1.6081 1.6061 16.0097 144.9765 0.00025208 -85.4248 0.36195
2.466 0.98805 5.51e-005 3.8182 0.012016 3.2387e-005 0.0011552 0.20635 0.00065907 0.20701 0.19033 0 0.033676 0.0389 0 1.0181 0.30426 0.086582 0.011671 5.1122 0.072836 8.9014e-005 0.81725 0.006013 0.0067741 0.0014394 0.98625 0.99125 3.1108e-006 1.2443e-005 0.13796 0.83558 0.86099 0.0014249 0.93461 0.5183 0.0019186 0.42472 1.6092 1.6072 16.0097 144.9765 0.00025166 -85.4265 0.36295
2.467 0.98805 5.51e-005 3.8182 0.012016 3.24e-005 0.0011552 0.20638 0.00065907 0.20703 0.19035 0 0.033675 0.0389 0 1.0182 0.30431 0.086598 0.011673 5.1132 0.072847 8.9028e-005 0.81724 0.0060137 0.0067748 0.001439 0.98626 0.99126 3.1099e-006 1.244e-005 0.13796 0.83605 0.86126 0.0014247 0.93501 0.51846 0.0019183 0.42473 1.6103 1.6083 16.0097 144.9765 0.00025124 -85.4282 0.36395
2.468 0.98805 5.51e-005 3.8182 0.012016 3.2413e-005 0.0011552 0.2064 0.00065907 0.20705 0.19037 0 0.033674 0.0389 0 1.0183 0.30435 0.086614 0.011675 5.1141 0.072858 8.9043e-005 0.81723 0.0060144 0.0067755 0.0014386 0.98626 0.99126 3.109e-006 1.2436e-005 0.13797 0.8365 0.86152 0.0014245 0.93541 0.51863 0.0019181 0.42474 1.6114 1.6095 16.0097 144.9765 0.00025082 -85.4298 0.36495
2.469 0.98805 5.51e-005 3.8182 0.012016 3.2426e-005 0.0011552 0.20642 0.00065907 0.20708 0.19039 0 0.033672 0.0389 0 1.0184 0.30439 0.08663 0.011676 5.115 0.072869 8.9058e-005 0.81722 0.006015 0.0067763 0.0014382 0.98627 0.99127 3.1081e-006 1.2432e-005 0.13797 0.83696 0.86179 0.0014243 0.9358 0.5188 0.0019178 0.42475 1.6125 1.6106 16.0097 144.9766 0.00025041 -85.4315 0.36595
2.47 0.98805 5.5099e-005 3.8182 0.012016 3.2439e-005 0.0011552 0.20644 0.00065907 0.2071 0.19042 0 0.033671 0.0389 0 1.0185 0.30444 0.086645 0.011678 5.116 0.07288 8.9073e-005 0.81721 0.0060157 0.006777 0.0014378 0.98628 0.99127 3.1072e-006 1.2429e-005 0.13798 0.83742 0.86205 0.0014241 0.93619 0.51896 0.0019175 0.42476 1.6137 1.6117 16.0097 144.9766 0.00024999 -85.4331 0.36695
2.471 0.98805 5.5099e-005 3.8182 0.012016 3.2452e-005 0.0011552 0.20647 0.00065907 0.20712 0.19044 0 0.03367 0.0389 0 1.0186 0.30448 0.086661 0.01168 5.1169 0.072892 8.9088e-005 0.8172 0.0060164 0.0067777 0.0014374 0.98628 0.99127 3.1063e-006 1.2425e-005 0.13798 0.83788 0.86231 0.0014239 0.93658 0.51913 0.0019173 0.42478 1.6148 1.6128 16.0097 144.9766 0.00024958 -85.4347 0.36795
2.472 0.98805 5.5099e-005 3.8182 0.012016 3.2465e-005 0.0011552 0.20649 0.00065907 0.20715 0.19046 0 0.033669 0.0389 0 1.0187 0.30453 0.086677 0.011682 5.1178 0.072903 8.9103e-005 0.81719 0.0060171 0.0067784 0.001437 0.98629 0.99128 3.1054e-006 1.2422e-005 0.13799 0.83833 0.86257 0.0014237 0.93696 0.51929 0.001917 0.42479 1.6159 1.6139 16.0097 144.9766 0.00024917 -85.4364 0.36895
2.473 0.98805 5.5099e-005 3.8182 0.012016 3.2479e-005 0.0011552 0.20651 0.00065907 0.20717 0.19048 0 0.033667 0.0389 0 1.0188 0.30457 0.086693 0.011684 5.1188 0.072914 8.9118e-005 0.81718 0.0060178 0.0067791 0.0014366 0.98629 0.99128 3.1045e-006 1.2418e-005 0.138 0.83878 0.86283 0.0014234 0.93735 0.51946 0.0019167 0.4248 1.617 1.615 16.0097 144.9766 0.00024876 -85.438 0.36995
2.474 0.98805 5.5099e-005 3.8182 0.012016 3.2492e-005 0.0011552 0.20654 0.00065907 0.20719 0.1905 0 0.033666 0.0389 0 1.0189 0.30461 0.086708 0.011685 5.1197 0.072925 8.9133e-005 0.81716 0.0060185 0.0067799 0.0014363 0.9863 0.99128 3.1037e-006 1.2415e-005 0.138 0.83923 0.86309 0.0014232 0.93773 0.51963 0.0019165 0.42481 1.6181 1.6162 16.0097 144.9766 0.00024836 -85.4395 0.37095
2.475 0.98805 5.5099e-005 3.8182 0.012016 3.2505e-005 0.0011552 0.20656 0.00065907 0.20721 0.19053 0 0.033665 0.0389 0 1.019 0.30466 0.086724 0.011687 5.1207 0.072936 8.9148e-005 0.81715 0.0060192 0.0067806 0.0014359 0.9863 0.99128 3.1028e-006 1.2411e-005 0.13801 0.83968 0.86334 0.001423 0.93811 0.51979 0.0019162 0.42483 1.6192 1.6173 16.0097 144.9767 0.00024795 -85.4411 0.37195
2.476 0.98805 5.5099e-005 3.8182 0.012016 3.2518e-005 0.0011552 0.20658 0.00065907 0.20724 0.19055 0 0.033664 0.0389 0 1.0191 0.3047 0.08674 0.011689 5.1216 0.072948 8.9162e-005 0.81714 0.0060198 0.0067813 0.0014355 0.9863 0.99129 3.1019e-006 1.2408e-005 0.13801 0.84013 0.8636 0.0014229 0.93848 0.51996 0.001916 0.42484 1.6203 1.6184 16.0097 144.9767 0.00024755 -85.4427 0.37295
2.477 0.98805 5.5099e-005 3.8182 0.012016 3.2531e-005 0.0011552 0.20661 0.00065907 0.20726 0.19057 0 0.033662 0.0389 0 1.0192 0.30475 0.086755 0.011691 5.1226 0.072959 8.9177e-005 0.81713 0.0060205 0.006782 0.0014351 0.98631 0.99129 3.1011e-006 1.2404e-005 0.13802 0.84058 0.86385 0.0014227 0.93886 0.52012 0.0019157 0.42485 1.6214 1.6195 16.0097 144.9767 0.00024715 -85.4443 0.37395
2.478 0.98805 5.5099e-005 3.8182 0.012016 3.2544e-005 0.0011552 0.20663 0.00065907 0.20728 0.19059 0 0.033661 0.0389 0 1.0193 0.30479 0.086771 0.011692 5.1235 0.07297 8.9192e-005 0.81712 0.0060212 0.0067827 0.0014348 0.98631 0.99129 3.1002e-006 1.2401e-005 0.13802 0.84102 0.86411 0.0014225 0.93923 0.52029 0.0019155 0.42486 1.6225 1.6206 16.0097 144.9767 0.00024675 -85.4458 0.37495
2.479 0.98805 5.5099e-005 3.8182 0.012016 3.2557e-005 0.0011552 0.20665 0.00065907 0.20731 0.19061 0 0.03366 0.0389 0 1.0194 0.30483 0.086787 0.011694 5.1244 0.072981 8.9207e-005 0.81711 0.0060219 0.0067835 0.0014344 0.98632 0.9913 3.0994e-006 1.2398e-005 0.13803 0.84147 0.86436 0.0014223 0.9396 0.52046 0.0019152 0.42487 1.6235 1.6217 16.0097 144.9767 0.00024635 -85.4473 0.37595
2.48 0.98805 5.5099e-005 3.8182 0.012016 3.257e-005 0.0011552 0.20668 0.00065907 0.20733 0.19063 0 0.033659 0.0389 0 1.0195 0.30488 0.086803 0.011696 5.1254 0.072992 8.9222e-005 0.8171 0.0060226 0.0067842 0.001434 0.98632 0.9913 3.0985e-006 1.2394e-005 0.13803 0.84191 0.86461 0.0014221 0.93997 0.52062 0.001915 0.42489 1.6246 1.6227 16.0097 144.9768 0.00024595 -85.4489 0.37695
2.481 0.98805 5.5099e-005 3.8182 0.012016 3.2583e-005 0.0011552 0.2067 0.00065907 0.20735 0.19066 0 0.033657 0.0389 0 1.0196 0.30492 0.086818 0.011698 5.1263 0.073003 8.9237e-005 0.81709 0.0060233 0.0067849 0.0014337 0.98633 0.9913 3.0977e-006 1.2391e-005 0.13804 0.84235 0.86486 0.0014219 0.94033 0.52079 0.0019147 0.4249 1.6257 1.6238 16.0097 144.9768 0.00024556 -85.4504 0.37795
2.482 0.98805 5.5099e-005 3.8182 0.012016 3.2596e-005 0.0011552 0.20672 0.00065907 0.20738 0.19068 0 0.033656 0.0389 0 1.0197 0.30497 0.086834 0.0117 5.1273 0.073015 8.9252e-005 0.81707 0.006024 0.0067856 0.0014333 0.98633 0.99131 3.0969e-006 1.2388e-005 0.13805 0.84279 0.86511 0.0014218 0.94069 0.52095 0.0019145 0.42491 1.6268 1.6249 16.0097 144.9768 0.00024516 -85.4519 0.37895
2.483 0.98805 5.5099e-005 3.8182 0.012016 3.2609e-005 0.0011552 0.20674 0.00065907 0.2074 0.1907 0 0.033655 0.0389 0 1.0198 0.30501 0.08685 0.011701 5.1282 0.073026 8.9267e-005 0.81706 0.0060247 0.0067864 0.001433 0.98634 0.99131 3.0961e-006 1.2384e-005 0.13805 0.84323 0.86536 0.0014216 0.94105 0.52112 0.0019142 0.42492 1.6279 1.626 16.0097 144.9768 0.00024477 -85.4534 0.37995
2.484 0.98805 5.5099e-005 3.8182 0.012016 3.2622e-005 0.0011552 0.20677 0.00065907 0.20742 0.19072 0 0.033654 0.0389 0 1.0199 0.30506 0.086866 0.011703 5.1292 0.073037 8.9282e-005 0.81705 0.0060253 0.0067871 0.0014326 0.98634 0.99131 3.0953e-006 1.2381e-005 0.13806 0.84367 0.8656 0.0014214 0.94141 0.52129 0.001914 0.42493 1.6289 1.6271 16.0097 144.9768 0.00024438 -85.4548 0.38095
2.485 0.98805 5.5098e-005 3.8182 0.012016 3.2635e-005 0.0011552 0.20679 0.00065907 0.20744 0.19074 0 0.033653 0.0389 0 1.02 0.3051 0.086881 0.011705 5.1301 0.073048 8.9296e-005 0.81704 0.006026 0.0067878 0.0014323 0.98635 0.99132 3.0944e-006 1.2378e-005 0.13806 0.84411 0.86585 0.0014212 0.94177 0.52145 0.0019138 0.42495 1.63 1.6282 16.0097 144.9769 0.000244 -85.4563 0.38195
2.486 0.98805 5.5098e-005 3.8182 0.012016 3.2649e-005 0.0011552 0.20681 0.00065907 0.20747 0.19076 0 0.033651 0.0389 0 1.0201 0.30514 0.086897 0.011707 5.1311 0.073059 8.9311e-005 0.81703 0.0060267 0.0067885 0.0014319 0.98635 0.99132 3.0936e-006 1.2375e-005 0.13807 0.84454 0.86609 0.001421 0.94212 0.52162 0.0019135 0.42496 1.6311 1.6292 16.0097 144.9769 0.00024361 -85.4578 0.38295
2.487 0.98805 5.5098e-005 3.8182 0.012016 3.2662e-005 0.0011552 0.20684 0.00065907 0.20749 0.19079 0 0.03365 0.0389 0 1.0202 0.30519 0.086913 0.011709 5.132 0.073071 8.9326e-005 0.81702 0.0060274 0.0067892 0.0014316 0.98636 0.99132 3.0929e-006 1.2371e-005 0.13807 0.84497 0.86634 0.0014209 0.94247 0.52178 0.0019133 0.42497 1.6321 1.6303 16.0097 144.9769 0.00024322 -85.4592 0.38395
2.488 0.98805 5.5098e-005 3.8182 0.012016 3.2675e-005 0.0011552 0.20686 0.00065907 0.20751 0.19081 0 0.033649 0.0389 0 1.0203 0.30523 0.086929 0.01171 5.133 0.073082 8.9341e-005 0.81701 0.0060281 0.00679 0.0014312 0.98636 0.99132 3.0921e-006 1.2368e-005 0.13808 0.84541 0.86658 0.0014207 0.94282 0.52195 0.0019131 0.42498 1.6332 1.6314 16.0097 144.9769 0.00024284 -85.4607 0.38495
2.489 0.98805 5.5098e-005 3.8182 0.012016 3.2688e-005 0.0011552 0.20688 0.00065907 0.20754 0.19083 0 0.033648 0.0389 0 1.0204 0.30528 0.086944 0.011712 5.1339 0.073093 8.9356e-005 0.817 0.0060288 0.0067907 0.0014309 0.98637 0.99133 3.0913e-006 1.2365e-005 0.13809 0.84584 0.86682 0.0014205 0.94317 0.52211 0.0019128 0.425 1.6343 1.6324 16.0097 144.9769 0.00024246 -85.4621 0.38595
2.49 0.98805 5.5098e-005 3.8182 0.012016 3.2701e-005 0.0011552 0.2069 0.00065907 0.20756 0.19085 0 0.033646 0.0389 0 1.0205 0.30532 0.08696 0.011714 5.1348 0.073104 8.9371e-005 0.81699 0.0060295 0.0067914 0.0014305 0.98637 0.99133 3.0905e-006 1.2362e-005 0.13809 0.84627 0.86706 0.0014203 0.94351 0.52228 0.0019126 0.42501 1.6353 1.6335 16.0097 144.9769 0.00024208 -85.4635 0.38695
2.491 0.98805 5.5098e-005 3.8182 0.012016 3.2714e-005 0.0011552 0.20693 0.00065907 0.20758 0.19087 0 0.033645 0.0389 0 1.0206 0.30536 0.086976 0.011716 5.1358 0.073115 8.9386e-005 0.81697 0.0060302 0.0067921 0.0014302 0.98637 0.99133 3.0897e-006 1.2359e-005 0.1381 0.84669 0.8673 0.0014201 0.94385 0.52244 0.0019124 0.42502 1.6364 1.6345 16.0097 144.977 0.0002417 -85.4649 0.38795
2.492 0.98805 5.5098e-005 3.8182 0.012016 3.2727e-005 0.0011552 0.20695 0.00065907 0.2076 0.19089 0 0.033644 0.0389 0 1.0207 0.30541 0.086992 0.011717 5.1367 0.073126 8.9401e-005 0.81696 0.0060308 0.0067929 0.0014299 0.98638 0.99134 3.089e-006 1.2356e-005 0.1381 0.84712 0.86754 0.0014199 0.94419 0.52261 0.0019121 0.42503 1.6374 1.6356 16.0097 144.977 0.00024132 -85.4663 0.38895
2.493 0.98805 5.5098e-005 3.8182 0.012016 3.274e-005 0.0011552 0.20697 0.00065907 0.20763 0.19092 0 0.033643 0.0389 0 1.0207 0.30545 0.087007 0.011719 5.1377 0.073138 8.9416e-005 0.81695 0.0060315 0.0067936 0.0014295 0.98638 0.99134 3.0882e-006 1.2353e-005 0.13811 0.84755 0.86778 0.0014198 0.94453 0.52277 0.0019119 0.42504 1.6385 1.6367 16.0097 144.977 0.00024095 -85.4677 0.38995
2.494 0.98805 5.5098e-005 3.8182 0.012016 3.2753e-005 0.0011552 0.207 0.00065907 0.20765 0.19094 0 0.033641 0.0389 0 1.0208 0.3055 0.087023 0.011721 5.1386 0.073149 8.943e-005 0.81694 0.0060322 0.0067943 0.0014292 0.98639 0.99134 3.0875e-006 1.235e-005 0.13811 0.84797 0.86802 0.0014196 0.94487 0.52294 0.0019117 0.42506 1.6395 1.6377 16.0097 144.977 0.00024057 -85.4691 0.39095
2.495 0.98805 5.5098e-005 3.8182 0.012016 3.2766e-005 0.0011552 0.20702 0.00065907 0.20767 0.19096 0 0.03364 0.0389 0 1.0209 0.30554 0.087039 0.011723 5.1396 0.07316 8.9445e-005 0.81693 0.0060329 0.006795 0.0014289 0.98639 0.99134 3.0867e-006 1.2347e-005 0.13812 0.84839 0.86825 0.0014194 0.9452 0.5231 0.0019115 0.42507 1.6406 1.6388 16.0097 144.977 0.0002402 -85.4705 0.39195
2.496 0.98805 5.5098e-005 3.8182 0.012016 3.2779e-005 0.0011552 0.20704 0.00065907 0.2077 0.19098 0 0.033639 0.0389 0 1.021 0.30558 0.087055 0.011725 5.1405 0.073171 8.946e-005 0.81692 0.0060336 0.0067957 0.0014286 0.9864 0.99135 3.086e-006 1.2344e-005 0.13813 0.84881 0.86849 0.0014192 0.94553 0.52327 0.0019112 0.42508 1.6416 1.6398 16.0097 144.9771 0.00023983 -85.4718 0.39295
2.497 0.98805 5.5098e-005 3.8182 0.012016 3.2792e-005 0.0011552 0.20706 0.00065907 0.20772 0.191 0 0.033638 0.0389 0 1.0211 0.30563 0.08707 0.011726 5.1415 0.073182 8.9475e-005 0.81691 0.0060343 0.0067965 0.0014282 0.9864 0.99135 3.0852e-006 1.2341e-005 0.13813 0.84924 0.86872 0.0014191 0.94586 0.52343 0.001911 0.42509 1.6426 1.6408 16.0097 144.9771 0.00023946 -85.4732 0.39395
2.498 0.98805 5.5098e-005 3.8182 0.012016 3.2805e-005 0.0011552 0.20709 0.00065907 0.20774 0.19102 0 0.033637 0.0389 0 1.0212 0.30567 0.087086 0.011728 5.1424 0.073194 8.949e-005 0.8169 0.006035 0.0067972 0.0014279 0.9864 0.99135 3.0845e-006 1.2338e-005 0.13814 0.84965 0.86896 0.0014189 0.94619 0.5236 0.0019108 0.42511 1.6437 1.6419 16.0097 144.9771 0.0002391 -85.4745 0.39495
2.499 0.98805 5.5098e-005 3.8182 0.012016 3.2819e-005 0.0011552 0.20711 0.00065907 0.20776 0.19104 0 0.033635 0.0389 0 1.0213 0.30572 0.087102 0.01173 5.1434 0.073205 8.9505e-005 0.81688 0.0060357 0.0067979 0.0014276 0.98641 0.99136 3.0838e-006 1.2335e-005 0.13814 0.85007 0.86919 0.0014188 0.94652 0.52376 0.0019106 0.42512 1.6447 1.6429 16.0097 144.9771 0.00023873 -85.4759 0.39595
2.5 0.98805 5.5097e-005 3.8182 0.012016 3.2832e-005 0.0011552 0.20713 0.00065907 0.20779 0.19107 0 0.033634 0.0389 0 1.0214 0.30576 0.087118 0.011732 5.1444 0.073216 8.952e-005 0.81687 0.0060364 0.0067986 0.0014273 0.98641 0.99136 3.083e-006 1.2332e-005 0.13815 0.85049 0.86942 0.0014186 0.94684 0.52393 0.0019104 0.42513 1.6457 1.6439 16.0097 144.9771 0.00023837 -85.4772 0.39695
2.501 0.98805 5.5097e-005 3.8182 0.012016 3.2845e-005 0.0011552 0.20715 0.00065907 0.20781 0.19109 0 0.033633 0.0389 0 1.0215 0.30581 0.087133 0.011734 5.1453 0.073227 8.9535e-005 0.81686 0.006037 0.0067994 0.001427 0.98642 0.99136 3.0823e-006 1.2329e-005 0.13815 0.8509 0.86965 0.0014184 0.94716 0.52409 0.0019102 0.42514 1.6467 1.645 16.0097 144.9772 0.000238 -85.4785 0.39795
2.502 0.98805 5.5097e-005 3.8182 0.012016 3.2858e-005 0.0011552 0.20718 0.00065907 0.20783 0.19111 0 0.033632 0.0389 0 1.0216 0.30585 0.087149 0.011735 5.1463 0.073238 8.955e-005 0.81685 0.0060377 0.0068001 0.0014267 0.98642 0.99136 3.0816e-006 1.2326e-005 0.13816 0.85132 0.86988 0.0014183 0.94748 0.52426 0.0019099 0.42516 1.6478 1.646 16.0097 144.9772 0.00023764 -85.4798 0.39895
2.503 0.98805 5.5097e-005 3.8182 0.012016 3.2871e-005 0.0011552 0.2072 0.00065907 0.20785 0.19113 0 0.033631 0.0389 0 1.0217 0.30589 0.087165 0.011737 5.1472 0.073249 8.9564e-005 0.81684 0.0060384 0.0068008 0.0014264 0.98642 0.99137 3.0809e-006 1.2324e-005 0.13816 0.85173 0.87011 0.0014181 0.9478 0.52442 0.0019097 0.42517 1.6488 1.647 16.0097 144.9772 0.00023728 -85.4811 0.39995
2.504 0.98805 5.5097e-005 3.8182 0.012016 3.2884e-005 0.0011552 0.20722 0.00065907 0.20788 0.19115 0 0.033629 0.0389 0 1.0218 0.30594 0.087181 0.011739 5.1482 0.073261 8.9579e-005 0.81683 0.0060391 0.0068015 0.0014261 0.98643 0.99137 3.0802e-006 1.2321e-005 0.13817 0.85214 0.87034 0.001418 0.94812 0.52459 0.0019095 0.42518 1.6498 1.6481 16.0097 144.9772 0.00023692 -85.4824 0.40095
2.505 0.98805 5.5097e-005 3.8182 0.012016 3.2897e-005 0.0011552 0.20724 0.00065907 0.2079 0.19117 0 0.033628 0.0389 0 1.0219 0.30598 0.087196 0.011741 5.1491 0.073272 8.9594e-005 0.81682 0.0060398 0.0068023 0.0014258 0.98643 0.99137 3.0795e-006 1.2318e-005 0.13818 0.85255 0.87056 0.0014178 0.94843 0.52475 0.0019093 0.42519 1.6508 1.6491 16.0097 144.9772 0.00023657 -85.4837 0.40195
2.506 0.98805 5.5097e-005 3.8182 0.012016 3.291e-005 0.0011552 0.20727 0.00065907 0.20792 0.19119 0 0.033627 0.0389 0 1.022 0.30603 0.087212 0.011743 5.1501 0.073283 8.9609e-005 0.81681 0.0060405 0.006803 0.0014254 0.98644 0.99137 3.0788e-006 1.2315e-005 0.13818 0.85296 0.87079 0.0014177 0.94874 0.52492 0.0019091 0.4252 1.6518 1.6501 16.0097 144.9773 0.00023621 -85.4849 0.40295
2.507 0.98805 5.5097e-005 3.8182 0.012016 3.2923e-005 0.0011553 0.20729 0.00065908 0.20794 0.19121 0 0.033626 0.0389 0 1.0221 0.30607 0.087228 0.011744 5.151 0.073294 8.9624e-005 0.8168 0.0060412 0.0068037 0.0014251 0.98644 0.99138 3.0781e-006 1.2312e-005 0.13819 0.85336 0.87101 0.0014175 0.94905 0.52508 0.0019089 0.42522 1.6528 1.6511 16.0097 144.9773 0.00023586 -85.4862 0.40395
2.508 0.98805 5.5097e-005 3.8182 0.012016 3.2936e-005 0.0011553 0.20731 0.00065908 0.20797 0.19124 0 0.033624 0.0389 0 1.0222 0.30612 0.087244 0.011746 5.152 0.073305 8.9639e-005 0.81678 0.0060419 0.0068044 0.0014248 0.98644 0.99138 3.0774e-006 1.231e-005 0.13819 0.85377 0.87124 0.0014173 0.94936 0.52525 0.0019087 0.42523 1.6538 1.6521 16.0097 144.9773 0.0002355 -85.4875 0.40495
2.509 0.98805 5.5097e-005 3.8182 0.012016 3.2949e-005 0.0011553 0.20733 0.00065908 0.20799 0.19126 0 0.033623 0.0389 0 1.0223 0.30616 0.087259 0.011748 5.1529 0.073317 8.9654e-005 0.81677 0.0060426 0.0068052 0.0014245 0.98645 0.99138 3.0768e-006 1.2307e-005 0.1382 0.85418 0.87146 0.0014172 0.94967 0.52541 0.0019085 0.42524 1.6548 1.6531 16.0097 144.9773 0.00023515 -85.4887 0.40595
2.51 0.98805 5.5097e-005 3.8182 0.012016 3.2962e-005 0.0011553 0.20736 0.00065908 0.20801 0.19128 0 0.033622 0.0389 0 1.0224 0.3062 0.087275 0.01175 5.1539 0.073328 8.9669e-005 0.81676 0.0060433 0.0068059 0.0014243 0.98645 0.99138 3.0761e-006 1.2304e-005 0.1382 0.85458 0.87168 0.001417 0.94997 0.52558 0.0019083 0.42525 1.6558 1.6541 16.0097 144.9773 0.0002348 -85.4899 0.40695
2.511 0.98805 5.5097e-005 3.8182 0.012016 3.2975e-005 0.0011553 0.20738 0.00065908 0.20803 0.1913 0 0.033621 0.0389 0 1.0225 0.30625 0.087291 0.011751 5.1549 0.073339 8.9684e-005 0.81675 0.0060439 0.0068066 0.001424 0.98646 0.99139 3.0754e-006 1.2302e-005 0.13821 0.85498 0.8719 0.0014169 0.95027 0.52574 0.0019081 0.42527 1.6568 1.6551 16.0097 144.9773 0.00023446 -85.4912 0.40795
2.512 0.98805 5.5097e-005 3.8182 0.012016 3.2989e-005 0.0011553 0.2074 0.00065908 0.20806 0.19132 0 0.03362 0.0389 0 1.0226 0.30629 0.087307 0.011753 5.1558 0.07335 8.9699e-005 0.81674 0.0060446 0.0068073 0.0014237 0.98646 0.99139 3.0748e-006 1.2299e-005 0.13822 0.85538 0.87212 0.0014167 0.95057 0.5259 0.0019079 0.42528 1.6578 1.6561 16.0097 144.9774 0.00023411 -85.4924 0.40895
2.513 0.98805 5.5097e-005 3.8182 0.012016 3.3002e-005 0.0011553 0.20742 0.00065908 0.20808 0.19134 0 0.033618 0.0389 0 1.0227 0.30634 0.087322 0.011755 5.1568 0.073361 8.9713e-005 0.81673 0.0060453 0.0068081 0.0014234 0.98646 0.99139 3.0741e-006 1.2296e-005 0.13822 0.85578 0.87234 0.0014166 0.95087 0.52607 0.0019077 0.42529 1.6588 1.6571 16.0097 144.9774 0.00023376 -85.4936 0.40995
2.514 0.98805 5.5097e-005 3.8182 0.012016 3.3015e-005 0.0011553 0.20745 0.00065908 0.2081 0.19136 0 0.033617 0.0389 0 1.0228 0.30638 0.087338 0.011757 5.1577 0.073372 8.9728e-005 0.81672 0.006046 0.0068088 0.0014231 0.98647 0.99139 3.0734e-006 1.2294e-005 0.13823 0.85618 0.87256 0.0014164 0.95117 0.52623 0.0019075 0.4253 1.6598 1.6581 16.0097 144.9774 0.00023342 -85.4948 0.41095
2.515 0.98805 5.5096e-005 3.8182 0.012016 3.3028e-005 0.0011553 0.20747 0.00065908 0.20812 0.19138 0 0.033616 0.0389 0 1.0229 0.30642 0.087354 0.011759 5.1587 0.073384 8.9743e-005 0.81671 0.0060467 0.0068095 0.0014228 0.98647 0.9914 3.0728e-006 1.2291e-005 0.13823 0.85658 0.87278 0.0014163 0.95146 0.5264 0.0019073 0.42532 1.6608 1.6591 16.0096 144.9774 0.00023308 -85.496 0.41195
2.516 0.98805 5.5096e-005 3.8182 0.012016 3.3041e-005 0.0011553 0.20749 0.00065908 0.20815 0.19141 0 0.033615 0.0389 0 1.023 0.30647 0.08737 0.01176 5.1596 0.073395 8.9758e-005 0.81669 0.0060474 0.0068102 0.0014225 0.98647 0.9914 3.0722e-006 1.2289e-005 0.13824 0.85697 0.87299 0.0014161 0.95175 0.52656 0.0019071 0.42533 1.6618 1.6601 16.0096 144.9774 0.00023274 -85.4972 0.41295
2.517 0.98805 5.5096e-005 3.8182 0.012016 3.3054e-005 0.0011553 0.20751 0.00065908 0.20817 0.19143 0 0.033614 0.0389 0 1.0231 0.30651 0.087386 0.011762 5.1606 0.073406 8.9773e-005 0.81668 0.0060481 0.006811 0.0014223 0.98648 0.9914 3.0715e-006 1.2286e-005 0.13824 0.85737 0.87321 0.001416 0.95204 0.52672 0.0019069 0.42534 1.6628 1.6611 16.0096 144.9775 0.0002324 -85.4983 0.41395
2.518 0.98805 5.5096e-005 3.8182 0.012016 3.3067e-005 0.0011553 0.20754 0.00065908 0.20819 0.19145 0 0.033612 0.0389 0 1.0232 0.30656 0.087401 0.011764 5.1616 0.073417 8.9788e-005 0.81667 0.0060488 0.0068117 0.001422 0.98648 0.9914 3.0709e-006 1.2283e-005 0.13825 0.85776 0.87342 0.0014158 0.95233 0.52689 0.0019067 0.42535 1.6637 1.6621 16.0096 144.9775 0.00023206 -85.4995 0.41495
2.519 0.98805 5.5096e-005 3.8182 0.012016 3.308e-005 0.0011553 0.20756 0.00065908 0.20821 0.19147 0 0.033611 0.0389 0 1.0233 0.3066 0.087417 0.011766 5.1625 0.073428 8.9803e-005 0.81666 0.0060495 0.0068124 0.0014217 0.98649 0.99141 3.0703e-006 1.2281e-005 0.13826 0.85815 0.87364 0.0014157 0.95262 0.52705 0.0019066 0.42537 1.6647 1.6631 16.0096 144.9775 0.00023172 -85.5007 0.41595
2.52 0.98805 5.5096e-005 3.8182 0.012016 3.3093e-005 0.0011553 0.20758 0.00065908 0.20823 0.19149 0 0.03361 0.0389 0 1.0234 0.30665 0.087433 0.011768 5.1635 0.07344 8.9818e-005 0.81665 0.0060502 0.0068131 0.0014214 0.98649 0.99141 3.0696e-006 1.2278e-005 0.13826 0.85855 0.87385 0.0014155 0.95291 0.52722 0.0019064 0.42538 1.6657 1.664 16.0096 144.9775 0.00023139 -85.5018 0.41695
2.521 0.98805 5.5096e-005 3.8182 0.012016 3.3106e-005 0.0011553 0.2076 0.00065908 0.20826 0.19151 0 0.033609 0.0389 0 1.0235 0.30669 0.087449 0.011769 5.1644 0.073451 8.9833e-005 0.81664 0.0060509 0.0068139 0.0014212 0.98649 0.99141 3.069e-006 1.2276e-005 0.13827 0.85894 0.87406 0.0014154 0.95319 0.52738 0.0019062 0.42539 1.6667 1.665 16.0096 144.9775 0.00023105 -85.503 0.41795
2.522 0.98805 5.5096e-005 3.8182 0.012016 3.3119e-005 0.0011553 0.20762 0.00065908 0.20828 0.19153 0 0.033608 0.0389 0 1.0236 0.30673 0.087464 0.011771 5.1654 0.073462 8.9848e-005 0.81663 0.0060515 0.0068146 0.0014209 0.9865 0.99141 3.0684e-006 1.2274e-005 0.13827 0.85932 0.87427 0.0014153 0.95347 0.52754 0.001906 0.4254 1.6676 1.666 16.0096 144.9776 0.00023072 -85.5041 0.41895
2.523 0.98805 5.5096e-005 3.8182 0.012016 3.3132e-005 0.0011553 0.20765 0.00065908 0.2083 0.19155 0 0.033606 0.0389 0 1.0237 0.30678 0.08748 0.011773 5.1664 0.073473 8.9862e-005 0.81662 0.0060522 0.0068153 0.0014206 0.9865 0.99142 3.0678e-006 1.2271e-005 0.13828 0.85971 0.87448 0.0014151 0.95375 0.52771 0.0019058 0.42542 1.6686 1.667 16.0096 144.9776 0.00023039 -85.5052 0.41995
2.524 0.98805 5.5096e-005 3.8182 0.012016 3.3145e-005 0.0011553 0.20767 0.00065908 0.20832 0.19157 0 0.033605 0.0389 0 1.0238 0.30682 0.087496 0.011775 5.1673 0.073484 8.9877e-005 0.81661 0.0060529 0.006816 0.0014204 0.9865 0.99142 3.0672e-006 1.2269e-005 0.13828 0.8601 0.87469 0.001415 0.95403 0.52787 0.0019056 0.42543 1.6696 1.6679 16.0096 144.9776 0.00023006 -85.5064 0.42095
2.525 0.98805 5.5096e-005 3.8182 0.012016 3.3159e-005 0.0011553 0.20769 0.00065908 0.20835 0.1916 0 0.033604 0.0389 0 1.0239 0.30687 0.087512 0.011776 5.1683 0.073495 8.9892e-005 0.81659 0.0060536 0.0068168 0.0014201 0.98651 0.99142 3.0666e-006 1.2266e-005 0.13829 0.86048 0.8749 0.0014149 0.95431 0.52803 0.0019055 0.42544 1.6705 1.6689 16.0096 144.9776 0.00022973 -85.5075 0.42195
2.526 0.98805 5.5096e-005 3.8182 0.012016 3.3172e-005 0.0011553 0.20771 0.00065908 0.20837 0.19162 0 0.033603 0.0389 0 1.024 0.30691 0.087527 0.011778 5.1693 0.073507 8.9907e-005 0.81658 0.0060543 0.0068175 0.0014198 0.98651 0.99142 3.066e-006 1.2264e-005 0.13829 0.86087 0.87511 0.0014147 0.95458 0.5282 0.0019053 0.42545 1.6715 1.6699 16.0096 144.9776 0.0002294 -85.5086 0.42295
2.527 0.98805 5.5096e-005 3.8182 0.012016 3.3185e-005 0.0011553 0.20774 0.00065908 0.20839 0.19164 0 0.033602 0.0389 0 1.024 0.30696 0.087543 0.01178 5.1702 0.073518 8.9922e-005 0.81657 0.006055 0.0068182 0.0014196 0.98651 0.99142 3.0654e-006 1.2261e-005 0.1383 0.86125 0.87532 0.0014146 0.95486 0.52836 0.0019051 0.42547 1.6724 1.6708 16.0096 144.9777 0.00022908 -85.5097 0.42395
2.528 0.98805 5.5096e-005 3.8182 0.012016 3.3198e-005 0.0011553 0.20776 0.00065908 0.20841 0.19166 0 0.0336 0.0389 0 1.0241 0.307 0.087559 0.011782 5.1712 0.073529 8.9937e-005 0.81656 0.0060557 0.0068189 0.0014193 0.98652 0.99143 3.0648e-006 1.2259e-005 0.13831 0.86163 0.87552 0.0014144 0.95513 0.52853 0.0019049 0.42548 1.6734 1.6718 16.0096 144.9777 0.00022875 -85.5108 0.42495
2.529 0.98805 5.5096e-005 3.8182 0.012016 3.3211e-005 0.0011553 0.20778 0.00065908 0.20843 0.19168 0 0.033599 0.0389 0 1.0242 0.30704 0.087575 0.011784 5.1721 0.07354 8.9952e-005 0.81655 0.0060564 0.0068197 0.0014191 0.98652 0.99143 3.0642e-006 1.2257e-005 0.13831 0.86201 0.87573 0.0014143 0.9554 0.52869 0.0019048 0.42549 1.6743 1.6727 16.0096 144.9777 0.00022843 -85.5118 0.42595
2.53 0.98805 5.5095e-005 3.8182 0.012015 3.3224e-005 0.0011553 0.2078 0.00065908 0.20846 0.1917 0 0.033598 0.0389 0 1.0243 0.30709 0.087591 0.011785 5.1731 0.073551 8.9967e-005 0.81654 0.0060571 0.0068204 0.0014188 0.98652 0.99143 3.0636e-006 1.2254e-005 0.13832 0.86239 0.87593 0.0014141 0.95566 0.52885 0.0019046 0.4255 1.6753 1.6737 16.0096 144.9777 0.00022811 -85.5129 0.42695
2.531 0.98805 5.5095e-005 3.8182 0.012015 3.3237e-005 0.0011553 0.20782 0.00065908 0.20848 0.19172 0 0.033597 0.0389 0 1.0244 0.30713 0.087606 0.011787 5.1741 0.073563 8.9982e-005 0.81653 0.0060578 0.0068211 0.0014186 0.98653 0.99143 3.063e-006 1.2252e-005 0.13832 0.86277 0.87614 0.001414 0.95593 0.52902 0.0019044 0.42552 1.6762 1.6746 16.0096 144.9777 0.00022779 -85.514 0.42795
2.532 0.98805 5.5095e-005 3.8182 0.012015 3.325e-005 0.0011553 0.20785 0.00065908 0.2085 0.19174 0 0.033596 0.0389 0 1.0245 0.30718 0.087622 0.011789 5.175 0.073574 8.9997e-005 0.81652 0.0060585 0.0068219 0.0014183 0.98653 0.99143 3.0625e-006 1.225e-005 0.13833 0.86314 0.87634 0.0014139 0.9562 0.52918 0.0019042 0.42553 1.6772 1.6756 16.0096 144.9778 0.00022747 -85.515 0.42895
2.533 0.98805 5.5095e-005 3.8182 0.012015 3.3263e-005 0.0011553 0.20787 0.00065908 0.20852 0.19176 0 0.033595 0.0389 0 1.0246 0.30722 0.087638 0.011791 5.176 0.073585 9.0012e-005 0.81651 0.0060592 0.0068226 0.0014181 0.98653 0.99144 3.0619e-006 1.2248e-005 0.13833 0.86352 0.87654 0.0014138 0.95646 0.52934 0.0019041 0.42554 1.6781 1.6765 16.0096 144.9778 0.00022715 -85.5161 0.42995
2.534 0.98805 5.5095e-005 3.8182 0.012015 3.3276e-005 0.0011553 0.20789 0.00065908 0.20854 0.19178 0 0.033593 0.0389 0 1.0247 0.30727 0.087654 0.011793 5.177 0.073596 9.0026e-005 0.81649 0.0060598 0.0068233 0.0014178 0.98654 0.99144 3.0613e-006 1.2245e-005 0.13834 0.86389 0.87674 0.0014136 0.95672 0.5295 0.0019039 0.42556 1.6791 1.6775 16.0096 144.9778 0.00022683 -85.5171 0.43095
2.535 0.98805 5.5095e-005 3.8182 0.012015 3.3289e-005 0.0011553 0.20791 0.00065908 0.20857 0.1918 0 0.033592 0.0389 0 1.0248 0.30731 0.08767 0.011794 5.1779 0.073607 9.0041e-005 0.81648 0.0060605 0.006824 0.0014176 0.98654 0.99144 3.0608e-006 1.2243e-005 0.13835 0.86427 0.87694 0.0014135 0.95698 0.52967 0.0019037 0.42557 1.68 1.6784 16.0095 144.9778 0.00022652 -85.5182 0.43195
2.536 0.98805 5.5095e-005 3.8182 0.012015 3.3302e-005 0.0011553 0.20793 0.00065908 0.20859 0.19182 0 0.033591 0.0389 0 1.0249 0.30735 0.087685 0.011796 5.1789 0.073618 9.0056e-005 0.81647 0.0060612 0.0068248 0.0014173 0.98654 0.99144 3.0602e-006 1.2241e-005 0.13835 0.86464 0.87714 0.0014134 0.95724 0.52983 0.0019036 0.42558 1.6809 1.6794 16.0095 144.9778 0.0002262 -85.5192 0.43295
2.537 0.98805 5.5095e-005 3.8182 0.012015 3.3315e-005 0.0011553 0.20796 0.00065908 0.20861 0.19185 0 0.03359 0.0389 0 1.025 0.3074 0.087701 0.011798 5.1799 0.07363 9.0071e-005 0.81646 0.0060619 0.0068255 0.0014171 0.98655 0.99145 3.0596e-006 1.2239e-005 0.13836 0.86501 0.87734 0.0014133 0.95749 0.52999 0.0019034 0.42559 1.6819 1.6803 16.0095 144.9779 0.00022589 -85.5202 0.43395
2.538 0.98805 5.5095e-005 3.8182 0.012015 3.3329e-005 0.0011553 0.20798 0.00065908 0.20863 0.19187 0 0.033589 0.0389 0 1.0251 0.30744 0.087717 0.0118 5.1808 0.073641 9.0086e-005 0.81645 0.0060626 0.0068262 0.0014168 0.98655 0.99145 3.0591e-006 1.2236e-005 0.13836 0.86538 0.87754 0.0014131 0.95775 0.53016 0.0019032 0.42561 1.6828 1.6812 16.0095 144.9779 0.00022558 -85.5212 0.43495
2.539 0.98805 5.5095e-005 3.8182 0.012015 3.3342e-005 0.0011553 0.208 0.00065908 0.20865 0.19189 0 0.033587 0.0389 0 1.0252 0.30749 0.087733 0.011802 5.1818 0.073652 9.0101e-005 0.81644 0.0060633 0.006827 0.0014166 0.98655 0.99145 3.0585e-006 1.2234e-005 0.13837 0.86575 0.87774 0.001413 0.958 0.53032 0.0019031 0.42562 1.6837 1.6821 16.0095 144.9779 0.00022527 -85.5223 0.43595
2.54 0.98805 5.5095e-005 3.8182 0.012015 3.3355e-005 0.0011553 0.20802 0.00065908 0.20868 0.19191 0 0.033586 0.0389 0 1.0253 0.30753 0.087748 0.011803 5.1828 0.073663 9.0116e-005 0.81643 0.006064 0.0068277 0.0014164 0.98655 0.99145 3.058e-006 1.2232e-005 0.13837 0.86612 0.87793 0.0014129 0.95825 0.53048 0.0019029 0.42563 1.6846 1.6831 16.0095 144.9779 0.00022496 -85.5233 0.43695
2.541 0.98805 5.5095e-005 3.8182 0.012015 3.3368e-005 0.0011553 0.20804 0.00065908 0.2087 0.19193 0 0.033585 0.0389 0 1.0254 0.30758 0.087764 0.011805 5.1838 0.073674 9.0131e-005 0.81642 0.0060647 0.0068284 0.0014161 0.98656 0.99145 3.0575e-006 1.223e-005 0.13838 0.86648 0.87813 0.0014128 0.9585 0.53065 0.0019027 0.42564 1.6856 1.684 16.0095 144.9779 0.00022465 -85.5243 0.43795
2.542 0.98805 5.5095e-005 3.8182 0.012015 3.3381e-005 0.0011553 0.20807 0.00065908 0.20872 0.19195 0 0.033584 0.0389 0 1.0255 0.30762 0.08778 0.011807 5.1847 0.073686 9.0146e-005 0.8164 0.0060654 0.0068291 0.0014159 0.98656 0.99146 3.0569e-006 1.2228e-005 0.13839 0.86685 0.87832 0.0014126 0.95875 0.53081 0.0019026 0.42566 1.6865 1.6849 16.0095 144.9779 0.00022434 -85.5252 0.43895
2.543 0.98805 5.5095e-005 3.8182 0.012015 3.3394e-005 0.0011553 0.20809 0.00065908 0.20874 0.19197 0 0.033583 0.0389 0 1.0256 0.30766 0.087796 0.011809 5.1857 0.073697 9.0161e-005 0.81639 0.0060661 0.0068299 0.0014157 0.98656 0.99146 3.0564e-006 1.2226e-005 0.13839 0.86721 0.87852 0.0014125 0.959 0.53097 0.0019024 0.42567 1.6874 1.6858 16.0095 144.978 0.00022404 -85.5262 0.43995
2.544 0.98805 5.5095e-005 3.8182 0.012015 3.3407e-005 0.0011553 0.20811 0.00065908 0.20876 0.19199 0 0.033582 0.0389 0 1.0257 0.30771 0.087812 0.01181 5.1867 0.073708 9.0176e-005 0.81638 0.0060668 0.0068306 0.0014154 0.98657 0.99146 3.0559e-006 1.2223e-005 0.1384 0.86758 0.87871 0.0014124 0.95924 0.53113 0.0019023 0.42568 1.6883 1.6868 16.0095 144.978 0.00022373 -85.5272 0.44095
2.545 0.98805 5.5094e-005 3.8182 0.012015 3.342e-005 0.0011553 0.20813 0.00065908 0.20879 0.19201 0 0.03358 0.0389 0 1.0258 0.30775 0.087827 0.011812 5.1876 0.073719 9.019e-005 0.81637 0.0060675 0.0068313 0.0014152 0.98657 0.99146 3.0553e-006 1.2221e-005 0.1384 0.86794 0.8789 0.0014123 0.95949 0.5313 0.0019021 0.42569 1.6892 1.6877 16.0095 144.978 0.00022343 -85.5282 0.44195
2.546 0.98805 5.5094e-005 3.8182 0.012015 3.3433e-005 0.0011553 0.20815 0.00065908 0.20881 0.19203 0 0.033579 0.0389 0 1.0259 0.3078 0.087843 0.011814 5.1886 0.07373 9.0205e-005 0.81636 0.0060682 0.0068321 0.001415 0.98657 0.99146 3.0548e-006 1.2219e-005 0.13841 0.8683 0.8791 0.0014122 0.95973 0.53146 0.001902 0.42571 1.6901 1.6886 16.0095 144.978 0.00022313 -85.5291 0.44295
2.547 0.98805 5.5094e-005 3.8182 0.012015 3.3446e-005 0.0011553 0.20817 0.00065908 0.20883 0.19205 0 0.033578 0.0389 0 1.026 0.30784 0.087859 0.011816 5.1896 0.073741 9.022e-005 0.81635 0.0060689 0.0068328 0.0014148 0.98658 0.99147 3.0543e-006 1.2217e-005 0.13841 0.86866 0.87929 0.0014121 0.95997 0.53162 0.0019018 0.42572 1.691 1.6895 16.0095 144.978 0.00022283 -85.5301 0.44395
2.548 0.98805 5.5094e-005 3.8182 0.012015 3.3459e-005 0.0011553 0.2082 0.00065908 0.20885 0.19207 0 0.033577 0.0389 0 1.0261 0.30789 0.087875 0.011818 5.1906 0.073753 9.0235e-005 0.81634 0.0060696 0.0068335 0.0014145 0.98658 0.99147 3.0538e-006 1.2215e-005 0.13842 0.86902 0.87948 0.001412 0.96021 0.53178 0.0019016 0.42573 1.6919 1.6904 16.0095 144.9781 0.00022253 -85.531 0.44495
2.549 0.98805 5.5094e-005 3.8182 0.012015 3.3472e-005 0.0011553 0.20822 0.00065908 0.20887 0.19209 0 0.033576 0.0389 0 1.0262 0.30793 0.087891 0.011819 5.1915 0.073764 9.025e-005 0.81633 0.0060702 0.0068342 0.0014143 0.98658 0.99147 3.0533e-006 1.2213e-005 0.13843 0.86937 0.87967 0.0014118 0.96045 0.53195 0.0019015 0.42574 1.6928 1.6913 16.0095 144.9781 0.00022223 -85.532 0.44595
2.55 0.98805 5.5094e-005 3.8182 0.012015 3.3485e-005 0.0011553 0.20824 0.00065908 0.20889 0.19211 0 0.033575 0.0389 0 1.0263 0.30798 0.087906 0.011821 5.1925 0.073775 9.0265e-005 0.81632 0.0060709 0.006835 0.0014141 0.98658 0.99147 3.0528e-006 1.2211e-005 0.13843 0.86973 0.87986 0.0014117 0.96068 0.53211 0.0019013 0.42576 1.6937 1.6922 16.0094 144.9781 0.00022194 -85.5329 0.44695
2.551 0.98805 5.5094e-005 3.8182 0.012015 3.3499e-005 0.0011553 0.20826 0.00065908 0.20892 0.19213 0 0.033573 0.0389 0 1.0264 0.30802 0.087922 0.011823 5.1935 0.073786 9.028e-005 0.8163 0.0060716 0.0068357 0.0014139 0.98659 0.99147 3.0523e-006 1.2209e-005 0.13844 0.87008 0.88004 0.0014116 0.96092 0.53227 0.0019012 0.42577 1.6946 1.6931 16.0094 144.9781 0.00022164 -85.5338 0.44795
2.552 0.98805 5.5094e-005 3.8182 0.012015 3.3512e-005 0.0011553 0.20828 0.00065909 0.20894 0.19216 0 0.033572 0.0389 0 1.0265 0.30806 0.087938 0.011825 5.1944 0.073797 9.0295e-005 0.81629 0.0060723 0.0068364 0.0014136 0.98659 0.99147 3.0518e-006 1.2207e-005 0.13844 0.87044 0.88023 0.0014114 0.96115 0.53243 0.001901 0.42578 1.6955 1.694 16.0094 144.9781 0.00022135 -85.5348 0.44895
2.553 0.98805 5.5094e-005 3.8182 0.012015 3.3525e-005 0.0011553 0.2083 0.00065909 0.20896 0.19218 0 0.033571 0.0389 0 1.0266 0.30811 0.087954 0.011827 5.1954 0.073808 9.031e-005 0.81628 0.006073 0.0068372 0.0014134 0.98659 0.99148 3.0513e-006 1.2205e-005 0.13845 0.87079 0.88042 0.0014113 0.96138 0.53259 0.0019009 0.4258 1.6964 1.6949 16.0094 144.9782 0.00022105 -85.5357 0.44995
2.554 0.98805 5.5094e-005 3.8182 0.012015 3.3538e-005 0.0011553 0.20833 0.00065909 0.20898 0.1922 0 0.03357 0.0389 0 1.0267 0.30815 0.08797 0.011828 5.1964 0.07382 9.0325e-005 0.81627 0.0060737 0.0068379 0.0014132 0.9866 0.99148 3.0508e-006 1.2203e-005 0.13845 0.87114 0.8806 0.0014112 0.96161 0.53276 0.0019007 0.42581 1.6973 1.6958 16.0094 144.9782 0.00022076 -85.5366 0.45095
2.555 0.98805 5.5094e-005 3.8182 0.012015 3.3551e-005 0.0011553 0.20835 0.00065909 0.209 0.19222 0 0.033569 0.0389 0 1.0268 0.3082 0.087985 0.01183 5.1974 0.073831 9.034e-005 0.81626 0.0060744 0.0068386 0.001413 0.9866 0.99148 3.0503e-006 1.2201e-005 0.13846 0.87149 0.88079 0.0014111 0.96184 0.53292 0.0019006 0.42582 1.6982 1.6967 16.0094 144.9782 0.00022047 -85.5375 0.45195
2.556 0.98805 5.5094e-005 3.8182 0.012015 3.3564e-005 0.0011553 0.20837 0.00065909 0.20902 0.19224 0 0.033568 0.0389 0 1.0269 0.30824 0.088001 0.011832 5.1983 0.073842 9.0354e-005 0.81625 0.0060751 0.0068393 0.0014128 0.9866 0.99148 3.0498e-006 1.2199e-005 0.13846 0.87184 0.88097 0.0014109 0.96207 0.53308 0.0019005 0.42583 1.6991 1.6976 16.0094 144.9782 0.00022018 -85.5384 0.45295
2.557 0.98805 5.5094e-005 3.8182 0.012015 3.3577e-005 0.0011553 0.20839 0.00065909 0.20905 0.19226 0 0.033566 0.0389 0 1.027 0.30829 0.088017 0.011834 5.1993 0.073853 9.0369e-005 0.81624 0.0060758 0.0068401 0.0014126 0.9866 0.99148 3.0493e-006 1.2197e-005 0.13847 0.87219 0.88116 0.0014108 0.9623 0.53324 0.0019003 0.42585 1.7 1.6985 16.0094 144.9782 0.00021989 -85.5393 0.45395
2.558 0.98805 5.5094e-005 3.8182 0.012015 3.359e-005 0.0011553 0.20841 0.00065909 0.20907 0.19228 0 0.033565 0.0389 0 1.0271 0.30833 0.088033 0.011835 5.2003 0.073864 9.0384e-005 0.81623 0.0060765 0.0068408 0.0014124 0.98661 0.99149 3.0489e-006 1.2195e-005 0.13848 0.87254 0.88134 0.0014107 0.96252 0.53341 0.0019002 0.42586 1.7008 1.6994 16.0094 144.9783 0.0002196 -85.5402 0.45495
2.559 0.98805 5.5094e-005 3.8182 0.012015 3.3603e-005 0.0011553 0.20843 0.00065909 0.20909 0.1923 0 0.033564 0.0389 0 1.0272 0.30837 0.088049 0.011837 5.2013 0.073876 9.0399e-005 0.81621 0.0060772 0.0068415 0.0014122 0.98661 0.99149 3.0484e-006 1.2194e-005 0.13848 0.87289 0.88152 0.0014106 0.96274 0.53357 0.0019 0.42587 1.7017 1.7003 16.0094 144.9783 0.00021932 -85.541 0.45595
2.56 0.98805 5.5093e-005 3.8182 0.012015 3.3616e-005 0.0011553 0.20846 0.00065909 0.20911 0.19232 0 0.033563 0.0389 0 1.0273 0.30842 0.088064 0.011839 5.2023 0.073887 9.0414e-005 0.8162 0.0060779 0.0068423 0.001412 0.98661 0.99149 3.0479e-006 1.2192e-005 0.13849 0.87323 0.8817 0.0014106 0.96296 0.53373 0.0018999 0.42588 1.7026 1.7011 16.0094 144.9783 0.00021903 -85.5419 0.45695
2.561 0.98805 5.5093e-005 3.8182 0.012015 3.3629e-005 0.0011553 0.20848 0.00065909 0.20913 0.19234 0 0.033562 0.0389 0 1.0274 0.30846 0.08808 0.011841 5.2032 0.073898 9.0429e-005 0.81619 0.0060786 0.006843 0.0014118 0.98661 0.99149 3.0475e-006 1.219e-005 0.13849 0.87358 0.88188 0.0014105 0.96318 0.53389 0.0018998 0.4259 1.7035 1.702 16.0093 144.9783 0.00021875 -85.5428 0.45795
2.562 0.98805 5.5093e-005 3.8182 0.012015 3.3642e-005 0.0011553 0.2085 0.00065909 0.20915 0.19236 0 0.033561 0.0389 0 1.0275 0.30851 0.088096 0.011843 5.2042 0.073909 9.0444e-005 0.81618 0.0060793 0.0068437 0.0014116 0.98662 0.99149 3.047e-006 1.2188e-005 0.1385 0.87392 0.88206 0.0014104 0.9634 0.53405 0.0018996 0.42591 1.7043 1.7029 16.0093 144.9783 0.00021846 -85.5437 0.45895
2.563 0.98805 5.5093e-005 3.8182 0.012015 3.3655e-005 0.0011553 0.20852 0.00065909 0.20917 0.19238 0 0.03356 0.0389 0 1.0275 0.30855 0.088112 0.011844 5.2052 0.07392 9.0459e-005 0.81617 0.00608 0.0068445 0.0014114 0.98662 0.99149 3.0465e-006 1.2186e-005 0.1385 0.87426 0.88224 0.0014103 0.96362 0.53421 0.0018995 0.42592 1.7052 1.7038 16.0093 144.9784 0.00021818 -85.5445 0.45995
2.564 0.98805 5.5093e-005 3.8182 0.012015 3.3668e-005 0.0011553 0.20854 0.00065909 0.2092 0.1924 0 0.033558 0.0389 0 1.0276 0.3086 0.088128 0.011846 5.2062 0.073931 9.0474e-005 0.81616 0.0060807 0.0068452 0.0014112 0.98662 0.9915 3.0461e-006 1.2184e-005 0.13851 0.8746 0.88242 0.0014102 0.96384 0.53438 0.0018993 0.42594 1.7061 1.7046 16.0093 144.9784 0.0002179 -85.5454 0.46095
2.565 0.98805 5.5093e-005 3.8182 0.012015 3.3682e-005 0.0011553 0.20856 0.00065909 0.20922 0.19242 0 0.033557 0.0389 0 1.0277 0.30864 0.088143 0.011848 5.2071 0.073943 9.0489e-005 0.81615 0.0060814 0.0068459 0.001411 0.98662 0.9915 3.0456e-006 1.2182e-005 0.13852 0.87494 0.8826 0.0014101 0.96405 0.53454 0.0018992 0.42595 1.7069 1.7055 16.0093 144.9784 0.00021762 -85.5462 0.46195
2.566 0.98805 5.5093e-005 3.8182 0.012015 3.3695e-005 0.0011553 0.20858 0.00065909 0.20924 0.19244 0 0.033556 0.0389 0 1.0278 0.30868 0.088159 0.01185 5.2081 0.073954 9.0504e-005 0.81614 0.0060821 0.0068467 0.0014108 0.98663 0.9915 3.0452e-006 1.2181e-005 0.13852 0.87528 0.88278 0.00141 0.96427 0.5347 0.0018991 0.42596 1.7078 1.7064 16.0093 144.9784 0.00021734 -85.547 0.46295
2.567 0.98805 5.5093e-005 3.8182 0.012015 3.3708e-005 0.0011553 0.20861 0.00065909 0.20926 0.19246 0 0.033555 0.0389 0 1.0279 0.30873 0.088175 0.011852 5.2091 0.073965 9.0519e-005 0.81613 0.0060828 0.0068474 0.0014106 0.98663 0.9915 3.0447e-006 1.2179e-005 0.13853 0.87562 0.88295 0.0014099 0.96448 0.53486 0.0018989 0.42597 1.7087 1.7072 16.0093 144.9784 0.00021707 -85.5479 0.46395
2.568 0.98805 5.5093e-005 3.8182 0.012015 3.3721e-005 0.0011553 0.20863 0.00065909 0.20928 0.19248 0 0.033554 0.0389 0 1.028 0.30877 0.088191 0.011853 5.2101 0.073976 9.0533e-005 0.81611 0.0060835 0.0068481 0.0014104 0.98663 0.9915 3.0443e-006 1.2177e-005 0.13853 0.87595 0.88313 0.0014098 0.96469 0.53502 0.0018988 0.42599 1.7095 1.7081 16.0093 144.9785 0.00021679 -85.5487 0.46495
2.569 0.98805 5.5093e-005 3.8182 0.012015 3.3734e-005 0.0011553 0.20865 0.00065909 0.2093 0.1925 0 0.033553 0.0389 0 1.0281 0.30882 0.088207 0.011855 5.2111 0.073987 9.0548e-005 0.8161 0.0060841 0.0068489 0.0014102 0.98663 0.9915 3.0438e-006 1.2175e-005 0.13854 0.87629 0.88331 0.0014097 0.9649 0.53518 0.0018987 0.426 1.7104 1.709 16.0093 144.9785 0.00021652 -85.5495 0.46595
2.57 0.98805 5.5093e-005 3.8182 0.012015 3.3747e-005 0.0011553 0.20867 0.00065909 0.20932 0.19252 0 0.033552 0.0389 0 1.0282 0.30886 0.088223 0.011857 5.2121 0.073999 9.0563e-005 0.81609 0.0060848 0.0068496 0.00141 0.98664 0.99151 3.0434e-006 1.2174e-005 0.13854 0.87663 0.88348 0.0014096 0.9651 0.53534 0.0018985 0.42601 1.7112 1.7098 16.0093 144.9785 0.00021624 -85.5503 0.46695
2.571 0.98805 5.5093e-005 3.8182 0.012015 3.376e-005 0.0011553 0.20869 0.00065909 0.20935 0.19254 0 0.03355 0.0389 0 1.0283 0.30891 0.088238 0.011859 5.213 0.07401 9.0578e-005 0.81608 0.0060855 0.0068503 0.0014098 0.98664 0.99151 3.043e-006 1.2172e-005 0.13855 0.87696 0.88365 0.0014095 0.96531 0.53551 0.0018984 0.42602 1.7121 1.7107 16.0093 144.9785 0.00021597 -85.5511 0.46795
2.572 0.98805 5.5093e-005 3.8182 0.012015 3.3773e-005 0.0011553 0.20871 0.00065909 0.20937 0.19256 0 0.033549 0.0389 0 1.0284 0.30895 0.088254 0.01186 5.214 0.074021 9.0593e-005 0.81607 0.0060862 0.006851 0.0014096 0.98664 0.99151 3.0425e-006 1.217e-005 0.13856 0.87729 0.88383 0.0014094 0.96552 0.53567 0.0018983 0.42604 1.7129 1.7115 16.0092 144.9785 0.0002157 -85.5519 0.46895
2.573 0.98805 5.5093e-005 3.8182 0.012015 3.3786e-005 0.0011553 0.20873 0.00065909 0.20939 0.19258 0 0.033548 0.0389 0 1.0285 0.309 0.08827 0.011862 5.215 0.074032 9.0608e-005 0.81606 0.0060869 0.0068518 0.0014094 0.98664 0.99151 3.0421e-006 1.2168e-005 0.13856 0.87762 0.884 0.0014093 0.96572 0.53583 0.0018981 0.42605 1.7138 1.7124 16.0092 144.9786 0.00021543 -85.5527 0.46995
2.574 0.98805 5.5093e-005 3.8182 0.012015 3.3799e-005 0.0011553 0.20876 0.00065909 0.20941 0.1926 0 0.033547 0.0389 0 1.0286 0.30904 0.088286 0.011864 5.216 0.074043 9.0623e-005 0.81605 0.0060876 0.0068525 0.0014092 0.98665 0.99151 3.0417e-006 1.2167e-005 0.13857 0.87795 0.88417 0.0014092 0.96592 0.53599 0.001898 0.42606 1.7146 1.7132 16.0092 144.9786 0.00021516 -85.5535 0.47095
2.575 0.98805 5.5092e-005 3.8182 0.012015 3.3812e-005 0.0011553 0.20878 0.00065909 0.20943 0.19262 0 0.033546 0.0389 0 1.0287 0.30908 0.088302 0.011866 5.217 0.074054 9.0638e-005 0.81604 0.0060883 0.0068532 0.001409 0.98665 0.99151 3.0412e-006 1.2165e-005 0.13857 0.87828 0.88434 0.0014091 0.96612 0.53615 0.0018979 0.42608 1.7155 1.7141 16.0092 144.9786 0.00021489 -85.5543 0.47195
2.576 0.98805 5.5092e-005 3.8182 0.012015 3.3825e-005 0.0011553 0.2088 0.00065909 0.20945 0.19264 0 0.033545 0.0389 0 1.0288 0.30913 0.088317 0.011868 5.218 0.074066 9.0653e-005 0.81603 0.006089 0.006854 0.0014089 0.98665 0.99151 3.0408e-006 1.2163e-005 0.13858 0.87861 0.88451 0.001409 0.96632 0.53631 0.0018978 0.42609 1.7163 1.7149 16.0092 144.9786 0.00021462 -85.5551 0.47295
2.577 0.98805 5.5092e-005 3.8182 0.012015 3.3838e-005 0.0011553 0.20882 0.00065909 0.20947 0.19266 0 0.033544 0.0389 0 1.0289 0.30917 0.088333 0.011869 5.2189 0.074077 9.0668e-005 0.81601 0.0060897 0.0068547 0.0014087 0.98665 0.99152 3.0404e-006 1.2162e-005 0.13858 0.87894 0.88468 0.0014089 0.96652 0.53647 0.0018976 0.4261 1.7171 1.7157 16.0092 144.9786 0.00021435 -85.5559 0.47395
2.578 0.98805 5.5092e-005 3.8182 0.012015 3.3852e-005 0.0011553 0.20884 0.00065909 0.2095 0.19268 0 0.033542 0.0389 0 1.029 0.30922 0.088349 0.011871 5.2199 0.074088 9.0683e-005 0.816 0.0060904 0.0068554 0.0014085 0.98666 0.99152 3.04e-006 1.216e-005 0.13859 0.87927 0.88485 0.0014088 0.96672 0.53663 0.0018975 0.42611 1.718 1.7166 16.0092 144.9787 0.00021409 -85.5567 0.47495
2.579 0.98805 5.5092e-005 3.8182 0.012015 3.3865e-005 0.0011553 0.20886 0.00065909 0.20952 0.1927 0 0.033541 0.0389 0 1.0291 0.30926 0.088365 0.011873 5.2209 0.074099 9.0698e-005 0.81599 0.0060911 0.0068562 0.0014083 0.98666 0.99152 3.0396e-006 1.2158e-005 0.1386 0.87959 0.88502 0.0014087 0.96692 0.53679 0.0018974 0.42613 1.7188 1.7174 16.0092 144.9787 0.00021382 -85.5574 0.47595
2.58 0.98805 5.5092e-005 3.8182 0.012015 3.3878e-005 0.0011553 0.20888 0.00065909 0.20954 0.19272 0 0.03354 0.0389 0 1.0292 0.30931 0.088381 0.011875 5.2219 0.07411 9.0712e-005 0.81598 0.0060918 0.0068569 0.0014081 0.98666 0.99152 3.0392e-006 1.2157e-005 0.1386 0.87992 0.88519 0.0014086 0.96711 0.53695 0.0018973 0.42614 1.7196 1.7183 16.0092 144.9787 0.00021356 -85.5582 0.47695
2.581 0.98805 5.5092e-005 3.8182 0.012015 3.3891e-005 0.0011553 0.2089 0.00065909 0.20956 0.19274 0 0.033539 0.0389 0 1.0293 0.30935 0.088397 0.011877 5.2229 0.074121 9.0727e-005 0.81597 0.0060925 0.0068576 0.001408 0.98666 0.99152 3.0388e-006 1.2155e-005 0.13861 0.88024 0.88535 0.0014085 0.96731 0.53712 0.0018971 0.42615 1.7205 1.7191 16.0091 144.9787 0.0002133 -85.5589 0.47795
2.582 0.98805 5.5092e-005 3.8182 0.012015 3.3904e-005 0.0011553 0.20893 0.00065909 0.20958 0.19276 0 0.033538 0.0389 0 1.0294 0.3094 0.088412 0.011878 5.2239 0.074133 9.0742e-005 0.81596 0.0060932 0.0068584 0.0014078 0.98667 0.99152 3.0384e-006 1.2153e-005 0.13861 0.88056 0.88552 0.0014084 0.9675 0.53728 0.001897 0.42617 1.7213 1.7199 16.0091 144.9787 0.00021304 -85.5597 0.47895
2.583 0.98805 5.5092e-005 3.8182 0.012015 3.3917e-005 0.0011553 0.20895 0.00065909 0.2096 0.19278 0 0.033537 0.0389 0 1.0295 0.30944 0.088428 0.01188 5.2249 0.074144 9.0757e-005 0.81595 0.0060939 0.0068591 0.0014076 0.98667 0.99153 3.038e-006 1.2152e-005 0.13862 0.88088 0.88569 0.0014083 0.96769 0.53744 0.0018969 0.42618 1.7221 1.7208 16.0091 144.9788 0.00021278 -85.5604 0.47995
2.584 0.98805 5.5092e-005 3.8182 0.012015 3.393e-005 0.0011553 0.20897 0.00065909 0.20962 0.1928 0 0.033536 0.0389 0 1.0296 0.30948 0.088444 0.011882 5.2258 0.074155 9.0772e-005 0.81594 0.0060946 0.0068598 0.0014074 0.98667 0.99153 3.0376e-006 1.215e-005 0.13862 0.8812 0.88585 0.0014082 0.96788 0.5376 0.0018968 0.42619 1.7229 1.7216 16.0091 144.9788 0.00021252 -85.5612 0.48095
2.585 0.98805 5.5092e-005 3.8182 0.012015 3.3943e-005 0.0011553 0.20899 0.00065909 0.20964 0.19282 0 0.033534 0.0389 0 1.0297 0.30953 0.08846 0.011884 5.2268 0.074166 9.0787e-005 0.81592 0.0060953 0.0068606 0.0014073 0.98667 0.99153 3.0372e-006 1.2149e-005 0.13863 0.88152 0.88602 0.0014081 0.96807 0.53776 0.0018967 0.4262 1.7238 1.7224 16.0091 144.9788 0.00021226 -85.5619 0.48195
2.586 0.98805 5.5092e-005 3.8182 0.012015 3.3956e-005 0.0011553 0.20901 0.00065909 0.20966 0.19284 0 0.033533 0.0389 0 1.0298 0.30957 0.088476 0.011886 5.2278 0.074177 9.0802e-005 0.81591 0.006096 0.0068613 0.0014071 0.98667 0.99153 3.0368e-006 1.2147e-005 0.13864 0.88184 0.88618 0.001408 0.96826 0.53792 0.0018965 0.42622 1.7246 1.7232 16.0091 144.9788 0.000212 -85.5626 0.48295
2.587 0.98805 5.5092e-005 3.8182 0.012015 3.3969e-005 0.0011554 0.20903 0.00065909 0.20969 0.19286 0 0.033532 0.0389 0 1.0299 0.30962 0.088492 0.011887 5.2288 0.074189 9.0817e-005 0.8159 0.0060967 0.006862 0.0014069 0.98668 0.99153 3.0364e-006 1.2145e-005 0.13864 0.88216 0.88634 0.001408 0.96844 0.53808 0.0018964 0.42623 1.7254 1.724 16.0091 144.9788 0.00021174 -85.5634 0.48395
2.588 0.98805 5.5092e-005 3.8182 0.012015 3.3982e-005 0.0011554 0.20905 0.00065909 0.20971 0.19288 0 0.033531 0.0389 0 1.03 0.30966 0.088507 0.011889 5.2298 0.0742 9.0832e-005 0.81589 0.0060974 0.0068628 0.0014067 0.98668 0.99153 3.036e-006 1.2144e-005 0.13865 0.88247 0.88651 0.0014079 0.96863 0.53824 0.0018963 0.42624 1.7262 1.7249 16.0091 144.9788 0.00021149 -85.5641 0.48495
2.589 0.98805 5.5092e-005 3.8182 0.012015 3.3995e-005 0.0011554 0.20907 0.00065909 0.20973 0.1929 0 0.03353 0.0389 0 1.0301 0.30971 0.088523 0.011891 5.2308 0.074211 9.0847e-005 0.81588 0.0060981 0.0068635 0.0014066 0.98668 0.99153 3.0356e-006 1.2142e-005 0.13865 0.88279 0.88667 0.0014078 0.96881 0.5384 0.0018962 0.42625 1.727 1.7257 16.0091 144.9789 0.00021123 -85.5648 0.48595
2.59 0.98805 5.5091e-005 3.8182 0.012015 3.4008e-005 0.0011554 0.20909 0.00065909 0.20975 0.19292 0 0.033529 0.0389 0 1.0302 0.30975 0.088539 0.011893 5.2318 0.074222 9.0862e-005 0.81587 0.0060988 0.0068642 0.0014064 0.98668 0.99154 3.0352e-006 1.2141e-005 0.13866 0.8831 0.88683 0.0014077 0.969 0.53856 0.0018961 0.42627 1.7278 1.7265 16.009 144.9789 0.00021098 -85.5655 0.48695
2.591 0.98805 5.5091e-005 3.8182 0.012015 3.4021e-005 0.0011554 0.20912 0.00065909 0.20977 0.19294 0 0.033528 0.0389 0 1.0303 0.3098 0.088555 0.011894 5.2328 0.074233 9.0877e-005 0.81586 0.0060995 0.006865 0.0014062 0.98669 0.99154 3.0348e-006 1.2139e-005 0.13866 0.88342 0.88699 0.0014076 0.96918 0.53872 0.001896 0.42628 1.7286 1.7273 16.009 144.9789 0.00021073 -85.5662 0.48795
2.592 0.98805 5.5091e-005 3.8182 0.012015 3.4035e-005 0.0011554 0.20914 0.00065909 0.20979 0.19296 0 0.033527 0.0389 0 1.0304 0.30984 0.088571 0.011896 5.2338 0.074244 9.0892e-005 0.81585 0.0061002 0.0068657 0.0014061 0.98669 0.99154 3.0345e-006 1.2138e-005 0.13867 0.88373 0.88715 0.0014075 0.96936 0.53888 0.0018959 0.42629 1.7294 1.7281 16.009 144.9789 0.00021048 -85.5669 0.48895
2.593 0.98805 5.5091e-005 3.8182 0.012015 3.4048e-005 0.0011554 0.20916 0.00065909 0.20981 0.19298 0 0.033525 0.0389 0 1.0305 0.30988 0.088587 0.011898 5.2348 0.074256 9.0906e-005 0.81584 0.0061009 0.0068664 0.0014059 0.98669 0.99154 3.0341e-006 1.2136e-005 0.13868 0.88404 0.88731 0.0014074 0.96954 0.53904 0.0018957 0.42631 1.7302 1.7289 16.009 144.9789 0.00021023 -85.5676 0.48995
2.594 0.98805 5.5091e-005 3.8182 0.012015 3.4061e-005 0.0011554 0.20918 0.00065909 0.20983 0.193 0 0.033524 0.0389 0 1.0306 0.30993 0.088602 0.0119 5.2357 0.074267 9.0921e-005 0.81582 0.0061016 0.0068672 0.0014058 0.98669 0.99154 3.0337e-006 1.2135e-005 0.13868 0.88435 0.88747 0.0014073 0.96972 0.5392 0.0018956 0.42632 1.731 1.7297 16.009 144.979 0.00020998 -85.5683 0.49095
2.595 0.98805 5.5091e-005 3.8182 0.012015 3.4074e-005 0.0011554 0.2092 0.00065909 0.20985 0.19302 0 0.033523 0.0389 0 1.0307 0.30997 0.088618 0.011902 5.2367 0.074278 9.0936e-005 0.81581 0.0061023 0.0068679 0.0014056 0.98669 0.99154 3.0334e-006 1.2133e-005 0.13869 0.88466 0.88763 0.0014073 0.96989 0.53936 0.0018955 0.42633 1.7318 1.7305 16.009 144.979 0.00020973 -85.569 0.49195
2.596 0.98805 5.5091e-005 3.8182 0.012015 3.4087e-005 0.0011554 0.20922 0.00065909 0.20987 0.19304 0 0.033522 0.0389 0 1.0308 0.31002 0.088634 0.011903 5.2377 0.074289 9.0951e-005 0.8158 0.006103 0.0068686 0.0014054 0.9867 0.99154 3.033e-006 1.2132e-005 0.13869 0.88497 0.88778 0.0014072 0.97007 0.53952 0.0018954 0.42634 1.7326 1.7313 16.009 144.979 0.00020948 -85.5697 0.49295
2.597 0.98805 5.5091e-005 3.8182 0.012015 3.41e-005 0.0011554 0.20924 0.00065909 0.2099 0.19306 0 0.033521 0.0389 0 1.0309 0.31006 0.08865 0.011905 5.2387 0.0743 9.0966e-005 0.81579 0.0061037 0.0068694 0.0014053 0.9867 0.99154 3.0326e-006 1.213e-005 0.1387 0.88528 0.88794 0.0014071 0.97024 0.53968 0.0018953 0.42636 1.7334 1.7321 16.009 144.979 0.00020924 -85.5704 0.49395
2.598 0.98805 5.5091e-005 3.8182 0.012015 3.4113e-005 0.0011554 0.20926 0.00065909 0.20992 0.19308 0 0.03352 0.0389 0 1.031 0.31011 0.088666 0.011907 5.2397 0.074311 9.0981e-005 0.81578 0.0061044 0.0068701 0.0014051 0.9867 0.99155 3.0323e-006 1.2129e-005 0.1387 0.88558 0.8881 0.001407 0.97042 0.53984 0.0018952 0.42637 1.7342 1.7329 16.0089 144.979 0.00020899 -85.571 0.49495
2.599 0.98805 5.5091e-005 3.8182 0.012015 3.4126e-005 0.0011554 0.20928 0.0006591 0.20994 0.1931 0 0.033519 0.0389 0 1.0311 0.31015 0.088682 0.011909 5.2407 0.074323 9.0996e-005 0.81577 0.0061051 0.0068709 0.001405 0.9867 0.99155 3.0319e-006 1.2128e-005 0.13871 0.88589 0.88825 0.0014069 0.97059 0.54 0.0018951 0.42638 1.735 1.7337 16.0089 144.9791 0.00020875 -85.5717 0.49595
2.6 0.98805 5.5091e-005 3.8182 0.012014 3.4139e-005 0.0011554 0.2093 0.0006591 0.20996 0.19312 0 0.033518 0.0389 0 1.0312 0.3102 0.088697 0.011911 5.2417 0.074334 9.1011e-005 0.81576 0.0061058 0.0068716 0.0014048 0.9867 0.99155 3.0315e-006 1.2126e-005 0.13872 0.8862 0.88841 0.0014068 0.97076 0.54016 0.001895 0.4264 1.7358 1.7345 16.0089 144.9791 0.0002085 -85.5724 0.49695
2.601 0.98805 5.5091e-005 3.8182 0.012014 3.4152e-005 0.0011554 0.20932 0.0006591 0.20998 0.19314 0 0.033516 0.0389 0 1.0312 0.31024 0.088713 0.011912 5.2427 0.074345 9.1026e-005 0.81575 0.0061065 0.0068723 0.0014046 0.98671 0.99155 3.0312e-006 1.2125e-005 0.13872 0.8865 0.88856 0.0014068 0.97093 0.54032 0.0018949 0.42641 1.7366 1.7353 16.0089 144.9791 0.00020826 -85.573 0.49795
2.602 0.98805 5.5091e-005 3.8182 0.012014 3.4165e-005 0.0011554 0.20935 0.0006591 0.21 0.19316 0 0.033515 0.0389 0 1.0313 0.31029 0.088729 0.011914 5.2437 0.074356 9.1041e-005 0.81573 0.0061072 0.0068731 0.0014045 0.98671 0.99155 3.0308e-006 1.2123e-005 0.13873 0.8868 0.88872 0.0014067 0.9711 0.54048 0.0018948 0.42642 1.7374 1.7361 16.0089 144.9791 0.00020802 -85.5737 0.49895
2.603 0.98805 5.5091e-005 3.8182 0.012014 3.4178e-005 0.0011554 0.20937 0.0006591 0.21002 0.19318 0 0.033514 0.0389 0 1.0314 0.31033 0.088745 0.011916 5.2447 0.074367 9.1056e-005 0.81572 0.0061079 0.0068738 0.0014043 0.98671 0.99155 3.0305e-006 1.2122e-005 0.13873 0.8871 0.88887 0.0014066 0.97127 0.54064 0.0018947 0.42643 1.7382 1.7369 16.0089 144.9791 0.00020778 -85.5743 0.49995
2.604 0.98805 5.5091e-005 3.8182 0.012014 3.4191e-005 0.0011554 0.20939 0.0006591 0.21004 0.1932 0 0.033513 0.0389 0 1.0315 0.31037 0.088761 0.011918 5.2457 0.074379 9.1071e-005 0.81571 0.0061086 0.0068745 0.0014042 0.98671 0.99155 3.0301e-006 1.2121e-005 0.13874 0.88741 0.88902 0.0014065 0.97144 0.5408 0.0018946 0.42645 1.739 1.7377 16.0089 144.9792 0.00020754 -85.575 0.50095
2.605 0.98805 5.509e-005 3.8182 0.012014 3.4205e-005 0.0011554 0.20941 0.0006591 0.21006 0.19322 0 0.033512 0.0389 0 1.0316 0.31042 0.088777 0.011919 5.2467 0.07439 9.1086e-005 0.8157 0.0061093 0.0068753 0.001404 0.98671 0.99156 3.0298e-006 1.2119e-005 0.13874 0.88771 0.88918 0.0014064 0.9716 0.54096 0.0018945 0.42646 1.7397 1.7385 16.0089 144.9792 0.0002073 -85.5756 0.50195
2.606 0.98805 5.509e-005 3.8182 0.012014 3.4218e-005 0.0011554 0.20943 0.0006591 0.21008 0.19324 0 0.033511 0.0389 0 1.0317 0.31046 0.088792 0.011921 5.2477 0.074401 9.11e-005 0.81569 0.00611 0.006876 0.0014039 0.98672 0.99156 3.0295e-006 1.2118e-005 0.13875 0.888 0.88933 0.0014064 0.97177 0.54112 0.0018944 0.42647 1.7405 1.7392 16.0088 144.9792 0.00020706 -85.5763 0.50295
2.607 0.98805 5.509e-005 3.8182 0.012014 3.4231e-005 0.0011554 0.20945 0.0006591 0.2101 0.19326 0 0.03351 0.0389 0 1.0318 0.31051 0.088808 0.011923 5.2487 0.074412 9.1115e-005 0.81568 0.0061107 0.0068767 0.0014037 0.98672 0.99156 3.0291e-006 1.2116e-005 0.13876 0.8883 0.88948 0.0014063 0.97193 0.54128 0.0018943 0.42649 1.7413 1.74 16.0088 144.9792 0.00020682 -85.5769 0.50395
2.608 0.98805 5.509e-005 3.8182 0.012014 3.4244e-005 0.0011554 0.20947 0.0006591 0.21012 0.19328 0 0.033509 0.0389 0 1.0319 0.31055 0.088824 0.011925 5.2497 0.074423 9.113e-005 0.81567 0.0061114 0.0068775 0.0014036 0.98672 0.99156 3.0288e-006 1.2115e-005 0.13876 0.8886 0.88963 0.0014062 0.9721 0.54144 0.0018942 0.4265 1.7421 1.7408 16.0088 144.9792 0.00020659 -85.5775 0.50495
2.609 0.98805 5.509e-005 3.8182 0.012014 3.4257e-005 0.0011554 0.20949 0.0006591 0.21014 0.1933 0 0.033508 0.0389 0 1.032 0.3106 0.08884 0.011927 5.2507 0.074434 9.1145e-005 0.81566 0.0061121 0.0068782 0.0014034 0.98672 0.99156 3.0284e-006 1.2114e-005 0.13877 0.8889 0.88978 0.0014061 0.97226 0.54159 0.0018941 0.42651 1.7428 1.7416 16.0088 144.9793 0.00020635 -85.5781 0.50595
2.61 0.98805 5.509e-005 3.8182 0.012014 3.427e-005 0.0011554 0.20951 0.0006591 0.21017 0.19332 0 0.033507 0.0389 0 1.0321 0.31064 0.088856 0.011928 5.2517 0.074446 9.116e-005 0.81565 0.0061128 0.0068789 0.0014033 0.98672 0.99156 3.0281e-006 1.2112e-005 0.13877 0.88919 0.88993 0.001406 0.97242 0.54175 0.001894 0.42652 1.7436 1.7423 16.0088 144.9793 0.00020612 -85.5788 0.50695
2.611 0.98805 5.509e-005 3.8182 0.012014 3.4283e-005 0.0011554 0.20953 0.0006591 0.21019 0.19334 0 0.033505 0.0389 0 1.0322 0.31069 0.088872 0.01193 5.2527 0.074457 9.1175e-005 0.81563 0.0061135 0.0068797 0.0014032 0.98673 0.99156 3.0278e-006 1.2111e-005 0.13878 0.88949 0.89008 0.001406 0.97258 0.54191 0.0018939 0.42654 1.7444 1.7431 16.0088 144.9793 0.00020588 -85.5794 0.50795
2.612 0.98805 5.509e-005 3.8182 0.012014 3.4296e-005 0.0011554 0.20955 0.0006591 0.21021 0.19336 0 0.033504 0.0389 0 1.0323 0.31073 0.088888 0.011932 5.2537 0.074468 9.119e-005 0.81562 0.0061142 0.0068804 0.001403 0.98673 0.99156 3.0275e-006 1.211e-005 0.13878 0.88978 0.89023 0.0014059 0.97274 0.54207 0.0018938 0.42655 1.7451 1.7439 16.0088 144.9793 0.00020565 -85.58 0.50895
2.613 0.98805 5.509e-005 3.8182 0.012014 3.4309e-005 0.0011554 0.20957 0.0006591 0.21023 0.19338 0 0.033503 0.0389 0 1.0324 0.31078 0.088903 0.011934 5.2547 0.074479 9.1205e-005 0.81561 0.0061149 0.0068812 0.0014029 0.98673 0.99157 3.0271e-006 1.2108e-005 0.13879 0.89007 0.89037 0.0014058 0.9729 0.54223 0.0018937 0.42656 1.7459 1.7446 16.0087 144.9793 0.00020542 -85.5806 0.50995
2.614 0.98805 5.509e-005 3.8182 0.012014 3.4322e-005 0.0011554 0.20959 0.0006591 0.21025 0.1934 0 0.033502 0.0389 0 1.0325 0.31082 0.088919 0.011936 5.2557 0.07449 9.122e-005 0.8156 0.0061156 0.0068819 0.0014027 0.98673 0.99157 3.0268e-006 1.2107e-005 0.1388 0.89036 0.89052 0.0014057 0.97305 0.54239 0.0018936 0.42658 1.7467 1.7454 16.0087 144.9794 0.00020519 -85.5812 0.51095
2.615 0.98805 5.509e-005 3.8182 0.012014 3.4335e-005 0.0011554 0.20961 0.0006591 0.21027 0.19342 0 0.033501 0.0389 0 1.0326 0.31086 0.088935 0.011937 5.2567 0.074501 9.1235e-005 0.81559 0.0061163 0.0068826 0.0014026 0.98673 0.99157 3.0265e-006 1.2106e-005 0.1388 0.89066 0.89067 0.0014057 0.97321 0.54255 0.0018935 0.42659 1.7474 1.7462 16.0087 144.9794 0.00020496 -85.5818 0.51195
2.616 0.98805 5.509e-005 3.8182 0.012014 3.4348e-005 0.0011554 0.20963 0.0006591 0.21029 0.19343 0 0.0335 0.0389 0 1.0327 0.31091 0.088951 0.011939 5.2577 0.074513 9.125e-005 0.81558 0.006117 0.0068834 0.0014025 0.98673 0.99157 3.0262e-006 1.2105e-005 0.13881 0.89094 0.89081 0.0014056 0.97336 0.54271 0.0018934 0.4266 1.7482 1.7469 16.0087 144.9794 0.00020473 -85.5824 0.51295
2.617 0.98805 5.509e-005 3.8182 0.012014 3.4361e-005 0.0011554 0.20966 0.0006591 0.21031 0.19345 0 0.033499 0.0389 0 1.0328 0.31095 0.088967 0.011941 5.2587 0.074524 9.1265e-005 0.81557 0.0061177 0.0068841 0.0014023 0.98674 0.99157 3.0259e-006 1.2103e-005 0.13881 0.89123 0.89096 0.0014055 0.97352 0.54287 0.0018933 0.42661 1.7489 1.7477 16.0087 144.9794 0.0002045 -85.583 0.51395
2.618 0.98805 5.509e-005 3.8182 0.012014 3.4374e-005 0.0011554 0.20968 0.0006591 0.21033 0.19347 0 0.033498 0.0389 0 1.0329 0.311 0.088983 0.011943 5.2597 0.074535 9.128e-005 0.81556 0.0061184 0.0068848 0.0014022 0.98674 0.99157 3.0255e-006 1.2102e-005 0.13882 0.89152 0.8911 0.0014054 0.97367 0.54303 0.0018932 0.42663 1.7497 1.7485 16.0087 144.9794 0.00020427 -85.5836 0.51495
2.619 0.98805 5.509e-005 3.8182 0.012014 3.4388e-005 0.0011554 0.2097 0.0006591 0.21035 0.19349 0 0.033497 0.0389 0 1.033 0.31104 0.088998 0.011944 5.2607 0.074546 9.1295e-005 0.81555 0.0061191 0.0068856 0.001402 0.98674 0.99157 3.0252e-006 1.2101e-005 0.13882 0.89181 0.89125 0.0014054 0.97382 0.54318 0.0018931 0.42664 1.7504 1.7492 16.0087 144.9795 0.00020405 -85.5842 0.51595
2.62 0.98805 5.5089e-005 3.8182 0.012014 3.4401e-005 0.0011554 0.20972 0.0006591 0.21037 0.19351 0 0.033496 0.0389 0 1.0331 0.31109 0.089014 0.011946 5.2617 0.074557 9.1309e-005 0.81553 0.0061198 0.0068863 0.0014019 0.98674 0.99157 3.0249e-006 1.21e-005 0.13883 0.8921 0.89139 0.0014053 0.97397 0.54334 0.001893 0.42665 1.7512 1.75 16.0086 144.9795 0.00020382 -85.5847 0.51695
2.621 0.98805 5.5089e-005 3.8182 0.012014 3.4414e-005 0.0011554 0.20974 0.0006591 0.21039 0.19353 0 0.033494 0.0389 0 1.0332 0.31113 0.08903 0.011948 5.2627 0.074568 9.1324e-005 0.81552 0.0061205 0.006887 0.0014018 0.98674 0.99157 3.0246e-006 1.2098e-005 0.13884 0.89238 0.89154 0.0014052 0.97412 0.5435 0.0018929 0.42667 1.7519 1.7507 16.0086 144.9795 0.0002036 -85.5853 0.51795
2.622 0.98805 5.5089e-005 3.8182 0.012014 3.4427e-005 0.0011554 0.20976 0.0006591 0.21041 0.19355 0 0.033493 0.0389 0 1.0333 0.31118 0.089046 0.01195 5.2637 0.07458 9.1339e-005 0.81551 0.0061212 0.0068878 0.0014016 0.98675 0.99158 3.0243e-006 1.2097e-005 0.13884 0.89267 0.89168 0.0014052 0.97427 0.54366 0.0018928 0.42668 1.7527 1.7515 16.0086 144.9795 0.00020337 -85.5859 0.51895
2.623 0.98805 5.5089e-005 3.8182 0.012014 3.444e-005 0.0011554 0.20978 0.0006591 0.21043 0.19357 0 0.033492 0.0389 0 1.0334 0.31122 0.089062 0.011952 5.2647 0.074591 9.1354e-005 0.8155 0.0061219 0.0068885 0.0014015 0.98675 0.99158 3.024e-006 1.2096e-005 0.13885 0.89295 0.89182 0.0014051 0.97442 0.54382 0.0018927 0.42669 1.7534 1.7522 16.0086 144.9795 0.00020315 -85.5865 0.51995
2.624 0.98805 5.5089e-005 3.8182 0.012014 3.4453e-005 0.0011554 0.2098 0.0006591 0.21045 0.19359 0 0.033491 0.0389 0 1.0335 0.31127 0.089078 0.011953 5.2657 0.074602 9.1369e-005 0.81549 0.0061226 0.0068893 0.0014014 0.98675 0.99158 3.0237e-006 1.2095e-005 0.13885 0.89323 0.89196 0.001405 0.97457 0.54398 0.0018926 0.4267 1.7542 1.753 16.0086 144.9796 0.00020293 -85.587 0.52095
2.625 0.98805 5.5089e-005 3.8182 0.012014 3.4466e-005 0.0011554 0.20982 0.0006591 0.21047 0.19361 0 0.03349 0.0389 0 1.0336 0.31131 0.089094 0.011955 5.2667 0.074613 9.1384e-005 0.81548 0.0061233 0.00689 0.0014012 0.98675 0.99158 3.0234e-006 1.2094e-005 0.13886 0.89351 0.8921 0.001405 0.97471 0.54414 0.0018925 0.42672 1.7549 1.7537 16.0086 144.9796 0.00020271 -85.5876 0.52195
2.626 0.98805 5.5089e-005 3.8182 0.012014 3.4479e-005 0.0011554 0.20984 0.0006591 0.21049 0.19363 0 0.033489 0.0389 0 1.0337 0.31135 0.089109 0.011957 5.2677 0.074624 9.1399e-005 0.81547 0.006124 0.0068907 0.0014011 0.98675 0.99158 3.0231e-006 1.2092e-005 0.13886 0.8938 0.89224 0.0014049 0.97486 0.54429 0.0018924 0.42673 1.7556 1.7544 16.0086 144.9796 0.00020249 -85.5881 0.52295
2.627 0.98805 5.5089e-005 3.8182 0.012014 3.4492e-005 0.0011554 0.20986 0.0006591 0.21051 0.19365 0 0.033488 0.0389 0 1.0338 0.3114 0.089125 0.011959 5.2687 0.074635 9.1414e-005 0.81546 0.0061247 0.0068915 0.001401 0.98675 0.99158 3.0228e-006 1.2091e-005 0.13887 0.89408 0.89238 0.0014048 0.975 0.54445 0.0018924 0.42674 1.7564 1.7552 16.0085 144.9796 0.00020227 -85.5887 0.52395
2.628 0.98805 5.5089e-005 3.8182 0.012014 3.4505e-005 0.0011554 0.20988 0.0006591 0.21054 0.19367 0 0.033487 0.0389 0 1.0339 0.31144 0.089141 0.011961 5.2697 0.074647 9.1429e-005 0.81544 0.0061254 0.0068922 0.0014009 0.98676 0.99158 3.0225e-006 1.209e-005 0.13888 0.89435 0.89252 0.0014048 0.97515 0.54461 0.0018923 0.42676 1.7571 1.7559 16.0085 144.9796 0.00020205 -85.5892 0.52495
2.629 0.98805 5.5089e-005 3.8182 0.012014 3.4518e-005 0.0011554 0.2099 0.0006591 0.21056 0.19369 0 0.033486 0.0389 0 1.034 0.31149 0.089157 0.011962 5.2707 0.074658 9.1444e-005 0.81543 0.0061261 0.006893 0.0014007 0.98676 0.99158 3.0222e-006 1.2089e-005 0.13888 0.89463 0.89266 0.0014047 0.97529 0.54477 0.0018922 0.42677 1.7579 1.7567 16.0085 144.9797 0.00020183 -85.5898 0.52595
2.63 0.98805 5.5089e-005 3.8182 0.012014 3.4531e-005 0.0011554 0.20992 0.0006591 0.21058 0.19371 0 0.033485 0.0389 0 1.0341 0.31153 0.089173 0.011964 5.2717 0.074669 9.1459e-005 0.81542 0.0061268 0.0068937 0.0014006 0.98676 0.99158 3.0219e-006 1.2088e-005 0.13889 0.89491 0.8928 0.0014046 0.97543 0.54493 0.0018921 0.42678 1.7586 1.7574 16.0085 144.9797 0.00020161 -85.5903 0.52695
2.631 0.98805 5.5089e-005 3.8182 0.012014 3.4544e-005 0.0011554 0.20994 0.0006591 0.2106 0.19373 0 0.033484 0.0389 0 1.0342 0.31158 0.089189 0.011966 5.2727 0.07468 9.1474e-005 0.81541 0.0061275 0.0068944 0.0014005 0.98676 0.99159 3.0216e-006 1.2086e-005 0.13889 0.89519 0.89294 0.0014046 0.97557 0.54509 0.001892 0.42679 1.7593 1.7581 16.0085 144.9797 0.0002014 -85.5909 0.52795
2.632 0.98805 5.5089e-005 3.8182 0.012014 3.4557e-005 0.0011554 0.20996 0.0006591 0.21062 0.19374 0 0.033482 0.0389 0 1.0343 0.31162 0.089205 0.011968 5.2737 0.074691 9.1489e-005 0.8154 0.0061282 0.0068952 0.0014004 0.98676 0.99159 3.0214e-006 1.2085e-005 0.1389 0.89546 0.89308 0.0014045 0.97571 0.54524 0.0018919 0.42681 1.76 1.7589 16.0085 144.9797 0.00020118 -85.5914 0.52895
2.633 0.98805 5.5089e-005 3.8182 0.012014 3.4571e-005 0.0011554 0.20998 0.0006591 0.21064 0.19376 0 0.033481 0.0389 0 1.0344 0.31167 0.089221 0.011969 5.2748 0.074702 9.1504e-005 0.81539 0.0061289 0.0068959 0.0014002 0.98676 0.99159 3.0211e-006 1.2084e-005 0.1389 0.89574 0.89321 0.0014045 0.97585 0.5454 0.0018918 0.42682 1.7608 1.7596 16.0084 144.9797 0.00020097 -85.5919 0.52995
2.634 0.98805 5.5089e-005 3.8182 0.012014 3.4584e-005 0.0011554 0.21 0.0006591 0.21066 0.19378 0 0.03348 0.0389 0 1.0345 0.31171 0.089236 0.011971 5.2758 0.074714 9.1518e-005 0.81538 0.0061296 0.0068966 0.0014001 0.98677 0.99159 3.0208e-006 1.2083e-005 0.13891 0.89601 0.89335 0.0014044 0.97599 0.54556 0.0018918 0.42683 1.7615 1.7603 16.0084 144.9798 0.00020075 -85.5925 0.53095
2.635 0.98805 5.5088e-005 3.8182 0.012014 3.4597e-005 0.0011554 0.21002 0.0006591 0.21068 0.1938 0 0.033479 0.0389 0 1.0346 0.31176 0.089252 0.011973 5.2768 0.074725 9.1533e-005 0.81537 0.0061303 0.0068974 0.0014 0.98677 0.99159 3.0205e-006 1.2082e-005 0.13892 0.89629 0.89349 0.0014043 0.97613 0.54572 0.0018917 0.42685 1.7622 1.761 16.0084 144.9798 0.00020054 -85.593 0.53195
2.636 0.98805 5.5088e-005 3.8182 0.012014 3.461e-005 0.0011554 0.21004 0.0006591 0.2107 0.19382 0 0.033478 0.0389 0 1.0347 0.3118 0.089268 0.011975 5.2778 0.074736 9.1548e-005 0.81536 0.006131 0.0068981 0.0013999 0.98677 0.99159 3.0202e-006 1.2081e-005 0.13892 0.89656 0.89362 0.0014042 0.97626 0.54588 0.0018916 0.42686 1.7629 1.7618 16.0084 144.9798 0.00020033 -85.5935 0.53295
2.637 0.98805 5.5088e-005 3.8182 0.012014 3.4623e-005 0.0011554 0.21006 0.0006591 0.21072 0.19384 0 0.033477 0.0389 0 1.0348 0.31185 0.089284 0.011977 5.2788 0.074747 9.1563e-005 0.81534 0.0061317 0.0068989 0.0013997 0.98677 0.99159 3.0199e-006 1.208e-005 0.13893 0.89683 0.89376 0.0014042 0.9764 0.54603 0.0018915 0.42687 1.7637 1.7625 16.0084 144.9798 0.00020012 -85.594 0.53395
2.638 0.98805 5.5088e-005 3.8182 0.012014 3.4636e-005 0.0011554 0.21008 0.0006591 0.21074 0.19386 0 0.033476 0.0389 0 1.0349 0.31189 0.0893 0.011978 5.2798 0.074758 9.1578e-005 0.81533 0.0061324 0.0068996 0.0013996 0.98677 0.99159 3.0197e-006 1.2079e-005 0.13893 0.8971 0.89389 0.0014041 0.97653 0.54619 0.0018914 0.42688 1.7644 1.7632 16.0084 144.9798 0.00019991 -85.5945 0.53495
2.639 0.98805 5.5088e-005 3.8182 0.012014 3.4649e-005 0.0011554 0.2101 0.0006591 0.21076 0.19388 0 0.033475 0.0389 0 1.035 0.31193 0.089316 0.01198 5.2808 0.074769 9.1593e-005 0.81532 0.0061331 0.0069003 0.0013995 0.98677 0.99159 3.0194e-006 1.2078e-005 0.13894 0.89737 0.89402 0.001404 0.97667 0.54635 0.0018913 0.4269 1.7651 1.7639 16.0083 144.9799 0.0001997 -85.595 0.53595
2.64 0.98805 5.5088e-005 3.8182 0.012014 3.4662e-005 0.0011554 0.21012 0.0006591 0.21078 0.1939 0 0.033474 0.0389 0 1.0351 0.31198 0.089332 0.011982 5.2818 0.074781 9.1608e-005 0.81531 0.0061338 0.0069011 0.0013994 0.98677 0.99159 3.0191e-006 1.2076e-005 0.13894 0.89764 0.89416 0.001404 0.9768 0.54651 0.0018913 0.42691 1.7658 1.7647 16.0083 144.9799 0.00019949 -85.5955 0.53695
2.641 0.98805 5.5088e-005 3.8182 0.012014 3.4675e-005 0.0011554 0.21014 0.0006591 0.2108 0.19392 0 0.033473 0.0389 0 1.0352 0.31202 0.089347 0.011984 5.2828 0.074792 9.1623e-005 0.8153 0.0061345 0.0069018 0.0013993 0.98678 0.9916 3.0189e-006 1.2075e-005 0.13895 0.89791 0.89429 0.0014039 0.97693 0.54666 0.0018912 0.42692 1.7665 1.7654 16.0083 144.9799 0.00019928 -85.596 0.53795
2.642 0.98805 5.5088e-005 3.8182 0.012014 3.4688e-005 0.0011554 0.21016 0.0006591 0.21082 0.19394 0 0.033472 0.0389 0 1.0353 0.31207 0.089363 0.011986 5.2838 0.074803 9.1638e-005 0.81529 0.0061352 0.0069026 0.0013992 0.98678 0.9916 3.0186e-006 1.2074e-005 0.13896 0.89817 0.89442 0.0014039 0.97706 0.54682 0.0018911 0.42694 1.7672 1.7661 16.0083 144.9799 0.00019907 -85.5965 0.53895
2.643 0.98805 5.5088e-005 3.8182 0.012014 3.4701e-005 0.0011554 0.21018 0.0006591 0.21084 0.19396 0 0.033471 0.0389 0 1.0353 0.31211 0.089379 0.011987 5.2849 0.074814 9.1653e-005 0.81528 0.0061359 0.0069033 0.001399 0.98678 0.9916 3.0183e-006 1.2073e-005 0.13896 0.89844 0.89455 0.0014039 0.97719 0.54698 0.001891 0.42695 1.7679 1.7668 16.0083 144.9799 0.00019887 -85.597 0.53995
2.644 0.98805 5.5088e-005 3.8182 0.012014 3.4714e-005 0.0011554 0.2102 0.0006591 0.21086 0.19397 0 0.033469 0.0389 0 1.0354 0.31216 0.089395 0.011989 5.2859 0.074825 9.1668e-005 0.81527 0.0061366 0.006904 0.0013989 0.98678 0.9916 3.0181e-006 1.2072e-005 0.13897 0.89871 0.89469 0.0014038 0.97732 0.54714 0.0018909 0.42696 1.7686 1.7675 16.0083 144.98 0.00019866 -85.5975 0.54095
2.645 0.98805 5.5088e-005 3.8182 0.012014 3.4727e-005 0.0011554 0.21022 0.0006591 0.21088 0.19399 0 0.033468 0.0389 0 1.0355 0.3122 0.089411 0.011991 5.2869 0.074836 9.1683e-005 0.81526 0.0061373 0.0069048 0.0013988 0.98678 0.9916 3.0178e-006 1.2071e-005 0.13897 0.89897 0.89482 0.0014037 0.97745 0.54729 0.0018909 0.42697 1.7693 1.7682 16.0082 144.98 0.00019845 -85.598 0.54195
2.646 0.98805 5.5088e-005 3.8182 0.012014 3.474e-005 0.0011554 0.21024 0.0006591 0.2109 0.19401 0 0.033467 0.0389 0 1.0356 0.31225 0.089427 0.011993 5.2879 0.074848 9.1698e-005 0.81524 0.006138 0.0069055 0.0013987 0.98678 0.9916 3.0175e-006 1.207e-005 0.13898 0.89924 0.89495 0.0014036 0.97758 0.54745 0.0018908 0.42699 1.77 1.7689 16.0082 144.98 0.00019825 -85.5985 0.54295
2.647 0.98805 5.5088e-005 3.8182 0.012014 3.4754e-005 0.0011554 0.21026 0.0006591 0.21092 0.19403 0 0.033466 0.0389 0 1.0357 0.31229 0.089443 0.011994 5.2889 0.074859 9.1713e-005 0.81523 0.0061387 0.0069063 0.0013986 0.98678 0.9916 3.0173e-006 1.2069e-005 0.13898 0.8995 0.89508 0.0014035 0.9777 0.54761 0.0018907 0.427 1.7707 1.7696 16.0082 144.98 0.00019805 -85.599 0.54395
2.648 0.98805 5.5088e-005 3.8182 0.012014 3.4767e-005 0.0011554 0.21029 0.0006591 0.21094 0.19405 0 0.033465 0.0389 0 1.0358 0.31234 0.089459 0.011996 5.2899 0.07487 9.1728e-005 0.81522 0.0061394 0.006907 0.0013984 0.98679 0.9916 3.017e-006 1.2068e-005 0.13899 0.89976 0.89521 0.0014034 0.97783 0.54777 0.0018906 0.42701 1.7714 1.7703 16.0082 144.98 0.00019784 -85.5995 0.54495
2.649 0.98805 5.5088e-005 3.8182 0.012014 3.478e-005 0.0011554 0.21031 0.00065911 0.21096 0.19407 0 0.033464 0.0389 0 1.0359 0.31238 0.089474 0.011998 5.2909 0.074881 9.1742e-005 0.81521 0.0061401 0.0069077 0.0013983 0.98679 0.9916 3.0168e-006 1.2067e-005 0.139 0.90002 0.89534 0.0014034 0.97796 0.54792 0.0018905 0.42703 1.7721 1.771 16.0082 144.9801 0.00019764 -85.6 0.54595
2.65 0.98805 5.5087e-005 3.8182 0.012014 3.4793e-005 0.0011554 0.21033 0.00065911 0.21098 0.19409 0 0.033463 0.0389 0 1.036 0.31243 0.08949 0.012 5.292 0.074892 9.1757e-005 0.8152 0.0061408 0.0069085 0.0013982 0.98679 0.9916 3.0165e-006 1.2066e-005 0.139 0.90028 0.89546 0.0014034 0.97808 0.54808 0.0018905 0.42704 1.7728 1.7717 16.0082 144.9801 0.00019744 -85.6004 0.54695
2.651 0.98805 5.5087e-005 3.8182 0.012014 3.4806e-005 0.0011554 0.21035 0.00065911 0.211 0.19411 0 0.033462 0.0389 0 1.0361 0.31247 0.089506 0.012002 5.293 0.074903 9.1772e-005 0.81519 0.0061415 0.0069092 0.0013981 0.98679 0.9916 3.0163e-006 1.2065e-005 0.13901 0.90054 0.89559 0.0014034 0.9782 0.54824 0.0018904 0.42705 1.7735 1.7724 16.0081 144.9801 0.00019724 -85.6009 0.54795
2.652 0.98805 5.5087e-005 3.8182 0.012014 3.4819e-005 0.0011554 0.21037 0.00065911 0.21102 0.19413 0 0.033461 0.0389 0 1.0362 0.31251 0.089522 0.012003 5.294 0.074915 9.1787e-005 0.81518 0.0061422 0.00691 0.001398 0.98679 0.99161 3.0161e-006 1.2064e-005 0.13901 0.9008 0.89572 0.0014035 0.97833 0.54839 0.0018903 0.42706 1.7742 1.7731 16.0081 144.9801 0.00019704 -85.6014 0.54895
2.653 0.98805 5.5087e-005 3.8182 0.012014 3.4832e-005 0.0011554 0.21039 0.00065911 0.21104 0.19414 0 0.03346 0.0389 0 1.0363 0.31256 0.089538 0.012005 5.295 0.074926 9.1802e-005 0.81517 0.0061429 0.0069107 0.0013979 0.98679 0.99161 3.0158e-006 1.2063e-005 0.13902 0.90106 0.89585 0.0014035 0.97845 0.54855 0.0018902 0.42708 1.7749 1.7738 16.0081 144.9801 0.00019684 -85.6018 0.54995
2.654 0.98805 5.5087e-005 3.8182 0.012014 3.4845e-005 0.0011554 0.21041 0.00065911 0.21106 0.19416 0 0.033459 0.0389 0 1.0364 0.3126 0.089554 0.012007 5.296 0.074937 9.1817e-005 0.81515 0.0061436 0.0069114 0.0013978 0.98679 0.99161 3.0156e-006 1.2062e-005 0.13902 0.90132 0.89597 0.0014034 0.97857 0.54871 0.0018902 0.42709 1.7756 1.7745 16.0081 144.9802 0.00019664 -85.6023 0.55095
2.655 0.98805 5.5087e-005 3.8182 0.012014 3.4858e-005 0.0011554 0.21043 0.00065911 0.21108 0.19418 0 0.033458 0.0389 0 1.0365 0.31265 0.08957 0.012009 5.297 0.074948 9.1832e-005 0.81514 0.0061443 0.0069122 0.0013977 0.9868 0.99161 3.0153e-006 1.2061e-005 0.13903 0.90158 0.8961 0.0014033 0.97869 0.54886 0.0018901 0.4271 1.7763 1.7752 16.0081 144.9802 0.00019645 -85.6027 0.55195
2.656 0.98805 5.5087e-005 3.8182 0.012014 3.4871e-005 0.0011554 0.21044 0.00065911 0.2111 0.1942 0 0.033457 0.0389 0 1.0366 0.31269 0.089586 0.012011 5.2981 0.074959 9.1847e-005 0.81513 0.006145 0.0069129 0.0013976 0.9868 0.99161 3.0151e-006 1.206e-005 0.13904 0.90183 0.89622 0.0014032 0.97881 0.54902 0.00189 0.42712 1.777 1.7759 16.0081 144.9802 0.00019625 -85.6032 0.55295
2.657 0.98805 5.5087e-005 3.8182 0.012014 3.4884e-005 0.0011554 0.21046 0.00065911 0.21112 0.19422 0 0.033456 0.0389 0 1.0367 0.31274 0.089602 0.012012 5.2991 0.07497 9.1862e-005 0.81512 0.0061457 0.0069137 0.0013975 0.9868 0.99161 3.0148e-006 1.2059e-005 0.13904 0.90209 0.89635 0.001403 0.97893 0.54918 0.00189 0.42713 1.7777 1.7766 16.008 144.9802 0.00019605 -85.6036 0.55395
2.658 0.98805 5.5087e-005 3.8182 0.012014 3.4897e-005 0.0011554 0.21048 0.00065911 0.21114 0.19424 0 0.033455 0.0389 0 1.0368 0.31278 0.089617 0.012014 5.3001 0.074982 9.1877e-005 0.81511 0.0061464 0.0069144 0.0013974 0.9868 0.99161 3.0146e-006 1.2058e-005 0.13905 0.90234 0.89647 0.0014028 0.97905 0.54933 0.0018899 0.42714 1.7784 1.7773 16.008 144.9802 0.00019586 -85.6041 0.55495
2.659 0.98805 5.5087e-005 3.8182 0.012014 3.491e-005 0.0011554 0.2105 0.00065911 0.21116 0.19426 0 0.033453 0.0389 0 1.0369 0.31283 0.089633 0.012016 5.3011 0.074993 9.1892e-005 0.8151 0.0061471 0.0069151 0.0013973 0.9868 0.99161 3.0143e-006 1.2057e-005 0.13905 0.90259 0.8966 0.0014028 0.97916 0.54949 0.0018898 0.42715 1.779 1.7779 16.008 144.9803 0.00019566 -85.6045 0.55595
2.66 0.98805 5.5087e-005 3.8182 0.012014 3.4923e-005 0.0011554 0.21052 0.00065911 0.21118 0.19428 0 0.033452 0.0389 0 1.037 0.31287 0.089649 0.012018 5.3021 0.075004 9.1907e-005 0.81509 0.0061478 0.0069159 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.13906 0.90285 0.89672 0.0014028 0.97928 0.54965 0.0018897 0.42717 1.7797 1.7786 16.008 144.9803 0.00019547 -85.605 0.55695
2.661 0.98805 5.5087e-005 3.8182 0.012014 3.4937e-005 0.0011554 0.21054 0.00065911 0.2112 0.1943 0 0.033451 0.0389 0 1.0371 0.31292 0.089665 0.012019 5.3031 0.075015 9.1922e-005 0.81508 0.0061485 0.0069166 0.0013971 0.9868 0.99161 3.0139e-006 1.2055e-005 0.13907 0.9031 0.89684 0.0014028 0.9794 0.5498 0.0018897 0.42718 1.7804 1.7793 16.008 144.9803 0.00019528 -85.6054 0.55795
2.662 0.98805 5.5087e-005 3.8182 0.012014 3.495e-005 0.0011554 0.21056 0.00065911 0.21122 0.19431 0 0.03345 0.0389 0 1.0372 0.31296 0.089681 0.012021 5.3042 0.075026 9.1937e-005 0.81507 0.0061492 0.0069174 0.001397 0.98681 0.99161 3.0136e-006 1.2054e-005 0.13907 0.90335 0.89697 0.0014028 0.97951 0.54996 0.0018896 0.42719 1.7811 1.78 16.008 144.9803 0.00019508 -85.6059 0.55895
2.663 0.98805 5.5087e-005 3.8182 0.012014 3.4963e-005 0.0011555 0.21058 0.00065911 0.21124 0.19433 0 0.033449 0.0389 0 1.0373 0.31301 0.089697 0.012023 5.3052 0.075037 9.1952e-005 0.81505 0.0061499 0.0069181 0.0013969 0.98681 0.99162 3.0134e-006 1.2054e-005 0.13908 0.9036 0.89709 0.0014028 0.97963 0.55012 0.0018895 0.42721 1.7817 1.7807 16.0079 144.9803 0.00019489 -85.6063 0.55995
2.664 0.98805 5.5087e-005 3.8182 0.012014 3.4976e-005 0.0011555 0.2106 0.00065911 0.21126 0.19435 0 0.033448 0.0389 0 1.0374 0.31305 0.089713 0.012025 5.3062 0.075049 9.1966e-005 0.81504 0.0061506 0.0069188 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.13908 0.90385 0.89721 0.0014027 0.97974 0.55027 0.0018895 0.42722 1.7824 1.7813 16.0079 144.9804 0.0001947 -85.6067 0.56095
2.665 0.98805 5.5086e-005 3.8182 0.012014 3.4989e-005 0.0011555 0.21062 0.00065911 0.21128 0.19437 0 0.033447 0.0389 0 1.0375 0.3131 0.089729 0.012027 5.3072 0.07506 9.1981e-005 0.81503 0.0061513 0.0069196 0.0013967 0.98681 0.99162 3.0129e-006 1.2052e-005 0.13909 0.9041 0.89733 0.0014027 0.97985 0.55043 0.0018894 0.42723 1.7831 1.782 16.0079 144.9804 0.00019451 -85.6071 0.56195
2.666 0.98805 5.5086e-005 3.8182 0.012014 3.5002e-005 0.0011555 0.21064 0.00065911 0.2113 0.19439 0 0.033446 0.0389 0 1.0376 0.31314 0.089744 0.012028 5.3083 0.075071 9.1996e-005 0.81502 0.0061521 0.0069203 0.0013966 0.98681 0.99162 3.0127e-006 1.2051e-005 0.13909 0.90435 0.89745 0.0014027 0.97997 0.55059 0.0018893 0.42724 1.7838 1.7827 16.0079 144.9804 0.00019432 -85.6076 0.56295
2.667 0.98805 5.5086e-005 3.8182 0.012014 3.5015e-005 0.0011555 0.21066 0.00065911 0.21132 0.19441 0 0.033445 0.0389 0 1.0377 0.31318 0.08976 0.01203 5.3093 0.075082 9.2011e-005 0.81501 0.0061528 0.0069211 0.0013965 0.98681 0.99162 3.0125e-006 1.205e-005 0.1391 0.9046 0.89757 0.0014026 0.98008 0.55074 0.0018893 0.42726 1.7844 1.7834 16.0079 144.9804 0.00019413 -85.608 0.56395
2.668 0.98805 5.5086e-005 3.8182 0.012014 3.5028e-005 0.0011555 0.21068 0.00065911 0.21134 0.19443 0 0.033444 0.0389 0 1.0378 0.31323 0.089776 0.012032 5.3103 0.075093 9.2026e-005 0.815 0.0061535 0.0069218 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.13911 0.90484 0.89769 0.0014026 0.98019 0.5509 0.0018892 0.42727 1.7851 1.784 16.0078 144.9804 0.00019394 -85.6084 0.56495
2.669 0.98805 5.5086e-005 3.8182 0.012014 3.5041e-005 0.0011555 0.2107 0.00065911 0.21136 0.19445 0 0.033443 0.0389 0 1.0379 0.31327 0.089792 0.012034 5.3113 0.075104 9.2041e-005 0.81499 0.0061542 0.0069226 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.13911 0.90509 0.89781 0.0014025 0.9803 0.55106 0.0018891 0.42728 1.7858 1.7847 16.0078 144.9805 0.00019376 -85.6088 0.56595
2.67 0.98805 5.5086e-005 3.8182 0.012013 3.5054e-005 0.0011555 0.21072 0.00065911 0.21138 0.19446 0 0.033442 0.0389 0 1.038 0.31332 0.089808 0.012036 5.3123 0.075116 9.2056e-005 0.81498 0.0061549 0.0069233 0.0013962 0.98682 0.99162 3.0118e-006 1.2047e-005 0.13912 0.90533 0.89793 0.0014024 0.98041 0.55121 0.0018891 0.4273 1.7864 1.7854 16.0078 144.9805 0.00019357 -85.6092 0.56695
2.671 0.98805 5.5086e-005 3.8182 0.012013 3.5067e-005 0.0011555 0.21074 0.00065911 0.2114 0.19448 0 0.033441 0.0389 0 1.0381 0.31336 0.089824 0.012037 5.3134 0.075127 9.2071e-005 0.81497 0.0061556 0.006924 0.0013961 0.98682 0.99162 3.0116e-006 1.2046e-005 0.13912 0.90558 0.89805 0.0014023 0.98052 0.55137 0.001889 0.42731 1.7871 1.786 16.0078 144.9805 0.00019338 -85.6097 0.56795
2.672 0.98805 5.5086e-005 3.8182 0.012013 3.508e-005 0.0011555 0.21076 0.00065911 0.21142 0.1945 0 0.03344 0.0389 0 1.0382 0.31341 0.08984 0.012039 5.3144 0.075138 9.2086e-005 0.81495 0.0061563 0.0069248 0.001396 0.98682 0.99162 3.0114e-006 1.2045e-005 0.13913 0.90582 0.89817 0.0014023 0.98062 0.55152 0.0018889 0.42732 1.7877 1.7867 16.0078 144.9805 0.0001932 -85.6101 0.56895
2.673 0.98805 5.5086e-005 3.8182 0.012013 3.5093e-005 0.0011555 0.21078 0.00065911 0.21144 0.19452 0 0.033439 0.0389 0 1.0383 0.31345 0.089856 0.012041 5.3154 0.075149 9.2101e-005 0.81494 0.006157 0.0069255 0.0013959 0.98682 0.99162 3.0112e-006 1.2045e-005 0.13913 0.90606 0.89829 0.0014022 0.98073 0.55168 0.0018889 0.42733 1.7884 1.7873 16.0078 144.9805 0.00019301 -85.6105 0.56995
2.674 0.98805 5.5086e-005 3.8182 0.012013 3.5106e-005 0.0011555 0.2108 0.00065911 0.21146 0.19454 0 0.033438 0.0389 0 1.0384 0.3135 0.089872 0.012043 5.3164 0.07516 9.2116e-005 0.81493 0.0061577 0.0069263 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.13914 0.9063 0.89841 0.0014021 0.98084 0.55184 0.0018888 0.42735 1.7891 1.788 16.0077 144.9806 0.00019283 -85.6109 0.57095
2.675 0.98805 5.5086e-005 3.8182 0.012013 3.512e-005 0.0011555 0.21082 0.00065911 0.21148 0.19456 0 0.033437 0.0389 0 1.0385 0.31354 0.089888 0.012044 5.3175 0.075171 9.2131e-005 0.81492 0.0061584 0.006927 0.0013957 0.98682 0.99163 3.0107e-006 1.2043e-005 0.13915 0.90655 0.89852 0.001402 0.98094 0.55199 0.0018887 0.42736 1.7897 1.7887 16.0077 144.9806 0.00019265 -85.6113 0.57195
2.676 0.98805 5.5086e-005 3.8182 0.012013 3.5133e-005 0.0011555 0.21084 0.00065911 0.21149 0.19458 0 0.033436 0.0389 0 1.0386 0.31359 0.089903 0.012046 5.3185 0.075183 9.2146e-005 0.81491 0.0061591 0.0069277 0.0013956 0.98682 0.99163 3.0105e-006 1.2042e-005 0.13915 0.90679 0.89864 0.001402 0.98105 0.55215 0.0018887 0.42737 1.7904 1.7893 16.0077 144.9806 0.00019246 -85.6117 0.57295
2.677 0.98805 5.5086e-005 3.8182 0.012013 3.5146e-005 0.0011555 0.21086 0.00065911 0.21151 0.19459 0 0.033435 0.0389 0 1.0387 0.31363 0.089919 0.012048 5.3195 0.075194 9.2161e-005 0.8149 0.0061598 0.0069285 0.0013955 0.98682 0.99163 3.0103e-006 1.2041e-005 0.13916 0.90703 0.89876 0.0014019 0.98115 0.5523 0.0018886 0.42739 1.791 1.79 16.0077 144.9806 0.00019228 -85.6121 0.57395
2.678 0.98805 5.5086e-005 3.8182 0.012013 3.5159e-005 0.0011555 0.21088 0.00065911 0.21153 0.19461 0 0.033434 0.0389 0 1.0388 0.31368 0.089935 0.01205 5.3206 0.075205 9.2176e-005 0.81489 0.0061605 0.0069292 0.0013954 0.98683 0.99163 3.0101e-006 1.204e-005 0.13916 0.90726 0.89887 0.0014019 0.98126 0.55246 0.0018885 0.4274 1.7917 1.7906 16.0077 144.9806 0.0001921 -85.6124 0.57495
2.679 0.98805 5.5086e-005 3.8182 0.012013 3.5172e-005 0.0011555 0.2109 0.00065911 0.21155 0.19463 0 0.033432 0.0389 0 1.0389 0.31372 0.089951 0.012052 5.3216 0.075216 9.2191e-005 0.81488 0.0061612 0.00693 0.0013953 0.98683 0.99163 3.0099e-006 1.204e-005 0.13917 0.9075 0.89899 0.0014018 0.98136 0.55261 0.0018885 0.42741 1.7923 1.7913 16.0076 144.9807 0.00019192 -85.6128 0.57595
2.68 0.98805 5.5085e-005 3.8182 0.012013 3.5185e-005 0.0011555 0.21092 0.00065911 0.21157 0.19465 0 0.033431 0.0389 0 1.039 0.31377 0.089967 0.012053 5.3226 0.075227 9.2205e-005 0.81487 0.0061619 0.0069307 0.0013953 0.98683 0.99163 3.0097e-006 1.2039e-005 0.13917 0.90774 0.8991 0.0014018 0.98146 0.55277 0.0018884 0.42742 1.793 1.7919 16.0076 144.9807 0.00019174 -85.6132 0.57695
2.681 0.98805 5.5085e-005 3.8182 0.012013 3.5198e-005 0.0011555 0.21094 0.00065911 0.21159 0.19467 0 0.03343 0.0389 0 1.0391 0.31381 0.089983 0.012055 5.3236 0.075238 9.222e-005 0.81485 0.0061626 0.0069315 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.13918 0.90798 0.89922 0.0014017 0.98157 0.55292 0.0018884 0.42744 1.7936 1.7926 16.0076 144.9807 0.00019156 -85.6136 0.57795
2.682 0.98805 5.5085e-005 3.8182 0.012013 3.5211e-005 0.0011555 0.21096 0.00065911 0.21161 0.19469 0 0.033429 0.0389 0 1.0392 0.31386 0.089999 0.012057 5.3247 0.07525 9.2235e-005 0.81484 0.0061633 0.0069322 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.13919 0.90821 0.89933 0.0014017 0.98167 0.55308 0.0018883 0.42745 1.7942 1.7932 16.0076 144.9807 0.00019138 -85.614 0.57895
2.683 0.98805 5.5085e-005 3.8182 0.012013 3.5224e-005 0.0011555 0.21098 0.00065911 0.21163 0.19471 0 0.033428 0.0389 0 1.0393 0.3139 0.090015 0.012059 5.3257 0.075261 9.225e-005 0.81483 0.006164 0.0069329 0.001395 0.98683 0.99163 3.0091e-006 1.2036e-005 0.13919 0.90845 0.89944 0.0014017 0.98177 0.55324 0.0018882 0.42746 1.7949 1.7939 16.0076 144.9807 0.0001912 -85.6144 0.57995
2.684 0.98805 5.5085e-005 3.8182 0.012013 3.5237e-005 0.0011555 0.211 0.00065911 0.21165 0.19472 0 0.033427 0.0389 0 1.0394 0.31394 0.090031 0.012061 5.3267 0.075272 9.2265e-005 0.81482 0.0061647 0.0069337 0.0013949 0.98683 0.99163 3.0089e-006 1.2036e-005 0.1392 0.90868 0.89956 0.0014016 0.98187 0.55339 0.0018882 0.42747 1.7955 1.7945 16.0075 144.9808 0.00019103 -85.6147 0.58095
2.685 0.98805 5.5085e-005 3.8182 0.012013 3.525e-005 0.0011555 0.21102 0.00065911 0.21167 0.19474 0 0.033426 0.0389 0 1.0395 0.31399 0.090047 0.012062 5.3278 0.075283 9.228e-005 0.81481 0.0061654 0.0069344 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.1392 0.90892 0.89967 0.0014016 0.98197 0.55355 0.0018881 0.42749 1.7962 1.7952 16.0075 144.9808 0.00019085 -85.6151 0.58195
2.686 0.98805 5.5085e-005 3.8182 0.012013 3.5263e-005 0.0011555 0.21104 0.00065911 0.21169 0.19476 0 0.033425 0.0389 0 1.0396 0.31403 0.090062 0.012064 5.3288 0.075294 9.2295e-005 0.8148 0.0061661 0.0069352 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.13921 0.90915 0.89978 0.0014016 0.98207 0.5537 0.0018881 0.4275 1.7968 1.7958 16.0075 144.9808 0.00019067 -85.6155 0.58295
2.687 0.98805 5.5085e-005 3.8182 0.012013 3.5276e-005 0.0011555 0.21105 0.00065911 0.21171 0.19478 0 0.033424 0.0389 0 1.0396 0.31408 0.090078 0.012066 5.3298 0.075305 9.231e-005 0.81479 0.0061669 0.0069359 0.0013946 0.98684 0.99163 3.0083e-006 1.2033e-005 0.13921 0.90938 0.89989 0.0014015 0.98216 0.55386 0.001888 0.42751 1.7974 1.7964 16.0075 144.9808 0.0001905 -85.6159 0.58395
2.688 0.98805 5.5085e-005 3.8182 0.012013 3.5289e-005 0.0011555 0.21107 0.00065911 0.21173 0.1948 0 0.033423 0.0389 0 1.0397 0.31412 0.090094 0.012068 5.3308 0.075316 9.2325e-005 0.81478 0.0061676 0.0069367 0.0013946 0.98684 0.99163 3.0081e-006 1.2032e-005 0.13922 0.90961 0.90001 0.0014015 0.98226 0.55401 0.0018879 0.42753 1.7981 1.7971 16.0075 144.9808 0.00019032 -85.6162 0.58495
2.689 0.98805 5.5085e-005 3.8182 0.012013 3.5302e-005 0.0011555 0.21109 0.00065911 0.21175 0.19482 0 0.033422 0.0389 0 1.0398 0.31417 0.09011 0.012069 5.3319 0.075328 9.234e-005 0.81476 0.0061683 0.0069374 0.0013945 0.98684 0.99164 3.0079e-006 1.2032e-005 0.13923 0.90984 0.90012 0.0014014 0.98236 0.55417 0.0018879 0.42754 1.7987 1.7977 16.0074 144.9809 0.00019015 -85.6166 0.58595
2.69 0.98805 5.5085e-005 3.8182 0.012013 3.5316e-005 0.0011555 0.21111 0.00065911 0.21177 0.19483 0 0.033421 0.0389 0 1.0399 0.31421 0.090126 0.012071 5.3329 0.075339 9.2355e-005 0.81475 0.006169 0.0069382 0.0013944 0.98684 0.99164 3.0077e-006 1.2031e-005 0.13923 0.91007 0.90023 0.0014014 0.98245 0.55432 0.0018878 0.42755 1.7993 1.7983 16.0074 144.9809 0.00018998 -85.6169 0.58695
2.691 0.98805 5.5085e-005 3.8182 0.012013 3.5329e-005 0.0011555 0.21113 0.00065911 0.21179 0.19485 0 0.03342 0.0389 0 1.04 0.31426 0.090142 0.012073 5.3339 0.07535 9.237e-005 0.81474 0.0061697 0.0069389 0.0013943 0.98684 0.99164 3.0075e-006 1.203e-005 0.13924 0.9103 0.90034 0.0014013 0.98255 0.55448 0.0018878 0.42756 1.8 1.799 16.0074 144.9809 0.0001898 -85.6173 0.58795
2.692 0.98805 5.5085e-005 3.8182 0.012013 3.5342e-005 0.0011555 0.21115 0.00065911 0.21181 0.19487 0 0.033419 0.0389 0 1.0401 0.3143 0.090158 0.012075 5.335 0.075361 9.2385e-005 0.81473 0.0061704 0.0069396 0.0013942 0.98684 0.99164 3.0073e-006 1.2029e-005 0.13924 0.91053 0.90045 0.0014013 0.98264 0.55463 0.0018877 0.42758 1.8006 1.7996 16.0074 144.9809 0.00018963 -85.6177 0.58895
2.693 0.98805 5.5085e-005 3.8182 0.012013 3.5355e-005 0.0011555 0.21117 0.00065911 0.21183 0.19489 0 0.033418 0.0389 0 1.0402 0.31435 0.090174 0.012077 5.336 0.075372 9.24e-005 0.81472 0.0061711 0.0069404 0.0013941 0.98684 0.99164 3.0072e-006 1.2029e-005 0.13925 0.91076 0.90056 0.0014012 0.98274 0.55479 0.0018876 0.42759 1.8012 1.8002 16.0074 144.9809 0.00018946 -85.618 0.58995
2.694 0.98805 5.5085e-005 3.8182 0.012013 3.5368e-005 0.0011555 0.21119 0.00065911 0.21185 0.19491 0 0.033417 0.0389 0 1.0403 0.31439 0.09019 0.012078 5.337 0.075383 9.2415e-005 0.81471 0.0061718 0.0069411 0.0013941 0.98684 0.99164 3.007e-006 1.2028e-005 0.13926 0.91099 0.90067 0.0014012 0.98283 0.55494 0.0018876 0.4276 1.8019 1.8009 16.0073 144.981 0.00018929 -85.6184 0.59095
2.695 0.98805 5.5084e-005 3.8182 0.012013 3.5381e-005 0.0011555 0.21121 0.00065911 0.21186 0.19493 0 0.033416 0.0389 0 1.0404 0.31444 0.090206 0.01208 5.3381 0.075395 9.243e-005 0.8147 0.0061725 0.0069419 0.001394 0.98684 0.99164 3.0068e-006 1.2027e-005 0.13926 0.91121 0.90078 0.0014012 0.98292 0.5551 0.0018875 0.42762 1.8025 1.8015 16.0073 144.981 0.00018912 -85.6187 0.59195
2.696 0.98805 5.5084e-005 3.8182 0.012013 3.5394e-005 0.0011555 0.21123 0.00065911 0.21188 0.19494 0 0.033415 0.0389 0 1.0405 0.31448 0.090221 0.012082 5.3391 0.075406 9.2444e-005 0.81469 0.0061732 0.0069426 0.0013939 0.98685 0.99164 3.0066e-006 1.2026e-005 0.13927 0.91144 0.90088 0.0014011 0.98302 0.55525 0.0018875 0.42763 1.8031 1.8021 16.0073 144.981 0.00018895 -85.6191 0.59295
2.697 0.98805 5.5084e-005 3.8182 0.012013 3.5407e-005 0.0011555 0.21125 0.00065911 0.2119 0.19496 0 0.033414 0.0389 0 1.0406 0.31453 0.090237 0.012084 5.3401 0.075417 9.2459e-005 0.81468 0.0061739 0.0069434 0.0013938 0.98685 0.99164 3.0064e-006 1.2026e-005 0.13927 0.91167 0.90099 0.0014011 0.98311 0.55541 0.0018874 0.42764 1.8037 1.8027 16.0073 144.981 0.00018878 -85.6194 0.59395
2.698 0.98805 5.5084e-005 3.8182 0.012013 3.542e-005 0.0011555 0.21127 0.00065911 0.21192 0.19498 0 0.033413 0.0389 0 1.0407 0.31457 0.090253 0.012085 5.3412 0.075428 9.2474e-005 0.81466 0.0061746 0.0069441 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.13928 0.91189 0.9011 0.001401 0.9832 0.55556 0.0018874 0.42765 1.8043 1.8034 16.0073 144.981 0.00018861 -85.6198 0.59495
2.699 0.98805 5.5084e-005 3.8182 0.012013 3.5433e-005 0.0011555 0.21129 0.00065911 0.21194 0.195 0 0.033412 0.0389 0 1.0408 0.31462 0.090269 0.012087 5.3422 0.075439 9.2489e-005 0.81465 0.0061753 0.0069449 0.0013937 0.98685 0.99164 3.0061e-006 1.2024e-005 0.13928 0.91211 0.90121 0.001401 0.98329 0.55572 0.0018873 0.42767 1.805 1.804 16.0072 144.9811 0.00018844 -85.6201 0.59595
2.7 0.98805 5.5084e-005 3.8182 0.012013 3.5446e-005 0.0011555 0.21131 0.00065911 0.21196 0.19502 0 0.033411 0.0389 0 1.0409 0.31466 0.090285 0.012089 5.3432 0.07545 9.2504e-005 0.81464 0.006176 0.0069456 0.0013936 0.98685 0.99164 3.0059e-006 1.2023e-005 0.13929 0.91234 0.90131 0.0014009 0.98338 0.55587 0.0018873 0.42768 1.8056 1.8046 16.0072 144.9811 0.00018828 -85.6204 0.59695
2.701 0.98805 5.5084e-005 3.8182 0.012013 3.5459e-005 0.0011555 0.21133 0.00065911 0.21198 0.19504 0 0.03341 0.0389 0 1.041 0.31471 0.090301 0.012091 5.3443 0.075462 9.2519e-005 0.81463 0.0061767 0.0069463 0.0013935 0.98685 0.99164 3.0057e-006 1.2023e-005 0.1393 0.91256 0.90142 0.0014009 0.98347 0.55602 0.0018872 0.42769 1.8062 1.8052 16.0072 144.9811 0.00018811 -85.6208 0.59795
2.702 0.98805 5.5084e-005 3.8182 0.012013 3.5472e-005 0.0011555 0.21134 0.00065912 0.212 0.19505 0 0.033409 0.0389 0 1.0411 0.31475 0.090317 0.012093 5.3453 0.075473 9.2534e-005 0.81462 0.0061774 0.0069471 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.1393 0.91278 0.90153 0.0014008 0.98356 0.55618 0.0018872 0.42771 1.8068 1.8058 16.0072 144.9811 0.00018794 -85.6211 0.59895
2.703 0.98805 5.5084e-005 3.8182 0.012013 3.5485e-005 0.0011555 0.21136 0.00065912 0.21202 0.19507 0 0.033408 0.0389 0 1.0412 0.3148 0.090333 0.012094 5.3464 0.075484 9.2549e-005 0.81461 0.0061781 0.0069478 0.0013933 0.98685 0.99164 3.0053e-006 1.2021e-005 0.13931 0.913 0.90163 0.0014008 0.98365 0.55633 0.0018871 0.42772 1.8074 1.8065 16.0072 144.9812 0.00018778 -85.6214 0.59995
2.704 0.98805 5.5084e-005 3.8182 0.012013 3.5499e-005 0.0011555 0.21138 0.00065912 0.21204 0.19509 0 0.033407 0.0389 0 1.0413 0.31484 0.090349 0.012096 5.3474 0.075495 9.2564e-005 0.8146 0.0061789 0.0069486 0.0013933 0.98685 0.99165 3.0052e-006 1.2021e-005 0.13931 0.91322 0.90174 0.0014008 0.98374 0.55649 0.001887 0.42773 1.808 1.8071 16.0071 144.9812 0.00018761 -85.6218 0.60095
2.705 0.98805 5.5084e-005 3.8182 0.012013 3.5512e-005 0.0011555 0.2114 0.00065912 0.21206 0.19511 0 0.033406 0.0389 0 1.0414 0.31489 0.090365 0.012098 5.3484 0.075506 9.2579e-005 0.81459 0.0061796 0.0069493 0.0013932 0.98685 0.99165 3.005e-006 1.202e-005 0.13932 0.91344 0.90184 0.0014007 0.98382 0.55664 0.001887 0.42774 1.8086 1.8077 16.0071 144.9812 0.00018745 -85.6221 0.60195
2.706 0.98805 5.5084e-005 3.8182 0.012013 3.5525e-005 0.0011555 0.21142 0.00065912 0.21208 0.19513 0 0.033405 0.0389 0 1.0415 0.31493 0.090381 0.0121 5.3495 0.075517 9.2594e-005 0.81458 0.0061803 0.0069501 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.13932 0.91366 0.90195 0.0014007 0.98391 0.5568 0.0018869 0.42776 1.8093 1.8083 16.0071 144.9812 0.00018729 -85.6224 0.60295
2.707 0.98805 5.5084e-005 3.8182 0.012013 3.5538e-005 0.0011555 0.21144 0.00065912 0.21209 0.19514 0 0.033404 0.0389 0 1.0416 0.31497 0.090397 0.012102 5.3505 0.075528 9.2609e-005 0.81456 0.006181 0.0069508 0.001393 0.98686 0.99165 3.0046e-006 1.2019e-005 0.13933 0.91388 0.90205 0.0014007 0.984 0.55695 0.0018869 0.42777 1.8099 1.8089 16.0071 144.9812 0.00018712 -85.6227 0.60395
2.708 0.98805 5.5084e-005 3.8182 0.012013 3.5551e-005 0.0011555 0.21146 0.00065912 0.21211 0.19516 0 0.033403 0.0389 0 1.0417 0.31502 0.090412 0.012103 5.3516 0.07554 9.2624e-005 0.81455 0.0061817 0.0069516 0.001393 0.98686 0.99165 3.0045e-006 1.2018e-005 0.13934 0.9141 0.90215 0.0014006 0.98408 0.5571 0.0018868 0.42778 1.8105 1.8095 16.0071 144.9813 0.00018696 -85.623 0.60495
2.709 0.98805 5.5084e-005 3.8182 0.012013 3.5564e-005 0.0011555 0.21148 0.00065912 0.21213 0.19518 0 0.033402 0.0389 0 1.0418 0.31506 0.090428 0.012105 5.3526 0.075551 9.2639e-005 0.81454 0.0061824 0.0069523 0.0013929 0.98686 0.99165 3.0043e-006 1.2017e-005 0.13934 0.91431 0.90226 0.0014006 0.98417 0.55726 0.0018868 0.42779 1.8111 1.8101 16.007 144.9813 0.0001868 -85.6234 0.60595
2.71 0.98805 5.5083e-005 3.8182 0.012013 3.5577e-005 0.0011555 0.2115 0.00065912 0.21215 0.1952 0 0.033401 0.0389 0 1.0419 0.31511 0.090444 0.012107 5.3536 0.075562 9.2654e-005 0.81453 0.0061831 0.006953 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.13935 0.91453 0.90236 0.0014005 0.98425 0.55741 0.0018867 0.42781 1.8117 1.8107 16.007 144.9813 0.00018664 -85.6237 0.60695
2.711 0.98805 5.5083e-005 3.8182 0.012013 3.559e-005 0.0011555 0.21152 0.00065912 0.21217 0.19522 0 0.0334 0.0389 0 1.042 0.31515 0.09046 0.012109 5.3547 0.075573 9.2669e-005 0.81452 0.0061838 0.0069538 0.0013928 0.98686 0.99165 3.004e-006 1.2016e-005 0.13935 0.91475 0.90246 0.0014005 0.98433 0.55757 0.0018867 0.42782 1.8123 1.8113 16.007 144.9813 0.00018648 -85.624 0.60795
2.712 0.98805 5.5083e-005 3.8182 0.012013 3.5603e-005 0.0011555 0.21154 0.00065912 0.21219 0.19523 0 0.033399 0.0389 0 1.0421 0.3152 0.090476 0.01211 5.3557 0.075584 9.2684e-005 0.81451 0.0061845 0.0069545 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.13936 0.91496 0.90256 0.0014005 0.98442 0.55772 0.0018866 0.42783 1.8129 1.8119 16.007 144.9813 0.00018632 -85.6243 0.60895
2.713 0.98805 5.5083e-005 3.8182 0.012013 3.5616e-005 0.0011555 0.21155 0.00065912 0.21221 0.19525 0 0.033398 0.0389 0 1.0422 0.31524 0.090492 0.012112 5.3568 0.075595 9.2698e-005 0.8145 0.0061852 0.0069553 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.13936 0.91517 0.90267 0.0014004 0.9845 0.55787 0.0018866 0.42785 1.8135 1.8125 16.007 144.9814 0.00018616 -85.6246 0.60995
2.714 0.98805 5.5083e-005 3.8182 0.012013 3.5629e-005 0.0011555 0.21157 0.00065912 0.21223 0.19527 0 0.033397 0.0389 0 1.0423 0.31529 0.090508 0.012114 5.3578 0.075606 9.2713e-005 0.81449 0.0061859 0.006956 0.0013925 0.98686 0.99165 3.0035e-006 1.2014e-005 0.13937 0.91539 0.90277 0.0014004 0.98458 0.55803 0.0018865 0.42786 1.8141 1.8131 16.0069 144.9814 0.000186 -85.6249 0.61095
2.715 0.98805 5.5083e-005 3.8182 0.012013 3.5642e-005 0.0011555 0.21159 0.00065912 0.21225 0.19529 0 0.033396 0.0389 0 1.0424 0.31533 0.090524 0.012116 5.3588 0.075618 9.2728e-005 0.81448 0.0061866 0.0069568 0.0013925 0.98686 0.99165 3.0033e-006 1.2013e-005 0.13938 0.9156 0.90287 0.0014003 0.98466 0.55818 0.0018865 0.42787 1.8147 1.8137 16.0069 144.9814 0.00018584 -85.6252 0.61195
2.716 0.98805 5.5083e-005 3.8182 0.012013 3.5655e-005 0.0011555 0.21161 0.00065912 0.21227 0.19531 0 0.033395 0.0389 0 1.0425 0.31538 0.09054 0.012118 5.3599 0.075629 9.2743e-005 0.81446 0.0061873 0.0069575 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.13938 0.91581 0.90297 0.0014003 0.98475 0.55833 0.0018864 0.42788 1.8153 1.8143 16.0069 144.9814 0.00018568 -85.6255 0.61295
2.717 0.98805 5.5083e-005 3.8182 0.012013 3.5668e-005 0.0011555 0.21163 0.00065912 0.21229 0.19532 0 0.033394 0.0389 0 1.0426 0.31542 0.090556 0.012119 5.3609 0.07564 9.2758e-005 0.81445 0.006188 0.0069583 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.13939 0.91602 0.90307 0.0014002 0.98483 0.55849 0.0018864 0.4279 1.8159 1.8149 16.0069 144.9814 0.00018553 -85.6258 0.61395
2.718 0.98805 5.5083e-005 3.8182 0.012013 3.5681e-005 0.0011555 0.21165 0.00065912 0.2123 0.19534 0 0.033393 0.0389 0 1.0427 0.31547 0.090572 0.012121 5.362 0.075651 9.2773e-005 0.81444 0.0061888 0.006959 0.0013923 0.98687 0.99165 3.0028e-006 1.2011e-005 0.13939 0.91624 0.90317 0.0014002 0.98491 0.55864 0.0018863 0.42791 1.8164 1.8155 16.0068 144.9815 0.00018537 -85.6261 0.61495
2.719 0.98805 5.5083e-005 3.8182 0.012013 3.5695e-005 0.0011555 0.21167 0.00065912 0.21232 0.19536 0 0.033392 0.0389 0 1.0428 0.31551 0.090588 0.012123 5.363 0.075662 9.2788e-005 0.81443 0.0061895 0.0069598 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.1394 0.91645 0.90327 0.0014002 0.98499 0.5588 0.0018863 0.42792 1.817 1.8161 16.0068 144.9815 0.00018521 -85.6264 0.61595
2.72 0.98805 5.5083e-005 3.8182 0.012013 3.5708e-005 0.0011555 0.21169 0.00065912 0.21234 0.19538 0 0.033391 0.0389 0 1.0429 0.31556 0.090604 0.012125 5.3641 0.075673 9.2803e-005 0.81442 0.0061902 0.0069605 0.0013921 0.98687 0.99166 3.0025e-006 1.201e-005 0.13941 0.91666 0.90337 0.0014001 0.98507 0.55895 0.0018863 0.42793 1.8176 1.8167 16.0068 144.9815 0.00018506 -85.6267 0.61695
2.721 0.98805 5.5083e-005 3.8182 0.012013 3.5721e-005 0.0011555 0.21171 0.00065912 0.21236 0.1954 0 0.03339 0.0389 0 1.043 0.3156 0.090619 0.012126 5.3651 0.075685 9.2818e-005 0.81441 0.0061909 0.0069613 0.0013921 0.98687 0.99166 3.0024e-006 1.2009e-005 0.13941 0.91686 0.90347 0.0014001 0.98514 0.5591 0.0018862 0.42795 1.8182 1.8173 16.0068 144.9815 0.0001849 -85.627 0.61795
2.722 0.98805 5.5083e-005 3.8182 0.012013 3.5734e-005 0.0011555 0.21173 0.00065912 0.21238 0.19541 0 0.033389 0.0389 0 1.0431 0.31565 0.090635 0.012128 5.3661 0.075696 9.2833e-005 0.8144 0.0061916 0.006962 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.13942 0.91707 0.90357 0.0014001 0.98522 0.55926 0.0018862 0.42796 1.8188 1.8179 16.0068 144.9815 0.00018475 -85.6273 0.61895
2.723 0.98805 5.5083e-005 3.8182 0.012013 3.5747e-005 0.0011555 0.21174 0.00065912 0.2124 0.19543 0 0.033388 0.0389 0 1.0432 0.31569 0.090651 0.01213 5.3672 0.075707 9.2848e-005 0.81439 0.0061923 0.0069628 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.13942 0.91728 0.90366 0.0014 0.9853 0.55941 0.0018861 0.42797 1.8194 1.8185 16.0067 144.9816 0.00018459 -85.6276 0.61995
2.724 0.98805 5.5083e-005 3.8182 0.012013 3.576e-005 0.0011555 0.21176 0.00065912 0.21242 0.19545 0 0.033387 0.0389 0 1.0433 0.31574 0.090667 0.012132 5.3682 0.075718 9.2863e-005 0.81437 0.006193 0.0069635 0.0013918 0.98687 0.99166 3.0019e-006 1.2008e-005 0.13943 0.91749 0.90376 0.0014 0.98538 0.55956 0.0018861 0.42799 1.82 1.8191 16.0067 144.9816 0.00018444 -85.6279 0.62095
2.725 0.98805 5.5082e-005 3.8182 0.012013 3.5773e-005 0.0011555 0.21178 0.00065912 0.21244 0.19547 0 0.033386 0.0389 0 1.0434 0.31578 0.090683 0.012134 5.3693 0.075729 9.2878e-005 0.81436 0.0061937 0.0069642 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.13943 0.91769 0.90386 0.0014 0.98545 0.55972 0.001886 0.428 1.8206 1.8196 16.0067 144.9816 0.00018429 -85.6282 0.62195
2.726 0.98805 5.5082e-005 3.8182 0.012013 3.5786e-005 0.0011555 0.2118 0.00065912 0.21246 0.19549 0 0.033385 0.0389 0 1.0435 0.31583 0.090699 0.012135 5.3703 0.07574 9.2893e-005 0.81435 0.0061944 0.006965 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.13944 0.9179 0.90396 0.0013999 0.98553 0.55987 0.001886 0.42801 1.8211 1.8202 16.0067 144.9816 0.00018414 -85.6285 0.62295
2.727 0.98805 5.5082e-005 3.8182 0.012013 3.5799e-005 0.0011555 0.21182 0.00065912 0.21247 0.1955 0 0.033384 0.0389 0 1.0436 0.31587 0.090715 0.012137 5.3714 0.075751 9.2908e-005 0.81434 0.0061951 0.0069657 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.13945 0.9181 0.90405 0.0013999 0.98561 0.56002 0.0018859 0.42802 1.8217 1.8208 16.0066 144.9816 0.00018398 -85.6287 0.62395
2.728 0.98805 5.5082e-005 3.8182 0.012013 3.5812e-005 0.0011555 0.21184 0.00065912 0.21249 0.19552 0 0.033383 0.0389 0 1.0437 0.31592 0.090731 0.012139 5.3724 0.075763 9.2923e-005 0.81433 0.0061958 0.0069665 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.13945 0.91831 0.90415 0.0013999 0.98568 0.56017 0.0018859 0.42804 1.8223 1.8214 16.0066 144.9817 0.00018383 -85.629 0.62495
2.729 0.98805 5.5082e-005 3.8182 0.012013 3.5825e-005 0.0011555 0.21186 0.00065912 0.21251 0.19554 0 0.033382 0.0389 0 1.0438 0.31596 0.090747 0.012141 5.3735 0.075774 9.2938e-005 0.81432 0.0061965 0.0069672 0.0013915 0.98688 0.99166 3.0012e-006 1.2005e-005 0.13946 0.91851 0.90425 0.0013998 0.98576 0.56033 0.0018858 0.42805 1.8229 1.822 16.0066 144.9817 0.00018368 -85.6293 0.62595
2.73 0.98805 5.5082e-005 3.8182 0.012013 3.5838e-005 0.0011555 0.21188 0.00065912 0.21253 0.19556 0 0.033381 0.0389 0 1.0439 0.31601 0.090763 0.012143 5.3745 0.075785 9.2952e-005 0.81431 0.0061972 0.006968 0.0013915 0.98688 0.99166 3.001e-006 1.2004e-005 0.13946 0.91872 0.90434 0.0013998 0.98583 0.56048 0.0018858 0.42806 1.8234 1.8225 16.0066 144.9817 0.00018353 -85.6296 0.62695
2.731 0.98805 5.5082e-005 3.8182 0.012013 3.5851e-005 0.0011555 0.21189 0.00065912 0.21255 0.19557 0 0.03338 0.0389 0 1.044 0.31605 0.090779 0.012144 5.3756 0.075796 9.2967e-005 0.8143 0.006198 0.0069687 0.0013914 0.98688 0.99166 3.0009e-006 1.2003e-005 0.13947 0.91892 0.90444 0.0013998 0.9859 0.56063 0.0018858 0.42807 1.824 1.8231 16.0066 144.9817 0.00018338 -85.6298 0.62795
2.732 0.98805 5.5082e-005 3.8182 0.012013 3.5864e-005 0.0011555 0.21191 0.00065912 0.21257 0.19559 0 0.033379 0.0389 0 1.0441 0.3161 0.090795 0.012146 5.3766 0.075807 9.2982e-005 0.81429 0.0061987 0.0069695 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.13947 0.91912 0.90453 0.0013997 0.98598 0.56079 0.0018857 0.42809 1.8246 1.8237 16.0065 144.9817 0.00018323 -85.6301 0.62895
2.733 0.98805 5.5082e-005 3.8182 0.012013 3.5878e-005 0.0011555 0.21193 0.00065912 0.21259 0.19561 0 0.033378 0.0389 0 1.0442 0.31614 0.090811 0.012148 5.3777 0.075818 9.2997e-005 0.81427 0.0061994 0.0069702 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.13948 0.91932 0.90463 0.0013997 0.98605 0.56094 0.0018857 0.4281 1.8252 1.8243 16.0065 144.9818 0.00018309 -85.6304 0.62995
2.734 0.98805 5.5082e-005 3.8182 0.012013 3.5891e-005 0.0011555 0.21195 0.00065912 0.21261 0.19563 0 0.033377 0.0389 0 1.0443 0.31619 0.090827 0.01215 5.3787 0.075829 9.3012e-005 0.81426 0.0062001 0.006971 0.0013912 0.98688 0.99166 3.0004e-006 1.2002e-005 0.13949 0.91952 0.90472 0.0013997 0.98612 0.56109 0.0018856 0.42811 1.8257 1.8248 16.0065 144.9818 0.00018294 -85.6307 0.63095
2.735 0.98805 5.5082e-005 3.8182 0.012013 3.5904e-005 0.0011555 0.21197 0.00065912 0.21262 0.19565 0 0.033376 0.0389 0 1.0443 0.31623 0.090842 0.012151 5.3798 0.075841 9.3027e-005 0.81425 0.0062008 0.0069717 0.0013911 0.98688 0.99166 3.0003e-006 1.2001e-005 0.13949 0.91972 0.90481 0.0013996 0.98619 0.56124 0.0018856 0.42813 1.8263 1.8254 16.0065 144.9818 0.00018279 -85.6309 0.63195
2.736 0.98805 5.5082e-005 3.8182 0.012013 3.5917e-005 0.0011555 0.21199 0.00065912 0.21264 0.19566 0 0.033375 0.0389 0 1.0444 0.31628 0.090858 0.012153 5.3808 0.075852 9.3042e-005 0.81424 0.0062015 0.0069725 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.1395 0.91992 0.90491 0.0013996 0.98626 0.5614 0.0018855 0.42814 1.8269 1.826 16.0064 144.9818 0.00018264 -85.6312 0.63295
2.737 0.98805 5.5082e-005 3.8182 0.012013 3.593e-005 0.0011556 0.21201 0.00065912 0.21266 0.19568 0 0.033374 0.0389 0 1.0445 0.31632 0.090874 0.012155 5.3819 0.075863 9.3057e-005 0.81423 0.0062022 0.0069732 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.1395 0.92012 0.905 0.0013996 0.98634 0.56155 0.0018855 0.42815 1.8274 1.8265 16.0064 144.9818 0.0001825 -85.6315 0.63395
2.738 0.98805 5.5082e-005 3.8182 0.012013 3.5943e-005 0.0011556 0.21203 0.00065912 0.21268 0.1957 0 0.033373 0.0389 0 1.0446 0.31637 0.09089 0.012157 5.3829 0.075874 9.3072e-005 0.81422 0.0062029 0.006974 0.001391 0.98688 0.99166 2.9999e-006 1.1999e-005 0.13951 0.92032 0.90509 0.0013995 0.98641 0.5617 0.0018855 0.42816 1.828 1.8271 16.0064 144.9819 0.00018235 -85.6317 0.63495
2.739 0.98805 5.5081e-005 3.8182 0.012012 3.5956e-005 0.0011556 0.21204 0.00065912 0.2127 0.19572 0 0.033372 0.0389 0 1.0447 0.31641 0.090906 0.012159 5.384 0.075885 9.3087e-005 0.81421 0.0062036 0.0069747 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.13952 0.92052 0.90519 0.0013995 0.98648 0.56186 0.0018854 0.42818 1.8286 1.8277 16.0064 144.9819 0.00018221 -85.632 0.63595
2.74 0.98805 5.5081e-005 3.8182 0.012012 3.5969e-005 0.0011556 0.21206 0.00065912 0.21272 0.19573 0 0.033371 0.0389 0 1.0448 0.31645 0.090922 0.01216 5.385 0.075896 9.3102e-005 0.8142 0.0062043 0.0069755 0.0013908 0.98688 0.99167 2.9996e-006 1.1998e-005 0.13952 0.92071 0.90528 0.0013995 0.98655 0.56201 0.0018854 0.42819 1.8291 1.8282 16.0064 144.9819 0.00018206 -85.6322 0.63695
2.741 0.98805 5.5081e-005 3.8182 0.012012 3.5982e-005 0.0011556 0.21208 0.00065912 0.21274 0.19575 0 0.03337 0.0389 0 1.0449 0.3165 0.090938 0.012162 5.3861 0.075907 9.3117e-005 0.81419 0.006205 0.0069762 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.13953 0.92091 0.90537 0.0013995 0.98661 0.56216 0.0018853 0.4282 1.8297 1.8288 16.0063 144.9819 0.00018192 -85.6325 0.63795
2.742 0.98805 5.5081e-005 3.8182 0.012012 3.5995e-005 0.0011556 0.2121 0.00065912 0.21275 0.19577 0 0.033369 0.0389 0 1.045 0.31654 0.090954 0.012164 5.3871 0.075919 9.3132e-005 0.81417 0.0062058 0.006977 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.13953 0.9211 0.90546 0.0013994 0.98668 0.56231 0.0018853 0.42821 1.8302 1.8294 16.0063 144.9819 0.00018177 -85.6327 0.63895
2.743 0.98805 5.5081e-005 3.8182 0.012012 3.6008e-005 0.0011556 0.21212 0.00065912 0.21277 0.19579 0 0.033368 0.0389 0 1.0451 0.31659 0.09097 0.012166 5.3882 0.07593 9.3147e-005 0.81416 0.0062065 0.0069777 0.0013907 0.98689 0.99167 2.9992e-006 1.1997e-005 0.13954 0.9213 0.90555 0.0013994 0.98675 0.56246 0.0018852 0.42823 1.8308 1.8299 16.0063 144.982 0.00018163 -85.633 0.63995
2.744 0.98805 5.5081e-005 3.8182 0.012012 3.6021e-005 0.0011556 0.21214 0.00065912 0.21279 0.1958 0 0.033367 0.0389 0 1.0452 0.31663 0.090986 0.012167 5.3892 0.075941 9.3162e-005 0.81415 0.0062072 0.0069785 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.13954 0.92149 0.90565 0.0013994 0.98682 0.56262 0.0018852 0.42824 1.8314 1.8305 16.0063 144.982 0.00018149 -85.6332 0.64095
2.745 0.98805 5.5081e-005 3.8182 0.012012 3.6034e-005 0.0011556 0.21216 0.00065912 0.21281 0.19582 0 0.033366 0.0389 0 1.0453 0.31668 0.091002 0.012169 5.3903 0.075952 9.3177e-005 0.81414 0.0062079 0.0069792 0.0013905 0.98689 0.99167 2.9989e-006 1.1996e-005 0.13955 0.92169 0.90574 0.0013993 0.98689 0.56277 0.0018852 0.42825 1.8319 1.8311 16.0062 144.982 0.00018135 -85.6335 0.64195
2.746 0.98805 5.5081e-005 3.8182 0.012012 3.6047e-005 0.0011556 0.21217 0.00065912 0.21283 0.19584 0 0.033365 0.0389 0 1.0454 0.31672 0.091018 0.012171 5.3914 0.075963 9.3192e-005 0.81413 0.0062086 0.0069799 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.13956 0.92188 0.90583 0.0013993 0.98695 0.56292 0.0018851 0.42826 1.8325 1.8316 16.0062 144.982 0.00018121 -85.6337 0.64295
2.747 0.98805 5.5081e-005 3.8182 0.012012 3.606e-005 0.0011556 0.21219 0.00065912 0.21285 0.19586 0 0.033364 0.0389 0 1.0455 0.31677 0.091034 0.012173 5.3924 0.075974 9.3206e-005 0.81412 0.0062093 0.0069807 0.0013904 0.98689 0.99167 2.9987e-006 1.1995e-005 0.13956 0.92207 0.90592 0.0013993 0.98702 0.56307 0.0018851 0.42828 1.833 1.8322 16.0062 144.982 0.00018106 -85.634 0.64395
2.748 0.98805 5.5081e-005 3.8182 0.012012 3.6074e-005 0.0011556 0.21221 0.00065912 0.21287 0.19587 0 0.033363 0.0389 0 1.0456 0.31681 0.09105 0.012175 5.3935 0.075985 9.3221e-005 0.81411 0.00621 0.0069814 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.13957 0.92227 0.90601 0.0013992 0.98709 0.56323 0.0018851 0.42829 1.8336 1.8327 16.0062 144.9821 0.00018092 -85.6342 0.64495
2.749 0.98805 5.5081e-005 3.8182 0.012012 3.6087e-005 0.0011556 0.21223 0.00065912 0.21288 0.19589 0 0.033362 0.0389 0 1.0457 0.31686 0.091066 0.012176 5.3945 0.075997 9.3236e-005 0.8141 0.0062107 0.0069822 0.0013903 0.98689 0.99167 2.9984e-006 1.1994e-005 0.13957 0.92246 0.9061 0.0013992 0.98715 0.56338 0.001885 0.4283 1.8341 1.8333 16.0061 144.9821 0.00018078 -85.6345 0.64595
2.75 0.98805 5.5081e-005 3.8182 0.012012 3.61e-005 0.0011556 0.21225 0.00065912 0.2129 0.19591 0 0.033361 0.0389 0 1.0458 0.3169 0.091082 0.012178 5.3956 0.076008 9.3251e-005 0.81409 0.0062114 0.0069829 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.13958 0.92265 0.90618 0.0013992 0.98722 0.56353 0.001885 0.42831 1.8347 1.8338 16.0061 144.9821 0.00018064 -85.6347 0.64695
2.751 0.98805 5.5081e-005 3.8182 0.012012 3.6113e-005 0.0011556 0.21227 0.00065912 0.21292 0.19593 0 0.03336 0.0389 0 1.0459 0.31695 0.091097 0.01218 5.3966 0.076019 9.3266e-005 0.81407 0.0062121 0.0069837 0.0013902 0.98689 0.99167 2.9981e-006 1.1993e-005 0.13958 0.92284 0.90627 0.0013991 0.98728 0.56368 0.0018849 0.42833 1.8352 1.8344 16.0061 144.9821 0.0001805 -85.635 0.64795
2.752 0.98805 5.5081e-005 3.8182 0.012012 3.6126e-005 0.0011556 0.21229 0.00065912 0.21294 0.19594 0 0.033359 0.0389 0 1.046 0.31699 0.091113 0.012182 5.3977 0.07603 9.3281e-005 0.81406 0.0062128 0.0069844 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.13959 0.92303 0.90636 0.0013991 0.98734 0.56383 0.0018849 0.42834 1.8358 1.8349 16.0061 144.9821 0.00018037 -85.6352 0.64895
2.753 0.98805 5.5081e-005 3.8182 0.012012 3.6139e-005 0.0011556 0.2123 0.00065912 0.21296 0.19596 0 0.033358 0.0389 0 1.0461 0.31704 0.091129 0.012184 5.3988 0.076041 9.3296e-005 0.81405 0.0062136 0.0069852 0.0013901 0.98689 0.99167 2.9979e-006 1.1992e-005 0.1396 0.92322 0.90645 0.0013991 0.98741 0.56398 0.0018849 0.42835 1.8363 1.8355 16.0061 144.9822 0.00018023 -85.6354 0.64995
2.754 0.98805 5.508e-005 3.8182 0.012012 3.6152e-005 0.0011556 0.21232 0.00065912 0.21298 0.19598 0 0.033357 0.0389 0 1.0462 0.31708 0.091145 0.012185 5.3998 0.076052 9.3311e-005 0.81404 0.0062143 0.0069859 0.00139 0.9869 0.99167 2.9978e-006 1.1991e-005 0.1396 0.9234 0.90654 0.0013991 0.98747 0.56414 0.0018848 0.42837 1.8369 1.836 16.006 144.9822 0.00018009 -85.6357 0.65095
2.755 0.98805 5.508e-005 3.8182 0.012012 3.6165e-005 0.0011556 0.21234 0.00065912 0.213 0.196 0 0.033356 0.0389 0 1.0463 0.31713 0.091161 0.012187 5.4009 0.076063 9.3326e-005 0.81403 0.006215 0.0069867 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.13961 0.92359 0.90663 0.001399 0.98754 0.56429 0.0018848 0.42838 1.8374 1.8366 16.006 144.9822 0.00017995 -85.6359 0.65195
2.756 0.98805 5.508e-005 3.8182 0.012012 3.6178e-005 0.0011556 0.21236 0.00065912 0.21301 0.19601 0 0.033355 0.0389 0 1.0464 0.31717 0.091177 0.012189 5.4019 0.076075 9.3341e-005 0.81402 0.0062157 0.0069874 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.13961 0.92378 0.90671 0.001399 0.9876 0.56444 0.0018847 0.42839 1.838 1.8371 16.006 144.9822 0.00017982 -85.6361 0.65295
2.757 0.98805 5.508e-005 3.8182 0.012012 3.6191e-005 0.0011556 0.21238 0.00065912 0.21303 0.19603 0 0.033354 0.0389 0 1.0465 0.31722 0.091193 0.012191 5.403 0.076086 9.3356e-005 0.81401 0.0062164 0.0069882 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.13962 0.92397 0.9068 0.001399 0.98766 0.56459 0.0018847 0.4284 1.8385 1.8377 16.006 144.9822 0.00017968 -85.6364 0.65395
2.758 0.98805 5.508e-005 3.8182 0.012012 3.6204e-005 0.0011556 0.2124 0.00065913 0.21305 0.19605 0 0.033353 0.0389 0 1.0466 0.31726 0.091209 0.012192 5.4041 0.076097 9.3371e-005 0.814 0.0062171 0.0069889 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.13963 0.92415 0.90689 0.001399 0.98772 0.56474 0.0018847 0.42842 1.839 1.8382 16.0059 144.9823 0.00017954 -85.6366 0.65495
2.759 0.98805 5.508e-005 3.8182 0.012012 3.6217e-005 0.0011556 0.21241 0.00065913 0.21307 0.19607 0 0.033352 0.0389 0 1.0467 0.31731 0.091225 0.012194 5.4051 0.076108 9.3386e-005 0.81399 0.0062178 0.0069897 0.0013898 0.9869 0.99167 2.9972e-006 1.1989e-005 0.13963 0.92434 0.90697 0.0013989 0.98778 0.56489 0.0018846 0.42843 1.8396 1.8387 16.0059 144.9823 0.00017941 -85.6368 0.65595
2.76 0.98805 5.508e-005 3.8182 0.012012 3.623e-005 0.0011556 0.21243 0.00065913 0.21309 0.19608 0 0.033351 0.0389 0 1.0468 0.31735 0.091241 0.012196 5.4062 0.076119 9.3401e-005 0.81397 0.0062185 0.0069904 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.13964 0.92452 0.90706 0.0013989 0.98784 0.56505 0.0018846 0.42844 1.8401 1.8393 16.0059 144.9823 0.00017927 -85.637 0.65695
2.761 0.98805 5.508e-005 3.8182 0.012012 3.6243e-005 0.0011556 0.21245 0.00065913 0.21311 0.1961 0 0.03335 0.0389 0 1.0469 0.3174 0.091257 0.012198 5.4072 0.07613 9.3416e-005 0.81396 0.0062192 0.0069912 0.0013897 0.9869 0.99168 2.9969e-006 1.1988e-005 0.13964 0.92471 0.90714 0.0013989 0.98791 0.5652 0.0018846 0.42845 1.8407 1.8398 16.0059 144.9823 0.00017914 -85.6373 0.65795
2.762 0.98805 5.508e-005 3.8182 0.012012 3.6256e-005 0.0011556 0.21247 0.00065913 0.21312 0.19612 0 0.033349 0.0389 0 1.047 0.31744 0.091273 0.0122 5.4083 0.076141 9.3431e-005 0.81395 0.0062199 0.0069919 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.13965 0.92489 0.90723 0.0013988 0.98797 0.56535 0.0018845 0.42847 1.8412 1.8404 16.0058 144.9823 0.00017901 -85.6375 0.65895
2.763 0.98805 5.508e-005 3.8182 0.012012 3.627e-005 0.0011556 0.21249 0.00065913 0.21314 0.19614 0 0.033348 0.0389 0 1.0471 0.31749 0.091289 0.012201 5.4094 0.076153 9.3446e-005 0.81394 0.0062207 0.0069927 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.13965 0.92507 0.90731 0.0013988 0.98803 0.5655 0.0018845 0.42848 1.8417 1.8409 16.0058 144.9824 0.00017887 -85.6377 0.65995
2.764 0.98805 5.508e-005 3.8182 0.012012 3.6283e-005 0.0011556 0.21251 0.00065913 0.21316 0.19615 0 0.033347 0.0389 0 1.0472 0.31753 0.091305 0.012203 5.4104 0.076164 9.346e-005 0.81393 0.0062214 0.0069934 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.13966 0.92526 0.9074 0.0013988 0.98808 0.56565 0.0018845 0.42849 1.8423 1.8414 16.0058 144.9824 0.00017874 -85.6379 0.66095
2.765 0.98805 5.508e-005 3.8182 0.012012 3.6296e-005 0.0011556 0.21252 0.00065913 0.21318 0.19617 0 0.033346 0.0389 0 1.0473 0.31758 0.091321 0.012205 5.4115 0.076175 9.3475e-005 0.81392 0.0062221 0.0069942 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.13967 0.92544 0.90748 0.0013988 0.98814 0.5658 0.0018844 0.4285 1.8428 1.842 16.0058 144.9824 0.00017861 -85.6381 0.66195
2.766 0.98805 5.508e-005 3.8182 0.012012 3.6309e-005 0.0011556 0.21254 0.00065913 0.2132 0.19619 0 0.033345 0.0389 0 1.0474 0.31762 0.091337 0.012207 5.4125 0.076186 9.349e-005 0.81391 0.0062228 0.0069949 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.13967 0.92562 0.90757 0.0013987 0.9882 0.56595 0.0018844 0.42852 1.8433 1.8425 16.0057 144.9824 0.00017848 -85.6384 0.66295
2.767 0.98805 5.508e-005 3.8182 0.012012 3.6322e-005 0.0011556 0.21256 0.00065913 0.21321 0.1962 0 0.033344 0.0389 0 1.0475 0.31767 0.091353 0.012208 5.4136 0.076197 9.3505e-005 0.8139 0.0062235 0.0069957 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.13968 0.9258 0.90765 0.0013987 0.98826 0.5661 0.0018844 0.42853 1.8439 1.843 16.0057 144.9824 0.00017834 -85.6386 0.66395
2.768 0.98805 5.508e-005 3.8182 0.012012 3.6335e-005 0.0011556 0.21258 0.00065913 0.21323 0.19622 0 0.033343 0.0389 0 1.0476 0.31771 0.091369 0.01221 5.4147 0.076208 9.352e-005 0.81389 0.0062242 0.0069964 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.13968 0.92598 0.90774 0.0013987 0.98832 0.56625 0.0018843 0.42854 1.8444 1.8436 16.0057 144.9825 0.00017821 -85.6388 0.66495
2.769 0.98805 5.5079e-005 3.8182 0.012012 3.6348e-005 0.0011556 0.2126 0.00065913 0.21325 0.19624 0 0.033342 0.0389 0 1.0477 0.31776 0.091385 0.012212 5.4157 0.076219 9.3535e-005 0.81387 0.0062249 0.0069972 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.13969 0.92616 0.90782 0.0013987 0.98838 0.56641 0.0018843 0.42855 1.8449 1.8441 16.0057 144.9825 0.00017808 -85.639 0.66595
2.77 0.98805 5.5079e-005 3.8182 0.012012 3.6361e-005 0.0011556 0.21261 0.00065913 0.21327 0.19626 0 0.033341 0.0389 0 1.0478 0.3178 0.091401 0.012214 5.4168 0.076231 9.355e-005 0.81386 0.0062256 0.0069979 0.0013892 0.98691 0.99168 2.9959e-006 1.1983e-005 0.13969 0.92634 0.9079 0.0013986 0.98843 0.56656 0.0018843 0.42857 1.8454 1.8446 16.0056 144.9825 0.00017795 -85.6392 0.66695
2.771 0.98805 5.5079e-005 3.8182 0.012012 3.6374e-005 0.0011556 0.21263 0.00065913 0.21329 0.19627 0 0.03334 0.0389 0 1.0479 0.31785 0.091417 0.012216 5.4179 0.076242 9.3565e-005 0.81385 0.0062263 0.0069987 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.1397 0.92652 0.90798 0.0013986 0.98849 0.56671 0.0018842 0.42858 1.846 1.8451 16.0056 144.9825 0.00017782 -85.6394 0.66795
2.772 0.98805 5.5079e-005 3.8182 0.012012 3.6387e-005 0.0011556 0.21265 0.00065913 0.21331 0.19629 0 0.033339 0.0389 0 1.048 0.31789 0.091432 0.012217 5.4189 0.076253 9.358e-005 0.81384 0.0062271 0.0069994 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.13971 0.9267 0.90807 0.0013986 0.98855 0.56686 0.0018842 0.42859 1.8465 1.8457 16.0056 144.9826 0.00017769 -85.6396 0.66895
2.773 0.98805 5.5079e-005 3.8182 0.012012 3.64e-005 0.0011556 0.21267 0.00065913 0.21332 0.19631 0 0.033339 0.0389 0 1.0481 0.31794 0.091448 0.012219 5.42 0.076264 9.3595e-005 0.81383 0.0062278 0.0070002 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.13971 0.92688 0.90815 0.0013985 0.9886 0.56701 0.0018842 0.4286 1.847 1.8462 16.0056 144.9826 0.00017757 -85.6398 0.66995
2.774 0.98805 5.5079e-005 3.8182 0.012012 3.6413e-005 0.0011556 0.21269 0.00065913 0.21334 0.19632 0 0.033338 0.0389 0 1.0482 0.31798 0.091464 0.012221 5.4211 0.076275 9.361e-005 0.81382 0.0062285 0.0070009 0.001389 0.98691 0.99168 2.9955e-006 1.1982e-005 0.13972 0.92705 0.90823 0.0013985 0.98866 0.56716 0.0018841 0.42862 1.8475 1.8467 16.0055 144.9826 0.00017744 -85.64 0.67095
2.775 0.98805 5.5079e-005 3.8182 0.012012 3.6426e-005 0.0011556 0.21271 0.00065913 0.21336 0.19634 0 0.033337 0.0389 0 1.0483 0.31803 0.09148 0.012223 5.4221 0.076286 9.3625e-005 0.81381 0.0062292 0.0070017 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.13972 0.92723 0.90831 0.0013985 0.98871 0.56731 0.0018841 0.42863 1.848 1.8472 16.0055 144.9826 0.00017731 -85.6402 0.67195
2.776 0.98805 5.5079e-005 3.8182 0.012012 3.6439e-005 0.0011556 0.21272 0.00065913 0.21338 0.19636 0 0.033336 0.0389 0 1.0484 0.31807 0.091496 0.012225 5.4232 0.076297 9.364e-005 0.8138 0.0062299 0.0070024 0.0013889 0.98691 0.99168 2.9953e-006 1.1981e-005 0.13973 0.92741 0.90839 0.0013985 0.98877 0.56746 0.0018841 0.42864 1.8486 1.8478 16.0055 144.9826 0.00017718 -85.6404 0.67295
2.777 0.98805 5.5079e-005 3.8182 0.012012 3.6452e-005 0.0011556 0.21274 0.00065913 0.2134 0.19638 0 0.033335 0.0389 0 1.0485 0.31812 0.091512 0.012226 5.4243 0.076308 9.3655e-005 0.81379 0.0062306 0.0070032 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.13974 0.92758 0.90847 0.0013984 0.98882 0.56761 0.001884 0.42865 1.8491 1.8483 16.0055 144.9827 0.00017705 -85.6406 0.67395
2.778 0.98805 5.5079e-005 3.8182 0.012012 3.6465e-005 0.0011556 0.21276 0.00065913 0.21341 0.19639 0 0.033334 0.0389 0 1.0486 0.31816 0.091528 0.012228 5.4253 0.07632 9.367e-005 0.81377 0.0062313 0.0070039 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.13974 0.92776 0.90856 0.0013984 0.98888 0.56776 0.001884 0.42867 1.8496 1.8488 16.0054 144.9827 0.00017693 -85.6408 0.67495
2.779 0.98805 5.5079e-005 3.8182 0.012012 3.6479e-005 0.0011556 0.21278 0.00065913 0.21343 0.19641 0 0.033333 0.0389 0 1.0487 0.31821 0.091544 0.01223 5.4264 0.076331 9.3685e-005 0.81376 0.006232 0.0070047 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.13975 0.92793 0.90864 0.0013984 0.98893 0.56791 0.001884 0.42868 1.8501 1.8493 16.0054 144.9827 0.0001768 -85.641 0.67595
2.78 0.98805 5.5079e-005 3.8182 0.012012 3.6492e-005 0.0011556 0.2128 0.00065913 0.21345 0.19643 0 0.033332 0.0389 0 1.0488 0.31825 0.09156 0.012232 5.4275 0.076342 9.37e-005 0.81375 0.0062327 0.0070054 0.0013888 0.98691 0.99168 2.9948e-006 1.1979e-005 0.13975 0.9281 0.90872 0.0013984 0.98899 0.56806 0.0018839 0.42869 1.8506 1.8498 16.0054 144.9827 0.00017668 -85.6412 0.67695
2.781 0.98805 5.5079e-005 3.8182 0.012012 3.6505e-005 0.0011556 0.21281 0.00065913 0.21347 0.19644 0 0.033331 0.0389 0 1.0489 0.3183 0.091576 0.012233 5.4285 0.076353 9.3714e-005 0.81374 0.0062335 0.0070062 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.13976 0.92828 0.9088 0.0013984 0.98904 0.56821 0.0018839 0.42871 1.8511 1.8504 16.0054 144.9827 0.00017655 -85.6414 0.67795
2.782 0.98805 5.5079e-005 3.8182 0.012012 3.6518e-005 0.0011556 0.21283 0.00065913 0.21349 0.19646 0 0.03333 0.0389 0 1.049 0.31834 0.091592 0.012235 5.4296 0.076364 9.3729e-005 0.81373 0.0062342 0.007007 0.0013887 0.98691 0.99168 2.9946e-006 1.1978e-005 0.13976 0.92845 0.90888 0.0013983 0.98909 0.56836 0.0018839 0.42872 1.8517 1.8509 16.0054 144.9828 0.00017643 -85.6416 0.67895
2.783 0.98805 5.5079e-005 3.8182 0.012012 3.6531e-005 0.0011556 0.21285 0.00065913 0.2135 0.19648 0 0.033329 0.0389 0 1.0491 0.31839 0.091608 0.012237 5.4307 0.076375 9.3744e-005 0.81372 0.0062349 0.0070077 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.13977 0.92862 0.90895 0.0013983 0.98914 0.56851 0.0018838 0.42873 1.8522 1.8514 16.0053 144.9828 0.0001763 -85.6418 0.67995
2.784 0.98805 5.5078e-005 3.8182 0.012012 3.6544e-005 0.0011556 0.21287 0.00065913 0.21352 0.1965 0 0.033328 0.0389 0 1.0492 0.31843 0.091624 0.012239 5.4318 0.076386 9.3759e-005 0.81371 0.0062356 0.0070085 0.0013886 0.98691 0.99168 2.9944e-006 1.1978e-005 0.13978 0.92879 0.90903 0.0013983 0.9892 0.56866 0.0018838 0.42874 1.8527 1.8519 16.0053 144.9828 0.00017618 -85.642 0.68095
2.785 0.98805 5.5078e-005 3.8182 0.012012 3.6557e-005 0.0011556 0.21289 0.00065913 0.21354 0.19651 0 0.033327 0.0389 0 1.0493 0.31848 0.09164 0.012241 5.4328 0.076398 9.3774e-005 0.8137 0.0062363 0.0070092 0.0013885 0.98691 0.99168 2.9943e-006 1.1977e-005 0.13978 0.92896 0.90911 0.0013983 0.98925 0.56881 0.0018838 0.42876 1.8532 1.8524 16.0053 144.9828 0.00017606 -85.6422 0.68195
2.786 0.98805 5.5078e-005 3.8182 0.012012 3.657e-005 0.0011556 0.2129 0.00065913 0.21356 0.19653 0 0.033326 0.0389 0 1.0494 0.31852 0.091656 0.012242 5.4339 0.076409 9.3789e-005 0.81369 0.006237 0.00701 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.13979 0.92913 0.90919 0.0013982 0.9893 0.56896 0.0018837 0.42877 1.8537 1.8529 16.0053 144.9828 0.00017593 -85.6424 0.68295
2.787 0.98805 5.5078e-005 3.8182 0.012012 3.6583e-005 0.0011556 0.21292 0.00065913 0.21358 0.19655 0 0.033325 0.0389 0 1.0495 0.31857 0.091672 0.012244 5.435 0.07642 9.3804e-005 0.81367 0.0062377 0.0070107 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.13979 0.9293 0.90927 0.0013982 0.98935 0.56911 0.0018837 0.42878 1.8542 1.8534 16.0052 144.9829 0.00017581 -85.6426 0.68395
2.788 0.98805 5.5078e-005 3.8182 0.012012 3.6596e-005 0.0011556 0.21294 0.00065913 0.21359 0.19656 0 0.033324 0.0389 0 1.0495 0.31861 0.091688 0.012246 5.436 0.076431 9.3819e-005 0.81366 0.0062384 0.0070115 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.1398 0.92947 0.90935 0.0013982 0.9894 0.56926 0.0018837 0.42879 1.8547 1.8539 16.0052 144.9829 0.00017569 -85.6428 0.68495
2.789 0.98805 5.5078e-005 3.8182 0.012012 3.6609e-005 0.0011556 0.21296 0.00065913 0.21361 0.19658 0 0.033323 0.0389 0 1.0496 0.31866 0.091704 0.012248 5.4371 0.076442 9.3834e-005 0.81365 0.0062391 0.0070122 0.0013884 0.98692 0.99169 2.9939e-006 1.1976e-005 0.1398 0.92964 0.90942 0.0013982 0.98945 0.56941 0.0018837 0.42881 1.8552 1.8544 16.0052 144.9829 0.00017557 -85.643 0.68595
2.79 0.98805 5.5078e-005 3.8182 0.012012 3.6622e-005 0.0011556 0.21297 0.00065913 0.21363 0.1966 0 0.033322 0.0389 0 1.0497 0.3187 0.09172 0.012249 5.4382 0.076453 9.3849e-005 0.81364 0.0062399 0.007013 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.13981 0.92981 0.9095 0.0013982 0.9895 0.56956 0.0018836 0.42882 1.8557 1.8549 16.0051 144.9829 0.00017545 -85.6431 0.68695
2.791 0.98805 5.5078e-005 3.8182 0.012012 3.6635e-005 0.0011556 0.21299 0.00065913 0.21365 0.19661 0 0.033321 0.0389 0 1.0498 0.31875 0.091736 0.012251 5.4393 0.076464 9.3864e-005 0.81363 0.0062406 0.0070137 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.13982 0.92998 0.90958 0.0013981 0.98955 0.56971 0.0018836 0.42883 1.8562 1.8554 16.0051 144.9829 0.00017532 -85.6433 0.68795
2.792 0.98805 5.5078e-005 3.8182 0.012012 3.6648e-005 0.0011556 0.21301 0.00065913 0.21367 0.19663 0 0.03332 0.0389 0 1.0499 0.31879 0.091752 0.012253 5.4403 0.076475 9.3879e-005 0.81362 0.0062413 0.0070145 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.13982 0.93015 0.90966 0.0013981 0.9896 0.56986 0.0018836 0.42884 1.8567 1.856 16.0051 144.983 0.0001752 -85.6435 0.68895
2.793 0.98805 5.5078e-005 3.8182 0.012012 3.6661e-005 0.0011556 0.21303 0.00065913 0.21368 0.19665 0 0.033319 0.0389 0 1.05 0.31884 0.091768 0.012255 5.4414 0.076487 9.3894e-005 0.81361 0.006242 0.0070152 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.13983 0.93031 0.90973 0.0013981 0.98965 0.57001 0.0018835 0.42886 1.8572 1.8565 16.0051 144.983 0.00017508 -85.6437 0.68995
2.794 0.98805 5.5078e-005 3.8182 0.012012 3.6675e-005 0.0011556 0.21305 0.00065913 0.2137 0.19666 0 0.033319 0.0389 0 1.0501 0.31888 0.091784 0.012257 5.4425 0.076498 9.3909e-005 0.8136 0.0062427 0.007016 0.0013881 0.98692 0.99169 2.9934e-006 1.1974e-005 0.13983 0.93048 0.90981 0.0013981 0.9897 0.57016 0.0018835 0.42887 1.8577 1.857 16.005 144.983 0.00017496 -85.6439 0.69095
2.795 0.98805 5.5078e-005 3.8182 0.012012 3.6688e-005 0.0011556 0.21306 0.00065913 0.21372 0.19668 0 0.033318 0.0389 0 1.0502 0.31893 0.0918 0.012258 5.4436 0.076509 9.3924e-005 0.81359 0.0062434 0.0070167 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.13984 0.93065 0.90988 0.0013981 0.98975 0.57031 0.0018835 0.42888 1.8582 1.8575 16.005 144.983 0.00017485 -85.644 0.69195
2.796 0.98805 5.5078e-005 3.8182 0.012012 3.6701e-005 0.0011556 0.21308 0.00065913 0.21374 0.1967 0 0.033317 0.0389 0 1.0503 0.31897 0.091816 0.01226 5.4446 0.07652 9.3939e-005 0.81357 0.0062441 0.0070175 0.0013881 0.98692 0.99169 2.9932e-006 1.1973e-005 0.13985 0.93081 0.90996 0.001398 0.9898 0.57046 0.0018835 0.42889 1.8587 1.858 16.005 144.983 0.00017473 -85.6442 0.69295
2.797 0.98805 5.5078e-005 3.8182 0.012012 3.6714e-005 0.0011556 0.2131 0.00065913 0.21375 0.19672 0 0.033316 0.0389 0 1.0504 0.31902 0.091832 0.012262 5.4457 0.076531 9.3954e-005 0.81356 0.0062448 0.0070182 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.13985 0.93098 0.91004 0.001398 0.98985 0.57061 0.0018834 0.4289 1.8592 1.8585 16.005 144.9831 0.00017461 -85.6444 0.69395
2.798 0.98805 5.5078e-005 3.8182 0.012012 3.6727e-005 0.0011556 0.21312 0.00065913 0.21377 0.19673 0 0.033315 0.0389 0 1.0505 0.31906 0.091848 0.012264 5.4468 0.076542 9.3968e-005 0.81355 0.0062456 0.007019 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.13986 0.93114 0.91011 0.001398 0.98989 0.57076 0.0018834 0.42892 1.8597 1.859 16.0049 144.9831 0.00017449 -85.6446 0.69495
2.799 0.98805 5.5077e-005 3.8182 0.012012 3.674e-005 0.0011556 0.21314 0.00065913 0.21379 0.19675 0 0.033314 0.0389 0 1.0506 0.31911 0.091864 0.012265 5.4479 0.076553 9.3983e-005 0.81354 0.0062463 0.0070197 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.13986 0.9313 0.91019 0.001398 0.98994 0.57091 0.0018834 0.42893 1.8602 1.8594 16.0049 144.9831 0.00017437 -85.6447 0.69595
2.8 0.98805 5.5077e-005 3.8182 0.012012 3.6753e-005 0.0011556 0.21315 0.00065913 0.21381 0.19677 0 0.033313 0.0389 0 1.0507 0.31915 0.091879 0.012267 5.4489 0.076564 9.3998e-005 0.81353 0.006247 0.0070205 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.13987 0.93147 0.91026 0.0013979 0.98999 0.57106 0.0018833 0.42894 1.8607 1.8599 16.0049 144.9831 0.00017426 -85.6449 0.69695
2.801 0.98805 5.5077e-005 3.8182 0.012012 3.6766e-005 0.0011556 0.21317 0.00065913 0.21383 0.19678 0 0.033312 0.0389 0 1.0508 0.3192 0.091895 0.012269 5.45 0.076576 9.4013e-005 0.81352 0.0062477 0.0070212 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.13987 0.93163 0.91033 0.0013979 0.99003 0.57121 0.0018833 0.42895 1.8612 1.8604 16.0049 144.9831 0.00017414 -85.6451 0.69795
2.802 0.98805 5.5077e-005 3.8182 0.012012 3.6779e-005 0.0011556 0.21319 0.00065913 0.21384 0.1968 0 0.033311 0.0389 0 1.0509 0.31924 0.091911 0.012271 5.4511 0.076587 9.4028e-005 0.81351 0.0062484 0.007022 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.13988 0.93179 0.91041 0.0013979 0.99008 0.57136 0.0018833 0.42897 1.8617 1.8609 16.0048 144.9832 0.00017402 -85.6453 0.69895
2.803 0.98805 5.5077e-005 3.8182 0.012012 3.6792e-005 0.0011556 0.21321 0.00065913 0.21386 0.19682 0 0.03331 0.0389 0 1.051 0.31929 0.091927 0.012273 5.4522 0.076598 9.4043e-005 0.8135 0.0062491 0.0070227 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.13989 0.93195 0.91048 0.0013979 0.99013 0.57151 0.0018833 0.42898 1.8622 1.8614 16.0048 144.9832 0.00017391 -85.6454 0.69995
2.804 0.98805 5.5077e-005 3.8182 0.012012 3.6805e-005 0.0011556 0.21322 0.00065913 0.21388 0.19683 0 0.033309 0.0389 0 1.0511 0.31933 0.091943 0.012274 5.4533 0.076609 9.4058e-005 0.81349 0.0062498 0.0070235 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.13989 0.93211 0.91056 0.0013979 0.99017 0.57166 0.0018832 0.42899 1.8627 1.8619 16.0048 144.9832 0.00017379 -85.6456 0.70095
2.805 0.98805 5.5077e-005 3.8182 0.012012 3.6818e-005 0.0011556 0.21324 0.00065913 0.2139 0.19685 0 0.033308 0.0389 0 1.0512 0.31938 0.091959 0.012276 5.4543 0.07662 9.4073e-005 0.81347 0.0062505 0.0070243 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.1399 0.93228 0.91063 0.0013978 0.99022 0.5718 0.0018832 0.429 1.8632 1.8624 16.0048 144.9832 0.00017368 -85.6458 0.70195
2.806 0.98805 5.5077e-005 3.8182 0.012012 3.6831e-005 0.0011556 0.21326 0.00065913 0.21391 0.19687 0 0.033307 0.0389 0 1.0513 0.31942 0.091975 0.012278 5.4554 0.076631 9.4088e-005 0.81346 0.0062513 0.007025 0.0013877 0.98693 0.99169 2.9923e-006 1.1969e-005 0.1399 0.93244 0.9107 0.0013978 0.99026 0.57195 0.0018832 0.42902 1.8636 1.8629 16.0047 144.9832 0.00017356 -85.6459 0.70295
2.807 0.98805 5.5077e-005 3.8182 0.012012 3.6844e-005 0.0011557 0.21328 0.00065913 0.21393 0.19688 0 0.033306 0.0389 0 1.0514 0.31947 0.091991 0.01228 5.4565 0.076642 9.4103e-005 0.81345 0.006252 0.0070258 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.13991 0.93259 0.91078 0.0013978 0.99031 0.5721 0.0018832 0.42903 1.8641 1.8634 16.0047 144.9833 0.00017345 -85.6461 0.70395
2.808 0.98805 5.5077e-005 3.8182 0.012011 3.6857e-005 0.0011557 0.21329 0.00065913 0.21395 0.1969 0 0.033305 0.0389 0 1.0515 0.31951 0.092007 0.012281 5.4576 0.076653 9.4118e-005 0.81344 0.0062527 0.0070265 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.13992 0.93275 0.91085 0.0013978 0.99035 0.57225 0.0018831 0.42904 1.8646 1.8639 16.0047 144.9833 0.00017333 -85.6463 0.70495
2.809 0.98805 5.5077e-005 3.8182 0.012011 3.687e-005 0.0011557 0.21331 0.00065913 0.21397 0.19692 0 0.033304 0.0389 0 1.0516 0.31956 0.092023 0.012283 5.4587 0.076665 9.4133e-005 0.81343 0.0062534 0.0070273 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.13992 0.93291 0.91092 0.0013978 0.9904 0.5724 0.0018831 0.42905 1.8651 1.8644 16.0047 144.9833 0.00017322 -85.6464 0.70595
2.81 0.98805 5.5077e-005 3.8182 0.012011 3.6884e-005 0.0011557 0.21333 0.00065913 0.21398 0.19693 0 0.033304 0.0389 0 1.0517 0.3196 0.092039 0.012285 5.4597 0.076676 9.4148e-005 0.81342 0.0062541 0.007028 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.13993 0.93307 0.91099 0.0013977 0.99044 0.57255 0.0018831 0.42907 1.8656 1.8648 16.0046 144.9833 0.00017311 -85.6466 0.70695
2.811 0.98805 5.5077e-005 3.8182 0.012011 3.6897e-005 0.0011557 0.21335 0.00065913 0.214 0.19695 0 0.033303 0.0389 0 1.0518 0.31965 0.092055 0.012287 5.4608 0.076687 9.4163e-005 0.81341 0.0062548 0.0070288 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.13993 0.93323 0.91106 0.0013977 0.99049 0.5727 0.0018831 0.42908 1.8661 1.8653 16.0046 144.9833 0.00017299 -85.6467 0.70795
2.812 0.98805 5.5077e-005 3.8182 0.012011 3.691e-005 0.0011557 0.21336 0.00065913 0.21402 0.19697 0 0.033302 0.0389 0 1.0519 0.31969 0.092071 0.012289 5.4619 0.076698 9.4178e-005 0.8134 0.0062555 0.0070295 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.13994 0.93339 0.91114 0.0013977 0.99053 0.57285 0.001883 0.42909 1.8665 1.8658 16.0046 144.9834 0.00017288 -85.6469 0.70895
2.813 0.98805 5.5077e-005 3.8182 0.012011 3.6923e-005 0.0011557 0.21338 0.00065913 0.21404 0.19698 0 0.033301 0.0389 0 1.052 0.31974 0.092087 0.01229 5.463 0.076709 9.4193e-005 0.81339 0.0062563 0.0070303 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.13994 0.93354 0.91121 0.0013977 0.99057 0.57299 0.001883 0.4291 1.867 1.8663 16.0046 144.9834 0.00017277 -85.647 0.70995
2.814 0.98805 5.5076e-005 3.8182 0.012011 3.6936e-005 0.0011557 0.2134 0.00065913 0.21405 0.197 0 0.0333 0.0389 0 1.0521 0.31978 0.092103 0.012292 5.4641 0.07672 9.4208e-005 0.81337 0.006257 0.007031 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.13995 0.9337 0.91128 0.0013977 0.99061 0.57314 0.001883 0.42912 1.8675 1.8668 16.0045 144.9834 0.00017266 -85.6472 0.71095
2.815 0.98805 5.5076e-005 3.8182 0.012011 3.6949e-005 0.0011557 0.21342 0.00065913 0.21407 0.19702 0 0.033299 0.0389 0 1.0522 0.31983 0.092119 0.012294 5.4652 0.076731 9.4222e-005 0.81336 0.0062577 0.0070318 0.0013873 0.98693 0.99169 2.9916e-006 1.1966e-005 0.13996 0.93385 0.91135 0.0013976 0.99066 0.57329 0.0018829 0.42913 1.868 1.8672 16.0045 144.9834 0.00017255 -85.6474 0.71195
2.816 0.98805 5.5076e-005 3.8182 0.012011 3.6962e-005 0.0011557 0.21343 0.00065914 0.21409 0.19703 0 0.033298 0.0389 0 1.0523 0.31987 0.092135 0.012296 5.4662 0.076742 9.4237e-005 0.81335 0.0062584 0.0070325 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.13996 0.93401 0.91142 0.0013976 0.9907 0.57344 0.0018829 0.42914 1.8685 1.8677 16.0045 144.9834 0.00017244 -85.6475 0.71295
2.817 0.98805 5.5076e-005 3.8182 0.012011 3.6975e-005 0.0011557 0.21345 0.00065914 0.21411 0.19705 0 0.033297 0.0389 0 1.0524 0.31992 0.092151 0.012297 5.4673 0.076754 9.4252e-005 0.81334 0.0062591 0.0070333 0.0013873 0.98693 0.9917 2.9914e-006 1.1966e-005 0.13997 0.93416 0.91149 0.0013976 0.99074 0.57359 0.0018829 0.42915 1.8689 1.8682 16.0044 144.9835 0.00017233 -85.6477 0.71395
2.818 0.98805 5.5076e-005 3.8182 0.012011 3.6988e-005 0.0011557 0.21347 0.00065914 0.21412 0.19707 0 0.033296 0.0389 0 1.0525 0.31996 0.092167 0.012299 5.4684 0.076765 9.4267e-005 0.81333 0.0062598 0.0070341 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.13997 0.93432 0.91156 0.0013976 0.99078 0.57374 0.0018829 0.42917 1.8694 1.8687 16.0044 144.9835 0.00017222 -85.6478 0.71495
2.819 0.98805 5.5076e-005 3.8182 0.012011 3.7001e-005 0.0011557 0.21349 0.00065914 0.21414 0.19708 0 0.033295 0.0389 0 1.0526 0.32001 0.092183 0.012301 5.4695 0.076776 9.4282e-005 0.81332 0.0062605 0.0070348 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.13998 0.93447 0.91163 0.0013976 0.99083 0.57389 0.0018829 0.42918 1.8699 1.8692 16.0044 144.9835 0.00017211 -85.648 0.71595
2.82 0.98805 5.5076e-005 3.8182 0.012011 3.7014e-005 0.0011557 0.2135 0.00065914 0.21416 0.1971 0 0.033294 0.0389 0 1.0527 0.32005 0.092199 0.012303 5.4706 0.076787 9.4297e-005 0.81331 0.0062612 0.0070356 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.13999 0.93463 0.9117 0.0013975 0.99087 0.57403 0.0018828 0.42919 1.8704 1.8696 16.0044 144.9835 0.000172 -85.6481 0.71695
2.821 0.98805 5.5076e-005 3.8182 0.012011 3.7027e-005 0.0011557 0.21352 0.00065914 0.21418 0.19712 0 0.033293 0.0389 0 1.0528 0.3201 0.092215 0.012305 5.4717 0.076798 9.4312e-005 0.8133 0.006262 0.0070363 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.13999 0.93478 0.91177 0.0013975 0.99091 0.57418 0.0018828 0.4292 1.8708 1.8701 16.0043 144.9836 0.00017189 -85.6483 0.71795
2.822 0.98805 5.5076e-005 3.8182 0.012011 3.704e-005 0.0011557 0.21354 0.00065914 0.21419 0.19713 0 0.033292 0.0389 0 1.0529 0.32014 0.092231 0.012306 5.4728 0.076809 9.4327e-005 0.81329 0.0062627 0.0070371 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.14 0.93493 0.91184 0.0013975 0.99095 0.57433 0.0018828 0.42922 1.8713 1.8706 16.0043 144.9836 0.00017178 -85.6484 0.71895
2.823 0.98805 5.5076e-005 3.8182 0.012011 3.7053e-005 0.0011557 0.21356 0.00065914 0.21421 0.19715 0 0.033292 0.0389 0 1.053 0.32019 0.092247 0.012308 5.4738 0.07682 9.4342e-005 0.81327 0.0062634 0.0070378 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.14 0.93508 0.91191 0.0013975 0.99099 0.57448 0.0018828 0.42923 1.8718 1.871 16.0043 144.9836 0.00017167 -85.6486 0.71995
2.824 0.98805 5.5076e-005 3.8182 0.012011 3.7066e-005 0.0011557 0.21357 0.00065914 0.21423 0.19716 0 0.033291 0.0389 0 1.0531 0.32023 0.092263 0.01231 5.4749 0.076831 9.4357e-005 0.81326 0.0062641 0.0070386 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.14001 0.93523 0.91198 0.0013975 0.99103 0.57463 0.0018827 0.42924 1.8722 1.8715 16.0043 144.9836 0.00017156 -85.6487 0.72095
2.825 0.98805 5.5076e-005 3.8182 0.012011 3.708e-005 0.0011557 0.21359 0.00065914 0.21425 0.19718 0 0.03329 0.0389 0 1.0532 0.32028 0.092279 0.012312 5.476 0.076842 9.4372e-005 0.81325 0.0062648 0.0070393 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.14001 0.93539 0.91204 0.0013974 0.99107 0.57477 0.0018827 0.42925 1.8727 1.872 16.0042 144.9836 0.00017146 -85.6489 0.72195
2.826 0.98805 5.5076e-005 3.8182 0.012011 3.7093e-005 0.0011557 0.21361 0.00065914 0.21426 0.1972 0 0.033289 0.0389 0 1.0533 0.32032 0.092295 0.012313 5.4771 0.076854 9.4387e-005 0.81324 0.0062655 0.0070401 0.0013869 0.98693 0.9917 2.9907e-006 1.1963e-005 0.14002 0.93554 0.91211 0.0013974 0.99111 0.57492 0.0018827 0.42926 1.8732 1.8725 16.0042 144.9837 0.00017135 -85.649 0.72295
2.827 0.98805 5.5076e-005 3.8182 0.012011 3.7106e-005 0.0011557 0.21363 0.00065914 0.21428 0.19721 0 0.033288 0.0389 0 1.0534 0.32037 0.092311 0.012315 5.4782 0.076865 9.4402e-005 0.81323 0.0062662 0.0070408 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.14003 0.93569 0.91218 0.0013974 0.99115 0.57507 0.0018827 0.42928 1.8736 1.8729 16.0042 144.9837 0.00017124 -85.6491 0.72395
2.828 0.98805 5.5075e-005 3.8182 0.012011 3.7119e-005 0.0011557 0.21364 0.00065914 0.2143 0.19723 0 0.033287 0.0389 0 1.0535 0.32042 0.092327 0.012317 5.4793 0.076876 9.4417e-005 0.81322 0.006267 0.0070416 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.14003 0.93584 0.91225 0.0013974 0.99119 0.57522 0.0018826 0.42929 1.8741 1.8734 16.0042 144.9837 0.00017114 -85.6493 0.72495
2.829 0.98805 5.5075e-005 3.8182 0.012011 3.7132e-005 0.0011557 0.21366 0.00065914 0.21432 0.19725 0 0.033286 0.0389 0 1.0536 0.32046 0.092343 0.012319 5.4804 0.076887 9.4432e-005 0.81321 0.0062677 0.0070424 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.14004 0.93598 0.91232 0.0013974 0.99123 0.57537 0.0018826 0.4293 1.8746 1.8739 16.0041 144.9837 0.00017103 -85.6494 0.72595
2.83 0.98805 5.5075e-005 3.8182 0.012011 3.7145e-005 0.0011557 0.21368 0.00065914 0.21433 0.19726 0 0.033285 0.0389 0 1.0537 0.32051 0.092359 0.012321 5.4815 0.076898 9.4447e-005 0.8132 0.0062684 0.0070431 0.0013868 0.98694 0.9917 2.9904e-006 1.1962e-005 0.14004 0.93613 0.91238 0.0013974 0.99127 0.57551 0.0018826 0.42931 1.875 1.8743 16.0041 144.9837 0.00017092 -85.6496 0.72695
2.831 0.98805 5.5075e-005 3.8182 0.012011 3.7158e-005 0.0011557 0.2137 0.00065914 0.21435 0.19728 0 0.033284 0.0389 0 1.0538 0.32055 0.092375 0.012322 5.4826 0.076909 9.4462e-005 0.81319 0.0062691 0.0070439 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.14005 0.93628 0.91245 0.0013973 0.9913 0.57566 0.0018826 0.42933 1.8755 1.8748 16.0041 144.9838 0.00017082 -85.6497 0.72795
2.832 0.98805 5.5075e-005 3.8182 0.012011 3.7171e-005 0.0011557 0.21371 0.00065914 0.21437 0.1973 0 0.033283 0.0389 0 1.0539 0.3206 0.092391 0.012324 5.4836 0.07692 9.4476e-005 0.81317 0.0062698 0.0070446 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.14006 0.93643 0.91252 0.0013973 0.99134 0.57581 0.0018826 0.42934 1.876 1.8752 16.004 144.9838 0.00017071 -85.6498 0.72895
2.833 0.98805 5.5075e-005 3.8182 0.012011 3.7184e-005 0.0011557 0.21373 0.00065914 0.21438 0.19731 0 0.033282 0.0389 0 1.054 0.32064 0.092407 0.012326 5.4847 0.076931 9.4491e-005 0.81316 0.0062705 0.0070454 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.14006 0.93658 0.91258 0.0013973 0.99138 0.57596 0.0018825 0.42935 1.8764 1.8757 16.004 144.9838 0.00017061 -85.65 0.72995
2.834 0.98805 5.5075e-005 3.8182 0.012011 3.7197e-005 0.0011557 0.21375 0.00065914 0.2144 0.19733 0 0.033281 0.0389 0 1.0541 0.32069 0.092423 0.012328 5.4858 0.076943 9.4506e-005 0.81315 0.0062712 0.0070461 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.14007 0.93672 0.91265 0.0013973 0.99142 0.5761 0.0018825 0.42936 1.8769 1.8762 16.004 144.9838 0.00017051 -85.6501 0.73095
2.835 0.98805 5.5075e-005 3.8182 0.012011 3.721e-005 0.0011557 0.21376 0.00065914 0.21442 0.19735 0 0.033281 0.0389 0 1.0542 0.32073 0.092439 0.012329 5.4869 0.076954 9.4521e-005 0.81314 0.006272 0.0070469 0.0013867 0.98694 0.9917 2.99e-006 1.196e-005 0.14007 0.93687 0.91272 0.0013973 0.99146 0.57625 0.0018825 0.42938 1.8773 1.8766 16.004 144.9838 0.0001704 -85.6503 0.73195
2.836 0.98805 5.5075e-005 3.8182 0.012011 3.7223e-005 0.0011557 0.21378 0.00065914 0.21444 0.19736 0 0.03328 0.0389 0 1.0543 0.32078 0.092455 0.012331 5.488 0.076965 9.4536e-005 0.81313 0.0062727 0.0070476 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.14008 0.93701 0.91278 0.0013973 0.99149 0.5764 0.0018825 0.42939 1.8778 1.8771 16.0039 144.9839 0.0001703 -85.6504 0.73295
2.837 0.98805 5.5075e-005 3.8182 0.012011 3.7236e-005 0.0011557 0.2138 0.00065914 0.21445 0.19738 0 0.033279 0.0389 0 1.0544 0.32082 0.092471 0.012333 5.4891 0.076976 9.4551e-005 0.81312 0.0062734 0.0070484 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.14008 0.93716 0.91285 0.0013973 0.99153 0.57655 0.0018824 0.4294 1.8782 1.8775 16.0039 144.9839 0.0001702 -85.6505 0.73395
2.838 0.98805 5.5075e-005 3.8182 0.012011 3.7249e-005 0.0011557 0.21382 0.00065914 0.21447 0.19739 0 0.033278 0.0389 0 1.0545 0.32087 0.092487 0.012335 5.4902 0.076987 9.4566e-005 0.81311 0.0062741 0.0070491 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.14009 0.93731 0.91291 0.0013972 0.99157 0.57669 0.0018824 0.42941 1.8787 1.878 16.0039 144.9839 0.00017009 -85.6507 0.73495
2.839 0.98805 5.5075e-005 3.8182 0.012011 3.7262e-005 0.0011557 0.21383 0.00065914 0.21449 0.19741 0 0.033277 0.0389 0 1.0546 0.32091 0.092503 0.012337 5.4913 0.076998 9.4581e-005 0.8131 0.0062748 0.0070499 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.1401 0.93745 0.91298 0.0013972 0.9916 0.57684 0.0018824 0.42942 1.8792 1.8785 16.0039 144.9839 0.00016999 -85.6508 0.73595
2.84 0.98805 5.5075e-005 3.8182 0.012011 3.7275e-005 0.0011557 0.21385 0.00065914 0.21451 0.19743 0 0.033276 0.0389 0 1.0547 0.32096 0.092519 0.012338 5.4924 0.077009 9.4596e-005 0.81309 0.0062755 0.0070507 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.1401 0.93759 0.91304 0.0013972 0.99164 0.57699 0.0018824 0.42944 1.8796 1.8789 16.0038 144.9839 0.00016989 -85.6509 0.73695
2.841 0.98805 5.5075e-005 3.8182 0.012011 3.7289e-005 0.0011557 0.21387 0.00065914 0.21452 0.19744 0 0.033275 0.0389 0 1.0548 0.321 0.092535 0.01234 5.4935 0.07702 9.4611e-005 0.81307 0.0062762 0.0070514 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.14011 0.93774 0.91311 0.0013972 0.99167 0.57714 0.0018824 0.42945 1.8801 1.8794 16.0038 144.984 0.00016979 -85.651 0.73795
2.842 0.98805 5.5075e-005 3.8182 0.012011 3.7302e-005 0.0011557 0.21388 0.00065914 0.21454 0.19746 0 0.033274 0.0389 0 1.0549 0.32105 0.092551 0.012342 5.4946 0.077031 9.4626e-005 0.81306 0.006277 0.0070522 0.0013864 0.98694 0.9917 2.9896e-006 1.1958e-005 0.14011 0.93788 0.91317 0.0013972 0.99171 0.57728 0.0018823 0.42946 1.8805 1.8798 16.0038 144.984 0.00016969 -85.6512 0.73895
2.843 0.98805 5.5074e-005 3.8182 0.012011 3.7315e-005 0.0011557 0.2139 0.00065914 0.21456 0.19748 0 0.033273 0.0389 0 1.055 0.32109 0.092567 0.012344 5.4957 0.077043 9.4641e-005 0.81305 0.0062777 0.0070529 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.14012 0.93802 0.91324 0.0013972 0.99175 0.57743 0.0018823 0.42947 1.881 1.8803 16.0037 144.984 0.00016959 -85.6513 0.73995
2.844 0.98805 5.5074e-005 3.8182 0.012011 3.7328e-005 0.0011557 0.21392 0.00065914 0.21457 0.19749 0 0.033272 0.0389 0 1.0551 0.32114 0.092583 0.012345 5.4968 0.077054 9.4656e-005 0.81304 0.0062784 0.0070537 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.14012 0.93817 0.9133 0.0013971 0.99178 0.57758 0.0018823 0.42949 1.8814 1.8807 16.0037 144.984 0.00016948 -85.6514 0.74095
2.845 0.98805 5.5074e-005 3.8182 0.012011 3.7341e-005 0.0011557 0.21394 0.00065914 0.21459 0.19751 0 0.033272 0.0389 0 1.0552 0.32118 0.092599 0.012347 5.4979 0.077065 9.4671e-005 0.81303 0.0062791 0.0070544 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.14013 0.93831 0.91337 0.0013971 0.99182 0.57773 0.0018823 0.4295 1.8819 1.8812 16.0037 144.984 0.00016938 -85.6516 0.74195
2.846 0.98805 5.5074e-005 3.8182 0.012011 3.7354e-005 0.0011557 0.21395 0.00065914 0.21461 0.19752 0 0.033271 0.0389 0 1.0552 0.32123 0.092615 0.012349 5.499 0.077076 9.4686e-005 0.81302 0.0062798 0.0070552 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.14014 0.93845 0.91343 0.0013971 0.99185 0.57787 0.0018823 0.42951 1.8823 1.8816 16.0037 144.9841 0.00016928 -85.6517 0.74295
2.847 0.98805 5.5074e-005 3.8182 0.012011 3.7367e-005 0.0011557 0.21397 0.00065914 0.21462 0.19754 0 0.03327 0.0389 0 1.0553 0.32127 0.092631 0.012351 5.5 0.077087 9.4701e-005 0.81301 0.0062805 0.0070559 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.14014 0.93859 0.91349 0.0013971 0.99189 0.57802 0.0018822 0.42952 1.8828 1.8821 16.0036 144.9841 0.00016918 -85.6518 0.74395
2.848 0.98805 5.5074e-005 3.8182 0.012011 3.738e-005 0.0011557 0.21399 0.00065914 0.21464 0.19756 0 0.033269 0.0389 0 1.0554 0.32132 0.092647 0.012353 5.5011 0.077098 9.4715e-005 0.813 0.0062812 0.0070567 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.14015 0.93873 0.91356 0.0013971 0.99192 0.57817 0.0018822 0.42954 1.8832 1.8825 16.0036 144.9841 0.00016909 -85.6519 0.74495
2.849 0.98805 5.5074e-005 3.8182 0.012011 3.7393e-005 0.0011557 0.214 0.00065914 0.21466 0.19757 0 0.033268 0.0389 0 1.0555 0.32136 0.092663 0.012354 5.5022 0.077109 9.473e-005 0.81299 0.006282 0.0070575 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.14015 0.93887 0.91362 0.0013971 0.99195 0.57831 0.0018822 0.42955 1.8837 1.883 16.0036 144.9841 0.00016899 -85.6521 0.74595
2.85 0.98805 5.5074e-005 3.8182 0.012011 3.7406e-005 0.0011557 0.21402 0.00065914 0.21468 0.19759 0 0.033267 0.0389 0 1.0556 0.32141 0.092679 0.012356 5.5033 0.07712 9.4745e-005 0.81297 0.0062827 0.0070582 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.14016 0.93901 0.91368 0.0013971 0.99199 0.57846 0.0018822 0.42956 1.8841 1.8834 16.0036 144.9841 0.00016889 -85.6522 0.74695
2.851 0.98805 5.5074e-005 3.8182 0.012011 3.7419e-005 0.0011557 0.21404 0.00065914 0.21469 0.1976 0 0.033266 0.0389 0 1.0557 0.32145 0.092695 0.012358 5.5044 0.077131 9.476e-005 0.81296 0.0062834 0.007059 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.14017 0.93915 0.91374 0.001397 0.99202 0.57861 0.0018822 0.42957 1.8845 1.8839 16.0035 144.9842 0.00016879 -85.6523 0.74795
2.852 0.98805 5.5074e-005 3.8182 0.012011 3.7432e-005 0.0011557 0.21406 0.00065914 0.21471 0.19762 0 0.033265 0.0389 0 1.0558 0.3215 0.092711 0.01236 5.5055 0.077142 9.4775e-005 0.81295 0.0062841 0.0070597 0.0013861 0.98695 0.9917 2.9889e-006 1.1955e-005 0.14017 0.93929 0.91381 0.001397 0.99206 0.57875 0.0018821 0.42958 1.885 1.8843 16.0035 144.9842 0.00016869 -85.6524 0.74895
2.853 0.98805 5.5074e-005 3.8182 0.012011 3.7445e-005 0.0011557 0.21407 0.00065914 0.21473 0.19764 0 0.033264 0.0389 0 1.0559 0.32154 0.092727 0.012361 5.5066 0.077154 9.479e-005 0.81294 0.0062848 0.0070605 0.0013861 0.98695 0.9917 2.9888e-006 1.1955e-005 0.14018 0.93943 0.91387 0.001397 0.99209 0.5789 0.0018821 0.4296 1.8854 1.8848 16.0035 144.9842 0.00016859 -85.6525 0.74995
2.854 0.98805 5.5074e-005 3.8182 0.012011 3.7458e-005 0.0011557 0.21409 0.00065914 0.21474 0.19765 0 0.033263 0.0389 0 1.056 0.32159 0.092743 0.012363 5.5077 0.077165 9.4805e-005 0.81293 0.0062855 0.0070612 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.14018 0.93956 0.91393 0.001397 0.99212 0.57905 0.0018821 0.42961 1.8859 1.8852 16.0034 144.9842 0.0001685 -85.6527 0.75095
2.855 0.98805 5.5074e-005 3.8182 0.012011 3.7471e-005 0.0011557 0.21411 0.00065914 0.21476 0.19767 0 0.033263 0.0389 0 1.0561 0.32163 0.092759 0.012365 5.5088 0.077176 9.482e-005 0.81292 0.0062863 0.007062 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.14019 0.9397 0.91399 0.001397 0.99216 0.57919 0.0018821 0.42962 1.8863 1.8856 16.0034 144.9842 0.0001684 -85.6528 0.75195
2.856 0.98805 5.5074e-005 3.8182 0.012011 3.7484e-005 0.0011557 0.21412 0.00065914 0.21478 0.19769 0 0.033262 0.0389 0 1.0562 0.32168 0.092775 0.012367 5.5099 0.077187 9.4835e-005 0.81291 0.006287 0.0070628 0.001386 0.98695 0.99171 2.9887e-006 1.1954e-005 0.14019 0.93984 0.91405 0.001397 0.99219 0.57934 0.0018821 0.42963 1.8868 1.8861 16.0034 144.9843 0.0001683 -85.6529 0.75295
2.857 0.98805 5.5074e-005 3.8182 0.012011 3.7498e-005 0.0011557 0.21414 0.00065914 0.21479 0.1977 0 0.033261 0.0389 0 1.0563 0.32172 0.092791 0.012369 5.511 0.077198 9.485e-005 0.8129 0.0062877 0.0070635 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.1402 0.93997 0.91411 0.001397 0.99222 0.57949 0.001882 0.42965 1.8872 1.8865 16.0034 144.9843 0.00016821 -85.653 0.75395
2.858 0.98805 5.5073e-005 3.8182 0.012011 3.7511e-005 0.0011557 0.21416 0.00065914 0.21481 0.19772 0 0.03326 0.0389 0 1.0564 0.32177 0.092807 0.01237 5.5121 0.077209 9.4865e-005 0.81289 0.0062884 0.0070643 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.14021 0.94011 0.91418 0.001397 0.99225 0.57963 0.001882 0.42966 1.8876 1.887 16.0033 144.9843 0.00016811 -85.6531 0.75495
2.859 0.98805 5.5073e-005 3.8182 0.012011 3.7524e-005 0.0011557 0.21417 0.00065914 0.21483 0.19773 0 0.033259 0.0389 0 1.0565 0.32181 0.092823 0.012372 5.5132 0.07722 9.488e-005 0.81287 0.0062891 0.007065 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.14021 0.94025 0.91424 0.0013969 0.99228 0.57978 0.001882 0.42967 1.8881 1.8874 16.0033 144.9843 0.00016802 -85.6532 0.75595
2.86 0.98805 5.5073e-005 3.8182 0.012011 3.7537e-005 0.0011557 0.21419 0.00065914 0.21485 0.19775 0 0.033258 0.0389 0 1.0566 0.32186 0.092839 0.012374 5.5143 0.077231 9.4895e-005 0.81286 0.0062898 0.0070658 0.0013859 0.98695 0.99171 2.9884e-006 1.1954e-005 0.14022 0.94038 0.9143 0.0013969 0.99232 0.57992 0.001882 0.42968 1.8885 1.8878 16.0033 144.9843 0.00016792 -85.6534 0.75695
2.861 0.98805 5.5073e-005 3.8182 0.012011 3.755e-005 0.0011557 0.21421 0.00065914 0.21486 0.19777 0 0.033257 0.0389 0 1.0567 0.32191 0.092855 0.012376 5.5154 0.077242 9.491e-005 0.81285 0.0062905 0.0070665 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.14022 0.94052 0.91436 0.0013969 0.99235 0.58007 0.001882 0.42969 1.8889 1.8883 16.0032 144.9844 0.00016783 -85.6535 0.75795
2.862 0.98805 5.5073e-005 3.8182 0.012011 3.7563e-005 0.0011557 0.21422 0.00065914 0.21488 0.19778 0 0.033256 0.0389 0 1.0568 0.32195 0.092871 0.012377 5.5165 0.077254 9.4925e-005 0.81284 0.0062913 0.0070673 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.14023 0.94065 0.91442 0.0013969 0.99238 0.58022 0.001882 0.42971 1.8894 1.8887 16.0032 144.9844 0.00016773 -85.6536 0.75895
2.863 0.98805 5.5073e-005 3.8182 0.012011 3.7576e-005 0.0011557 0.21424 0.00065914 0.2149 0.1978 0 0.033255 0.0389 0 1.0569 0.322 0.092887 0.012379 5.5176 0.077265 9.494e-005 0.81283 0.006292 0.0070681 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.14024 0.94078 0.91448 0.0013969 0.99241 0.58036 0.0018819 0.42972 1.8898 1.8891 16.0032 144.9844 0.00016764 -85.6537 0.75995
2.864 0.98805 5.5073e-005 3.8182 0.012011 3.7589e-005 0.0011557 0.21426 0.00065914 0.21491 0.19781 0 0.033255 0.0389 0 1.057 0.32204 0.092903 0.012381 5.5188 0.077276 9.4954e-005 0.81282 0.0062927 0.0070688 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.14024 0.94092 0.91454 0.0013969 0.99244 0.58051 0.0018819 0.42973 1.8902 1.8896 16.0032 144.9844 0.00016754 -85.6538 0.76095
2.865 0.98805 5.5073e-005 3.8182 0.012011 3.7602e-005 0.0011557 0.21428 0.00065914 0.21493 0.19783 0 0.033254 0.0389 0 1.0571 0.32209 0.092919 0.012383 5.5199 0.077287 9.4969e-005 0.81281 0.0062934 0.0070696 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.14025 0.94105 0.9146 0.0013968 0.99247 0.58065 0.0018819 0.42974 1.8907 1.89 16.0031 144.9844 0.00016745 -85.6539 0.76195
2.866 0.98805 5.5073e-005 3.8182 0.012011 3.7615e-005 0.0011557 0.21429 0.00065914 0.21495 0.19784 0 0.033253 0.0389 0 1.0572 0.32213 0.092935 0.012385 5.521 0.077298 9.4984e-005 0.8128 0.0062941 0.0070703 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.14025 0.94118 0.91466 0.0013968 0.9925 0.5808 0.0018819 0.42976 1.8911 1.8904 16.0031 144.9845 0.00016736 -85.654 0.76295
2.867 0.98805 5.5073e-005 3.8182 0.012011 3.7628e-005 0.0011557 0.21431 0.00065914 0.21496 0.19786 0 0.033252 0.0389 0 1.0573 0.32218 0.092951 0.012386 5.5221 0.077309 9.4999e-005 0.81279 0.0062948 0.0070711 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.14026 0.94132 0.91472 0.0013968 0.99253 0.58095 0.0018819 0.42977 1.8915 1.8909 16.0031 144.9845 0.00016726 -85.6541 0.76395
2.868 0.98805 5.5073e-005 3.8182 0.012011 3.7641e-005 0.0011557 0.21433 0.00065914 0.21498 0.19788 0 0.033251 0.0389 0 1.0574 0.32222 0.092967 0.012388 5.5232 0.07732 9.5014e-005 0.81277 0.0062956 0.0070718 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.14026 0.94145 0.91478 0.0013968 0.99256 0.58109 0.0018818 0.42978 1.892 1.8913 16.003 144.9845 0.00016717 -85.6542 0.76495
2.869 0.98805 5.5073e-005 3.8182 0.012011 3.7654e-005 0.0011557 0.21434 0.00065914 0.215 0.19789 0 0.03325 0.0389 0 1.0575 0.32227 0.092983 0.01239 5.5243 0.077331 9.5029e-005 0.81276 0.0062963 0.0070726 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.14027 0.94158 0.91483 0.0013968 0.99259 0.58124 0.0018818 0.42979 1.8924 1.8917 16.003 144.9845 0.00016708 -85.6543 0.76595
2.87 0.98805 5.5073e-005 3.8182 0.012011 3.7667e-005 0.0011557 0.21436 0.00065914 0.21501 0.19791 0 0.033249 0.0389 0 1.0576 0.32231 0.092999 0.012392 5.5254 0.077342 9.5044e-005 0.81275 0.006297 0.0070734 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.14028 0.94171 0.91489 0.0013968 0.99262 0.58138 0.0018818 0.4298 1.8928 1.8922 16.003 144.9846 0.00016699 -85.6545 0.76695
2.871 0.98805 5.5073e-005 3.8182 0.012011 3.768e-005 0.0011557 0.21438 0.00065914 0.21503 0.19792 0 0.033248 0.0389 0 1.0577 0.32236 0.093015 0.012393 5.5265 0.077353 9.5059e-005 0.81274 0.0062977 0.0070741 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.14028 0.94184 0.91495 0.0013968 0.99265 0.58153 0.0018818 0.42982 1.8932 1.8926 16.003 144.9846 0.00016689 -85.6546 0.76795
2.872 0.98805 5.5073e-005 3.8182 0.012011 3.7693e-005 0.0011557 0.21439 0.00065914 0.21505 0.19794 0 0.033247 0.0389 0 1.0578 0.3224 0.093031 0.012395 5.5276 0.077365 9.5074e-005 0.81273 0.0062984 0.0070749 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.14029 0.94197 0.91501 0.0013967 0.99268 0.58168 0.0018818 0.42983 1.8937 1.893 16.0029 144.9846 0.0001668 -85.6547 0.76895
2.873 0.98805 5.5072e-005 3.8182 0.012011 3.7706e-005 0.0011557 0.21441 0.00065914 0.21506 0.19796 0 0.033247 0.0389 0 1.0579 0.32245 0.093047 0.012397 5.5287 0.077376 9.5089e-005 0.81272 0.0062991 0.0070756 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.14029 0.9421 0.91507 0.0013967 0.99271 0.58182 0.0018818 0.42984 1.8941 1.8934 16.0029 144.9846 0.00016671 -85.6548 0.76995
2.874 0.98805 5.5072e-005 3.8182 0.012011 3.772e-005 0.0011557 0.21443 0.00065914 0.21508 0.19797 0 0.033246 0.0389 0 1.058 0.32249 0.093063 0.012399 5.5298 0.077387 9.5104e-005 0.81271 0.0062998 0.0070764 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.1403 0.94223 0.91513 0.0013967 0.99274 0.58197 0.0018817 0.42985 1.8945 1.8939 16.0029 144.9846 0.00016662 -85.6549 0.77095
2.875 0.98805 5.5072e-005 3.8182 0.012011 3.7733e-005 0.0011557 0.21444 0.00065914 0.2151 0.19799 0 0.033245 0.0389 0 1.0581 0.32254 0.093079 0.012401 5.5309 0.077398 9.5119e-005 0.8127 0.0063006 0.0070771 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.14031 0.94236 0.91518 0.0013967 0.99277 0.58211 0.0018817 0.42986 1.8949 1.8943 16.0028 144.9847 0.00016653 -85.655 0.77195
2.876 0.98805 5.5072e-005 3.8182 0.012011 3.7746e-005 0.0011558 0.21446 0.00065914 0.21511 0.198 0 0.033244 0.0389 0 1.0582 0.32258 0.093095 0.012402 5.532 0.077409 9.5134e-005 0.81269 0.0063013 0.0070779 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.14031 0.94249 0.91524 0.0013967 0.9928 0.58226 0.0018817 0.42988 1.8954 1.8947 16.0028 144.9847 0.00016644 -85.6551 0.77295
2.877 0.98805 5.5072e-005 3.8182 0.01201 3.7759e-005 0.0011558 0.21448 0.00065914 0.21513 0.19802 0 0.033243 0.0389 0 1.0583 0.32263 0.093111 0.012404 5.5331 0.07742 9.5149e-005 0.81268 0.006302 0.0070787 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.14032 0.94262 0.9153 0.0013967 0.99283 0.5824 0.0018817 0.42989 1.8958 1.8951 16.0028 144.9847 0.00016635 -85.6552 0.77395
2.878 0.98805 5.5072e-005 3.8182 0.01201 3.7772e-005 0.0011558 0.21449 0.00065914 0.21515 0.19803 0 0.033242 0.0389 0 1.0584 0.32267 0.093127 0.012406 5.5342 0.077431 9.5164e-005 0.81266 0.0063027 0.0070794 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.14032 0.94275 0.91535 0.0013967 0.99286 0.58255 0.0018817 0.4299 1.8962 1.8956 16.0028 144.9847 0.00016626 -85.6553 0.77495
2.879 0.98805 5.5072e-005 3.8182 0.01201 3.7785e-005 0.0011558 0.21451 0.00065915 0.21516 0.19805 0 0.033241 0.0389 0 1.0585 0.32272 0.093143 0.012408 5.5354 0.077442 9.5178e-005 0.81265 0.0063034 0.0070802 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.14033 0.94287 0.91541 0.0013967 0.99288 0.58269 0.0018817 0.42991 1.8966 1.896 16.0027 144.9847 0.00016617 -85.6554 0.77595
2.88 0.98805 5.5072e-005 3.8182 0.01201 3.7798e-005 0.0011558 0.21453 0.00065915 0.21518 0.19807 0 0.03324 0.0389 0 1.0586 0.32276 0.093159 0.012409 5.5365 0.077453 9.5193e-005 0.81264 0.0063041 0.0070809 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.14033 0.943 0.91547 0.0013967 0.99291 0.58284 0.0018817 0.42993 1.897 1.8964 16.0027 144.9848 0.00016608 -85.6555 0.77695
2.881 0.98805 5.5072e-005 3.8182 0.01201 3.7811e-005 0.0011558 0.21454 0.00065915 0.2152 0.19808 0 0.03324 0.0389 0 1.0587 0.32281 0.093175 0.012411 5.5376 0.077464 9.5208e-005 0.81263 0.0063049 0.0070817 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.14034 0.94313 0.91552 0.0013967 0.99294 0.58298 0.0018816 0.42994 1.8975 1.8968 16.0027 144.9848 0.00016599 -85.6556 0.77795
2.882 0.98805 5.5072e-005 3.8182 0.01201 3.7824e-005 0.0011558 0.21456 0.00065915 0.21521 0.1981 0 0.033239 0.0389 0 1.0588 0.32285 0.093191 0.012413 5.5387 0.077476 9.5223e-005 0.81262 0.0063056 0.0070824 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.14035 0.94325 0.91558 0.0013966 0.99297 0.58313 0.0018816 0.42995 1.8979 1.8973 16.0026 144.9848 0.0001659 -85.6557 0.77895
2.883 0.98805 5.5072e-005 3.8182 0.01201 3.7837e-005 0.0011558 0.21458 0.00065915 0.21523 0.19811 0 0.033238 0.0389 0 1.0589 0.3229 0.093207 0.012415 5.5398 0.077487 9.5238e-005 0.81261 0.0063063 0.0070832 0.0013854 0.98695 0.99171 2.9871e-006 1.1948e-005 0.14035 0.94338 0.91564 0.0013966 0.99299 0.58327 0.0018816 0.42996 1.8983 1.8977 16.0026 144.9848 0.00016582 -85.6558 0.77995
2.884 0.98805 5.5072e-005 3.8182 0.01201 3.785e-005 0.0011558 0.21459 0.00065915 0.21525 0.19813 0 0.033237 0.0389 0 1.059 0.32294 0.093223 0.012417 5.5409 0.077498 9.5253e-005 0.8126 0.006307 0.007084 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.14036 0.9435 0.91569 0.0013966 0.99302 0.58342 0.0018816 0.42997 1.8987 1.8981 16.0026 144.9848 0.00016573 -85.6559 0.78095
2.885 0.98805 5.5072e-005 3.8182 0.01201 3.7863e-005 0.0011558 0.21461 0.00065915 0.21526 0.19814 0 0.033236 0.0389 0 1.0591 0.32299 0.093239 0.012418 5.542 0.077509 9.5268e-005 0.81259 0.0063077 0.0070847 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.14036 0.94363 0.91575 0.0013966 0.99305 0.58356 0.0018816 0.42999 1.8991 1.8985 16.0026 144.9849 0.00016564 -85.656 0.78195
2.886 0.98805 5.5072e-005 3.8182 0.01201 3.7876e-005 0.0011558 0.21463 0.00065915 0.21528 0.19816 0 0.033235 0.0389 0 1.0592 0.32304 0.093255 0.01242 5.5431 0.07752 9.5283e-005 0.81258 0.0063084 0.0070855 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.14037 0.94375 0.9158 0.0013966 0.99308 0.58371 0.0018816 0.43 1.8995 1.8989 16.0025 144.9849 0.00016555 -85.6561 0.78295
2.887 0.98805 5.5072e-005 3.8182 0.01201 3.7889e-005 0.0011558 0.21464 0.00065915 0.2153 0.19818 0 0.033234 0.0389 0 1.0593 0.32308 0.093271 0.012422 5.5442 0.077531 9.5298e-005 0.81256 0.0063092 0.0070862 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.14038 0.94388 0.91586 0.0013966 0.9931 0.58385 0.0018815 0.43001 1.9 1.8993 16.0025 144.9849 0.00016547 -85.6562 0.78395
2.888 0.98805 5.5071e-005 3.8182 0.01201 3.7902e-005 0.0011558 0.21466 0.00065915 0.21531 0.19819 0 0.033233 0.0389 0 1.0594 0.32313 0.093287 0.012424 5.5454 0.077542 9.5313e-005 0.81255 0.0063099 0.007087 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.14038 0.944 0.91591 0.0013966 0.99313 0.584 0.0018815 0.43002 1.9004 1.8997 16.0025 144.9849 0.00016538 -85.6562 0.78495
2.889 0.98805 5.5071e-005 3.8182 0.01201 3.7915e-005 0.0011558 0.21467 0.00065915 0.21533 0.19821 0 0.033233 0.0389 0 1.0595 0.32317 0.093303 0.012425 5.5465 0.077553 9.5328e-005 0.81254 0.0063106 0.0070878 0.0013853 0.98696 0.99171 2.9868e-006 1.1947e-005 0.14039 0.94413 0.91597 0.0013965 0.99315 0.58414 0.0018815 0.43003 1.9008 1.9002 16.0024 144.9849 0.00016529 -85.6563 0.78595
2.89 0.98805 5.5071e-005 3.8182 0.01201 3.7929e-005 0.0011558 0.21469 0.00065915 0.21535 0.19822 0 0.033232 0.0389 0 1.0596 0.32322 0.093319 0.012427 5.5476 0.077564 9.5343e-005 0.81253 0.0063113 0.0070885 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.14039 0.94425 0.91602 0.0013965 0.99318 0.58429 0.0018815 0.43005 1.9012 1.9006 16.0024 144.985 0.00016521 -85.6564 0.78695
2.891 0.98805 5.5071e-005 3.8182 0.01201 3.7942e-005 0.0011558 0.21471 0.00065915 0.21536 0.19824 0 0.033231 0.0389 0 1.0597 0.32326 0.093335 0.012429 5.5487 0.077575 9.5358e-005 0.81252 0.006312 0.0070893 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.1404 0.94437 0.91608 0.0013965 0.99321 0.58443 0.0018815 0.43006 1.9016 1.901 16.0024 144.985 0.00016512 -85.6565 0.78795
2.892 0.98805 5.5071e-005 3.8182 0.01201 3.7955e-005 0.0011558 0.21472 0.00065915 0.21538 0.19825 0 0.03323 0.0389 0 1.0598 0.32331 0.093351 0.012431 5.5498 0.077586 9.5373e-005 0.81251 0.0063127 0.00709 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.1404 0.94449 0.91613 0.0013965 0.99323 0.58458 0.0018815 0.43007 1.902 1.9014 16.0024 144.985 0.00016504 -85.6566 0.78895
2.893 0.98805 5.5071e-005 3.8182 0.01201 3.7968e-005 0.0011558 0.21474 0.00065915 0.2154 0.19827 0 0.033229 0.0389 0 1.0599 0.32335 0.093367 0.012432 5.5509 0.077598 9.5388e-005 0.8125 0.0063135 0.0070908 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.14041 0.94462 0.91619 0.0013965 0.99326 0.58472 0.0018815 0.43008 1.9024 1.9018 16.0023 144.985 0.00016495 -85.6567 0.78995
2.894 0.98805 5.5071e-005 3.8182 0.01201 3.7981e-005 0.0011558 0.21476 0.00065915 0.21541 0.19829 0 0.033228 0.0389 0 1.06 0.3234 0.093383 0.012434 5.552 0.077609 9.5402e-005 0.81249 0.0063142 0.0070915 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.14042 0.94474 0.91624 0.0013965 0.99328 0.58487 0.0018814 0.43009 1.9028 1.9022 16.0023 144.985 0.00016487 -85.6568 0.79095
2.895 0.98805 5.5071e-005 3.8182 0.01201 3.7994e-005 0.0011558 0.21477 0.00065915 0.21543 0.1983 0 0.033227 0.0389 0 1.0601 0.32344 0.093399 0.012436 5.5532 0.07762 9.5417e-005 0.81248 0.0063149 0.0070923 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.14042 0.94486 0.9163 0.0013965 0.99331 0.58501 0.0018814 0.43011 1.9032 1.9026 16.0023 144.9851 0.00016478 -85.6569 0.79195
2.896 0.98805 5.5071e-005 3.8182 0.01201 3.8007e-005 0.0011558 0.21479 0.00065915 0.21544 0.19832 0 0.033227 0.0389 0 1.0602 0.32349 0.093415 0.012438 5.5543 0.077631 9.5432e-005 0.81246 0.0063156 0.0070931 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.14043 0.94498 0.91635 0.0013965 0.99333 0.58516 0.0018814 0.43012 1.9037 1.903 16.0022 144.9851 0.0001647 -85.657 0.79295
2.897 0.98805 5.5071e-005 3.8182 0.01201 3.802e-005 0.0011558 0.21481 0.00065915 0.21546 0.19833 0 0.033226 0.0389 0 1.0603 0.32353 0.093431 0.01244 5.5554 0.077642 9.5447e-005 0.81245 0.0063163 0.0070938 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.14043 0.9451 0.9164 0.0013964 0.99336 0.5853 0.0018814 0.43013 1.9041 1.9034 16.0022 144.9851 0.00016461 -85.6571 0.79395
2.898 0.98805 5.5071e-005 3.8182 0.01201 3.8033e-005 0.0011558 0.21482 0.00065915 0.21548 0.19835 0 0.033225 0.0389 0 1.0604 0.32358 0.093447 0.012441 5.5565 0.077653 9.5462e-005 0.81244 0.006317 0.0070946 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.14044 0.94522 0.91646 0.0013964 0.99338 0.58544 0.0018814 0.43014 1.9045 1.9038 16.0022 144.9851 0.00016453 -85.6571 0.79495
2.899 0.98805 5.5071e-005 3.8182 0.01201 3.8046e-005 0.0011558 0.21484 0.00065915 0.21549 0.19836 0 0.033224 0.0389 0 1.0605 0.32362 0.093463 0.012443 5.5576 0.077664 9.5477e-005 0.81243 0.0063178 0.0070953 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.14045 0.94534 0.91651 0.0013964 0.99341 0.58559 0.0018814 0.43015 1.9049 1.9043 16.0021 144.9851 0.00016445 -85.6572 0.79595
2.9 0.98805 5.5071e-005 3.8182 0.01201 3.8059e-005 0.0011558 0.21486 0.00065915 0.21551 0.19838 0 0.033223 0.0389 0 1.0606 0.32367 0.093479 0.012445 5.5588 0.077675 9.5492e-005 0.81242 0.0063185 0.0070961 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.14045 0.94546 0.91656 0.0013964 0.99343 0.58573 0.0018814 0.43017 1.9053 1.9047 16.0021 144.9852 0.00016436 -85.6573 0.79695
2.901 0.98805 5.5071e-005 3.8182 0.01201 3.8072e-005 0.0011558 0.21487 0.00065915 0.21553 0.19839 0 0.033222 0.0389 0 1.0607 0.32371 0.093495 0.012447 5.5599 0.077686 9.5507e-005 0.81241 0.0063192 0.0070969 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.14046 0.94558 0.91661 0.0013964 0.99346 0.58588 0.0018813 0.43018 1.9057 1.9051 16.0021 144.9852 0.00016428 -85.6574 0.79795
2.902 0.98805 5.507e-005 3.8182 0.01201 3.8085e-005 0.0011558 0.21489 0.00065915 0.21554 0.19841 0 0.033221 0.0389 0 1.0608 0.32376 0.093511 0.012448 5.561 0.077697 9.5522e-005 0.8124 0.0063199 0.0070976 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.14046 0.9457 0.91667 0.0013964 0.99348 0.58602 0.0018813 0.43019 1.9061 1.9055 16.0021 144.9852 0.0001642 -85.6575 0.79895
2.903 0.98805 5.507e-005 3.8182 0.01201 3.8098e-005 0.0011558 0.2149 0.00065915 0.21556 0.19843 0 0.033221 0.0389 0 1.0609 0.3238 0.093527 0.01245 5.5621 0.077708 9.5537e-005 0.81239 0.0063206 0.0070984 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.14047 0.94582 0.91672 0.0013964 0.99351 0.58617 0.0018813 0.4302 1.9065 1.9059 16.002 144.9852 0.00016412 -85.6576 0.79995
2.904 0.98805 5.507e-005 3.8182 0.01201 3.8111e-005 0.0011558 0.21492 0.00065915 0.21558 0.19844 0 0.03322 0.0389 0 1.061 0.32385 0.093543 0.012452 5.5632 0.07772 9.5552e-005 0.81238 0.0063214 0.0070991 0.001385 0.98696 0.99171 2.9861e-006 1.1944e-005 0.14047 0.94593 0.91677 0.0013964 0.99353 0.58631 0.0018813 0.43021 1.9069 1.9063 16.002 144.9852 0.00016403 -85.6577 0.80095
2.905 0.98805 5.507e-005 3.8182 0.01201 3.8124e-005 0.0011558 0.21494 0.00065915 0.21559 0.19846 0 0.033219 0.0389 0 1.0611 0.3239 0.093559 0.012454 5.5644 0.077731 9.5567e-005 0.81236 0.0063221 0.0070999 0.0013849 0.98696 0.99171 2.9861e-006 1.1944e-005 0.14048 0.94605 0.91682 0.0013964 0.99355 0.58645 0.0018813 0.43023 1.9073 1.9067 16.002 144.9853 0.00016395 -85.6577 0.80195
2.906 0.98805 5.507e-005 3.8182 0.01201 3.8137e-005 0.0011558 0.21495 0.00065915 0.21561 0.19847 0 0.033218 0.0389 0 1.0612 0.32394 0.093575 0.012456 5.5655 0.077742 9.5582e-005 0.81235 0.0063228 0.0071007 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.14049 0.94617 0.91688 0.0013964 0.99358 0.5866 0.0018813 0.43024 1.9077 1.9071 16.0019 144.9853 0.00016387 -85.6578 0.80295
2.907 0.98805 5.507e-005 3.8182 0.01201 3.8151e-005 0.0011558 0.21497 0.00065915 0.21562 0.19849 0 0.033217 0.0389 0 1.0613 0.32399 0.093591 0.012457 5.5666 0.077753 9.5597e-005 0.81234 0.0063235 0.0071014 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.14049 0.94629 0.91693 0.0013963 0.9936 0.58674 0.0018813 0.43025 1.9081 1.9075 16.0019 144.9853 0.00016379 -85.6579 0.80395
2.908 0.98805 5.507e-005 3.8182 0.01201 3.8164e-005 0.0011558 0.21499 0.00065915 0.21564 0.1985 0 0.033216 0.0389 0 1.0614 0.32403 0.093608 0.012459 5.5677 0.077764 9.5611e-005 0.81233 0.0063242 0.0071022 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.1405 0.9464 0.91698 0.0013963 0.99362 0.58689 0.0018813 0.43026 1.9085 1.9079 16.0019 144.9853 0.00016371 -85.658 0.80495
2.909 0.98805 5.507e-005 3.8182 0.01201 3.8177e-005 0.0011558 0.215 0.00065915 0.21566 0.19852 0 0.033215 0.0389 0 1.0614 0.32408 0.093624 0.012461 5.5688 0.077775 9.5626e-005 0.81232 0.0063249 0.0071029 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.1405 0.94652 0.91703 0.0013963 0.99365 0.58703 0.0018812 0.43027 1.9089 1.9083 16.0019 144.9854 0.00016363 -85.6581 0.80595
2.91 0.98805 5.507e-005 3.8182 0.01201 3.819e-005 0.0011558 0.21502 0.00065915 0.21567 0.19853 0 0.033215 0.0389 0 1.0615 0.32412 0.09364 0.012463 5.57 0.077786 9.5641e-005 0.81231 0.0063257 0.0071037 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.14051 0.94663 0.91708 0.0013963 0.99367 0.58717 0.0018812 0.43029 1.9093 1.9087 16.0018 144.9854 0.00016355 -85.6581 0.80695
2.911 0.98805 5.507e-005 3.8182 0.01201 3.8203e-005 0.0011558 0.21503 0.00065915 0.21569 0.19855 0 0.033214 0.0389 0 1.0616 0.32417 0.093656 0.012464 5.5711 0.077797 9.5656e-005 0.8123 0.0063264 0.0071045 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.14052 0.94675 0.91713 0.0013963 0.99369 0.58732 0.0018812 0.4303 1.9097 1.9091 16.0018 144.9854 0.00016347 -85.6582 0.80795
2.912 0.98805 5.507e-005 3.8182 0.01201 3.8216e-005 0.0011558 0.21505 0.00065915 0.21571 0.19856 0 0.033213 0.0389 0 1.0617 0.32421 0.093672 0.012466 5.5722 0.077808 9.5671e-005 0.81229 0.0063271 0.0071052 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.14052 0.94686 0.91718 0.0013963 0.99372 0.58746 0.0018812 0.43031 1.9101 1.9095 16.0018 144.9854 0.00016339 -85.6583 0.80895
2.913 0.98805 5.507e-005 3.8182 0.01201 3.8229e-005 0.0011558 0.21507 0.00065915 0.21572 0.19858 0 0.033212 0.0389 0 1.0618 0.32426 0.093688 0.012468 5.5733 0.077819 9.5686e-005 0.81228 0.0063278 0.007106 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.14053 0.94698 0.91723 0.0013963 0.99374 0.5876 0.0018812 0.43032 1.9105 1.9099 16.0017 144.9854 0.00016331 -85.6584 0.80995
2.914 0.98805 5.507e-005 3.8182 0.01201 3.8242e-005 0.0011558 0.21508 0.00065915 0.21574 0.19859 0 0.033211 0.0389 0 1.0619 0.3243 0.093704 0.01247 5.5745 0.07783 9.5701e-005 0.81227 0.0063285 0.0071067 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.14053 0.94709 0.91728 0.0013963 0.99376 0.58775 0.0018812 0.43033 1.9108 1.9103 16.0017 144.9855 0.00016323 -85.6585 0.81095
2.915 0.98805 5.507e-005 3.8182 0.01201 3.8255e-005 0.0011558 0.2151 0.00065915 0.21575 0.19861 0 0.03321 0.0389 0 1.062 0.32435 0.09372 0.012472 5.5756 0.077841 9.5716e-005 0.81225 0.0063292 0.0071075 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.14054 0.94721 0.91734 0.0013963 0.99378 0.58789 0.0018812 0.43035 1.9112 1.9106 16.0017 144.9855 0.00016315 -85.6585 0.81195
2.916 0.98805 5.507e-005 3.8182 0.01201 3.8268e-005 0.0011558 0.21512 0.00065915 0.21577 0.19862 0 0.033209 0.0389 0 1.0621 0.32439 0.093736 0.012473 5.5767 0.077853 9.5731e-005 0.81224 0.00633 0.0071083 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.14055 0.94732 0.91739 0.0013963 0.9938 0.58803 0.0018811 0.43036 1.9116 1.911 16.0016 144.9855 0.00016307 -85.6586 0.81295
2.917 0.98805 5.5069e-005 3.8182 0.01201 3.8281e-005 0.0011558 0.21513 0.00065915 0.21579 0.19864 0 0.033209 0.0389 0 1.0622 0.32444 0.093752 0.012475 5.5778 0.077864 9.5746e-005 0.81223 0.0063307 0.007109 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.14055 0.94743 0.91744 0.0013963 0.99383 0.58818 0.0018811 0.43037 1.912 1.9114 16.0016 144.9855 0.00016299 -85.6587 0.81395
2.918 0.98805 5.5069e-005 3.8182 0.01201 3.8294e-005 0.0011558 0.21515 0.00065915 0.2158 0.19866 0 0.033208 0.0389 0 1.0623 0.32448 0.093768 0.012477 5.579 0.077875 9.5761e-005 0.81222 0.0063314 0.0071098 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.14056 0.94755 0.91749 0.0013962 0.99385 0.58832 0.0018811 0.43038 1.9124 1.9118 16.0016 144.9855 0.00016291 -85.6588 0.81495
2.919 0.98805 5.5069e-005 3.8182 0.01201 3.8307e-005 0.0011558 0.21516 0.00065915 0.21582 0.19867 0 0.033207 0.0389 0 1.0624 0.32453 0.093784 0.012479 5.5801 0.077886 9.5776e-005 0.81221 0.0063321 0.0071105 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.14056 0.94766 0.91753 0.0013962 0.99387 0.58846 0.0018811 0.43039 1.9128 1.9122 16.0016 144.9856 0.00016283 -85.6588 0.81595
2.92 0.98805 5.5069e-005 3.8182 0.01201 3.832e-005 0.0011558 0.21518 0.00065915 0.21583 0.19869 0 0.033206 0.0389 0 1.0625 0.32457 0.0938 0.01248 5.5812 0.077897 9.5791e-005 0.8122 0.0063328 0.0071113 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.14057 0.94777 0.91758 0.0013962 0.99389 0.58861 0.0018811 0.43041 1.9132 1.9126 16.0015 144.9856 0.00016276 -85.6589 0.81695
2.921 0.98805 5.5069e-005 3.8182 0.01201 3.8333e-005 0.0011558 0.2152 0.00065915 0.21585 0.1987 0 0.033205 0.0389 0 1.0626 0.32462 0.093816 0.012482 5.5823 0.077908 9.5806e-005 0.81219 0.0063336 0.0071121 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.14057 0.94788 0.91763 0.0013962 0.99391 0.58875 0.0018811 0.43042 1.9136 1.913 16.0015 144.9856 0.00016268 -85.659 0.81795
2.922 0.98805 5.5069e-005 3.8182 0.01201 3.8346e-005 0.0011558 0.21521 0.00065915 0.21587 0.19872 0 0.033204 0.0389 0 1.0627 0.32467 0.093832 0.012484 5.5835 0.077919 9.582e-005 0.81218 0.0063343 0.0071128 0.0013846 0.98696 0.99172 2.9854e-006 1.1941e-005 0.14058 0.94799 0.91768 0.0013962 0.99393 0.58889 0.0018811 0.43043 1.914 1.9134 16.0015 144.9856 0.0001626 -85.6591 0.81895
2.923 0.98805 5.5069e-005 3.8182 0.01201 3.8359e-005 0.0011558 0.21523 0.00065915 0.21588 0.19873 0 0.033204 0.0389 0 1.0628 0.32471 0.093848 0.012486 5.5846 0.07793 9.5835e-005 0.81217 0.006335 0.0071136 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.14059 0.94811 0.91773 0.0013962 0.99395 0.58904 0.0018811 0.43044 1.9144 1.9138 16.0014 144.9856 0.00016252 -85.6591 0.81995
2.924 0.98805 5.5069e-005 3.8182 0.01201 3.8373e-005 0.0011558 0.21524 0.00065915 0.2159 0.19875 0 0.033203 0.0389 0 1.0629 0.32476 0.093864 0.012487 5.5857 0.077941 9.585e-005 0.81215 0.0063357 0.0071143 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.14059 0.94822 0.91778 0.0013962 0.99398 0.58918 0.0018811 0.43045 1.9147 1.9142 16.0014 144.9857 0.00016245 -85.6592 0.82095
2.925 0.98805 5.5069e-005 3.8182 0.01201 3.8386e-005 0.0011558 0.21526 0.00065915 0.21591 0.19876 0 0.033202 0.0389 0 1.063 0.3248 0.09388 0.012489 5.5868 0.077952 9.5865e-005 0.81214 0.0063364 0.0071151 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.1406 0.94833 0.91783 0.0013962 0.994 0.58932 0.001881 0.43047 1.9151 1.9145 16.0014 144.9857 0.00016237 -85.6593 0.82195
2.926 0.98805 5.5069e-005 3.8182 0.01201 3.8399e-005 0.0011558 0.21528 0.00065915 0.21593 0.19878 0 0.033201 0.0389 0 1.0631 0.32485 0.093896 0.012491 5.588 0.077963 9.588e-005 0.81213 0.0063371 0.0071159 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1406 0.94844 0.91788 0.0013962 0.99402 0.58947 0.001881 0.43048 1.9155 1.9149 16.0013 144.9857 0.0001623 -85.6594 0.82295
2.927 0.98805 5.5069e-005 3.8182 0.01201 3.8412e-005 0.0011558 0.21529 0.00065915 0.21595 0.19879 0 0.0332 0.0389 0 1.0632 0.32489 0.093912 0.012493 5.5891 0.077974 9.5895e-005 0.81212 0.0063379 0.0071166 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.14061 0.94855 0.91793 0.0013962 0.99404 0.58961 0.001881 0.43049 1.9159 1.9153 16.0013 144.9857 0.00016222 -85.6594 0.82395
2.928 0.98805 5.5069e-005 3.8182 0.01201 3.8425e-005 0.0011558 0.21531 0.00065915 0.21596 0.19881 0 0.033199 0.0389 0 1.0633 0.32494 0.093928 0.012495 5.5902 0.077985 9.591e-005 0.81211 0.0063386 0.0071174 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.14062 0.94866 0.91797 0.0013962 0.99406 0.58975 0.001881 0.4305 1.9163 1.9157 16.0013 144.9857 0.00016214 -85.6595 0.82495
2.929 0.98805 5.5069e-005 3.8182 0.01201 3.8438e-005 0.0011558 0.21532 0.00065915 0.21598 0.19882 0 0.033198 0.0389 0 1.0634 0.32498 0.093944 0.012496 5.5914 0.077997 9.5925e-005 0.8121 0.0063393 0.0071181 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.14062 0.94876 0.91802 0.0013962 0.99408 0.58989 0.001881 0.43051 1.9167 1.9161 16.0013 144.9858 0.00016207 -85.6596 0.82595
2.93 0.98805 5.5069e-005 3.8182 0.01201 3.8451e-005 0.0011558 0.21534 0.00065915 0.21599 0.19884 0 0.033198 0.0389 0 1.0635 0.32503 0.09396 0.012498 5.5925 0.078008 9.594e-005 0.81209 0.00634 0.0071189 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.14063 0.94887 0.91807 0.0013962 0.9941 0.59004 0.001881 0.43052 1.917 1.9165 16.0012 144.9858 0.00016199 -85.6596 0.82695
2.931 0.98805 5.5069e-005 3.8182 0.01201 3.8464e-005 0.0011558 0.21536 0.00065915 0.21601 0.19885 0 0.033197 0.0389 0 1.0636 0.32507 0.093976 0.0125 5.5936 0.078019 9.5955e-005 0.81208 0.0063407 0.0071197 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.14063 0.94898 0.91812 0.0013961 0.99412 0.59018 0.001881 0.43054 1.9174 1.9169 16.0012 144.9858 0.00016192 -85.6597 0.82795
2.932 0.98805 5.5068e-005 3.8182 0.01201 3.8477e-005 0.0011558 0.21537 0.00065915 0.21603 0.19887 0 0.033196 0.0389 0 1.0637 0.32512 0.093992 0.012502 5.5948 0.07803 9.597e-005 0.81207 0.0063415 0.0071204 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.14064 0.94909 0.91817 0.0013961 0.99414 0.59032 0.001881 0.43055 1.9178 1.9172 16.0012 144.9858 0.00016184 -85.6598 0.82895
2.933 0.98805 5.5068e-005 3.8182 0.01201 3.849e-005 0.0011558 0.21539 0.00065915 0.21604 0.19888 0 0.033195 0.0389 0 1.0638 0.32516 0.094008 0.012503 5.5959 0.078041 9.5985e-005 0.81206 0.0063422 0.0071212 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.14064 0.9492 0.91821 0.0013961 0.99416 0.59047 0.001881 0.43056 1.9182 1.9176 16.0011 144.9858 0.00016177 -85.6598 0.82995
2.934 0.98805 5.5068e-005 3.8182 0.01201 3.8503e-005 0.0011558 0.2154 0.00065915 0.21606 0.1989 0 0.033194 0.0389 0 1.0639 0.32521 0.094024 0.012505 5.597 0.078052 9.6e-005 0.81204 0.0063429 0.0071219 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.14065 0.9493 0.91826 0.0013961 0.99418 0.59061 0.0018809 0.43057 1.9186 1.918 16.0011 144.9859 0.00016169 -85.6599 0.83095
2.935 0.98805 5.5068e-005 3.8182 0.01201 3.8516e-005 0.0011558 0.21542 0.00065915 0.21607 0.19891 0 0.033193 0.0389 0 1.064 0.32525 0.09404 0.012507 5.5981 0.078063 9.6014e-005 0.81203 0.0063436 0.0071227 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.14066 0.94941 0.91831 0.0013961 0.9942 0.59075 0.0018809 0.43058 1.9189 1.9184 16.0011 144.9859 0.00016162 -85.66 0.83195
2.936 0.98805 5.5068e-005 3.8182 0.01201 3.8529e-005 0.0011558 0.21544 0.00065915 0.21609 0.19893 0 0.033193 0.0389 0 1.0641 0.3253 0.094056 0.012509 5.5993 0.078074 9.6029e-005 0.81202 0.0063443 0.0071235 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.14066 0.94952 0.91835 0.0013961 0.99422 0.59089 0.0018809 0.4306 1.9193 1.9188 16.001 144.9859 0.00016155 -85.66 0.83295
2.937 0.98805 5.5068e-005 3.8182 0.01201 3.8542e-005 0.0011558 0.21545 0.00065915 0.21611 0.19894 0 0.033192 0.0389 0 1.0642 0.32535 0.094072 0.012511 5.6004 0.078085 9.6044e-005 0.81201 0.006345 0.0071242 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.14067 0.94962 0.9184 0.0013961 0.99424 0.59104 0.0018809 0.43061 1.9197 1.9191 16.001 144.9859 0.00016147 -85.6601 0.83395
2.938 0.98805 5.5068e-005 3.8182 0.01201 3.8555e-005 0.0011558 0.21547 0.00065915 0.21612 0.19896 0 0.033191 0.0389 0 1.0643 0.32539 0.094088 0.012512 5.6015 0.078096 9.6059e-005 0.812 0.0063458 0.007125 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.14067 0.94973 0.91845 0.0013961 0.99426 0.59118 0.0018809 0.43062 1.9201 1.9195 16.001 144.9859 0.0001614 -85.6602 0.83495
2.939 0.98805 5.5068e-005 3.8182 0.01201 3.8568e-005 0.0011558 0.21548 0.00065915 0.21614 0.19897 0 0.03319 0.0389 0 1.0644 0.32544 0.094105 0.012514 5.6027 0.078107 9.6074e-005 0.81199 0.0063465 0.0071258 0.0013843 0.98697 0.99172 2.9848e-006 1.1939e-005 0.14068 0.94984 0.91849 0.0013961 0.99427 0.59132 0.0018809 0.43063 1.9204 1.9199 16.0009 144.986 0.00016133 -85.6602 0.83595
2.94 0.98805 5.5068e-005 3.8182 0.01201 3.8581e-005 0.0011558 0.2155 0.00065915 0.21615 0.19899 0 0.033189 0.0389 0 1.0645 0.32548 0.094121 0.012516 5.6038 0.078118 9.6089e-005 0.81198 0.0063472 0.0071265 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.14069 0.94994 0.91854 0.0013961 0.99429 0.59146 0.0018809 0.43064 1.9208 1.9203 16.0009 144.986 0.00016125 -85.6603 0.83695
2.941 0.98805 5.5068e-005 3.8182 0.01201 3.8595e-005 0.0011558 0.21551 0.00065915 0.21617 0.199 0 0.033188 0.0389 0 1.0646 0.32553 0.094137 0.012518 5.605 0.078129 9.6104e-005 0.81197 0.0063479 0.0071273 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.14069 0.95005 0.91859 0.0013961 0.99431 0.5916 0.0018809 0.43065 1.9212 1.9206 16.0009 144.986 0.00016118 -85.6604 0.83795
2.942 0.98805 5.5068e-005 3.8182 0.01201 3.8608e-005 0.0011559 0.21553 0.00065915 0.21618 0.19902 0 0.033188 0.0389 0 1.0647 0.32557 0.094153 0.012519 5.6061 0.07814 9.6119e-005 0.81196 0.0063486 0.007128 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.1407 0.95015 0.91863 0.001396 0.99433 0.59175 0.0018809 0.43067 1.9216 1.921 16.0009 144.986 0.00016111 -85.6604 0.83895
2.943 0.98805 5.5068e-005 3.8182 0.01201 3.8621e-005 0.0011559 0.21555 0.00065915 0.2162 0.19903 0 0.033187 0.0389 0 1.0648 0.32562 0.094169 0.012521 5.6072 0.078152 9.6134e-005 0.81194 0.0063494 0.0071288 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.1407 0.95026 0.91868 0.001396 0.99435 0.59189 0.0018808 0.43068 1.9219 1.9214 16.0008 144.986 0.00016104 -85.6605 0.83995
2.944 0.98805 5.5068e-005 3.8182 0.01201 3.8634e-005 0.0011559 0.21556 0.00065915 0.21622 0.19905 0 0.033186 0.0389 0 1.0649 0.32566 0.094185 0.012523 5.6084 0.078163 9.6149e-005 0.81193 0.0063501 0.0071296 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.14071 0.95036 0.91872 0.001396 0.99437 0.59203 0.0018808 0.43069 1.9223 1.9218 16.0008 144.9861 0.00016096 -85.6606 0.84095
2.945 0.98805 5.5068e-005 3.8182 0.012009 3.8647e-005 0.0011559 0.21558 0.00065916 0.21623 0.19906 0 0.033185 0.0389 0 1.065 0.32571 0.094201 0.012525 5.6095 0.078174 9.6164e-005 0.81192 0.0063508 0.0071303 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.14071 0.95046 0.91877 0.001396 0.99439 0.59217 0.0018808 0.4307 1.9227 1.9221 16.0008 144.9861 0.00016089 -85.6606 0.84195
2.946 0.98805 5.5068e-005 3.8182 0.012009 3.866e-005 0.0011559 0.21559 0.00065916 0.21625 0.19908 0 0.033184 0.0389 0 1.0651 0.32575 0.094217 0.012526 5.6106 0.078185 9.6179e-005 0.81191 0.0063515 0.0071311 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14072 0.95057 0.91881 0.001396 0.9944 0.59231 0.0018808 0.43071 1.9231 1.9225 16.0007 144.9861 0.00016082 -85.6607 0.84295
2.947 0.98805 5.5067e-005 3.8182 0.012009 3.8673e-005 0.0011559 0.21561 0.00065916 0.21626 0.19909 0 0.033184 0.0389 0 1.0652 0.3258 0.094233 0.012528 5.6118 0.078196 9.6194e-005 0.8119 0.0063522 0.0071318 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14073 0.95067 0.91886 0.001396 0.99442 0.59246 0.0018808 0.43073 1.9234 1.9229 16.0007 144.9861 0.00016075 -85.6607 0.84395
2.948 0.98805 5.5067e-005 3.8182 0.012009 3.8686e-005 0.0011559 0.21562 0.00065916 0.21628 0.19911 0 0.033183 0.0389 0 1.0653 0.32584 0.094249 0.01253 5.6129 0.078207 9.6208e-005 0.81189 0.006353 0.0071326 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14073 0.95077 0.9189 0.001396 0.99444 0.5926 0.0018808 0.43074 1.9238 1.9232 16.0007 144.9862 0.00016068 -85.6608 0.84495
2.949 0.98805 5.5067e-005 3.8182 0.012009 3.8699e-005 0.0011559 0.21564 0.00065916 0.2163 0.19912 0 0.033182 0.0389 0 1.0654 0.32589 0.094265 0.012532 5.614 0.078218 9.6223e-005 0.81188 0.0063537 0.0071334 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.14074 0.95088 0.91895 0.001396 0.99446 0.59274 0.0018808 0.43075 1.9242 1.9236 16.0006 144.9862 0.00016061 -85.6609 0.84595
2.95 0.98805 5.5067e-005 3.8182 0.012009 3.8712e-005 0.0011559 0.21566 0.00065916 0.21631 0.19914 0 0.033181 0.0389 0 1.0655 0.32594 0.094281 0.012534 5.6152 0.078229 9.6238e-005 0.81187 0.0063544 0.0071341 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.14074 0.95098 0.91899 0.001396 0.99448 0.59288 0.0018808 0.43076 1.9245 1.924 16.0006 144.9862 0.00016054 -85.6609 0.84695
2.951 0.98805 5.5067e-005 3.8182 0.012009 3.8725e-005 0.0011559 0.21567 0.00065916 0.21633 0.19915 0 0.03318 0.0389 0 1.0656 0.32598 0.094297 0.012535 5.6163 0.07824 9.6253e-005 0.81186 0.0063551 0.0071349 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.14075 0.95108 0.91904 0.001396 0.99449 0.59302 0.0018808 0.43077 1.9249 1.9244 16.0006 144.9862 0.00016047 -85.661 0.84795
2.952 0.98805 5.5067e-005 3.8182 0.012009 3.8738e-005 0.0011559 0.21569 0.00065916 0.21634 0.19917 0 0.033179 0.0389 0 1.0657 0.32603 0.094313 0.012537 5.6175 0.078251 9.6268e-005 0.81185 0.0063558 0.0071357 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.14076 0.95118 0.91908 0.001396 0.99451 0.59317 0.0018808 0.43078 1.9253 1.9247 16.0005 144.9862 0.0001604 -85.661 0.84895
2.953 0.98805 5.5067e-005 3.8182 0.012009 3.8751e-005 0.0011559 0.2157 0.00065916 0.21636 0.19918 0 0.033179 0.0389 0 1.0658 0.32607 0.094329 0.012539 5.6186 0.078262 9.6283e-005 0.81183 0.0063566 0.0071364 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.14076 0.95128 0.91913 0.001396 0.99453 0.59331 0.0018808 0.4308 1.9256 1.9251 16.0005 144.9863 0.00016033 -85.6611 0.84995
2.954 0.98805 5.5067e-005 3.8182 0.012009 3.8764e-005 0.0011559 0.21572 0.00065916 0.21637 0.1992 0 0.033178 0.0389 0 1.0659 0.32612 0.094345 0.012541 5.6197 0.078273 9.6298e-005 0.81182 0.0063573 0.0071372 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.14077 0.95138 0.91917 0.001396 0.99454 0.59345 0.0018807 0.43081 1.926 1.9255 16.0005 144.9863 0.00016026 -85.6612 0.85095
2.955 0.98805 5.5067e-005 3.8182 0.012009 3.8777e-005 0.0011559 0.21573 0.00065916 0.21639 0.19921 0 0.033177 0.0389 0 1.066 0.32616 0.094361 0.012542 5.6209 0.078284 9.6313e-005 0.81181 0.006358 0.0071379 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.14077 0.95148 0.91922 0.001396 0.99456 0.59359 0.0018807 0.43082 1.9264 1.9258 16.0005 144.9863 0.00016019 -85.6612 0.85195
2.956 0.98805 5.5067e-005 3.8182 0.012009 3.879e-005 0.0011559 0.21575 0.00065916 0.2164 0.19923 0 0.033176 0.0389 0 1.0661 0.32621 0.094377 0.012544 5.622 0.078295 9.6328e-005 0.8118 0.0063587 0.0071387 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14078 0.95158 0.91926 0.001396 0.99458 0.59373 0.0018807 0.43083 1.9267 1.9262 16.0004 144.9863 0.00016012 -85.6613 0.85295
2.957 0.98805 5.5067e-005 3.8182 0.012009 3.8803e-005 0.0011559 0.21577 0.00065916 0.21642 0.19924 0 0.033175 0.0389 0 1.0662 0.32625 0.094393 0.012546 5.6232 0.078306 9.6343e-005 0.81179 0.0063594 0.0071395 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14078 0.95168 0.9193 0.0013959 0.9946 0.59387 0.0018807 0.43084 1.9271 1.9266 16.0004 144.9863 0.00016005 -85.6613 0.85395
2.958 0.98805 5.5067e-005 3.8182 0.012009 3.8817e-005 0.0011559 0.21578 0.00065916 0.21644 0.19926 0 0.033174 0.0389 0 1.0663 0.3263 0.094409 0.012548 5.6243 0.078317 9.6358e-005 0.81178 0.0063601 0.0071402 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14079 0.95178 0.91935 0.0013959 0.99461 0.59401 0.0018807 0.43085 1.9275 1.9269 16.0004 144.9864 0.00015998 -85.6614 0.85495
2.959 0.98805 5.5067e-005 3.8182 0.012009 3.883e-005 0.0011559 0.2158 0.00065916 0.21645 0.19927 0 0.033174 0.0389 0 1.0664 0.32634 0.094425 0.012549 5.6254 0.078329 9.6373e-005 0.81177 0.0063609 0.007141 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.1408 0.95188 0.91939 0.0013959 0.99463 0.59416 0.0018807 0.43087 1.9278 1.9273 16.0003 144.9864 0.00015992 -85.6614 0.85595
2.96 0.98805 5.5067e-005 3.8182 0.012009 3.8843e-005 0.0011559 0.21581 0.00065916 0.21647 0.19929 0 0.033173 0.0389 0 1.0665 0.32639 0.094441 0.012551 5.6266 0.07834 9.6388e-005 0.81176 0.0063616 0.0071418 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.1408 0.95198 0.91943 0.0013959 0.99465 0.5943 0.0018807 0.43088 1.9282 1.9277 16.0003 144.9864 0.00015985 -85.6615 0.85695
2.961 0.98805 5.5066e-005 3.8182 0.012009 3.8856e-005 0.0011559 0.21583 0.00065916 0.21648 0.1993 0 0.033172 0.0389 0 1.0666 0.32643 0.094457 0.012553 5.6277 0.078351 9.6402e-005 0.81175 0.0063623 0.0071425 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.14081 0.95208 0.91948 0.0013959 0.99466 0.59444 0.0018807 0.43089 1.9286 1.928 16.0003 144.9864 0.00015978 -85.6616 0.85795
2.962 0.98805 5.5066e-005 3.8182 0.012009 3.8869e-005 0.0011559 0.21584 0.00065916 0.2165 0.19931 0 0.033171 0.0389 0 1.0667 0.32648 0.094473 0.012555 5.6289 0.078362 9.6417e-005 0.81173 0.006363 0.0071433 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14081 0.95218 0.91952 0.0013959 0.99468 0.59458 0.0018807 0.4309 1.9289 1.9284 16.0002 144.9864 0.00015971 -85.6616 0.85895
2.963 0.98805 5.5066e-005 3.8182 0.012009 3.8882e-005 0.0011559 0.21586 0.00065916 0.21651 0.19933 0 0.03317 0.0389 0 1.0668 0.32653 0.09449 0.012557 5.63 0.078373 9.6432e-005 0.81172 0.0063637 0.007144 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14082 0.95228 0.91956 0.0013959 0.99469 0.59472 0.0018807 0.43091 1.9293 1.9287 16.0002 144.9865 0.00015964 -85.6617 0.85995
2.964 0.98805 5.5066e-005 3.8182 0.012009 3.8895e-005 0.0011559 0.21587 0.00065916 0.21653 0.19934 0 0.03317 0.0389 0 1.0669 0.32657 0.094506 0.012558 5.6312 0.078384 9.6447e-005 0.81171 0.0063645 0.0071448 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14083 0.95237 0.91961 0.0013959 0.99471 0.59486 0.0018807 0.43093 1.9296 1.9291 16.0002 144.9865 0.00015958 -85.6617 0.86095
2.965 0.98805 5.5066e-005 3.8182 0.012009 3.8908e-005 0.0011559 0.21589 0.00065916 0.21654 0.19936 0 0.033169 0.0389 0 1.067 0.32662 0.094522 0.01256 5.6323 0.078395 9.6462e-005 0.8117 0.0063652 0.0071456 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14083 0.95247 0.91965 0.0013959 0.99473 0.595 0.0018806 0.43094 1.93 1.9295 16.0001 144.9865 0.00015951 -85.6618 0.86195
2.966 0.98805 5.5066e-005 3.8182 0.012009 3.8921e-005 0.0011559 0.21591 0.00065916 0.21656 0.19937 0 0.033168 0.0389 0 1.0671 0.32666 0.094538 0.012562 5.6335 0.078406 9.6477e-005 0.81169 0.0063659 0.0071463 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.14084 0.95257 0.91969 0.0013959 0.99474 0.59514 0.0018806 0.43095 1.9304 1.9298 16.0001 144.9865 0.00015944 -85.6618 0.86295
2.967 0.98805 5.5066e-005 3.8182 0.012009 3.8934e-005 0.0011559 0.21592 0.00065916 0.21658 0.19939 0 0.033167 0.0389 0 1.0672 0.32671 0.094554 0.012564 5.6346 0.078417 9.6492e-005 0.81168 0.0063666 0.0071471 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.14084 0.95266 0.91973 0.0013959 0.99476 0.59528 0.0018806 0.43096 1.9307 1.9302 16.0001 144.9865 0.00015938 -85.6619 0.86395
2.968 0.98805 5.5066e-005 3.8182 0.012009 3.8947e-005 0.0011559 0.21594 0.00065916 0.21659 0.1994 0 0.033166 0.0389 0 1.0673 0.32675 0.09457 0.012565 5.6357 0.078428 9.6507e-005 0.81167 0.0063673 0.0071479 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.14085 0.95276 0.91978 0.0013959 0.99477 0.59543 0.0018806 0.43097 1.9311 1.9305 16 144.9866 0.00015931 -85.6619 0.86495
2.969 0.98805 5.5066e-005 3.8182 0.012009 3.896e-005 0.0011559 0.21595 0.00065916 0.21661 0.19942 0 0.033166 0.0389 0 1.0674 0.3268 0.094586 0.012567 5.6369 0.078439 9.6522e-005 0.81166 0.0063681 0.0071486 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14086 0.95286 0.91982 0.0013959 0.99479 0.59557 0.0018806 0.43098 1.9314 1.9309 16 144.9866 0.00015924 -85.662 0.86595
2.97 0.98805 5.5066e-005 3.8182 0.012009 3.8973e-005 0.0011559 0.21597 0.00065916 0.21662 0.19943 0 0.033165 0.0389 0 1.0675 0.32684 0.094602 0.012569 5.638 0.07845 9.6537e-005 0.81165 0.0063688 0.0071494 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14086 0.95295 0.91986 0.0013958 0.99481 0.59571 0.0018806 0.431 1.9318 1.9312 16 144.9866 0.00015918 -85.662 0.86695
2.971 0.98805 5.5066e-005 3.8182 0.012009 3.8986e-005 0.0011559 0.21598 0.00065916 0.21664 0.19945 0 0.033164 0.0389 0 1.0676 0.32689 0.094618 0.012571 5.6392 0.078461 9.6552e-005 0.81164 0.0063695 0.0071501 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14087 0.95305 0.9199 0.0013958 0.99482 0.59585 0.0018806 0.43101 1.9321 1.9316 16 144.9866 0.00015911 -85.6621 0.86795
2.972 0.98805 5.5066e-005 3.8182 0.012009 3.8999e-005 0.0011559 0.216 0.00065916 0.21665 0.19946 0 0.033163 0.0389 0 1.0677 0.32693 0.094634 0.012572 5.6403 0.078472 9.6567e-005 0.81162 0.0063702 0.0071509 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14087 0.95314 0.91994 0.0013958 0.99484 0.59599 0.0018806 0.43102 1.9325 1.932 15.9999 144.9866 0.00015905 -85.6621 0.86895
2.973 0.98805 5.5066e-005 3.8182 0.012009 3.9012e-005 0.0011559 0.21601 0.00065916 0.21667 0.19948 0 0.033162 0.0389 0 1.0678 0.32698 0.09465 0.012574 5.6415 0.078483 9.6581e-005 0.81161 0.0063709 0.0071517 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14088 0.95324 0.91998 0.0013958 0.99485 0.59613 0.0018806 0.43103 1.9328 1.9323 15.9999 144.9867 0.00015898 -85.6622 0.86995
2.974 0.98805 5.5066e-005 3.8182 0.012009 3.9025e-005 0.0011559 0.21603 0.00065916 0.21668 0.19949 0 0.033161 0.0389 0 1.0679 0.32702 0.094666 0.012576 5.6426 0.078494 9.6596e-005 0.8116 0.0063717 0.0071524 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14088 0.95333 0.92003 0.0013958 0.99487 0.59627 0.0018806 0.43104 1.9332 1.9327 15.9999 144.9867 0.00015892 -85.6622 0.87095
2.975 0.98805 5.5066e-005 3.8182 0.012009 3.9038e-005 0.0011559 0.21604 0.00065916 0.2167 0.19951 0 0.033161 0.0389 0 1.068 0.32707 0.094682 0.012578 5.6438 0.078505 9.6611e-005 0.81159 0.0063724 0.0071532 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14089 0.95343 0.92007 0.0013958 0.99488 0.59641 0.0018806 0.43105 1.9336 1.933 15.9998 144.9867 0.00015885 -85.6623 0.87195
2.976 0.98805 5.5065e-005 3.8182 0.012009 3.9052e-005 0.0011559 0.21606 0.00065916 0.21671 0.19952 0 0.03316 0.0389 0 1.0681 0.32712 0.094698 0.01258 5.6449 0.078517 9.6626e-005 0.81158 0.0063731 0.007154 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.1409 0.95352 0.92011 0.0013958 0.9949 0.59655 0.0018806 0.43107 1.9339 1.9334 15.9998 144.9867 0.00015879 -85.6623 0.87295
2.977 0.98805 5.5065e-005 3.8182 0.012009 3.9065e-005 0.0011559 0.21608 0.00065916 0.21673 0.19953 0 0.033159 0.0389 0 1.0682 0.32716 0.094714 0.012581 5.6461 0.078528 9.6641e-005 0.81157 0.0063738 0.0071547 0.0013839 0.98697 0.99172 2.9836e-006 1.1934e-005 0.1409 0.95362 0.92015 0.0013958 0.99491 0.59669 0.0018805 0.43108 1.9343 1.9337 15.9998 144.9867 0.00015872 -85.6624 0.87395
2.978 0.98805 5.5065e-005 3.8182 0.012009 3.9078e-005 0.0011559 0.21609 0.00065916 0.21675 0.19955 0 0.033158 0.0389 0 1.0683 0.32721 0.09473 0.012583 5.6472 0.078539 9.6656e-005 0.81156 0.0063745 0.0071555 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.14091 0.95371 0.92019 0.0013958 0.99493 0.59683 0.0018805 0.43109 1.9346 1.9341 15.9997 144.9868 0.00015866 -85.6624 0.87495
2.979 0.98805 5.5065e-005 3.8182 0.012009 3.9091e-005 0.0011559 0.21611 0.00065916 0.21676 0.19956 0 0.033157 0.0389 0 1.0684 0.32725 0.094746 0.012585 5.6484 0.07855 9.6671e-005 0.81155 0.0063753 0.0071562 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.14091 0.9538 0.92023 0.0013958 0.99494 0.59697 0.0018805 0.4311 1.935 1.9344 15.9997 144.9868 0.0001586 -85.6625 0.87595
2.98 0.98805 5.5065e-005 3.8182 0.012009 3.9104e-005 0.0011559 0.21612 0.00065916 0.21678 0.19958 0 0.033157 0.0389 0 1.0684 0.3273 0.094762 0.012587 5.6495 0.078561 9.6686e-005 0.81154 0.006376 0.007157 0.0013838 0.98698 0.99172 2.9836e-006 1.1934e-005 0.14092 0.9539 0.92027 0.0013958 0.99496 0.59711 0.0018805 0.43111 1.9353 1.9348 15.9997 144.9868 0.00015853 -85.6625 0.87695
2.981 0.98805 5.5065e-005 3.8182 0.012009 3.9117e-005 0.0011559 0.21614 0.00065916 0.21679 0.19959 0 0.033156 0.0389 0 1.0685 0.32734 0.094778 0.012588 5.6507 0.078572 9.6701e-005 0.81152 0.0063767 0.0071578 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14093 0.95399 0.92031 0.0013958 0.99497 0.59725 0.0018805 0.43112 1.9357 1.9351 15.9996 144.9868 0.00015847 -85.6626 0.87795
2.982 0.98805 5.5065e-005 3.8182 0.012009 3.913e-005 0.0011559 0.21615 0.00065916 0.21681 0.19961 0 0.033155 0.0389 0 1.0686 0.32739 0.094795 0.01259 5.6518 0.078583 9.6716e-005 0.81151 0.0063774 0.0071585 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14093 0.95408 0.92035 0.0013958 0.99498 0.59739 0.0018805 0.43114 1.936 1.9355 15.9996 144.9868 0.0001584 -85.6626 0.87895
2.983 0.98805 5.5065e-005 3.8182 0.012009 3.9143e-005 0.0011559 0.21617 0.00065916 0.21682 0.19962 0 0.033154 0.0389 0 1.0687 0.32743 0.094811 0.012592 5.653 0.078594 9.6731e-005 0.8115 0.0063781 0.0071593 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14094 0.95417 0.92039 0.0013958 0.995 0.59753 0.0018805 0.43115 1.9364 1.9358 15.9996 144.9869 0.00015834 -85.6627 0.87995
2.984 0.98805 5.5065e-005 3.8182 0.012009 3.9156e-005 0.0011559 0.21618 0.00065916 0.21684 0.19964 0 0.033153 0.0389 0 1.0688 0.32748 0.094827 0.012594 5.6541 0.078605 9.6745e-005 0.81149 0.0063789 0.0071601 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14094 0.95426 0.92043 0.0013958 0.99501 0.59767 0.0018805 0.43116 1.9367 1.9362 15.9995 144.9869 0.00015828 -85.6627 0.88095
2.985 0.98805 5.5065e-005 3.8182 0.012009 3.9169e-005 0.0011559 0.2162 0.00065916 0.21685 0.19965 0 0.033153 0.0389 0 1.0689 0.32752 0.094843 0.012595 5.6553 0.078616 9.676e-005 0.81148 0.0063796 0.0071608 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.14095 0.95436 0.92047 0.0013958 0.99503 0.59781 0.0018805 0.43117 1.937 1.9365 15.9995 144.9869 0.00015822 -85.6628 0.88195
2.986 0.98805 5.5065e-005 3.8182 0.012009 3.9182e-005 0.0011559 0.21621 0.00065916 0.21687 0.19966 0 0.033152 0.0389 0 1.069 0.32757 0.094859 0.012597 5.6564 0.078627 9.6775e-005 0.81147 0.0063803 0.0071616 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.14095 0.95445 0.92051 0.0013957 0.99504 0.59795 0.0018805 0.43118 1.9374 1.9369 15.9995 144.9869 0.00015815 -85.6628 0.88295
2.987 0.98805 5.5065e-005 3.8182 0.012009 3.9195e-005 0.0011559 0.21623 0.00065916 0.21688 0.19968 0 0.033151 0.0389 0 1.0691 0.32762 0.094875 0.012599 5.6576 0.078638 9.679e-005 0.81146 0.006381 0.0071624 0.0013837 0.98698 0.99172 2.9834e-006 1.1933e-005 0.14096 0.95454 0.92055 0.0013957 0.99505 0.59809 0.0018805 0.43119 1.9377 1.9372 15.9994 144.987 0.00015809 -85.6629 0.88395
2.988 0.98805 5.5065e-005 3.8182 0.012009 3.9208e-005 0.0011559 0.21624 0.00065916 0.2169 0.19969 0 0.03315 0.0389 0 1.0692 0.32766 0.094891 0.012601 5.6587 0.078649 9.6805e-005 0.81145 0.0063817 0.0071631 0.0013837 0.98698 0.99172 2.9834e-006 1.1933e-005 0.14097 0.95463 0.92059 0.0013957 0.99507 0.59823 0.0018805 0.4312 1.9381 1.9376 15.9994 144.987 0.00015803 -85.6629 0.88495
2.989 0.98805 5.5065e-005 3.8182 0.012009 3.9221e-005 0.0011559 0.21626 0.00065916 0.21691 0.19971 0 0.033149 0.0389 0 1.0693 0.32771 0.094907 0.012603 5.6599 0.07866 9.682e-005 0.81144 0.0063825 0.0071639 0.0013837 0.98698 0.99172 2.9833e-006 1.1933e-005 0.14097 0.95472 0.92063 0.0013957 0.99508 0.59837 0.0018805 0.43122 1.9384 1.9379 15.9994 144.987 0.00015797 -85.663 0.88595
2.99 0.98805 5.5065e-005 3.8182 0.012009 3.9234e-005 0.0011559 0.21627 0.00065916 0.21693 0.19972 0 0.033149 0.0389 0 1.0694 0.32775 0.094923 0.012604 5.6611 0.078671 9.6835e-005 0.81143 0.0063832 0.0071646 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14098 0.95481 0.92067 0.0013957 0.9951 0.59851 0.0018805 0.43123 1.9388 1.9383 15.9994 144.987 0.00015791 -85.663 0.88695
2.991 0.98805 5.5064e-005 3.8182 0.012009 3.9247e-005 0.0011559 0.21629 0.00065916 0.21694 0.19974 0 0.033148 0.0389 0 1.0695 0.3278 0.094939 0.012606 5.6622 0.078682 9.685e-005 0.81141 0.0063839 0.0071654 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14098 0.9549 0.92071 0.0013957 0.99511 0.59865 0.0018804 0.43124 1.9391 1.9386 15.9993 144.987 0.00015784 -85.663 0.88795
2.992 0.98805 5.5064e-005 3.8182 0.012009 3.926e-005 0.0011559 0.2163 0.00065916 0.21696 0.19975 0 0.033147 0.0389 0 1.0696 0.32784 0.094955 0.012608 5.6634 0.078693 9.6865e-005 0.8114 0.0063846 0.0071662 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14099 0.95499 0.92075 0.0013957 0.99512 0.59879 0.0018804 0.43125 1.9395 1.939 15.9993 144.9871 0.00015778 -85.6631 0.88895
2.993 0.98805 5.5064e-005 3.8182 0.012009 3.9273e-005 0.0011559 0.21632 0.00065916 0.21697 0.19977 0 0.033146 0.0389 0 1.0697 0.32789 0.094971 0.01261 5.6645 0.078704 9.688e-005 0.81139 0.0063853 0.0071669 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.141 0.95508 0.92079 0.0013957 0.99514 0.59893 0.0018804 0.43126 1.9398 1.9393 15.9993 144.9871 0.00015772 -85.6631 0.88995
2.994 0.98805 5.5064e-005 3.8182 0.012009 3.9287e-005 0.0011559 0.21633 0.00065916 0.21699 0.19978 0 0.033145 0.0389 0 1.0698 0.32793 0.094987 0.012611 5.6657 0.078715 9.6895e-005 0.81138 0.0063861 0.0071677 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.141 0.95517 0.92082 0.0013957 0.99515 0.59907 0.0018804 0.43127 1.9401 1.9396 15.9992 144.9871 0.00015766 -85.6632 0.89095
2.995 0.98805 5.5064e-005 3.8182 0.012009 3.93e-005 0.0011559 0.21635 0.00065916 0.217 0.19979 0 0.033145 0.0389 0 1.0699 0.32798 0.095003 0.012613 5.6668 0.078726 9.691e-005 0.81137 0.0063868 0.0071685 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14101 0.95526 0.92086 0.0013957 0.99516 0.59921 0.0018804 0.43129 1.9405 1.94 15.9992 144.9871 0.0001576 -85.6632 0.89195
2.996 0.98805 5.5064e-005 3.8182 0.012009 3.9313e-005 0.0011559 0.21636 0.00065916 0.21702 0.19981 0 0.033144 0.0389 0 1.07 0.32802 0.095019 0.012615 5.668 0.078737 9.6924e-005 0.81136 0.0063875 0.0071692 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14101 0.95534 0.9209 0.0013957 0.99518 0.59935 0.0018804 0.4313 1.9408 1.9403 15.9992 144.9871 0.00015754 -85.6633 0.89295
2.997 0.98805 5.5064e-005 3.8182 0.012009 3.9326e-005 0.0011559 0.21638 0.00065916 0.21703 0.19982 0 0.033143 0.0389 0 1.0701 0.32807 0.095035 0.012617 5.6691 0.078749 9.6939e-005 0.81135 0.0063882 0.00717 0.0013836 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14102 0.95543 0.92094 0.0013957 0.99519 0.59949 0.0018804 0.43131 1.9412 1.9407 15.9991 144.9872 0.00015748 -85.6633 0.89395
2.998 0.98805 5.5064e-005 3.8182 0.012009 3.9339e-005 0.0011559 0.21639 0.00065916 0.21705 0.19984 0 0.033142 0.0389 0 1.0702 0.32812 0.095051 0.012618 5.6703 0.07876 9.6954e-005 0.81134 0.0063889 0.0071708 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14103 0.95552 0.92098 0.0013957 0.9952 0.59963 0.0018804 0.43132 1.9415 1.941 15.9991 144.9872 0.00015742 -85.6633 0.89495
2.999 0.98805 5.5064e-005 3.8182 0.012009 3.9352e-005 0.0011559 0.21641 0.00065916 0.21706 0.19985 0 0.033142 0.0389 0 1.0703 0.32816 0.095067 0.01262 5.6715 0.078771 9.6969e-005 0.81133 0.0063897 0.0071715 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14103 0.95561 0.92102 0.0013957 0.99521 0.59977 0.0018804 0.43133 1.9418 1.9413 15.9991 144.9872 0.00015736 -85.6634 0.89595
3 0.98805 5.5064e-005 3.8182 0.012009 3.9365e-005 0.0011559 0.21642 0.00065916 0.21708 0.19987 0 0.033141 0.0389 0 1.0704 0.32821 0.095084 0.012622 5.6726 0.078782 9.6984e-005 0.81132 0.0063904 0.0071723 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14104 0.95569 0.92105 0.0013957 0.99523 0.59991 0.0018804 0.43134 1.9422 1.9417 15.999 144.9872 0.0001573 -85.6634 0.89695
3.001 0.98805 5.5064e-005 3.8182 0.012009 3.9378e-005 0.0011559 0.21644 0.00065916 0.21709 0.19988 0 0.03314 0.0389 0 1.0705 0.32825 0.0951 0.012624 5.6738 0.078793 9.6999e-005 0.8113 0.0063911 0.007173 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14104 0.95578 0.92109 0.0013957 0.99524 0.60005 0.0018804 0.43135 1.9425 1.942 15.999 144.9872 0.00015724 -85.6635 0.89795
3.002 0.98805 5.5064e-005 3.8182 0.012009 3.9391e-005 0.0011559 0.21646 0.00065916 0.21711 0.19989 0 0.033139 0.0389 0 1.0706 0.3283 0.095116 0.012626 5.6749 0.078804 9.7014e-005 0.81129 0.0063918 0.0071738 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14105 0.95587 0.92113 0.0013957 0.99525 0.60019 0.0018804 0.43137 1.9429 1.9424 15.999 144.9873 0.00015718 -85.6635 0.89895
3.003 0.98805 5.5064e-005 3.8182 0.012009 3.9404e-005 0.0011559 0.21647 0.00065916 0.21712 0.19991 0 0.033138 0.0389 0 1.0707 0.32834 0.095132 0.012627 5.6761 0.078815 9.7029e-005 0.81128 0.0063925 0.0071746 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14105 0.95596 0.92117 0.0013957 0.99526 0.60033 0.0018804 0.43138 1.9432 1.9427 15.9989 144.9873 0.00015712 -85.6635 0.89995
3.004 0.98805 5.5064e-005 3.8182 0.012009 3.9417e-005 0.0011559 0.21649 0.00065916 0.21714 0.19992 0 0.033138 0.0389 0 1.0708 0.32839 0.095148 0.012629 5.6773 0.078826 9.7044e-005 0.81127 0.0063933 0.0071753 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14106 0.95604 0.9212 0.0013957 0.99528 0.60046 0.0018804 0.43139 1.9435 1.943 15.9989 144.9873 0.00015706 -85.6636 0.90095
3.005 0.98805 5.5063e-005 3.8182 0.012009 3.943e-005 0.0011559 0.2165 0.00065916 0.21715 0.19994 0 0.033137 0.0389 0 1.0709 0.32843 0.095164 0.012631 5.6784 0.078837 9.7059e-005 0.81126 0.006394 0.0071761 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14107 0.95613 0.92124 0.0013957 0.99529 0.6006 0.0018804 0.4314 1.9439 1.9434 15.9989 144.9873 0.000157 -85.6636 0.90195
3.006 0.98805 5.5063e-005 3.8182 0.012009 3.9443e-005 0.0011559 0.21652 0.00065916 0.21717 0.19995 0 0.033136 0.0389 0 1.071 0.32848 0.09518 0.012633 5.6796 0.078848 9.7074e-005 0.81125 0.0063947 0.0071769 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14107 0.95621 0.92128 0.0013957 0.9953 0.60074 0.0018803 0.43141 1.9442 1.9437 15.9988 144.9873 0.00015694 -85.6637 0.90295
3.007 0.98805 5.5063e-005 3.8182 0.012009 3.9456e-005 0.001156 0.21653 0.00065916 0.21718 0.19997 0 0.033135 0.0389 0 1.0711 0.32852 0.095196 0.012634 5.6807 0.078859 9.7088e-005 0.81124 0.0063954 0.0071776 0.0013835 0.98698 0.99173 2.9829e-006 1.1932e-005 0.14108 0.9563 0.92132 0.0013957 0.99531 0.60088 0.0018803 0.43142 1.9445 1.944 15.9988 144.9874 0.00015689 -85.6637 0.90395
3.008 0.98805 5.5063e-005 3.8182 0.012009 3.9469e-005 0.001156 0.21655 0.00065916 0.2172 0.19998 0 0.033134 0.0389 0 1.0712 0.32857 0.095212 0.012636 5.6819 0.07887 9.7103e-005 0.81123 0.0063962 0.0071784 0.0013835 0.98698 0.99173 2.9829e-006 1.1932e-005 0.14108 0.95638 0.92135 0.0013956 0.99533 0.60102 0.0018803 0.43144 1.9449 1.9444 15.9988 144.9874 0.00015683 -85.6637 0.90495
3.009 0.98805 5.5063e-005 3.8182 0.012009 3.9482e-005 0.001156 0.21656 0.00065916 0.21721 0.19999 0 0.033134 0.0389 0 1.0713 0.32862 0.095228 0.012638 5.6831 0.078881 9.7118e-005 0.81122 0.0063969 0.0071792 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.14109 0.95647 0.92139 0.0013956 0.99534 0.60116 0.0018803 0.43145 1.9452 1.9447 15.9987 144.9874 0.00015677 -85.6638 0.90595
3.01 0.98805 5.5063e-005 3.8182 0.012009 3.9495e-005 0.001156 0.21657 0.00065916 0.21723 0.20001 0 0.033133 0.0389 0 1.0714 0.32866 0.095244 0.01264 5.6842 0.078892 9.7133e-005 0.81121 0.0063976 0.0071799 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.1411 0.95655 0.92143 0.0013956 0.99535 0.6013 0.0018803 0.43146 1.9455 1.9451 15.9987 144.9874 0.00015671 -85.6638 0.90695
3.011 0.98805 5.5063e-005 3.8182 0.012009 3.9508e-005 0.001156 0.21659 0.00065916 0.21724 0.20002 0 0.033132 0.0389 0 1.0715 0.32871 0.09526 0.012641 5.6854 0.078903 9.7148e-005 0.81119 0.0063983 0.0071807 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.1411 0.95664 0.92146 0.0013956 0.99536 0.60144 0.0018803 0.43147 1.9459 1.9454 15.9987 144.9874 0.00015666 -85.6639 0.90795
3.012 0.98805 5.5063e-005 3.8182 0.012009 3.9522e-005 0.001156 0.2166 0.00065916 0.21726 0.20004 0 0.033131 0.0389 0 1.0716 0.32875 0.095276 0.012643 5.6866 0.078914 9.7163e-005 0.81118 0.006399 0.0071815 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14111 0.95672 0.9215 0.0013956 0.99537 0.60158 0.0018803 0.43148 1.9462 1.9457 15.9986 144.9875 0.0001566 -85.6639 0.90895
3.013 0.98805 5.5063e-005 3.8182 0.012009 3.9535e-005 0.001156 0.21662 0.00065916 0.21727 0.20005 0 0.033131 0.0389 0 1.0717 0.3288 0.095292 0.012645 5.6877 0.078925 9.7178e-005 0.81117 0.0063998 0.0071822 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14111 0.95681 0.92154 0.0013956 0.99539 0.60171 0.0018803 0.43149 1.9465 1.946 15.9986 144.9875 0.00015654 -85.6639 0.90995
3.014 0.98805 5.5063e-005 3.8182 0.012008 3.9548e-005 0.001156 0.21663 0.00065916 0.21729 0.20006 0 0.03313 0.0389 0 1.0718 0.32884 0.095308 0.012647 5.6889 0.078936 9.7193e-005 0.81116 0.0064005 0.007183 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14112 0.95689 0.92157 0.0013956 0.9954 0.60185 0.0018803 0.4315 1.9469 1.9464 15.9986 144.9875 0.00015648 -85.664 0.91095
3.015 0.98805 5.5063e-005 3.8182 0.012008 3.9561e-005 0.001156 0.21665 0.00065916 0.2173 0.20008 0 0.033129 0.0389 0 1.0719 0.32889 0.095324 0.012648 5.6901 0.078947 9.7208e-005 0.81115 0.0064012 0.0071837 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14112 0.95697 0.92161 0.0013956 0.99541 0.60199 0.0018803 0.43152 1.9472 1.9467 15.9985 144.9875 0.00015643 -85.664 0.91195
3.016 0.98805 5.5063e-005 3.8182 0.012008 3.9574e-005 0.001156 0.21666 0.00065917 0.21732 0.20009 0 0.033128 0.0389 0 1.072 0.32893 0.095341 0.01265 5.6912 0.078958 9.7223e-005 0.81114 0.0064019 0.0071845 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14113 0.95706 0.92164 0.0013956 0.99542 0.60213 0.0018803 0.43153 1.9475 1.947 15.9985 144.9875 0.00015637 -85.664 0.91295
3.017 0.98805 5.5063e-005 3.8182 0.012008 3.9587e-005 0.001156 0.21668 0.00065917 0.21733 0.20011 0 0.033127 0.0389 0 1.0721 0.32898 0.095357 0.012652 5.6924 0.078969 9.7237e-005 0.81113 0.0064026 0.0071853 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14114 0.95714 0.92168 0.0013956 0.99543 0.60227 0.0018803 0.43154 1.9479 1.9474 15.9985 144.9876 0.00015631 -85.6641 0.91395
3.018 0.98805 5.5063e-005 3.8182 0.012008 3.96e-005 0.001156 0.21669 0.00065917 0.21735 0.20012 0 0.033127 0.0389 0 1.0722 0.32903 0.095373 0.012654 5.6935 0.07898 9.7252e-005 0.81112 0.0064034 0.007186 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14114 0.95722 0.92172 0.0013956 0.99544 0.60241 0.0018803 0.43155 1.9482 1.9477 15.9984 144.9876 0.00015626 -85.6641 0.91495
3.019 0.98805 5.5063e-005 3.8182 0.012008 3.9613e-005 0.001156 0.21671 0.00065917 0.21736 0.20013 0 0.033126 0.0389 0 1.0723 0.32907 0.095389 0.012656 5.6947 0.078991 9.7267e-005 0.81111 0.0064041 0.0071868 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14115 0.9573 0.92175 0.0013956 0.99545 0.60255 0.0018803 0.43156 1.9485 1.948 15.9984 144.9876 0.0001562 -85.6641 0.91595
3.02 0.98805 5.5062e-005 3.8182 0.012008 3.9626e-005 0.001156 0.21672 0.00065917 0.21738 0.20015 0 0.033125 0.0389 0 1.0724 0.32912 0.095405 0.012657 5.6959 0.079002 9.7282e-005 0.81109 0.0064048 0.0071876 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14115 0.95738 0.92179 0.0013956 0.99547 0.60268 0.0018803 0.43157 1.9488 1.9484 15.9984 144.9876 0.00015615 -85.6642 0.91695
3.021 0.98805 5.5062e-005 3.8182 0.012008 3.9639e-005 0.001156 0.21674 0.00065917 0.21739 0.20016 0 0.033124 0.0389 0 1.0725 0.32916 0.095421 0.012659 5.697 0.079013 9.7297e-005 0.81108 0.0064055 0.0071883 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14116 0.95747 0.92182 0.0013956 0.99548 0.60282 0.0018803 0.43158 1.9492 1.9487 15.9984 144.9876 0.00015609 -85.6642 0.91795
3.022 0.98805 5.5062e-005 3.8182 0.012008 3.9652e-005 0.001156 0.21675 0.00065917 0.21741 0.20018 0 0.033124 0.0389 0 1.0726 0.32921 0.095437 0.012661 5.6982 0.079024 9.7312e-005 0.81107 0.0064062 0.0071891 0.0013834 0.98698 0.99173 2.9827e-006 1.193e-005 0.14117 0.95755 0.92186 0.0013956 0.99549 0.60296 0.0018803 0.4316 1.9495 1.949 15.9983 144.9877 0.00015603 -85.6642 0.91895
3.023 0.98805 5.5062e-005 3.8182 0.012008 3.9665e-005 0.001156 0.21677 0.00065917 0.21742 0.20019 0 0.033123 0.0389 0 1.0727 0.32925 0.095453 0.012663 5.6994 0.079035 9.7327e-005 0.81106 0.006407 0.0071899 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14117 0.95763 0.92189 0.0013956 0.9955 0.6031 0.0018802 0.43161 1.9498 1.9493 15.9983 144.9877 0.00015598 -85.6643 0.91995
3.024 0.98805 5.5062e-005 3.8182 0.012008 3.9678e-005 0.001156 0.21678 0.00065917 0.21744 0.2002 0 0.033122 0.0389 0 1.0728 0.3293 0.095469 0.012664 5.7006 0.079046 9.7342e-005 0.81105 0.0064077 0.0071906 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14118 0.95771 0.92193 0.0013956 0.99551 0.60324 0.0018802 0.43162 1.9502 1.9497 15.9983 144.9877 0.00015592 -85.6643 0.92095
3.025 0.98805 5.5062e-005 3.8182 0.012008 3.9691e-005 0.001156 0.2168 0.00065917 0.21745 0.20022 0 0.033121 0.0389 0 1.0729 0.32934 0.095485 0.012666 5.7017 0.079058 9.7357e-005 0.81104 0.0064084 0.0071914 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14118 0.95779 0.92196 0.0013956 0.99552 0.60337 0.0018802 0.43163 1.9505 1.95 15.9982 144.9877 0.00015587 -85.6643 0.92195
3.026 0.98805 5.5062e-005 3.8182 0.012008 3.9704e-005 0.001156 0.21681 0.00065917 0.21747 0.20023 0 0.03312 0.0389 0 1.073 0.32939 0.095501 0.012668 5.7029 0.079069 9.7372e-005 0.81103 0.0064091 0.0071922 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14119 0.95787 0.922 0.0013956 0.99553 0.60351 0.0018802 0.43164 1.9508 1.9503 15.9982 144.9878 0.00015581 -85.6644 0.92295
3.027 0.98805 5.5062e-005 3.8182 0.012008 3.9717e-005 0.001156 0.21683 0.00065917 0.21748 0.20025 0 0.03312 0.0389 0 1.0731 0.32944 0.095517 0.01267 5.7041 0.07908 9.7386e-005 0.81102 0.0064099 0.0071929 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.1412 0.95795 0.92203 0.0013956 0.99554 0.60365 0.0018802 0.43165 1.9511 1.9506 15.9982 144.9878 0.00015576 -85.6644 0.92395
3.028 0.98805 5.5062e-005 3.8182 0.012008 3.973e-005 0.001156 0.21684 0.00065917 0.2175 0.20026 0 0.033119 0.0389 0 1.0732 0.32948 0.095533 0.012671 5.7052 0.079091 9.7401e-005 0.81101 0.0064106 0.0071937 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.1412 0.95803 0.92207 0.0013956 0.99555 0.60379 0.0018802 0.43166 1.9514 1.951 15.9981 144.9878 0.0001557 -85.6644 0.92495
3.029 0.98805 5.5062e-005 3.8182 0.012008 3.9743e-005 0.001156 0.21686 0.00065917 0.21751 0.20027 0 0.033118 0.0389 0 1.0733 0.32953 0.095549 0.012673 5.7064 0.079102 9.7416e-005 0.811 0.0064113 0.0071945 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14121 0.95811 0.9221 0.0013956 0.99556 0.60393 0.0018802 0.43168 1.9518 1.9513 15.9981 144.9878 0.00015565 -85.6645 0.92595
3.03 0.98805 5.5062e-005 3.8182 0.012008 3.9757e-005 0.001156 0.21687 0.00065917 0.21753 0.20029 0 0.033117 0.0389 0 1.0734 0.32957 0.095566 0.012675 5.7076 0.079113 9.7431e-005 0.81098 0.006412 0.0071952 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14121 0.95819 0.92214 0.0013956 0.99557 0.60406 0.0018802 0.43169 1.9521 1.9516 15.9981 144.9878 0.0001556 -85.6645 0.92695
3.031 0.98805 5.5062e-005 3.8182 0.012008 3.977e-005 0.001156 0.21689 0.00065917 0.21754 0.2003 0 0.033117 0.0389 0 1.0735 0.32962 0.095582 0.012677 5.7087 0.079124 9.7446e-005 0.81097 0.0064127 0.007196 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14122 0.95827 0.92217 0.0013956 0.99558 0.6042 0.0018802 0.4317 1.9524 1.9519 15.998 144.9879 0.00015554 -85.6645 0.92795
3.032 0.98805 5.5062e-005 3.8182 0.012008 3.9783e-005 0.001156 0.2169 0.00065917 0.21756 0.20032 0 0.033116 0.0389 0 1.0736 0.32966 0.095598 0.012679 5.7099 0.079135 9.7461e-005 0.81096 0.0064135 0.0071968 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14122 0.95835 0.9222 0.0013955 0.99559 0.60434 0.0018802 0.43171 1.9527 1.9523 15.998 144.9879 0.00015549 -85.6646 0.92895
3.033 0.98805 5.5062e-005 3.8182 0.012008 3.9796e-005 0.001156 0.21692 0.00065917 0.21757 0.20033 0 0.033115 0.0389 0 1.0737 0.32971 0.095614 0.01268 5.7111 0.079146 9.7476e-005 0.81095 0.0064142 0.0071975 0.0013833 0.98698 0.99173 2.9825e-006 1.193e-005 0.14123 0.95843 0.92224 0.0013955 0.9956 0.60448 0.0018802 0.43172 1.9531 1.9526 15.998 144.9879 0.00015543 -85.6646 0.92995
3.034 0.98805 5.5062e-005 3.8182 0.012008 3.9809e-005 0.001156 0.21693 0.00065917 0.21758 0.20034 0 0.033114 0.0389 0 1.0738 0.32975 0.09563 0.012682 5.7123 0.079157 9.7491e-005 0.81094 0.0064149 0.0071983 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.14124 0.95851 0.92227 0.0013955 0.99561 0.60462 0.0018802 0.43173 1.9534 1.9529 15.9979 144.9879 0.00015538 -85.6646 0.93095
3.035 0.98805 5.5061e-005 3.8182 0.012008 3.9822e-005 0.001156 0.21694 0.00065917 0.2176 0.20036 0 0.033114 0.0389 0 1.0739 0.3298 0.095646 0.012684 5.7134 0.079168 9.7506e-005 0.81093 0.0064156 0.0071991 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.14124 0.95858 0.92231 0.0013955 0.99562 0.60475 0.0018802 0.43174 1.9537 1.9532 15.9979 144.9879 0.00015533 -85.6647 0.93195
3.036 0.98805 5.5061e-005 3.8182 0.012008 3.9835e-005 0.001156 0.21696 0.00065917 0.21761 0.20037 0 0.033113 0.0389 0 1.074 0.32984 0.095662 0.012686 5.7146 0.079179 9.7521e-005 0.81092 0.0064163 0.0071998 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.14125 0.95866 0.92234 0.0013955 0.99563 0.60489 0.0018802 0.43175 1.954 1.9535 15.9979 144.988 0.00015528 -85.6647 0.93295
3.037 0.98805 5.5061e-005 3.8182 0.012008 3.9848e-005 0.001156 0.21697 0.00065917 0.21763 0.20039 0 0.033112 0.0389 0 1.0741 0.32989 0.095678 0.012687 5.7158 0.07919 9.7535e-005 0.81091 0.0064171 0.0072006 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.14125 0.95874 0.92237 0.0013955 0.99564 0.60503 0.0018802 0.43177 1.9543 1.9539 15.9978 144.988 0.00015522 -85.6647 0.93395
3.038 0.98805 5.5061e-005 3.8182 0.012008 3.9861e-005 0.001156 0.21699 0.00065917 0.21764 0.2004 0 0.033111 0.0389 0 1.0742 0.32994 0.095694 0.012689 5.717 0.079201 9.755e-005 0.8109 0.0064178 0.0072013 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14126 0.95882 0.92241 0.0013955 0.99565 0.60517 0.0018802 0.43178 1.9547 1.9542 15.9978 144.988 0.00015517 -85.6648 0.93495
3.039 0.98805 5.5061e-005 3.8182 0.012008 3.9874e-005 0.001156 0.217 0.00065917 0.21766 0.20041 0 0.033111 0.0389 0 1.0743 0.32998 0.09571 0.012691 5.7181 0.079212 9.7565e-005 0.81089 0.0064185 0.0072021 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14127 0.95889 0.92244 0.0013955 0.99566 0.6053 0.0018802 0.43179 1.955 1.9545 15.9978 144.988 0.00015512 -85.6648 0.93595
3.04 0.98805 5.5061e-005 3.8182 0.012008 3.9887e-005 0.001156 0.21702 0.00065917 0.21767 0.20043 0 0.03311 0.0389 0 1.0744 0.33003 0.095726 0.012693 5.7193 0.079223 9.758e-005 0.81087 0.0064192 0.0072029 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14127 0.95897 0.92247 0.0013955 0.99567 0.60544 0.0018802 0.4318 1.9553 1.9548 15.9977 144.988 0.00015506 -85.6648 0.93695
3.041 0.98805 5.5061e-005 3.8182 0.012008 3.99e-005 0.001156 0.21703 0.00065917 0.21769 0.20044 0 0.033109 0.0389 0 1.0745 0.33007 0.095742 0.012694 5.7205 0.079234 9.7595e-005 0.81086 0.00642 0.0072036 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14128 0.95905 0.92251 0.0013955 0.99568 0.60558 0.0018802 0.43181 1.9556 1.9551 15.9977 144.9881 0.00015501 -85.6648 0.93795
3.042 0.98805 5.5061e-005 3.8182 0.012008 3.9913e-005 0.001156 0.21705 0.00065917 0.2177 0.20046 0 0.033108 0.0389 0 1.0746 0.33012 0.095758 0.012696 5.7216 0.079245 9.761e-005 0.81085 0.0064207 0.0072044 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14128 0.95913 0.92254 0.0013955 0.99569 0.60571 0.0018801 0.43182 1.9559 1.9555 15.9977 144.9881 0.00015496 -85.6649 0.93895
3.043 0.98805 5.5061e-005 3.8182 0.012008 3.9926e-005 0.001156 0.21706 0.00065917 0.21772 0.20047 0 0.033107 0.0389 0 1.0747 0.33016 0.095774 0.012698 5.7228 0.079256 9.7625e-005 0.81084 0.0064214 0.0072052 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14129 0.9592 0.92257 0.0013955 0.9957 0.60585 0.0018801 0.43183 1.9562 1.9558 15.9976 144.9881 0.00015491 -85.6649 0.93995
3.044 0.98805 5.5061e-005 3.8182 0.012008 3.9939e-005 0.001156 0.21708 0.00065917 0.21773 0.20048 0 0.033107 0.0389 0 1.0748 0.33021 0.095791 0.0127 5.724 0.079267 9.764e-005 0.81083 0.0064221 0.0072059 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14129 0.95928 0.9226 0.0013955 0.99571 0.60599 0.0018801 0.43185 1.9566 1.9561 15.9976 144.9881 0.00015486 -85.6649 0.94095
3.045 0.98805 5.5061e-005 3.8182 0.012008 3.9952e-005 0.001156 0.21709 0.00065917 0.21775 0.2005 0 0.033106 0.0389 0 1.0749 0.33025 0.095807 0.012701 5.7252 0.079278 9.7655e-005 0.81082 0.0064228 0.0072067 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.1413 0.95935 0.92264 0.0013955 0.99572 0.60613 0.0018801 0.43186 1.9569 1.9564 15.9976 144.9881 0.00015481 -85.665 0.94195
3.046 0.98805 5.5061e-005 3.8182 0.012008 3.9965e-005 0.001156 0.21711 0.00065917 0.21776 0.20051 0 0.033105 0.0389 0 1.075 0.3303 0.095823 0.012703 5.7264 0.079289 9.767e-005 0.81081 0.0064236 0.0072075 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14131 0.95943 0.92267 0.0013955 0.99573 0.60626 0.0018801 0.43187 1.9572 1.9567 15.9975 144.9882 0.00015475 -85.665 0.94295
3.047 0.98805 5.5061e-005 3.8182 0.012008 3.9978e-005 0.001156 0.21712 0.00065917 0.21777 0.20052 0 0.033104 0.0389 0 1.0751 0.33035 0.095839 0.012705 5.7275 0.0793 9.7684e-005 0.8108 0.0064243 0.0072082 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.14131 0.9595 0.9227 0.0013955 0.99574 0.6064 0.0018801 0.43188 1.9575 1.957 15.9975 144.9882 0.0001547 -85.665 0.94395
3.048 0.98805 5.5061e-005 3.8182 0.012008 3.9991e-005 0.001156 0.21713 0.00065917 0.21779 0.20054 0 0.033104 0.0389 0 1.0752 0.33039 0.095855 0.012707 5.7287 0.079311 9.7699e-005 0.81079 0.006425 0.007209 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.14132 0.95958 0.92274 0.0013955 0.99575 0.60654 0.0018801 0.43189 1.9578 1.9574 15.9975 144.9882 0.00015465 -85.665 0.94495
3.049 0.98805 5.506e-005 3.8182 0.012008 4.0005e-005 0.001156 0.21715 0.00065917 0.2178 0.20055 0 0.033103 0.0389 0 1.0753 0.33044 0.095871 0.012708 5.7299 0.079322 9.7714e-005 0.81078 0.0064257 0.0072098 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.14132 0.95965 0.92277 0.0013955 0.99576 0.60667 0.0018801 0.4319 1.9581 1.9577 15.9974 144.9882 0.0001546 -85.6651 0.94595
3.05 0.98805 5.506e-005 3.8182 0.012008 4.0018e-005 0.001156 0.21716 0.00065917 0.21782 0.20057 0 0.033102 0.0389 0 1.0754 0.33048 0.095887 0.01271 5.7311 0.079333 9.7729e-005 0.81076 0.0064264 0.0072105 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.14133 0.95973 0.9228 0.0013955 0.99577 0.60681 0.0018801 0.43191 1.9584 1.958 15.9974 144.9882 0.00015455 -85.6651 0.94695
3.051 0.98805 5.506e-005 3.8182 0.012008 4.0031e-005 0.001156 0.21718 0.00065917 0.21783 0.20058 0 0.033101 0.0389 0 1.0755 0.33053 0.095903 0.012712 5.7322 0.079344 9.7744e-005 0.81075 0.0064272 0.0072113 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.14134 0.9598 0.92283 0.0013955 0.99578 0.60695 0.0018801 0.43192 1.9588 1.9583 15.9974 144.9883 0.0001545 -85.6651 0.94795
3.052 0.98805 5.506e-005 3.8182 0.012008 4.0044e-005 0.001156 0.21719 0.00065917 0.21785 0.20059 0 0.033101 0.0389 0 1.0756 0.33057 0.095919 0.012714 5.7334 0.079355 9.7759e-005 0.81074 0.0064279 0.0072121 0.0013832 0.98698 0.99173 2.9822e-006 1.1929e-005 0.14134 0.95988 0.92286 0.0013955 0.99579 0.60708 0.0018801 0.43194 1.9591 1.9586 15.9973 144.9883 0.00015445 -85.6652 0.94895
3.053 0.98805 5.506e-005 3.8182 0.012008 4.0057e-005 0.001156 0.21721 0.00065917 0.21786 0.20061 0 0.0331 0.0389 0 1.0757 0.33062 0.095935 0.012716 5.7346 0.079366 9.7774e-005 0.81073 0.0064286 0.0072128 0.0013832 0.98698 0.99173 2.9822e-006 1.1928e-005 0.14135 0.95995 0.9229 0.0013955 0.9958 0.60722 0.0018801 0.43195 1.9594 1.9589 15.9973 144.9883 0.0001544 -85.6652 0.94995
3.054 0.98805 5.506e-005 3.8182 0.012008 4.007e-005 0.001156 0.21722 0.00065917 0.21788 0.20062 0 0.033099 0.0389 0 1.0758 0.33066 0.095951 0.012717 5.7358 0.079377 9.7789e-005 0.81072 0.0064293 0.0072136 0.0013832 0.98698 0.99173 2.9822e-006 1.1928e-005 0.14135 0.96003 0.92293 0.0013955 0.99581 0.60736 0.0018801 0.43196 1.9597 1.9592 15.9973 144.9883 0.00015435 -85.6652 0.95095
3.055 0.98805 5.506e-005 3.8182 0.012008 4.0083e-005 0.001156 0.21724 0.00065917 0.21789 0.20063 0 0.033098 0.0389 0 1.0759 0.33071 0.095967 0.012719 5.737 0.079388 9.7804e-005 0.81071 0.0064301 0.0072144 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14136 0.9601 0.92296 0.0013955 0.99581 0.60749 0.0018801 0.43197 1.96 1.9595 15.9972 144.9883 0.0001543 -85.6652 0.95195
3.056 0.98805 5.506e-005 3.8182 0.012008 4.0096e-005 0.001156 0.21725 0.00065917 0.2179 0.20065 0 0.033098 0.0389 0 1.076 0.33076 0.095983 0.012721 5.7381 0.079399 9.7818e-005 0.8107 0.0064308 0.0072151 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14137 0.96017 0.92299 0.0013955 0.99582 0.60763 0.0018801 0.43198 1.9603 1.9599 15.9972 144.9884 0.00015425 -85.6653 0.95295
3.057 0.98805 5.506e-005 3.8182 0.012008 4.0109e-005 0.001156 0.21726 0.00065917 0.21792 0.20066 0 0.033097 0.0389 0 1.0761 0.3308 0.096 0.012723 5.7393 0.07941 9.7833e-005 0.81069 0.0064315 0.0072159 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14137 0.96025 0.92302 0.0013955 0.99583 0.60777 0.0018801 0.43199 1.9606 1.9602 15.9972 144.9884 0.0001542 -85.6653 0.95395
3.058 0.98805 5.506e-005 3.8182 0.012008 4.0122e-005 0.001156 0.21728 0.00065917 0.21793 0.20067 0 0.033096 0.0389 0 1.0762 0.33085 0.096016 0.012724 5.7405 0.079421 9.7848e-005 0.81068 0.0064322 0.0072167 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14138 0.96032 0.92305 0.0013955 0.99584 0.6079 0.0018801 0.432 1.9609 1.9605 15.9971 144.9884 0.00015415 -85.6653 0.95495
3.059 0.98805 5.506e-005 3.8182 0.012008 4.0135e-005 0.001156 0.21729 0.00065917 0.21795 0.20069 0 0.033095 0.0389 0 1.0762 0.33089 0.096032 0.012726 5.7417 0.079432 9.7863e-005 0.81067 0.0064329 0.0072174 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14138 0.96039 0.92308 0.0013955 0.99585 0.60804 0.0018801 0.43201 1.9612 1.9608 15.9971 144.9884 0.0001541 -85.6653 0.95595
3.06 0.98805 5.506e-005 3.8182 0.012008 4.0148e-005 0.001156 0.21731 0.00065917 0.21796 0.2007 0 0.033095 0.0389 0 1.0763 0.33094 0.096048 0.012728 5.7429 0.079443 9.7878e-005 0.81065 0.0064337 0.0072182 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14139 0.96046 0.92312 0.0013955 0.99586 0.60818 0.0018801 0.43203 1.9615 1.9611 15.9971 144.9885 0.00015405 -85.6654 0.95695
3.061 0.98805 5.506e-005 3.8182 0.012008 4.0161e-005 0.001156 0.21732 0.00065917 0.21798 0.20072 0 0.033094 0.0389 0 1.0764 0.33098 0.096064 0.01273 5.7441 0.079454 9.7893e-005 0.81064 0.0064344 0.007219 0.0013832 0.98698 0.99173 2.9821e-006 1.1928e-005 0.14139 0.96053 0.92315 0.0013954 0.99587 0.60831 0.0018801 0.43204 1.9619 1.9614 15.997 144.9885 0.000154 -85.6654 0.95795
3.062 0.98805 5.506e-005 3.8182 0.012008 4.0174e-005 0.001156 0.21734 0.00065917 0.21799 0.20073 0 0.033093 0.0389 0 1.0765 0.33103 0.09608 0.012731 5.7452 0.079465 9.7908e-005 0.81063 0.0064351 0.0072197 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.1414 0.96061 0.92318 0.0013954 0.99587 0.60845 0.0018801 0.43205 1.9622 1.9617 15.997 144.9885 0.00015395 -85.6654 0.95895
3.063 0.98805 5.506e-005 3.8182 0.012008 4.0187e-005 0.001156 0.21735 0.00065917 0.218 0.20074 0 0.033092 0.0389 0 1.0766 0.33108 0.096096 0.012733 5.7464 0.079476 9.7923e-005 0.81062 0.0064358 0.0072205 0.0013832 0.98698 0.99173 2.982e-006 1.1928e-005 0.14141 0.96068 0.92321 0.0013954 0.99588 0.60859 0.0018801 0.43206 1.9625 1.962 15.997 144.9885 0.00015391 -85.6654 0.95995
3.064 0.98805 5.5059e-005 3.8182 0.012008 4.02e-005 0.001156 0.21736 0.00065917 0.21802 0.20076 0 0.033092 0.0389 0 1.0767 0.33112 0.096112 0.012735 5.7476 0.079487 9.7938e-005 0.81061 0.0064366 0.0072213 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.14141 0.96075 0.92324 0.0013954 0.99589 0.60872 0.0018801 0.43207 1.9628 1.9623 15.9969 144.9885 0.00015386 -85.6655 0.96095
3.065 0.98805 5.5059e-005 3.8182 0.012008 4.0213e-005 0.001156 0.21738 0.00065917 0.21803 0.20077 0 0.033091 0.0389 0 1.0768 0.33117 0.096128 0.012737 5.7488 0.079498 9.7953e-005 0.8106 0.0064373 0.007222 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.14142 0.96082 0.92327 0.0013954 0.9959 0.60886 0.0018801 0.43208 1.9631 1.9626 15.9969 144.9886 0.00015381 -85.6655 0.96195
3.066 0.98805 5.5059e-005 3.8182 0.012008 4.0226e-005 0.001156 0.21739 0.00065917 0.21805 0.20078 0 0.03309 0.0389 0 1.0769 0.33121 0.096144 0.012738 5.75 0.079509 9.7967e-005 0.81059 0.006438 0.0072228 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.14142 0.96089 0.9233 0.0013954 0.99591 0.60899 0.00188 0.43209 1.9634 1.9629 15.9969 144.9886 0.00015376 -85.6655 0.96295
3.067 0.98805 5.5059e-005 3.8182 0.012008 4.0239e-005 0.001156 0.21741 0.00065917 0.21806 0.2008 0 0.033089 0.0389 0 1.077 0.33126 0.09616 0.01274 5.7512 0.07952 9.7982e-005 0.81058 0.0064387 0.0072236 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.14143 0.96096 0.92333 0.0013954 0.99592 0.60913 0.00188 0.4321 1.9637 1.9632 15.9968 144.9886 0.00015371 -85.6655 0.96395
3.068 0.98805 5.5059e-005 3.8182 0.012008 4.0253e-005 0.001156 0.21742 0.00065917 0.21808 0.20081 0 0.033089 0.0389 0 1.0771 0.3313 0.096176 0.012742 5.7524 0.079531 9.7997e-005 0.81057 0.0064394 0.0072243 0.0013831 0.98698 0.99173 2.982e-006 1.1928e-005 0.14144 0.96103 0.92336 0.0013954 0.99592 0.60927 0.00188 0.43212 1.964 1.9636 15.9968 144.9886 0.00015367 -85.6656 0.96495
3.069 0.98805 5.5059e-005 3.8182 0.012008 4.0266e-005 0.001156 0.21744 0.00065917 0.21809 0.20082 0 0.033088 0.0389 0 1.0772 0.33135 0.096192 0.012744 5.7535 0.079542 9.8012e-005 0.81056 0.0064402 0.0072251 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.14144 0.9611 0.92339 0.0013954 0.99593 0.6094 0.00188 0.43213 1.9643 1.9639 15.9968 144.9886 0.00015362 -85.6656 0.96595
3.07 0.98805 5.5059e-005 3.8182 0.012008 4.0279e-005 0.0011561 0.21745 0.00065917 0.2181 0.20084 0 0.033087 0.0389 0 1.0773 0.33139 0.096209 0.012746 5.7547 0.079553 9.8027e-005 0.81054 0.0064409 0.0072259 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.14145 0.96117 0.92342 0.0013954 0.99594 0.60954 0.00188 0.43214 1.9646 1.9642 15.9967 144.9887 0.00015357 -85.6656 0.96695
3.071 0.98805 5.5059e-005 3.8182 0.012008 4.0292e-005 0.0011561 0.21746 0.00065917 0.21812 0.20085 0 0.033086 0.0389 0 1.0774 0.33144 0.096225 0.012747 5.7559 0.079564 9.8042e-005 0.81053 0.0064416 0.0072266 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.14145 0.96124 0.92345 0.0013954 0.99595 0.60967 0.00188 0.43215 1.9649 1.9645 15.9967 144.9887 0.00015352 -85.6656 0.96795
3.072 0.98805 5.5059e-005 3.8182 0.012008 4.0305e-005 0.0011561 0.21748 0.00065917 0.21813 0.20086 0 0.033086 0.0389 0 1.0775 0.33149 0.096241 0.012749 5.7571 0.079575 9.8057e-005 0.81052 0.0064423 0.0072274 0.0013831 0.98698 0.99173 2.9819e-006 1.1928e-005 0.14146 0.96131 0.92348 0.0013954 0.99596 0.60981 0.00188 0.43216 1.9652 1.9648 15.9967 144.9887 0.00015348 -85.6656 0.96895
3.073 0.98805 5.5059e-005 3.8182 0.012008 4.0318e-005 0.0011561 0.21749 0.00065917 0.21815 0.20088 0 0.033085 0.0389 0 1.0776 0.33153 0.096257 0.012751 5.7583 0.079586 9.8072e-005 0.81051 0.0064431 0.0072282 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.14146 0.96138 0.92351 0.0013954 0.99596 0.60995 0.00188 0.43217 1.9655 1.9651 15.9966 144.9887 0.00015343 -85.6657 0.96995
3.074 0.98805 5.5059e-005 3.8182 0.012008 4.0331e-005 0.0011561 0.21751 0.00065917 0.21816 0.20089 0 0.033084 0.0389 0 1.0777 0.33158 0.096273 0.012753 5.7595 0.079597 9.8086e-005 0.8105 0.0064438 0.0072289 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.14147 0.96145 0.92354 0.0013954 0.99597 0.61008 0.00188 0.43218 1.9658 1.9654 15.9966 144.9887 0.00015338 -85.6657 0.97095
3.075 0.98805 5.5059e-005 3.8182 0.012008 4.0344e-005 0.0011561 0.21752 0.00065917 0.21818 0.2009 0 0.033083 0.0389 0 1.0778 0.33162 0.096289 0.012754 5.7607 0.079608 9.8101e-005 0.81049 0.0064445 0.0072297 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.14148 0.96152 0.92357 0.0013954 0.99598 0.61022 0.00188 0.43219 1.9661 1.9657 15.9966 144.9888 0.00015334 -85.6657 0.97195
3.076 0.98805 5.5059e-005 3.8182 0.012008 4.0357e-005 0.0011561 0.21754 0.00065917 0.21819 0.20092 0 0.033083 0.0389 0 1.0779 0.33167 0.096305 0.012756 5.7619 0.079619 9.8116e-005 0.81048 0.0064452 0.0072305 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.14148 0.96159 0.9236 0.0013954 0.99599 0.61035 0.00188 0.4322 1.9664 1.966 15.9965 144.9888 0.00015329 -85.6657 0.97295
3.077 0.98805 5.5059e-005 3.8182 0.012008 4.037e-005 0.0011561 0.21755 0.00065917 0.2182 0.20093 0 0.033082 0.0389 0 1.078 0.33171 0.096321 0.012758 5.763 0.07963 9.8131e-005 0.81047 0.0064459 0.0072312 0.0013831 0.98698 0.99173 2.9819e-006 1.1927e-005 0.14149 0.96166 0.92363 0.0013954 0.996 0.61049 0.00188 0.43222 1.9667 1.9663 15.9965 144.9888 0.00015324 -85.6658 0.97395
3.078 0.98805 5.5059e-005 3.8182 0.012008 4.0383e-005 0.0011561 0.21756 0.00065917 0.21822 0.20094 0 0.033081 0.0389 0 1.0781 0.33176 0.096337 0.01276 5.7642 0.079641 9.8146e-005 0.81046 0.0064467 0.007232 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.14149 0.96173 0.92366 0.0013954 0.996 0.61062 0.00188 0.43223 1.967 1.9666 15.9965 144.9888 0.0001532 -85.6658 0.97495
3.079 0.98805 5.5058e-005 3.8182 0.012008 4.0396e-005 0.0011561 0.21758 0.00065917 0.21823 0.20096 0 0.033081 0.0389 0 1.0782 0.3318 0.096353 0.012761 5.7654 0.079652 9.8161e-005 0.81045 0.0064474 0.0072328 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.1415 0.9618 0.92369 0.0013954 0.99601 0.61076 0.00188 0.43224 1.9673 1.9669 15.9964 144.9888 0.00015315 -85.6658 0.97595
3.08 0.98805 5.5058e-005 3.8182 0.012008 4.0409e-005 0.0011561 0.21759 0.00065917 0.21825 0.20097 0 0.03308 0.0389 0 1.0783 0.33185 0.096369 0.012763 5.7666 0.079663 9.8176e-005 0.81043 0.0064481 0.0072335 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.14151 0.96186 0.92372 0.0013954 0.99602 0.6109 0.00188 0.43225 1.9676 1.9672 15.9964 144.9889 0.0001531 -85.6658 0.97695
3.081 0.98805 5.5058e-005 3.8182 0.012008 4.0422e-005 0.0011561 0.21761 0.00065917 0.21826 0.20098 0 0.033079 0.0389 0 1.0784 0.3319 0.096385 0.012765 5.7678 0.079674 9.8191e-005 0.81042 0.0064488 0.0072343 0.0013831 0.98698 0.99173 2.9818e-006 1.1927e-005 0.14151 0.96193 0.92375 0.0013954 0.99603 0.61103 0.00188 0.43226 1.9679 1.9675 15.9964 144.9889 0.00015306 -85.6658 0.97795
3.082 0.98805 5.5058e-005 3.8182 0.012007 4.0435e-005 0.0011561 0.21762 0.00065917 0.21827 0.201 0 0.033078 0.0389 0 1.0785 0.33194 0.096402 0.012767 5.769 0.079685 9.8206e-005 0.81041 0.0064496 0.0072351 0.0013831 0.98699 0.99173 2.9818e-006 1.1927e-005 0.14152 0.962 0.92378 0.0013954 0.99603 0.61117 0.00188 0.43227 1.9682 1.9678 15.9963 144.9889 0.00015301 -85.6659 0.97895
3.083 0.98805 5.5058e-005 3.8182 0.012007 4.0448e-005 0.0011561 0.21763 0.00065917 0.21829 0.20101 0 0.033078 0.0389 0 1.0786 0.33199 0.096418 0.012768 5.7702 0.079696 9.822e-005 0.8104 0.0064503 0.0072358 0.0013831 0.98699 0.99173 2.9818e-006 1.1927e-005 0.14152 0.96207 0.92381 0.0013954 0.99604 0.6113 0.00188 0.43228 1.9685 1.9681 15.9963 144.9889 0.00015297 -85.6659 0.97995
3.084 0.98805 5.5058e-005 3.8182 0.012007 4.0461e-005 0.0011561 0.21765 0.00065917 0.2183 0.20102 0 0.033077 0.0389 0 1.0787 0.33203 0.096434 0.01277 5.7714 0.079707 9.8235e-005 0.81039 0.006451 0.0072366 0.001383 0.98699 0.99173 2.9818e-006 1.1927e-005 0.14153 0.96213 0.92383 0.0013954 0.99605 0.61144 0.00188 0.43229 1.9688 1.9684 15.9963 144.9889 0.00015292 -85.6659 0.98095
3.085 0.98805 5.5058e-005 3.8182 0.012007 4.0474e-005 0.0011561 0.21766 0.00065917 0.21832 0.20104 0 0.033076 0.0389 0 1.0788 0.33208 0.09645 0.012772 5.7726 0.079718 9.825e-005 0.81038 0.0064517 0.0072374 0.001383 0.98699 0.99173 2.9818e-006 1.1927e-005 0.14154 0.9622 0.92386 0.0013954 0.99606 0.61157 0.00188 0.4323 1.9691 1.9687 15.9962 144.989 0.00015288 -85.6659 0.98195
3.086 0.98805 5.5058e-005 3.8182 0.012007 4.0487e-005 0.0011561 0.21768 0.00065917 0.21833 0.20105 0 0.033075 0.0389 0 1.0789 0.33212 0.096466 0.012774 5.7738 0.079729 9.8265e-005 0.81037 0.0064524 0.0072381 0.001383 0.98699 0.99173 2.9818e-006 1.1927e-005 0.14154 0.96227 0.92389 0.0013954 0.99606 0.61171 0.00188 0.43232 1.9694 1.969 15.9962 144.989 0.00015283 -85.6659 0.98295
3.087 0.98805 5.5058e-005 3.8182 0.012007 4.0501e-005 0.0011561 0.21769 0.00065917 0.21834 0.20106 0 0.033075 0.0389 0 1.079 0.33217 0.096482 0.012775 5.775 0.07974 9.828e-005 0.81036 0.0064532 0.0072389 0.001383 0.98699 0.99173 2.9818e-006 1.1927e-005 0.14155 0.96233 0.92392 0.0013954 0.99607 0.61184 0.00188 0.43233 1.9697 1.9693 15.9962 144.989 0.00015279 -85.666 0.98395
3.088 0.98805 5.5058e-005 3.8182 0.012007 4.0514e-005 0.0011561 0.2177 0.00065917 0.21836 0.20108 0 0.033074 0.0389 0 1.0791 0.33222 0.096498 0.012777 5.7762 0.079751 9.8295e-005 0.81035 0.0064539 0.0072397 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14155 0.9624 0.92395 0.0013954 0.99608 0.61198 0.00188 0.43234 1.97 1.9696 15.9961 144.989 0.00015274 -85.666 0.98495
3.089 0.98805 5.5058e-005 3.8182 0.012007 4.0527e-005 0.0011561 0.21772 0.00065917 0.21837 0.20109 0 0.033073 0.0389 0 1.0792 0.33226 0.096514 0.012779 5.7774 0.079762 9.831e-005 0.81034 0.0064546 0.0072404 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14156 0.96247 0.92398 0.0013954 0.99608 0.61211 0.00188 0.43235 1.9703 1.9699 15.9961 144.989 0.0001527 -85.666 0.98595
3.09 0.98805 5.5058e-005 3.8182 0.012007 4.054e-005 0.0011561 0.21773 0.00065917 0.21839 0.2011 0 0.033072 0.0389 0 1.0793 0.33231 0.09653 0.012781 5.7785 0.079773 9.8325e-005 0.81033 0.0064553 0.0072412 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14156 0.96253 0.92401 0.0013954 0.99609 0.61225 0.00188 0.43236 1.9706 1.9702 15.9961 144.9891 0.00015265 -85.666 0.98695
3.091 0.98805 5.5058e-005 3.8182 0.012007 4.0553e-005 0.0011561 0.21775 0.00065917 0.2184 0.20112 0 0.033072 0.0389 0 1.0794 0.33235 0.096546 0.012782 5.7797 0.079784 9.834e-005 0.81031 0.0064561 0.007242 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14157 0.9626 0.92403 0.0013954 0.9961 0.61238 0.00188 0.43237 1.9709 1.9704 15.996 144.9891 0.00015261 -85.666 0.98795
3.092 0.98805 5.5058e-005 3.8182 0.012007 4.0566e-005 0.0011561 0.21776 0.00065918 0.21841 0.20113 0 0.033071 0.0389 0 1.0795 0.3324 0.096562 0.012784 5.7809 0.079795 9.8354e-005 0.8103 0.0064568 0.0072427 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14158 0.96266 0.92406 0.0013954 0.99611 0.61252 0.00188 0.43238 1.9712 1.9707 15.996 144.9891 0.00015256 -85.6661 0.98895
3.093 0.98805 5.5057e-005 3.8182 0.012007 4.0579e-005 0.0011561 0.21777 0.00065918 0.21843 0.20114 0 0.03307 0.0389 0 1.0796 0.33244 0.096579 0.012786 5.7821 0.079806 9.8369e-005 0.81029 0.0064575 0.0072435 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14158 0.96273 0.92409 0.0013954 0.99611 0.61265 0.00188 0.43239 1.9715 1.971 15.996 144.9891 0.00015252 -85.6661 0.98995
3.094 0.98805 5.5057e-005 3.8182 0.012007 4.0592e-005 0.0011561 0.21779 0.00065918 0.21844 0.20116 0 0.03307 0.0389 0 1.0797 0.33249 0.096595 0.012788 5.7833 0.079817 9.8384e-005 0.81028 0.0064582 0.0072443 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14159 0.96279 0.92412 0.0013954 0.99612 0.61279 0.00188 0.4324 1.9718 1.9713 15.9959 144.9891 0.00015248 -85.6661 0.99095
3.095 0.98805 5.5057e-005 3.8182 0.012007 4.0605e-005 0.0011561 0.2178 0.00065918 0.21846 0.20117 0 0.033069 0.0389 0 1.0798 0.33254 0.096611 0.01279 5.7845 0.079828 9.8399e-005 0.81027 0.0064589 0.007245 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14159 0.96286 0.92415 0.0013953 0.99613 0.61292 0.00188 0.43242 1.9721 1.9716 15.9959 144.9892 0.00015243 -85.6661 0.99195
3.096 0.98805 5.5057e-005 3.8182 0.012007 4.0618e-005 0.0011561 0.21782 0.00065918 0.21847 0.20118 0 0.033068 0.0389 0 1.0799 0.33258 0.096627 0.012791 5.7857 0.079839 9.8414e-005 0.81026 0.0064597 0.0072458 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.1416 0.96292 0.92417 0.0013953 0.99613 0.61306 0.0018799 0.43243 1.9723 1.9719 15.9959 144.9892 0.00015239 -85.6661 0.99295
3.097 0.98805 5.5057e-005 3.8182 0.012007 4.0631e-005 0.0011561 0.21783 0.00065918 0.21848 0.2012 0 0.033067 0.0389 0 1.08 0.33263 0.096643 0.012793 5.7869 0.07985 9.8429e-005 0.81025 0.0064604 0.0072466 0.001383 0.98699 0.99173 2.9817e-006 1.1927e-005 0.14161 0.96299 0.9242 0.0013953 0.99614 0.61319 0.0018799 0.43244 1.9726 1.9722 15.9958 144.9892 0.00015234 -85.6661 0.99395
3.098 0.98805 5.5057e-005 3.8182 0.012007 4.0644e-005 0.0011561 0.21784 0.00065918 0.2185 0.20121 0 0.033067 0.0389 0 1.0801 0.33267 0.096659 0.012795 5.7881 0.079861 9.8444e-005 0.81024 0.0064611 0.0072473 0.001383 0.98699 0.99173 2.9816e-006 1.1927e-005 0.14161 0.96305 0.92423 0.0013953 0.99615 0.61333 0.0018799 0.43245 1.9729 1.9725 15.9958 144.9892 0.0001523 -85.6662 0.99495
3.099 0.98805 5.5057e-005 3.8182 0.012007 4.0657e-005 0.0011561 0.21786 0.00065918 0.21851 0.20122 0 0.033066 0.0389 0 1.0802 0.33272 0.096675 0.012797 5.7893 0.079872 9.8459e-005 0.81023 0.0064618 0.0072481 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.14162 0.96311 0.92426 0.0013953 0.99615 0.61346 0.0018799 0.43246 1.9732 1.9728 15.9957 144.9893 0.00015226 -85.6662 0.99595
3.1 0.98805 5.5057e-005 3.8182 0.012007 4.067e-005 0.0011561 0.21787 0.00065918 0.21853 0.20124 0 0.033065 0.0389 0 1.0803 0.33276 0.096691 0.012798 5.7905 0.079883 9.8473e-005 0.81022 0.0064626 0.0072489 0.001383 0.98699 0.99173 2.9816e-006 1.1926e-005 0.14162 0.96318 0.92428 0.0013953 0.99616 0.6136 0.0018799 0.43247 1.9735 1.9731 15.9957 144.9893 0.00015222 -85.6656 0.99695
3.101 0.98805 5.5057e-005 3.8182 0.012007 4.0683e-005 0.0011561 0.21789 0.00065918 0.21854 0.20125 0 0.033064 0.0389 0 1.0804 0.33281 0.096707 0.0128 5.7917 0.079894 9.8488e-005 0.8102 0.0064633 0.0072497 0.0064697 0.98324 0.991 1.451e-005 5.3306e-005 0.14163 0.96319 0.92431 0.0027724 0.99615 0.61371 0.0023951 0.43243 1.9738 1.9734 15.9957 144.9893 0.00015218 -76.1643 0.99795
3.102 0.98805 5.5057e-005 3.8182 0.012007 4.0696e-005 0.0011561 0.2179 0.00065918 0.21855 0.20126 0 0.033064 0.0389 0 1.0805 0.33285 0.096723 0.012802 5.7929 0.079905 9.8503e-005 0.81019 0.006464 0.0072504 0.026207 0.97172 0.98767 6.5937e-005 0.00022936 0.14164 0.96298 0.92434 0.0052994 0.9961 0.61381 0.0033357 0.43231 1.9741 1.9737 15.9956 144.9892 0.00015217 -67.1503 0.99895
3.103 0.98805 5.5057e-005 3.8182 0.012007 4.0709e-005 0.0011561 0.21791 0.00065918 0.21857 0.20128 0 0.033063 0.0389 0 1.0806 0.3329 0.096739 0.012804 5.7941 0.079916 9.8518e-005 0.81018 0.0064647 0.0072512 0.094828 0.94724 0.97734 0.00028423 0.00091264 0.14164 0.96223 0.92436 0.0092457 0.99584 0.6139 0.0044245 0.43214 1.9744 1.974 15.9955 144.9892 0.00015218 -58.019 0.99995
3.104 0.98805 5.5057e-005 3.8182 0.012007 4.0722e-005 0.0011561 0.21793 0.00065918 0.21858 0.20129 0 0.033062 0.0389 0 1.0807 0.33295 0.096756 0.012805 5.7953 0.079927 9.8533e-005 0.81017 0.0064654 0.007252 0.48749 0.85656 0.93878 0.0021753 0.0054674 0.14165 0.96021 0.92438 0.015748 0.99173 0.61391 0.0056232 0.43195 1.9747 1.9742 15.9963 144.9892 0.00015222 -37.2482 0.15669
3.105 0.98805 5.5057e-005 3.8182 0.012007 4.0735e-005 0.0011561 0.21794 0.00065918 0.2186 0.2013 0 0.033062 0.0389 0 1.0808 0.33299 0.096772 0.012807 5.7965 0.079938 9.8548e-005 0.81016 0.0064662 0.0072527 0.9996 0.0021805 0.71221 0.93797 0.99597 0.14165 0.92671 0.92142 0.3328 0.96432 0.60044 0.044101 0.43175 1.931 0.95324 16.0002 144.9889 0.00023512 24.2056 0.0019526
3.106 0.98805 5.5057e-005 3.8182 0.012007 4.0749e-005 0.0011561 0.21795 0.00065918 0.21861 0.20132 0 0.033061 0.0389 0 1.0809 0.33304 0.096788 0.012809 5.7977 0.079949 9.8563e-005 0.81015 0.0064669 0.0072535 0.99935 1.4182e-006 0.52835 0.99688 0.99934 0.14166 0.88664 0.90353 0.60534 0.93716 0.58368 0.095721 0.43154 1.7451 0.58788 15.9998 144.9875 0.0003442 18.9585 0.0029526
3.107 0.98805 5.5057e-005 3.8182 0.012007 4.0762e-005 0.0011561 0.21797 0.00065918 0.21862 0.20133 0 0.03306 0.0389 0 1.081 0.33308 0.096804 0.012811 5.7989 0.07996 9.8578e-005 0.81014 0.0064676 0.0072543 0.9988 7.6157e-010 0.39239 0.99413 0.99829 0.14166 0.84924 0.88042 0.72127 0.91076 0.56771 0.1339 0.43134 1.5678 0.5623 15.9994 144.9859 0.00041276 13.297 0.0039526
3.108 0.98805 5.5056e-005 3.8182 0.012007 4.0775e-005 0.0011561 0.21798 0.00065918 0.21864 0.20134 0 0.033059 0.0389 0 1.0811 0.33313 0.09682 0.012812 5.8001 0.079971 9.8592e-005 0.81013 0.0064683 0.007255 0.99818 -9.9186e-011 0.29183 0.9887 0.99665 0.14167 0.81508 0.85484 0.77086 0.88512 0.55276 0.16322 0.43113 1.4198 0.59951 15.9991 144.9842 0.00046375 9.4896 0.0049526
3.109 0.98805 5.5056e-005 3.8182 0.012007 4.0788e-005 0.0011561 0.218 0.00065918 0.21865 0.20135 0 0.033059 0.0389 0 1.0812 0.33317 0.096836 0.012814 5.8013 0.079982 9.8607e-005 0.81012 0.0064691 0.0072558 0.99759 -1.5818e-011 0.21735 0.98205 0.99469 0.14168 0.78394 0.82808 0.79096 0.8602 0.53885 0.18734 0.43093 1.302 0.6567 15.9988 144.9825 0.00050275 6.9593 0.0059526
3.11 0.98805 5.5056e-005 3.8182 0.012007 4.0801e-005 0.0011561 0.21801 0.00065918 0.21866 0.20137 0 0.033058 0.0389 0 1.0813 0.33322 0.096852 0.012816 5.8025 0.079993 9.8622e-005 0.81011 0.0064698 0.0072566 0.99704 -4.974e-011 0.16208 0.97465 0.99252 0.14168 0.75536 0.80103 0.79626 0.83598 0.52591 0.20804 0.43072 1.2115 0.7186 15.9985 144.9809 0.0005325 5.0641 0.0069526
3.111 0.98805 5.5056e-005 3.8182 0.012007 4.0814e-005 0.0011561 0.21802 0.00065918 0.21868 0.20138 0 0.033057 0.0389 0 1.0814 0.33327 0.096868 0.012818 5.8037 0.080004 9.8637e-005 0.81009 0.0064705 0.0072573 0.99647 8.0079e-011 0.12101 0.9665 0.9901 0.14169 0.72902 0.77431 0.7933 0.81246 0.51386 0.22618 0.43052 1.1442 0.77742 15.9982 144.9793 0.00055506 3.4716 0.0079526
3.112 0.98805 5.5056e-005 3.8182 0.012007 4.0827e-005 0.0011561 0.21804 0.00065918 0.21869 0.20139 0 0.033057 0.0389 0 1.0815 0.33331 0.096884 0.012819 5.8049 0.080015 9.8652e-005 0.81008 0.0064712 0.0072581 0.99586 5.0531e-011 0.090461 0.95741 0.98734 0.14169 0.7047 0.74836 0.78526 0.7896 0.50268 0.24221 0.43031 1.0956 0.82898 15.9979 144.9778 0.00057219 2.0203 0.0089526
3.113 0.98805 5.5056e-005 3.8182 0.012007 4.084e-005 0.0011561 0.21805 0.00065918 0.21871 0.20141 0 0.033056 0.0389 0 1.0816 0.33336 0.0969 0.012821 5.8061 0.080026 9.8667e-005 0.81007 0.006472 0.0072589 0.99517 2.8596e-011 0.067713 0.94703 0.98409 0.1417 0.68225 0.72348 0.7738 0.76739 0.49234 0.25641 0.43011 1.0615 0.87155 15.9976 144.9765 0.00058532 0.62316 0.0099526
3.114 0.98805 5.5056e-005 3.8182 0.012007 4.0853e-005 0.0011561 0.21806 0.00065918 0.21872 0.20142 0 0.033055 0.0389 0 1.0817 0.3334 0.096916 0.012823 5.8073 0.080037 9.8682e-005 0.81006 0.0064727 0.0072596 0.99436 7.041e-011 0.05076 0.93493 0.98015 0.14171 0.66158 0.69992 0.75978 0.74582 0.48284 0.26895 0.4299 1.0385 0.90513 15.9973 144.9751 0.00059556 -0.77679 0.010953
3.115 0.98805 5.5056e-005 3.8182 0.012007 4.0866e-005 0.0011561 0.21808 0.00065918 0.21873 0.20143 0 0.033054 0.0389 0 1.0818 0.33345 0.096933 0.012825 5.8085 0.080048 9.8697e-005 0.81005 0.0064734 0.0072604 0.99338 4.1751e-011 0.038118 0.92055 0.97527 0.14171 0.64262 0.67785 0.74362 0.72486 0.47419 0.27995 0.4297 1.0235 0.93074 15.9971 144.9739 0.00060371 -2.2259 0.011953
3.116 0.98805 5.5056e-005 3.8182 0.012007 4.0879e-005 0.0011561 0.21809 0.00065918 0.21875 0.20145 0 0.033054 0.0389 0 1.0819 0.33349 0.096949 0.012826 5.8097 0.080059 9.8711e-005 0.81004 0.0064741 0.0072612 0.99215 -2.0712e-011 0.028684 0.90311 0.96907 0.14172 0.62533 0.65743 0.72544 0.7045 0.46641 0.28948 0.42949 1.0141 0.94985 15.9968 144.9728 0.00061033 -3.7715 0.012953
3.117 0.98805 5.5056e-005 3.8182 0.012007 4.0892e-005 0.0011561 0.21811 0.00065918 0.21876 0.20146 0 0.033053 0.0389 0 1.082 0.33354 0.096965 0.012828 5.811 0.08007 9.8726e-005 0.81003 0.0064748 0.0072619 0.99052 6.0807e-011 0.02164 0.88156 0.96096 0.14172 0.60971 0.6388 0.70517 0.68473 0.45954 0.29758 0.42929 1.0087 0.96397 15.9966 144.9717 0.00061577 -5.4701 0.013953
3.118 0.98805 5.5056e-005 3.8182 0.012007 4.0905e-005 0.0011561 0.21812 0.00065918 0.21877 0.20147 0 0.033052 0.0389 0 1.0821 0.33359 0.096981 0.01283 5.8122 0.080081 9.8741e-005 0.81002 0.0064756 0.0072627 0.98826 -1.9333e-011 0.016381 0.85434 0.95009 0.14173 0.59579 0.62214 0.68254 0.66555 0.45361 0.30426 0.42908 1.006 0.97442 15.9963 144.9708 0.00062024 -7.3971 0.014953
3.119 0.98805 5.5056e-005 3.8182 0.012007 4.0918e-005 0.0011561 0.21813 0.00065918 0.21879 0.20148 0 0.033052 0.0389 0 1.0822 0.33363 0.096997 0.012832 5.8134 0.080092 9.8756e-005 0.81001 0.0064763 0.0072635 0.9849 1.0743e-011 0.012457 0.81916 0.93496 0.14173 0.58362 0.60763 0.65717 0.64693 0.44866 0.30951 0.42888 1.0051 0.98226 15.9961 144.9699 0.00062383 -9.6584 0.015953
3.12 0.98805 5.5056e-005 3.8182 0.012007 4.0931e-005 0.0011561 0.21815 0.00065918 0.2188 0.2015 0 0.033051 0.0389 0 1.0823 0.33368 0.097013 0.012834 5.8146 0.080103 9.8771e-005 0.81 0.006477 0.0072642 0.97951 -1.0375e-011 0.0095354 0.77257 0.91319 0.14174 0.57329 0.59548 0.62856 0.6289 0.44473 0.31329 0.42868 1.0053 0.98829 15.9959 144.9691 0.00062656 -12.4021 0.016953
3.121 0.98805 5.5056e-005 3.8182 0.012007 4.0944e-005 0.0011561 0.21816 0.00065918 0.21882 0.20151 0 0.03305 0.0389 0 1.0824 0.33372 0.097029 0.012835 5.8158 0.080114 9.8786e-005 0.80999 0.0064777 0.007265 0.97 1.3605e-011 0.0073732 0.70945 0.88069 0.14175 0.56487 0.5859 0.59627 0.61149 0.44182 0.31557 0.42847 1.0064 0.99311 15.9957 144.9684 0.00062838 -15.8248 0.017953
3.122 0.98805 5.5056e-005 3.8182 0.012007 4.0957e-005 0.0011561 0.21817 0.00065918 0.21883 0.20152 0 0.033049 0.0389 0 1.0825 0.33377 0.097045 0.012837 5.817 0.080125 9.8801e-005 0.80997 0.0064785 0.0072658 0.95152 3.494e-013 0.0057947 0.6228 0.83076 0.14175 0.55837 0.57902 0.56007 0.59479 0.43985 0.3164 0.42827 1.0079 0.99718 15.9955 144.9677 0.00062918 -20.1377 0.018953
3.123 0.98805 5.5055e-005 3.8182 0.012007 4.097e-005 0.0011561 0.21819 0.00065918 0.21884 0.20154 0 0.033049 0.0389 0 1.0826 0.33381 0.097061 0.012839 5.8182 0.080136 9.8815e-005 0.80996 0.0064792 0.0072665 0.91304 -2.2218e-012 0.0046746 0.50535 0.75333 0.14176 0.55363 0.5747 0.52011 0.57909 0.43866 0.31589 0.42807 1.0098 1.0008 15.9953 144.9672 0.0006289 -25.4178 0.019953
3.124 0.98805 5.5055e-005 3.8182 0.012007 4.0983e-005 0.0011561 0.2182 0.00065918 0.21886 0.20155 0 0.033048 0.0389 0 1.0827 0.33386 0.097077 0.012841 5.8194 0.080147 9.883e-005 0.80995 0.0064799 0.0072673 0.83539 -6.4635e-013 0.0039166 0.35785 0.63763 0.14176 0.55027 0.57238 0.47606 0.56512 0.43802 0.31425 0.42786 1.012 1.004 15.9952 144.9668 0.00062775 -31.3192 0.020953
3.125 0.98805 5.5055e-005 3.8182 0.012007 4.0996e-005 0.0011561 0.21822 0.00065918 0.21887 0.20156 0 0.033047 0.0389 0 1.0828 0.33391 0.097093 0.012842 5.8206 0.080158 9.8845e-005 0.80994 0.0064806 0.0072681 0.70709 -1.7532e-013 0.0034271 0.20449 0.4839 0.14177 0.54785 0.57116 0.42586 0.55437 0.43773 0.3115 0.42766 1.0142 1.0068 15.9951 144.9665 0.00062611 -37.0238 0.021953
3.126 0.98805 5.5055e-005 3.8182 0.012007 4.101e-005 0.0011561 0.21823 0.00065918 0.21888 0.20158 0 0.033047 0.0389 0 1.0829 0.33395 0.09711 0.012844 5.8218 0.080169 9.886e-005 0.80993 0.0064814 0.0072689 0.55221 0.00016301 0.0031604 0.087927 0.31693 0.14178 0.54603 0.57051 0.36705 0.54827 0.43762 0.30741 0.42746 1.0166 1.0095 15.995 144.9662 0.00062429 -41.9044 0.022953
3.127 0.98805 5.5055e-005 3.8182 0.012007 4.1023e-005 0.0011561 0.21824 0.00065918 0.2189 0.20159 0 0.033046 0.0389 0 1.083 0.334 0.097126 0.012846 5.823 0.08018 9.8875e-005 0.80992 0.0064821 0.0072696 0.41099 0.00077363 0.0032304 0.027819 0.17483 0.14178 0.54468 0.57054 0.30032 0.54639 0.43763 0.30162 0.42727 1.0189 1.0121 15.9949 144.966 0.00062242 -45.8823 0.023953
3.128 0.98805 5.5055e-005 3.8182 0.012007 4.1036e-005 0.0011561 0.21826 0.00065918 0.21891 0.2016 0 0.033045 0.0389 0 1.0831 0.33404 0.097142 0.012848 5.8242 0.080191 9.889e-005 0.80991 0.0064828 0.0072704 0.30403 0.0017986 0.0036381 0.0071481 0.080912 0.14179 0.54369 0.57149 0.23082 0.54681 0.4377 0.29387 0.42707 1.0213 1.0147 15.9948 144.9658 0.00062051 -49.0754 0.024953
3.129 0.98805 5.5055e-005 3.8182 0.012007 4.1049e-005 0.0011561 0.21827 0.00065918 0.21892 0.20161 0 0.033044 0.0389 0 1.0832 0.33409 0.097158 0.012849 5.8255 0.080202 9.8905e-005 0.8099 0.0064835 0.0072712 0.23025 0.0033573 0.0043938 0.0021391 0.032317 0.14179 0.54303 0.5732 0.16619 0.54811 0.43779 0.28407 0.42688 1.0237 1.0172 15.9948 144.9657 0.00061858 -51.6237 0.025953
3.13 0.98805 5.5055e-005 3.8182 0.012007 4.1062e-005 0.0011561 0.21828 0.00065918 0.21894 0.20163 0 0.033044 0.0389 0 1.0833 0.33413 0.097174 0.012851 5.8267 0.080213 9.892e-005 0.80989 0.0064842 0.0072719 0.18039 0.0055312 0.0054951 0.0010528 0.012139 0.1418 0.54262 0.57533 0.11287 0.54964 0.43791 0.27236 0.42669 1.0262 1.0196 15.9948 144.9657 0.00061662 -53.6742 0.026953
3.131 0.98805 5.5055e-005 3.8182 0.012007 4.1075e-005 0.0011562 0.2183 0.00065918 0.21895 0.20164 0 0.033043 0.0389 0 1.0834 0.33418 0.09719 0.012853 5.8279 0.080223 9.8934e-005 0.80988 0.006485 0.0072727 0.14578 0.0083736 0.006933 0.00070987 0.0050603 0.14181 0.54243 0.57761 0.073547 0.5512 0.43803 0.259 0.42651 1.0286 1.0221 15.9948 144.9656 0.00061465 -55.3673 0.027953
3.132 0.98805 5.5055e-005 3.8182 0.012007 4.1088e-005 0.0011562 0.21831 0.00065918 0.21896 0.20165 0 0.033042 0.0389 0 1.0835 0.33423 0.097206 0.012855 5.8291 0.080234 9.8949e-005 0.80986 0.0064857 0.0072735 0.12057 0.011928 0.0087004 0.00053162 0.0027315 0.14181 0.54241 0.57993 0.047294 0.5527 0.43816 0.24429 0.42633 1.031 1.0246 15.9947 144.9656 0.00061267 -56.8208 0.028953
3.133 0.98805 5.5055e-005 3.8182 0.012007 4.1101e-005 0.0011562 0.21832 0.00065918 0.21898 0.20167 0 0.033042 0.0389 0 1.0836 0.33427 0.097222 0.012856 5.8303 0.080245 9.8964e-005 0.80985 0.0064864 0.0072742 0.10123 0.016249 0.010798 0.00041541 0.0018626 0.14182 0.54254 0.58224 0.031149 0.55413 0.43829 0.22853 0.42615 1.0334 1.027 15.9947 144.9655 0.00061068 -58.1222 0.029953
3.134 0.98805 5.5055e-005 3.8182 0.012007 4.1114e-005 0.0011562 0.21834 0.00065918 0.21899 0.20168 0 0.033041 0.0389 0 1.0837 0.33432 0.097238 0.012858 5.8315 0.080256 9.8979e-005 0.80984 0.0064871 0.007275 0.085755 0.021411 0.013235 0.00033181 0.0014242 0.14182 0.5428 0.58454 0.021807 0.55551 0.43843 0.21196 0.42598 1.0358 1.0295 15.9947 144.9655 0.00060869 -59.3292 0.030953
3.135 0.98805 5.5055e-005 3.8182 0.012007 4.1127e-005 0.0011562 0.21835 0.00065918 0.21901 0.20169 0 0.03304 0.0389 0 1.0838 0.33436 0.097254 0.01286 5.8327 0.080267 9.8994e-005 0.80983 0.0064879 0.0072758 0.073015 0.02751 0.016032 0.00026939 0.001136 0.14183 0.54317 0.58682 0.016553 0.55681 0.43856 0.19483 0.4258 1.0383 1.0319 15.9947 144.9655 0.00060669 -60.4764 0.031953
3.136 0.98805 5.5055e-005 3.8182 0.012007 4.114e-005 0.0011562 0.21836 0.00065918 0.21902 0.2017 0 0.03304 0.0389 0 1.0839 0.33441 0.097271 0.012862 5.8339 0.080278 9.9009e-005 0.80982 0.0064886 0.0072765 0.062357 0.034665 0.019213 0.00022012 0.00092144 0.14183 0.54365 0.58908 0.013536 0.55807 0.4387 0.17737 0.42563 1.0407 1.0343 15.9948 144.9654 0.00060469 -61.5828 0.032953
3.137 0.98805 5.5054e-005 3.8182 0.012007 4.1153e-005 0.0011562 0.21838 0.00065918 0.21903 0.20172 0 0.033039 0.0389 0 1.084 0.33445 0.097287 0.012863 5.8351 0.080289 9.9024e-005 0.80981 0.0064893 0.0072773 0.053367 0.043015 0.022809 0.00018121 0.00075418 0.14184 0.54422 0.59132 0.011656 0.55927 0.43884 0.15982 0.42547 1.0431 1.0368 15.9948 144.9654 0.00060268 -62.6581 0.033953
3.138 0.98805 5.5054e-005 3.8182 0.012007 4.1166e-005 0.0011562 0.21839 0.00065918 0.21905 0.20173 0 0.033038 0.0389 0 1.0841 0.3345 0.097303 0.012865 5.8364 0.0803 9.9038e-005 0.8098 0.00649 0.0072781 0.045755 0.05271 0.026855 0.00014999 0.00062132 0.14185 0.54488 0.59354 0.010336 0.56043 0.43898 0.14243 0.42531 1.0455 1.0392 15.9948 144.9654 0.00060067 -63.7069 0.034953
3.139 0.98805 5.5054e-005 3.8182 0.012007 4.1179e-005 0.0011562 0.2184 0.00065918 0.21906 0.20174 0 0.033037 0.0389 0 1.0842 0.33455 0.097319 0.012867 5.8376 0.080311 9.9053e-005 0.80979 0.0064908 0.0072788 0.039298 0.063911 0.031389 0.00012468 0.00051469 0.14185 0.54561 0.59573 0.0093037 0.56155 0.43912 0.12543 0.42515 1.0479 1.0416 15.9948 144.9654 0.00059866 -64.7313 0.035953
3.14 0.98805 5.5054e-005 3.8182 0.012007 4.1192e-005 0.0011562 0.21842 0.00065918 0.21907 0.20175 0 0.033037 0.0389 0 1.0843 0.33459 0.097335 0.012869 5.8388 0.080322 9.9068e-005 0.80978 0.0064915 0.0072796 0.033817 0.076786 0.036452 0.00010416 0.00042851 0.14186 0.54641 0.59791 0.0084392 0.56265 0.43926 0.10909 0.425 1.0503 1.0441 15.9948 144.9653 0.00059665 -65.7324 0.036953
3.141 0.98805 5.5054e-005 3.8182 0.012007 4.1205e-005 0.0011562 0.21843 0.00065918 0.21909 0.20177 0 0.033036 0.0389 0 1.0844 0.33464 0.097351 0.01287 5.84 0.080333 9.9083e-005 0.80977 0.0064922 0.0072804 0.02916 0.091505 0.042091 8.7382e-005 0.00035848 0.14186 0.54727 0.60006 0.00769 0.56373 0.4394 0.093639 0.42485 1.0527 1.0465 15.9949 144.9653 0.00059464 -66.7103 0.037953
3.142 0.98805 5.5054e-005 3.8182 0.012007 4.1218e-005 0.0011562 0.21844 0.00065918 0.2191 0.20178 0 0.033035 0.0389 0 1.0845 0.33468 0.097367 0.012872 5.8412 0.080344 9.9098e-005 0.80975 0.0064929 0.0072811 0.025202 0.10823 0.048356 7.3635e-005 0.00030132 0.14187 0.54819 0.60219 0.0070313 0.56479 0.43954 0.079277 0.4247 1.0551 1.0489 15.9949 144.9653 0.00059263 -67.6651 0.038953
3.143 0.98805 5.5054e-005 3.8182 0.012007 4.1231e-005 0.0011562 0.21846 0.00065918 0.21911 0.20179 0 0.033035 0.0389 0 1.0846 0.33473 0.097383 0.012874 5.8424 0.080355 9.9113e-005 0.80974 0.0064936 0.0072819 0.021837 0.12712 0.055301 6.2319e-005 0.00025446 0.14188 0.54915 0.60431 0.0064483 0.56584 0.43968 0.06618 0.42456 1.0575 1.0513 15.995 144.9653 0.00059061 -68.5962 0.039953
3.144 0.98805 5.5054e-005 3.8182 0.012007 4.1244e-005 0.0011562 0.21847 0.00065918 0.21913 0.20181 0 0.033034 0.0389 0 1.0847 0.33477 0.097399 0.012876 5.8437 0.080366 9.9128e-005 0.80973 0.0064944 0.0072827 0.018973 0.14831 0.06299 5.2986e-005 0.0002159 0.14188 0.55016 0.6064 0.0059304 0.56689 0.43982 0.054471 0.42443 1.0599 1.0537 15.995 144.9652 0.0005886 -69.5031 0.040953
3.145 0.98805 5.5054e-005 3.8182 0.012007 4.1257e-005 0.0011562 0.21848 0.00065918 0.21914 0.20182 0 0.033033 0.0389 0 1.0848 0.33482 0.097415 0.012877 5.8449 0.080377 9.9142e-005 0.80972 0.0064951 0.0072835 0.016535 0.17191 0.071489 4.5255e-005 0.00018408 0.14189 0.5512 0.60847 0.0054692 0.56795 0.43996 0.04422 0.4243 1.0623 1.0561 15.9951 144.9652 0.00058658 -70.3847 0.041953
3.146 0.98805 5.5054e-005 3.8182 0.012007 4.127e-005 0.0011562 0.2185 0.00065918 0.21915 0.20183 0 0.033033 0.0389 0 1.0849 0.33487 0.097432 0.012879 5.8461 0.080388 9.9157e-005 0.80971 0.0064958 0.0072842 0.014459 0.19798 0.080871 3.8841e-005 0.00015774 0.14189 0.55228 0.61052 0.005058 0.56901 0.44011 0.03544 0.42418 1.0647 1.0586 15.9951 144.9652 0.00058457 -71.24 0.042953
3.147 0.98805 5.5054e-005 3.8182 0.012007 4.1284e-005 0.0011562 0.21851 0.00065918 0.21917 0.20184 0 0.033032 0.0389 0 1.0849 0.33491 0.097448 0.012881 5.8473 0.080399 9.9172e-005 0.8097 0.0064965 0.007285 0.01269 0.22655 0.091215 3.3505e-005 0.00013586 0.1419 0.55338 0.61255 0.0046909 0.57008 0.44025 0.028091 0.42406 1.0671 1.061 15.9952 144.9651 0.00058256 -72.0676 0.043953
3.148 0.98805 5.5054e-005 3.8182 0.012007 4.1297e-005 0.0011562 0.21853 0.00065918 0.21918 0.20186 0 0.033031 0.0389 0 1.085 0.33496 0.097464 0.012883 5.8485 0.08041 9.9187e-005 0.80969 0.0064973 0.0072858 0.011182 0.25756 0.1026 2.9053e-005 0.00011766 0.14191 0.55451 0.61457 0.0043631 0.57117 0.4404 0.022081 0.42395 1.0695 1.0634 15.9952 144.9651 0.00058055 -72.8661 0.044953
3.149 0.98805 5.5054e-005 3.8182 0.012007 4.131e-005 0.0011562 0.21854 0.00065918 0.21919 0.20187 0 0.03303 0.0389 0 1.0851 0.335 0.09748 0.012884 5.8497 0.080421 9.9202e-005 0.80968 0.006498 0.0072865 0.0098956 0.29091 0.1151 2.5333e-005 0.00010247 0.14191 0.55566 0.61656 0.0040702 0.57229 0.44054 0.017282 0.42384 1.0719 1.0658 15.9953 144.9651 0.00057854 -73.6342 0.045953
3.15 0.98805 5.5054e-005 3.8182 0.012006 4.1323e-005 0.0011562 0.21855 0.00065918 0.21921 0.20188 0 0.03303 0.0389 0 1.0852 0.33505 0.097496 0.012886 5.851 0.080432 9.9217e-005 0.80967 0.0064987 0.0072873 0.0087976 0.32639 0.12878 2.2217e-005 8.9763e-005 0.14192 0.55683 0.61853 0.0038086 0.57343 0.44069 0.013539 0.42374 1.0742 1.0682 15.9954 144.9651 0.00057654 -74.3703 0.046953
3.151 0.98805 5.5054e-005 3.8182 0.012006 4.1336e-005 0.0011562 0.21857 0.00065918 0.21922 0.20189 0 0.033029 0.0389 0 1.0853 0.33509 0.097512 0.012888 5.8522 0.080443 9.9232e-005 0.80966 0.0064994 0.0072881 0.0078599 0.36375 0.1437 1.9599e-005 7.9111e-005 0.14192 0.55801 0.62049 0.0035749 0.5746 0.44084 0.010685 0.42365 1.0766 1.0706 15.9954 144.965 0.00057453 -75.0733 0.047953
3.152 0.98805 5.5053e-005 3.8182 0.012006 4.1349e-005 0.0011562 0.21858 0.00065918 0.21923 0.20191 0 0.033028 0.0389 0 1.0854 0.33514 0.097528 0.01289 5.8534 0.080454 9.9246e-005 0.80965 0.0065002 0.0072888 0.0070585 0.40263 0.15989 1.7397e-005 7.0157e-005 0.14193 0.55921 0.62242 0.0033664 0.57581 0.44099 0.0085543 0.42356 1.079 1.073 15.9955 144.965 0.00057253 -75.742 0.048953
3.153 0.98805 5.5053e-005 3.8182 0.012006 4.1362e-005 0.0011562 0.21859 0.00065918 0.21925 0.20192 0 0.033028 0.0389 0 1.0855 0.33519 0.097544 0.012891 5.8546 0.080465 9.9261e-005 0.80963 0.0065009 0.0072896 0.0063726 0.44261 0.17735 1.5542e-005 6.2614e-005 0.14193 0.56041 0.62434 0.0031803 0.57705 0.44115 0.0069917 0.42347 1.0814 1.0754 15.9956 144.965 0.00057054 -76.3755 0.049953
3.154 0.98805 5.5053e-005 3.8182 0.012006 4.1375e-005 0.0011562 0.2186 0.00065918 0.21926 0.20193 0 0.033027 0.0389 0 1.0856 0.33523 0.09756 0.012893 5.8558 0.080476 9.9276e-005 0.80962 0.0065016 0.0072904 0.0057849 0.48323 0.19605 1.3969e-005 5.6248e-005 0.14194 0.56163 0.62624 0.0030144 0.57833 0.4413 0.005862 0.4234 1.0837 1.0777 15.9957 144.9649 0.00056855 -76.9734 0.050953
3.155 0.98806 5.5053e-005 3.8182 0.012006 4.1388e-005 0.0011562 0.21862 0.00065918 0.21927 0.20194 0 0.033026 0.0389 0 1.0857 0.33528 0.097576 0.012895 5.8571 0.080487 9.9291e-005 0.80961 0.0065023 0.0072911 0.0052809 0.52398 0.21592 1.2638e-005 5.0857e-005 0.14195 0.56285 0.62812 0.0028666 0.57965 0.44146 0.0050519 0.42332 1.0861 1.0801 15.9958 144.9649 0.00056656 -77.5355 0.051953
3.156 0.98806 5.5053e-005 3.8182 0.012006 4.1401e-005 0.0011562 0.21863 0.00065918 0.21929 0.20196 0 0.033026 0.0389 0 1.0858 0.33532 0.097593 0.012897 5.8583 0.080498 9.9306e-005 0.8096 0.006503 0.0072919 0.0048479 0.56435 0.23687 1.1507e-005 4.628e-005 0.14195 0.56408 0.62998 0.0027349 0.58101 0.44161 0.004471 0.42325 1.0885 1.0825 15.9958 144.9649 0.00056458 -78.0617 0.052953
3.157 0.98806 5.5053e-005 3.8182 0.012006 4.1414e-005 0.0011562 0.21864 0.00065918 0.2193 0.20197 0 0.033025 0.0389 0 1.0859 0.33537 0.097609 0.012898 5.8595 0.080509 9.9321e-005 0.80959 0.0065038 0.0072927 0.004476 0.60384 0.25877 1.055e-005 4.2378e-005 0.14196 0.56531 0.63183 0.0026176 0.58241 0.44177 0.0040509 0.42319 1.0908 1.0849 15.9959 144.9649 0.0005626 -78.5526 0.053953
3.158 0.98806 5.5053e-005 3.8182 0.012006 4.1427e-005 0.0011562 0.21866 0.00065918 0.21931 0.20198 0 0.033024 0.0389 0 1.086 0.33541 0.097625 0.0129 5.8607 0.080519 9.9336e-005 0.80958 0.0065045 0.0072934 0.0041541 0.64198 0.28148 9.7218e-006 3.9057e-005 0.14196 0.56655 0.63366 0.0025132 0.58385 0.44193 0.0037418 0.42313 1.0932 1.0873 15.996 144.9649 0.00056063 -79.009 0.054953
3.159 0.98806 5.5053e-005 3.8182 0.012006 4.144e-005 0.0011562 0.21867 0.00065918 0.21933 0.20199 0 0.033024 0.0389 0 1.0861 0.33546 0.097641 0.012902 5.8619 0.08053 9.935e-005 0.80957 0.0065052 0.0072942 0.0038766 0.67837 0.30484 9.018e-006 3.6209e-005 0.14197 0.56779 0.63547 0.0024202 0.58534 0.44209 0.0035084 0.42308 1.0955 1.0896 15.9961 144.9648 0.00055867 -79.4317 0.055953
3.16 0.98806 5.5053e-005 3.8182 0.012006 4.1453e-005 0.0011562 0.21868 0.00065918 0.21934 0.20201 0 0.033023 0.0389 0 1.0862 0.33551 0.097657 0.012904 5.8632 0.080541 9.9365e-005 0.80956 0.0065059 0.007295 0.0036371 0.71267 0.32868 8.413e-006 3.3765e-005 0.14198 0.56903 0.63726 0.0023375 0.58687 0.44226 0.0033268 0.42303 1.0979 1.092 15.9962 144.9648 0.00055671 -79.8222 0.056953
3.161 0.98806 5.5053e-005 3.8182 0.012006 4.1466e-005 0.0011562 0.2187 0.00065918 0.21935 0.20202 0 0.033022 0.0389 0 1.0863 0.33555 0.097673 0.012906 5.8644 0.080552 9.938e-005 0.80955 0.0065067 0.0072958 0.0034284 0.74461 0.35284 7.8914e-006 3.1662e-005 0.14198 0.57028 0.63904 0.0022639 0.58843 0.44242 0.0031814 0.42298 1.1002 1.0944 15.9963 144.9648 0.00055477 -80.1817 0.057953
3.162 0.98806 5.5053e-005 3.8182 0.012006 4.1479e-005 0.0011562 0.21871 0.00065918 0.21937 0.20203 0 0.033021 0.0389 0 1.0864 0.3356 0.097689 0.012907 5.8656 0.080563 9.9395e-005 0.80954 0.0065074 0.0072965 0.0032475 0.77404 0.37715 7.4412e-006 2.9845e-005 0.14199 0.57152 0.6408 0.0021984 0.59003 0.44259 0.0030616 0.42294 1.1026 1.0967 15.9964 144.9648 0.00055282 -80.512 0.058953
3.163 0.98806 5.5053e-005 3.8182 0.012006 4.1492e-005 0.0011562 0.21872 0.00065918 0.21938 0.20204 0 0.033021 0.0389 0 1.0865 0.33564 0.097705 0.012909 5.8668 0.080574 9.941e-005 0.80953 0.0065081 0.0072973 0.0030901 0.80085 0.40147 7.0513e-006 2.8273e-005 0.14199 0.57276 0.64255 0.00214 0.59167 0.44276 0.0029608 0.4229 1.1049 1.0991 15.9965 144.9648 0.00055089 -80.8147 0.059953
3.164 0.98806 5.5053e-005 3.8182 0.012006 4.1505e-005 0.0011562 0.21874 0.00065918 0.21939 0.20206 0 0.03302 0.0389 0 1.0866 0.33569 0.097721 0.012911 5.8681 0.080585 9.9425e-005 0.80951 0.0065088 0.0072981 0.0029524 0.82503 0.42564 6.7126e-006 2.6909e-005 0.142 0.57401 0.64428 0.0020881 0.59335 0.44292 0.0028745 0.42286 1.1072 1.1014 15.9966 144.9648 0.00054897 -81.0915 0.060953
3.165 0.98806 5.5053e-005 3.8182 0.012006 4.1518e-005 0.0011562 0.21875 0.00065918 0.21941 0.20207 0 0.033019 0.0389 0 1.0867 0.33573 0.097737 0.012913 5.8693 0.080596 9.944e-005 0.8095 0.0065096 0.0072988 0.0028322 0.84664 0.44956 6.4177e-006 2.572e-005 0.14201 0.57525 0.64599 0.0020417 0.59505 0.44309 0.0027998 0.42283 1.1096 1.1038 15.9967 144.9648 0.00054705 -81.3441 0.061953
3.166 0.98806 5.5052e-005 3.8182 0.012006 4.1531e-005 0.0011562 0.21876 0.00065918 0.21942 0.20208 0 0.033019 0.0389 0 1.0868 0.33578 0.097754 0.012914 5.8705 0.080607 9.9454e-005 0.80949 0.0065103 0.0072996 0.0027266 0.86577 0.47311 6.1602e-006 2.4683e-005 0.14201 0.57649 0.64769 0.0020004 0.59678 0.44326 0.0027345 0.4228 1.1119 1.1061 15.9968 144.9648 0.00054514 -81.5744 0.062953
3.167 0.98806 5.5052e-005 3.8182 0.012006 4.1545e-005 0.0011562 0.21878 0.00065918 0.21943 0.20209 0 0.033018 0.0389 0 1.0869 0.33583 0.09777 0.012916 5.8717 0.080618 9.9469e-005 0.80948 0.006511 0.0073004 0.0026341 0.88258 0.49621 5.9349e-006 2.3776e-005 0.14202 0.57773 0.64938 0.0019636 0.59854 0.44344 0.0026771 0.42277 1.1142 1.1085 15.9969 144.9648 0.00054324 -81.784 0.063953
3.168 0.98806 5.5052e-005 3.8182 0.012006 4.1558e-005 0.0011562 0.21879 0.00065918 0.21944 0.20211 0 0.033017 0.0389 0 1.087 0.33587 0.097786 0.012918 5.873 0.080629 9.9484e-005 0.80947 0.0065117 0.0073011 0.0025523 0.89722 0.51876 5.7371e-006 2.298e-005 0.14202 0.57897 0.65104 0.0019307 0.60032 0.44361 0.0026264 0.42274 1.1165 1.1108 15.997 144.9648 0.00054135 -81.9746 0.064953
3.169 0.98806 5.5052e-005 3.8182 0.012006 4.1571e-005 0.0011562 0.2188 0.00065918 0.21946 0.20212 0 0.033017 0.0389 0 1.0871 0.33592 0.097802 0.01292 5.8742 0.08064 9.9499e-005 0.80946 0.0065125 0.0073019 0.0024805 0.9099 0.54072 5.5632e-006 2.228e-005 0.14203 0.58021 0.6527 0.0019012 0.60213 0.44378 0.0025816 0.42272 1.1189 1.1132 15.9971 144.9648 0.00053947 -82.1479 0.065953
3.17 0.98806 5.5052e-005 3.8182 0.012006 4.1584e-005 0.0011562 0.21882 0.00065918 0.21947 0.20213 0 0.033016 0.0389 0 1.0872 0.33596 0.097818 0.012921 5.8754 0.080651 9.9514e-005 0.80945 0.0065132 0.0073027 0.0024169 0.92081 0.56202 5.4098e-006 2.1663e-005 0.14203 0.58144 0.65434 0.0018749 0.60395 0.44396 0.0025418 0.4227 1.1212 1.1155 15.9972 144.9647 0.00053759 -82.3052 0.066953
3.171 0.98806 5.5052e-005 3.8182 0.012006 4.1597e-005 0.0011562 0.21883 0.00065918 0.21948 0.20214 0 0.033015 0.0389 0 1.0873 0.33601 0.097834 0.012923 5.8766 0.080662 9.9529e-005 0.80944 0.0065139 0.0073034 0.0023605 0.93014 0.58265 5.2743e-006 2.1118e-005 0.14204 0.58267 0.65596 0.0018514 0.60579 0.44413 0.0025064 0.42267 1.1235 1.1178 15.9972 144.9647 0.00053573 -82.448 0.067953
3.172 0.98806 5.5052e-005 3.8182 0.012006 4.161e-005 0.0011562 0.21884 0.00065918 0.2195 0.20216 0 0.033015 0.0389 0 1.0874 0.33605 0.09785 0.012925 5.8779 0.080673 9.9544e-005 0.80943 0.0065146 0.0073042 0.0023104 0.93808 0.60255 5.1541e-006 2.0635e-005 0.14205 0.5839 0.65757 0.0018302 0.60765 0.44431 0.0024748 0.42265 1.1258 1.1202 15.9973 144.9647 0.00053388 -82.5776 0.068953
3.173 0.98806 5.5052e-005 3.8182 0.012006 4.1623e-005 0.0011562 0.21886 0.00065918 0.21951 0.20217 0 0.033014 0.0389 0 1.0875 0.3361 0.097866 0.012927 5.8791 0.080684 9.9558e-005 0.80942 0.0065153 0.007305 0.0022658 0.94481 0.62173 5.0475e-006 2.0206e-005 0.14205 0.58513 0.65917 0.0018112 0.60952 0.44448 0.0024466 0.42264 1.1281 1.1225 15.9974 144.9647 0.00053203 -82.6953 0.069953
3.174 0.98806 5.5052e-005 3.8182 0.012006 4.1636e-005 0.0011562 0.21887 0.00065919 0.21952 0.20218 0 0.033013 0.0389 0 1.0876 0.33615 0.097882 0.012928 5.8803 0.080695 9.9573e-005 0.8094 0.0065161 0.0073058 0.0022261 0.95049 0.64017 4.9525e-006 1.9824e-005 0.14206 0.58635 0.66075 0.0017942 0.6114 0.44466 0.0024214 0.42262 1.1304 1.1248 15.9975 144.9647 0.0005302 -82.8022 0.070953
3.175 0.98806 5.5052e-005 3.8182 0.012006 4.1649e-005 0.0011562 0.21888 0.00065919 0.21954 0.20219 0 0.033013 0.0389 0 1.0877 0.33619 0.097899 0.01293 5.8816 0.080706 9.9588e-005 0.80939 0.0065168 0.0073065 0.0021905 0.95528 0.65786 4.8677e-006 1.9483e-005 0.14206 0.58757 0.66232 0.0017788 0.61329 0.44483 0.0023988 0.4226 1.1327 1.1271 15.9976 144.9647 0.00052837 -82.8994 0.071953
3.176 0.98806 5.5052e-005 3.8182 0.012006 4.1662e-005 0.0011562 0.21889 0.00065919 0.21955 0.20221 0 0.033012 0.0389 0 1.0878 0.33624 0.097915 0.012932 5.8828 0.080717 9.9603e-005 0.80938 0.0065175 0.0073073 0.0021587 0.95929 0.67481 4.7919e-006 1.9179e-005 0.14207 0.58879 0.66387 0.001765 0.61518 0.44501 0.0023785 0.42259 1.135 1.1294 15.9977 144.9647 0.00052656 -82.9878 0.072953
3.177 0.98806 5.5052e-005 3.8182 0.012006 4.1675e-005 0.0011562 0.21891 0.00065919 0.21956 0.20222 0 0.033011 0.0389 0 1.0879 0.33628 0.097931 0.012934 5.884 0.080727 9.9618e-005 0.80937 0.0065182 0.0073081 0.0021301 0.96266 0.69103 4.7238e-006 1.8905e-005 0.14208 0.59 0.66541 0.0017525 0.61709 0.44519 0.0023602 0.42257 1.1373 1.1317 15.9978 144.9647 0.00052475 -83.0683 0.073953
3.178 0.98806 5.5052e-005 3.8182 0.012006 4.1688e-005 0.0011562 0.21892 0.00065919 0.21958 0.20223 0 0.033011 0.0389 0 1.088 0.33633 0.097947 0.012935 5.8852 0.080738 9.9633e-005 0.80936 0.006519 0.0073088 0.0021043 0.96547 0.70653 4.6626e-006 1.8659e-005 0.14208 0.59121 0.66694 0.0017411 0.61899 0.44537 0.0023438 0.42256 1.1396 1.134 15.9979 144.9647 0.00052295 -83.1417 0.074953
3.179 0.98806 5.5052e-005 3.8182 0.012006 4.1701e-005 0.0011562 0.21893 0.00065919 0.21959 0.20224 0 0.03301 0.0389 0 1.0881 0.33638 0.097963 0.012937 5.8865 0.080749 9.9647e-005 0.80935 0.0065197 0.0073096 0.0020811 0.96783 0.72132 4.6074e-006 1.8438e-005 0.14209 0.59242 0.66845 0.0017308 0.6209 0.44555 0.0023289 0.42255 1.1419 1.1364 15.998 144.9648 0.00052117 -83.2087 0.075953
3.18 0.98806 5.5052e-005 3.8182 0.012006 4.1714e-005 0.0011562 0.21895 0.00065919 0.2196 0.20226 0 0.033009 0.0389 0 1.0882 0.33642 0.097979 0.012939 5.8877 0.08076 9.9662e-005 0.80934 0.0065204 0.0073104 0.0020602 0.9698 0.73543 4.5577e-006 1.8238e-005 0.14209 0.59363 0.66996 0.0017215 0.62282 0.44572 0.0023154 0.42254 1.1441 1.1387 15.9981 144.9648 0.00051939 -83.27 0.076953
3.181 0.98806 5.5051e-005 3.8182 0.012006 4.1727e-005 0.0011562 0.21896 0.00065919 0.21961 0.20227 0 0.033009 0.0389 0 1.0883 0.33647 0.097995 0.012941 5.8889 0.080771 9.9677e-005 0.80933 0.0065211 0.0073111 0.002041 0.97144 0.74887 4.5124e-006 1.8056e-005 0.1421 0.59483 0.67144 0.001713 0.62473 0.4459 0.0023032 0.42253 1.1464 1.1409 15.9982 144.9648 0.00051762 -83.3262 0.077953
3.182 0.98806 5.5051e-005 3.8182 0.012006 4.174e-005 0.0011562 0.21897 0.00065919 0.21963 0.20228 0 0.033008 0.0389 0 1.0884 0.33651 0.098011 0.012942 5.8902 0.080782 9.9692e-005 0.80932 0.0065219 0.0073119 0.0020232 0.97282 0.76166 4.471e-006 1.789e-005 0.1421 0.59603 0.67292 0.0017052 0.62664 0.44608 0.0022921 0.42252 1.1487 1.1432 15.9983 144.9648 0.00051586 -83.3777 0.078953
3.183 0.98806 5.5051e-005 3.8182 0.012006 4.1753e-005 0.0011562 0.21899 0.00065919 0.21964 0.20229 0 0.033007 0.0389 0 1.0885 0.33656 0.098027 0.012944 5.8914 0.080793 9.9707e-005 0.80931 0.0065226 0.0073127 0.0020074 0.97398 0.77383 4.4337e-006 1.774e-005 0.14211 0.59722 0.67438 0.0016981 0.62856 0.44626 0.0022819 0.42251 1.151 1.1455 15.9984 144.9648 0.00051411 -83.4251 0.079953
3.184 0.98806 5.5051e-005 3.8182 0.012006 4.1766e-005 0.0011562 0.219 0.00065919 0.21965 0.20231 0 0.033007 0.0389 0 1.0886 0.3366 0.098043 0.012946 5.8926 0.080804 9.9722e-005 0.8093 0.0065233 0.0073135 0.0019933 0.97494 0.78539 4.3996e-006 1.7603e-005 0.14212 0.59842 0.67584 0.0016916 0.63047 0.44644 0.0022726 0.4225 1.1532 1.1478 15.9985 144.9648 0.00051237 -83.4689 0.080953
3.185 0.98806 5.5051e-005 3.8182 0.012006 4.1779e-005 0.0011562 0.21901 0.00065919 0.21967 0.20232 0 0.033006 0.0389 0 1.0887 0.33665 0.09806 0.012948 5.8939 0.080815 9.9737e-005 0.80928 0.006524 0.0073142 0.0019802 0.97576 0.79638 4.3682e-006 1.7477e-005 0.14212 0.5996 0.67727 0.0016855 0.63238 0.44662 0.0022641 0.42249 1.1555 1.1501 15.9986 144.9648 0.00051064 -83.5093 0.081953
3.186 0.98806 5.5051e-005 3.8182 0.012006 4.1792e-005 0.0011562 0.21902 0.00065919 0.21968 0.20233 0 0.033005 0.0389 0 1.0888 0.3367 0.098076 0.012949 5.8951 0.080826 9.9751e-005 0.80927 0.0065248 0.007315 0.0019679 0.97644 0.80681 4.3392e-006 1.7361e-005 0.14213 0.60079 0.6787 0.00168 0.63429 0.4468 0.0022563 0.42248 1.1578 1.1524 15.9987 144.9648 0.00050892 -83.5468 0.082953
3.187 0.98806 5.5051e-005 3.8182 0.012006 4.1805e-005 0.0011562 0.21904 0.00065919 0.21969 0.20234 0 0.033005 0.0389 0 1.0889 0.33674 0.098092 0.012951 5.8963 0.080837 9.9766e-005 0.80926 0.0065255 0.0073158 0.0019562 0.97702 0.81671 4.3123e-006 1.7253e-005 0.14213 0.60197 0.68012 0.0016748 0.63619 0.44698 0.0022491 0.42247 1.16 1.1546 15.9988 144.9648 0.00050721 -83.5817 0.083953
3.188 0.98806 5.5051e-005 3.8182 0.012006 4.1819e-005 0.0011562 0.21905 0.00065919 0.2197 0.20235 0 0.033004 0.0389 0 1.089 0.33679 0.098108 0.012953 5.8976 0.080848 9.9781e-005 0.80925 0.0065262 0.0073165 0.0019455 0.97752 0.8261 4.2875e-006 1.7153e-005 0.14214 0.60315 0.68152 0.00167 0.63809 0.44716 0.0022424 0.42246 1.1623 1.1569 15.9989 144.9648 0.00050551 -83.6142 0.084953
3.189 0.98806 5.5051e-005 3.8182 0.012006 4.1832e-005 0.0011562 0.21906 0.00065919 0.21972 0.20237 0 0.033003 0.0389 0 1.0891 0.33683 0.098124 0.012955 5.8988 0.080859 9.9796e-005 0.80924 0.0065269 0.0073173 0.0019358 0.97794 0.835 4.2645e-006 1.7061e-005 0.14215 0.60433 0.68291 0.0016656 0.63999 0.44734 0.0022361 0.42246 1.1645 1.1592 15.999 144.9648 0.00050382 -83.6445 0.085953
3.19 0.98806 5.5051e-005 3.8182 0.012006 4.1845e-005 0.0011563 0.21908 0.00065919 0.21973 0.20238 0 0.033002 0.0389 0 1.0892 0.33688 0.09814 0.012956 5.9 0.08087 9.9811e-005 0.80923 0.0065276 0.0073181 0.0019268 0.97831 0.84344 4.2431e-006 1.6975e-005 0.14215 0.6055 0.68429 0.0016614 0.64188 0.44752 0.0022303 0.42245 1.1668 1.1614 15.999 144.9648 0.00050214 -83.673 0.086953
3.191 0.98806 5.5051e-005 3.8182 0.012006 4.1858e-005 0.0011563 0.21909 0.00065919 0.21974 0.20239 0 0.033002 0.0389 0 1.0893 0.33692 0.098156 0.012958 5.9013 0.080881 9.9826e-005 0.80922 0.0065284 0.0073188 0.0019186 0.97862 0.85143 4.2231e-006 1.6895e-005 0.14216 0.60666 0.68566 0.0016575 0.64377 0.4477 0.0022249 0.42244 1.169 1.1637 15.9991 144.9648 0.00050046 -83.6998 0.087953
3.192 0.98806 5.5051e-005 3.8182 0.012006 4.1871e-005 0.0011563 0.2191 0.00065919 0.21976 0.2024 0 0.033001 0.0389 0 1.0894 0.33697 0.098172 0.01296 5.9025 0.080892 9.984e-005 0.80921 0.0065291 0.0073196 0.0019107 0.97889 0.859 4.2042e-006 1.6819e-005 0.14216 0.60783 0.68702 0.0016538 0.64565 0.44788 0.0022198 0.42244 1.1712 1.166 15.9992 144.9648 0.0004988 -83.7251 0.088953
3.193 0.98806 5.5051e-005 3.8182 0.012006 4.1884e-005 0.0011563 0.21911 0.00065919 0.21977 0.20242 0 0.033 0.0389 0 1.0895 0.33702 0.098188 0.012962 5.9037 0.080902 9.9855e-005 0.8092 0.0065298 0.0073204 0.0019028 0.97913 0.86618 4.1863e-006 1.6748e-005 0.14217 0.60899 0.68836 0.0016503 0.64753 0.44806 0.0022151 0.42243 1.1735 1.1682 15.9993 144.9648 0.00049714 -83.749 0.089953
3.194 0.98806 5.5051e-005 3.8182 0.012006 4.1897e-005 0.0011563 0.21913 0.00065919 0.21978 0.20243 0 0.033 0.0389 0 1.0896 0.33706 0.098205 0.012963 5.905 0.080913 9.987e-005 0.80919 0.0065305 0.0073211 0.0018955 0.97934 0.87296 4.1694e-006 1.668e-005 0.14218 0.61015 0.6897 0.001647 0.6494 0.44824 0.0022106 0.42242 1.1757 1.1705 15.9994 144.9648 0.0004955 -83.7717 0.090953
3.195 0.98806 5.5051e-005 3.8182 0.012006 4.191e-005 0.0011563 0.21914 0.00065919 0.2198 0.20244 0 0.032999 0.0389 0 1.0897 0.33711 0.098221 0.012965 5.9062 0.080924 9.9885e-005 0.80918 0.0065313 0.0073219 0.0018886 0.97953 0.87939 4.1535e-006 1.6616e-005 0.14218 0.6113 0.69102 0.0016439 0.65127 0.44843 0.0022063 0.42242 1.1779 1.1727 15.9995 144.9648 0.00049386 -83.7933 0.091953
3.196 0.98806 5.505e-005 3.8182 0.012006 4.1923e-005 0.0011563 0.21915 0.00065919 0.21981 0.20245 0 0.032998 0.0389 0 1.0898 0.33715 0.098237 0.012967 5.9074 0.080935 9.99e-005 0.80916 0.006532 0.0073227 0.0018821 0.9797 0.88547 4.1384e-006 1.6555e-005 0.14219 0.61245 0.69234 0.0016409 0.65313 0.44861 0.0022023 0.42241 1.1801 1.1749 15.9996 144.9648 0.00049223 -83.8139 0.092953
3.197 0.98806 5.505e-005 3.8182 0.012006 4.1936e-005 0.0011563 0.21917 0.00065919 0.21982 0.20246 0 0.032998 0.0389 0 1.0899 0.3372 0.098253 0.012969 5.9087 0.080946 9.9915e-005 0.80915 0.0065327 0.0073235 0.0018763 0.97985 0.89122 4.124e-006 1.6498e-005 0.14219 0.6136 0.69364 0.0016381 0.65498 0.44879 0.0021984 0.42241 1.1824 1.1772 15.9997 144.9648 0.00049061 -83.8337 0.093953
3.198 0.98806 5.505e-005 3.8182 0.012006 4.1949e-005 0.0011563 0.21918 0.00065919 0.21983 0.20248 0 0.032997 0.0389 0 1.09 0.33725 0.098269 0.01297 5.9099 0.080957 9.9929e-005 0.80914 0.0065334 0.0073242 0.0018706 0.97998 0.89666 4.1102e-006 1.6443e-005 0.1422 0.61475 0.69493 0.0016354 0.65683 0.44897 0.0021947 0.4224 1.1846 1.1794 15.9998 144.9649 0.000489 -83.8526 0.094953
3.199 0.98806 5.505e-005 3.8182 0.012006 4.1962e-005 0.0011563 0.21919 0.00065919 0.21985 0.20249 0 0.032996 0.0389 0 1.0901 0.33729 0.098285 0.012972 5.9112 0.080968 9.9944e-005 0.80913 0.0065342 0.007325 0.0018649 0.98011 0.90181 4.0969e-006 1.6389e-005 0.1422 0.61589 0.69622 0.0016328 0.65867 0.44915 0.0021912 0.4224 1.1868 1.1816 15.9998 144.9649 0.0004874 -83.8708 0.095953
3.2 0.98806 5.505e-005 3.8182 0.012006 4.1975e-005 0.0011563 0.2192 0.00065919 0.21986 0.2025 0 0.032996 0.0389 0 1.0902 0.33734 0.098301 0.012974 5.9124 0.080979 9.9959e-005 0.80912 0.0065349 0.0073258 0.0018594 0.98022 0.90667 4.0842e-006 1.6338e-005 0.14221 0.61702 0.69749 0.0016303 0.6605 0.44933 0.0021878 0.42239 1.189 1.1839 15.9999 144.9649 0.00048581 -83.8884 0.096953
3.201 0.98806 5.505e-005 3.8182 0.012006 4.1988e-005 0.0011563 0.21922 0.00065919 0.21987 0.20251 0 0.032995 0.0389 0 1.0903 0.33738 0.098317 0.012976 5.9136 0.08099 9.9974e-005 0.80911 0.0065356 0.0073265 0.001854 0.98033 0.91127 4.0718e-006 1.6289e-005 0.14222 0.61816 0.69875 0.0016278 0.66233 0.44951 0.0021845 0.42239 1.1912 1.1861 16 144.9649 0.00048423 -83.9054 0.097953
3.202 0.98806 5.505e-005 3.8182 0.012006 4.2001e-005 0.0011563 0.21923 0.00065919 0.21988 0.20252 0 0.032994 0.0389 0 1.0904 0.33743 0.098333 0.012977 5.9149 0.081001 9.9989e-005 0.8091 0.0065363 0.0073273 0.0018488 0.98043 0.91562 4.06e-006 1.6241e-005 0.14222 0.61929 0.7 0.0016255 0.66415 0.44969 0.0021814 0.42239 1.1934 1.1883 16.0001 144.9649 0.00048265 -83.9218 0.098953
3.203 0.98806 5.505e-005 3.8182 0.012006 4.2014e-005 0.0011563 0.21924 0.00065919 0.2199 0.20254 0 0.032994 0.0389 0 1.0905 0.33747 0.09835 0.012979 5.9161 0.081012 0.0001 0.80909 0.0065371 0.0073281 0.0018439 0.98052 0.91973 4.0485e-006 1.6195e-005 0.14223 0.62041 0.70125 0.0016232 0.66596 0.44987 0.0021784 0.42238 1.1956 1.1905 16.0002 144.9649 0.00048109 -83.9378 0.099953
3.204 0.98806 5.505e-005 3.8182 0.012006 4.2027e-005 0.0011563 0.21926 0.00065919 0.21991 0.20255 0 0.032993 0.0389 0 1.0906 0.33752 0.098366 0.012981 5.9173 0.081023 0.00010002 0.80908 0.0065378 0.0073288 0.0018392 0.98061 0.92362 4.0374e-006 1.6151e-005 0.14223 0.62154 0.70248 0.001621 0.66776 0.45005 0.0021754 0.42238 1.1978 1.1927 16.0003 144.9649 0.00047953 -83.9533 0.10095
3.205 0.98806 5.505e-005 3.8182 0.012006 4.204e-005 0.0011563 0.21927 0.00065919 0.21992 0.20256 0 0.032993 0.0389 0 1.0907 0.33757 0.098382 0.012983 5.9186 0.081034 0.00010003 0.80907 0.0065385 0.0073296 0.0018346 0.98069 0.92729 4.0266e-006 1.6108e-005 0.14224 0.62266 0.7037 0.0016188 0.66956 0.45024 0.0021725 0.42238 1.2 1.1949 16.0003 144.9649 0.00047798 -83.9685 0.10195
3.206 0.98806 5.505e-005 3.8182 0.012006 4.2053e-005 0.0011563 0.21928 0.00065919 0.21994 0.20257 0 0.032992 0.0389 0 1.0908 0.33761 0.098398 0.012984 5.9198 0.081045 0.00010005 0.80906 0.0065392 0.0073304 0.0018302 0.98077 0.93076 4.0161e-006 1.6066e-005 0.14225 0.62377 0.70491 0.0016167 0.67135 0.45042 0.0021698 0.42237 1.2022 1.1971 16.0004 144.9649 0.00047644 -83.9833 0.10295
3.207 0.98806 5.505e-005 3.8182 0.012006 4.2066e-005 0.0011563 0.21929 0.00065919 0.21995 0.20259 0 0.032991 0.0389 0 1.0909 0.33766 0.098414 0.012986 5.9211 0.081055 0.00010006 0.80904 0.0065399 0.0073312 0.0018259 0.98084 0.93403 4.0058e-006 1.6025e-005 0.14225 0.62489 0.70612 0.0016147 0.67314 0.4506 0.002167 0.42237 1.2043 1.1993 16.0005 144.9649 0.00047491 -83.9977 0.10395
3.208 0.98806 5.505e-005 3.8182 0.012006 4.2079e-005 0.0011563 0.21931 0.00065919 0.21996 0.2026 0 0.032991 0.0389 0 1.091 0.3377 0.09843 0.012988 5.9223 0.081066 0.00010008 0.80903 0.0065407 0.0073319 0.0018216 0.98091 0.93713 3.9958e-006 1.5985e-005 0.14226 0.626 0.70731 0.0016127 0.67492 0.45078 0.0021644 0.42237 1.2065 1.2015 16.0006 144.9649 0.00047338 -84.0118 0.10495
3.209 0.98806 5.505e-005 3.8182 0.012006 4.2092e-005 0.0011563 0.21932 0.00065919 0.21997 0.20261 0 0.03299 0.0389 0 1.0911 0.33775 0.098446 0.01299 5.9236 0.081077 0.00010009 0.80902 0.0065414 0.0073327 0.0018174 0.98098 0.94005 3.986e-006 1.5945e-005 0.14226 0.6271 0.7085 0.0016107 0.67669 0.45096 0.0021618 0.42236 1.2087 1.2037 16.0007 144.9649 0.00047187 -84.0257 0.10595
3.21 0.98806 5.5049e-005 3.8182 0.012006 4.2106e-005 0.0011563 0.21933 0.00065919 0.21999 0.20262 0 0.032989 0.0389 0 1.0912 0.3378 0.098462 0.012991 5.9248 0.081088 0.00010011 0.80901 0.0065421 0.0073335 0.0018132 0.98105 0.94282 3.9764e-006 1.5907e-005 0.14227 0.62821 0.70967 0.0016088 0.67845 0.45114 0.0021593 0.42236 1.2108 1.2059 16.0008 144.9649 0.00047036 -84.0393 0.10695
3.211 0.98806 5.5049e-005 3.8182 0.012006 4.2119e-005 0.0011563 0.21934 0.00065919 0.22 0.20263 0 0.032989 0.0389 0 1.0913 0.33784 0.098478 0.012993 5.926 0.081099 0.00010012 0.809 0.0065428 0.0073342 0.0018091 0.98111 0.94543 3.967e-006 1.5869e-005 0.14228 0.62931 0.71084 0.0016069 0.6802 0.45132 0.0021568 0.42236 1.213 1.2081 16.0008 144.965 0.00046886 -84.0527 0.10795
3.212 0.98806 5.5049e-005 3.8182 0.012006 4.2132e-005 0.0011563 0.21936 0.00065919 0.22001 0.20265 0 0.032988 0.0389 0 1.0914 0.33789 0.098495 0.012995 5.9273 0.08111 0.00010014 0.80899 0.0065436 0.007335 0.0018052 0.98117 0.94789 3.9578e-006 1.5832e-005 0.14228 0.6304 0.712 0.0016051 0.68195 0.45151 0.0021544 0.42235 1.2152 1.2103 16.0009 144.965 0.00046737 -84.0658 0.10895
3.213 0.98806 5.5049e-005 3.8182 0.012006 4.2145e-005 0.0011563 0.21937 0.00065919 0.22002 0.20266 0 0.032987 0.0389 0 1.0915 0.33793 0.098511 0.012997 5.9285 0.081121 0.00010015 0.80898 0.0065443 0.0073358 0.0018013 0.98123 0.95022 3.9488e-006 1.5796e-005 0.14229 0.6315 0.71315 0.0016033 0.68369 0.45169 0.002152 0.42235 1.2173 1.2124 16.001 144.965 0.00046589 -84.0787 0.10995
3.214 0.98806 5.5049e-005 3.8182 0.012006 4.2158e-005 0.0011563 0.21938 0.00065919 0.22004 0.20267 0 0.032987 0.0389 0 1.0916 0.33798 0.098527 0.012998 5.9298 0.081132 0.00010017 0.80897 0.006545 0.0073365 0.0017976 0.98129 0.95242 3.9399e-006 1.5761e-005 0.14229 0.63259 0.71429 0.0016015 0.68543 0.45187 0.0021496 0.42235 1.2195 1.2146 16.0011 144.965 0.00046441 -84.0914 0.11095
3.215 0.98806 5.5049e-005 3.8182 0.012006 4.2171e-005 0.0011563 0.2194 0.00065919 0.22005 0.20268 0 0.032986 0.0389 0 1.0917 0.33802 0.098543 0.013 5.931 0.081143 0.00010018 0.80896 0.0065457 0.0073373 0.0017939 0.98135 0.95449 3.9312e-006 1.5726e-005 0.1423 0.63367 0.71542 0.0015997 0.68715 0.45205 0.0021473 0.42235 1.2216 1.2168 16.0011 144.965 0.00046294 -84.1039 0.11195
3.216 0.98806 5.5049e-005 3.8182 0.012006 4.2184e-005 0.0011563 0.21941 0.00065919 0.22006 0.20269 0 0.032985 0.0389 0 1.0918 0.33807 0.098559 0.013002 5.9323 0.081154 0.0001002 0.80895 0.0065465 0.0073381 0.0017902 0.98141 0.95645 3.9226e-006 1.5691e-005 0.1423 0.63476 0.71654 0.001598 0.68887 0.45223 0.002145 0.42235 1.2238 1.2189 16.0012 144.965 0.00046149 -84.1163 0.11295
3.217 0.98806 5.5049e-005 3.8182 0.012006 4.2197e-005 0.0011563 0.21942 0.00065919 0.22008 0.20271 0 0.032985 0.0389 0 1.0919 0.33812 0.098575 0.013004 5.9335 0.081165 0.00010021 0.80894 0.0065472 0.0073389 0.0017866 0.98146 0.9583 3.9141e-006 1.5658e-005 0.14231 0.63584 0.71766 0.0015963 0.69058 0.45241 0.0021428 0.42234 1.2259 1.2211 16.0013 144.965 0.00046003 -84.1285 0.11395
3.218 0.98806 5.5049e-005 3.8182 0.012005 4.221e-005 0.0011563 0.21943 0.00065919 0.22009 0.20272 0 0.032984 0.0389 0 1.092 0.33816 0.098591 0.013005 5.9347 0.081176 0.00010023 0.80892 0.0065479 0.0073396 0.001783 0.98151 0.96005 3.9058e-006 1.5624e-005 0.14232 0.63691 0.71877 0.0015946 0.69229 0.45259 0.0021406 0.42234 1.228 1.2232 16.0014 144.965 0.00045859 -84.1406 0.11495
3.219 0.98806 5.5049e-005 3.8182 0.012005 4.2223e-005 0.0011563 0.21945 0.00065919 0.2201 0.20273 0 0.032983 0.0389 0 1.0921 0.33821 0.098607 0.013007 5.936 0.081186 0.00010024 0.80891 0.0065486 0.0073404 0.0017795 0.98157 0.9617 3.8976e-006 1.5591e-005 0.14232 0.63799 0.71986 0.001593 0.69398 0.45277 0.0021384 0.42234 1.2302 1.2254 16.0015 144.965 0.00045716 -84.1525 0.11595
3.22 0.98806 5.5049e-005 3.8182 0.012005 4.2236e-005 0.0011563 0.21946 0.00065919 0.22011 0.20274 0 0.032983 0.0389 0 1.0922 0.33825 0.098623 0.013009 5.9372 0.081197 0.00010026 0.8089 0.0065494 0.0073412 0.001776 0.98162 0.96326 3.8895e-006 1.5559e-005 0.14233 0.63906 0.72095 0.0015913 0.69567 0.45296 0.0021363 0.42234 1.2323 1.2275 16.0015 144.965 0.00045573 -84.1642 0.11695
3.221 0.98806 5.5049e-005 3.8182 0.012005 4.2249e-005 0.0011563 0.21947 0.00065919 0.22013 0.20275 0 0.032982 0.0389 0 1.0923 0.3383 0.09864 0.013011 5.9385 0.081208 0.00010027 0.80889 0.0065501 0.0073419 0.0017725 0.98167 0.96473 3.8815e-006 1.5527e-005 0.14233 0.64012 0.72204 0.0015897 0.69735 0.45314 0.0021341 0.42234 1.2344 1.2297 16.0016 144.965 0.00045431 -84.1758 0.11795
3.222 0.98806 5.5049e-005 3.8182 0.012005 4.2262e-005 0.0011563 0.21948 0.00065919 0.22014 0.20276 0 0.032981 0.0389 0 1.0924 0.33835 0.098656 0.013012 5.9397 0.081219 0.00010029 0.80888 0.0065508 0.0073427 0.0017691 0.98172 0.96612 3.8736e-006 1.5495e-005 0.14234 0.64119 0.72311 0.0015881 0.69903 0.45332 0.002132 0.42234 1.2366 1.2318 16.0017 144.9651 0.0004529 -84.1873 0.11895
3.223 0.98806 5.5049e-005 3.8182 0.012005 4.2275e-005 0.0011563 0.2195 0.00065919 0.22015 0.20278 0 0.032981 0.0389 0 1.0925 0.33839 0.098672 0.013014 5.941 0.08123 0.0001003 0.80887 0.0065515 0.0073435 0.0017658 0.98177 0.96743 3.8658e-006 1.5464e-005 0.14235 0.64225 0.72418 0.0015865 0.70069 0.4535 0.00213 0.42234 1.2387 1.2339 16.0018 144.9651 0.00045149 -84.1987 0.11995
3.224 0.98806 5.5049e-005 3.8182 0.012005 4.2288e-005 0.0011563 0.21951 0.00065919 0.22016 0.20279 0 0.03298 0.0389 0 1.0926 0.33844 0.098688 0.013016 5.9422 0.081241 0.00010032 0.80886 0.0065522 0.0073442 0.0017625 0.98182 0.96867 3.8581e-006 1.5433e-005 0.14235 0.64331 0.72523 0.001585 0.70235 0.45368 0.0021279 0.42234 1.2408 1.2361 16.0018 144.9651 0.00045009 -84.21 0.12095
3.225 0.98806 5.5048e-005 3.8182 0.012005 4.2301e-005 0.0011563 0.21952 0.00065919 0.22018 0.2028 0 0.032979 0.0389 0 1.0927 0.33848 0.098704 0.013018 5.9435 0.081252 0.00010033 0.80885 0.006553 0.007345 0.0017592 0.98186 0.96984 3.8505e-006 1.5403e-005 0.14236 0.64436 0.72628 0.0015834 0.70401 0.45386 0.0021259 0.42234 1.2429 1.2382 16.0019 144.9651 0.0004487 -84.2211 0.12195
3.226 0.98806 5.5048e-005 3.8182 0.012005 4.2314e-005 0.0011563 0.21953 0.00065919 0.22019 0.20281 0 0.032979 0.0389 0 1.0928 0.33853 0.09872 0.013019 5.9447 0.081263 0.00010034 0.80884 0.0065537 0.0073458 0.0017561 0.98191 0.97094 3.843e-006 1.5373e-005 0.14236 0.64541 0.72733 0.0015819 0.70565 0.45404 0.0021239 0.42234 1.245 1.2403 16.002 144.9651 0.00044732 -84.2322 0.12295
3.227 0.98806 5.5048e-005 3.8182 0.012005 4.2327e-005 0.0011563 0.21955 0.00065919 0.2202 0.20282 0 0.032978 0.0389 0 1.0929 0.33857 0.098736 0.013021 5.946 0.081274 0.00010036 0.80883 0.0065544 0.0073466 0.0017529 0.98196 0.97198 3.8356e-006 1.5343e-005 0.14237 0.64646 0.72836 0.0015804 0.70729 0.45423 0.0021219 0.42233 1.2471 1.2424 16.002 144.9651 0.00044595 -84.2431 0.12395
3.228 0.98806 5.5048e-005 3.8182 0.012005 4.234e-005 0.0011563 0.21956 0.00065919 0.22021 0.20284 0 0.032977 0.0389 0 1.093 0.33862 0.098752 0.013023 5.9472 0.081285 0.00010037 0.80882 0.0065551 0.0073473 0.0017498 0.982 0.97297 3.8282e-006 1.5314e-005 0.14237 0.6475 0.72939 0.0015789 0.70892 0.45441 0.0021199 0.42233 1.2492 1.2445 16.0021 144.9651 0.00044458 -84.2539 0.12495
3.229 0.98806 5.5048e-005 3.8182 0.012005 4.2353e-005 0.0011563 0.21957 0.00065919 0.22023 0.20285 0 0.032977 0.0389 0 1.0931 0.33867 0.098769 0.013025 5.9485 0.081296 0.00010039 0.8088 0.0065559 0.0073481 0.0017467 0.98205 0.97389 3.821e-006 1.5285e-005 0.14238 0.64854 0.73041 0.0015774 0.71054 0.45459 0.002118 0.42233 1.2513 1.2466 16.0022 144.9651 0.00044322 -84.2646 0.12595
3.23 0.98806 5.5048e-005 3.8182 0.012005 4.2366e-005 0.0011563 0.21958 0.00065919 0.22024 0.20286 0 0.032976 0.0389 0 1.0932 0.33871 0.098785 0.013026 5.9497 0.081307 0.0001004 0.80879 0.0065566 0.0073489 0.0017436 0.98209 0.97477 3.8138e-006 1.5256e-005 0.14239 0.64958 0.73142 0.0015759 0.71215 0.45477 0.0021161 0.42233 1.2534 1.2487 16.0023 144.9651 0.00044187 -84.2752 0.12695
3.231 0.98806 5.5048e-005 3.8182 0.012005 4.2379e-005 0.0011563 0.2196 0.00065919 0.22025 0.20287 0 0.032976 0.0389 0 1.0933 0.33876 0.098801 0.013028 5.951 0.081317 0.00010042 0.80878 0.0065573 0.0073496 0.0017405 0.98214 0.9756 3.8067e-006 1.5228e-005 0.14239 0.65062 0.73243 0.0015745 0.71376 0.45495 0.0021142 0.42233 1.2554 1.2508 16.0023 144.9651 0.00044052 -84.2858 0.12795
3.232 0.98806 5.5048e-005 3.8182 0.012005 4.2393e-005 0.0011563 0.21961 0.00065919 0.22026 0.20288 0 0.032975 0.0389 0 1.0934 0.3388 0.098817 0.01303 5.9522 0.081328 0.00010043 0.80877 0.006558 0.0073504 0.0017375 0.98218 0.97638 3.7997e-006 1.52e-005 0.1424 0.65165 0.73343 0.0015731 0.71536 0.45513 0.0021123 0.42233 1.2575 1.2529 16.0024 144.9651 0.00043918 -84.2962 0.12895
3.233 0.98806 5.5048e-005 3.8182 0.012005 4.2406e-005 0.0011563 0.21962 0.00065919 0.22028 0.2029 0 0.032974 0.0389 0 1.0935 0.33885 0.098833 0.013032 5.9535 0.081339 0.00010045 0.80876 0.0065588 0.0073512 0.0017345 0.98222 0.97712 3.7927e-006 1.5172e-005 0.1424 0.65268 0.73442 0.0015716 0.71696 0.45532 0.0021105 0.42234 1.2596 1.255 16.0025 144.9652 0.00043785 -84.3065 0.12995
3.234 0.98806 5.5048e-005 3.8182 0.012005 4.2419e-005 0.0011563 0.21963 0.00065919 0.22029 0.20291 0 0.032974 0.0389 0 1.0936 0.3389 0.098849 0.013033 5.9547 0.08135 0.00010046 0.80875 0.0065595 0.007352 0.0017315 0.98226 0.97782 3.7859e-006 1.5144e-005 0.14241 0.6537 0.7354 0.0015702 0.71854 0.4555 0.0021086 0.42234 1.2617 1.2571 16.0025 144.9652 0.00043652 -84.3168 0.13095
3.235 0.98806 5.5048e-005 3.8182 0.012005 4.2432e-005 0.0011563 0.21965 0.00065919 0.2203 0.20292 0 0.032973 0.0389 0 1.0937 0.33894 0.098865 0.013035 5.956 0.081361 0.00010048 0.80874 0.0065602 0.0073527 0.0017285 0.98231 0.97847 3.7791e-006 1.5117e-005 0.14242 0.65472 0.73638 0.0015688 0.72012 0.45568 0.0021068 0.42234 1.2637 1.2592 16.0026 144.9652 0.00043521 -84.3269 0.13195
3.236 0.98806 5.5048e-005 3.8182 0.012005 4.2445e-005 0.0011563 0.21966 0.00065919 0.22031 0.20293 0 0.032972 0.0389 0 1.0938 0.33899 0.098881 0.013037 5.9572 0.081372 0.00010049 0.80873 0.0065609 0.0073535 0.0017256 0.98235 0.97909 3.7724e-006 1.509e-005 0.14242 0.65574 0.73735 0.0015674 0.72169 0.45586 0.002105 0.42234 1.2658 1.2613 16.0027 144.9652 0.0004339 -84.337 0.13295
3.237 0.98806 5.5048e-005 3.8182 0.012005 4.2458e-005 0.0011563 0.21967 0.00065919 0.22033 0.20294 0 0.032972 0.0389 0 1.0939 0.33903 0.098897 0.013039 5.9585 0.081383 0.00010051 0.80872 0.0065617 0.0073543 0.0017228 0.98239 0.97968 3.7657e-006 1.5064e-005 0.14243 0.65676 0.73831 0.0015661 0.72325 0.45604 0.0021032 0.42234 1.2679 1.2634 16.0027 144.9652 0.00043259 -84.347 0.13395
3.238 0.98806 5.5048e-005 3.8182 0.012005 4.2471e-005 0.0011563 0.21968 0.00065919 0.22034 0.20295 0 0.032971 0.0389 0 1.094 0.33908 0.098914 0.01304 5.9597 0.081394 0.00010052 0.80871 0.0065624 0.007355 0.00172 0.98243 0.98023 3.7591e-006 1.5037e-005 0.14243 0.65777 0.73927 0.0015647 0.72481 0.45622 0.0021014 0.42234 1.2699 1.2654 16.0028 144.9652 0.0004313 -84.3569 0.13495
3.239 0.98806 5.5047e-005 3.8182 0.012005 4.2484e-005 0.0011563 0.2197 0.00065919 0.22035 0.20297 0 0.03297 0.0389 0 1.0941 0.33913 0.09893 0.013042 5.961 0.081405 0.00010054 0.8087 0.0065631 0.0073558 0.0017172 0.98247 0.98076 3.7526e-006 1.5011e-005 0.14244 0.65878 0.74022 0.0015634 0.72636 0.4564 0.0020997 0.42234 1.272 1.2675 16.0029 144.9652 0.00043001 -84.3667 0.13595
3.24 0.98806 5.5047e-005 3.8182 0.012005 4.2497e-005 0.0011563 0.21971 0.00065919 0.22036 0.20298 0 0.03297 0.0389 0 1.0942 0.33917 0.098946 0.013044 5.9622 0.081416 0.00010055 0.80868 0.0065638 0.0073566 0.0017145 0.98251 0.98125 3.7461e-006 1.4985e-005 0.14245 0.65979 0.74116 0.001562 0.7279 0.45659 0.0020979 0.42234 1.274 1.2695 16.0029 144.9652 0.00042872 -84.3764 0.13695
3.241 0.98806 5.5047e-005 3.8182 0.012005 4.251e-005 0.0011563 0.21972 0.00065919 0.22038 0.20299 0 0.032969 0.0389 0 1.0943 0.33922 0.098962 0.013046 5.9635 0.081426 0.00010057 0.80867 0.0065645 0.0073573 0.0017118 0.98255 0.98172 3.7397e-006 1.496e-005 0.14245 0.66079 0.7421 0.0015607 0.72944 0.45677 0.0020962 0.42234 1.2761 1.2716 16.003 144.9652 0.00042745 -84.3861 0.13795
3.242 0.98806 5.5047e-005 3.8182 0.012005 4.2523e-005 0.0011563 0.21973 0.00065919 0.22039 0.203 0 0.032968 0.0389 0 1.0944 0.33926 0.098978 0.013047 5.9648 0.081437 0.00010058 0.80866 0.0065653 0.0073581 0.0017091 0.98258 0.98216 3.7334e-006 1.4934e-005 0.14246 0.66179 0.74303 0.0015594 0.73096 0.45695 0.0020945 0.42234 1.2781 1.2737 16.0031 144.9653 0.00042618 -84.3956 0.13895
3.243 0.98806 5.5047e-005 3.8182 0.012005 4.2536e-005 0.0011563 0.21975 0.00065919 0.2204 0.20301 0 0.032968 0.0389 0 1.0945 0.33931 0.098994 0.013049 5.966 0.081448 0.0001006 0.80865 0.006566 0.0073589 0.0017064 0.98262 0.98257 3.7271e-006 1.4909e-005 0.14246 0.66279 0.74395 0.0015581 0.73248 0.45713 0.0020928 0.42234 1.2801 1.2757 16.0031 144.9653 0.00042491 -84.4051 0.13995
3.244 0.98806 5.5047e-005 3.8182 0.012005 4.2549e-005 0.0011563 0.21976 0.00065919 0.22041 0.20302 0 0.032967 0.0389 0 1.0945 0.33935 0.09901 0.013051 5.9673 0.081459 0.00010061 0.80864 0.0065667 0.0073597 0.0017037 0.98266 0.98297 3.7209e-006 1.4884e-005 0.14247 0.66379 0.74487 0.0015568 0.734 0.45731 0.0020911 0.42235 1.2822 1.2778 16.0032 144.9653 0.00042366 -84.4146 0.14095
3.245 0.98806 5.5047e-005 3.8182 0.012005 4.2562e-005 0.0011563 0.21977 0.00065919 0.22042 0.20304 0 0.032966 0.0389 0 1.0946 0.3394 0.099026 0.013053 5.9685 0.08147 0.00010063 0.80863 0.0065674 0.0073604 0.001701 0.9827 0.98334 3.7148e-006 1.486e-005 0.14247 0.66478 0.74578 0.0015556 0.7355 0.45749 0.0020895 0.42235 1.2842 1.2798 16.0033 144.9653 0.00042241 -84.4239 0.14195
3.246 0.98806 5.5047e-005 3.8182 0.012005 4.2575e-005 0.0011563 0.21978 0.00065919 0.22044 0.20305 0 0.032966 0.0389 0 1.0947 0.33945 0.099042 0.013054 5.9698 0.081481 0.00010064 0.80862 0.0065682 0.0073612 0.0016983 0.98273 0.98369 3.7087e-006 1.4835e-005 0.14248 0.66577 0.74668 0.0015543 0.737 0.45767 0.0020878 0.42235 1.2862 1.2818 16.0033 144.9653 0.00042117 -84.4332 0.14295
3.247 0.98806 5.5047e-005 3.8182 0.012005 4.2588e-005 0.0011563 0.21979 0.00065919 0.22045 0.20306 0 0.032965 0.0389 0 1.0948 0.33949 0.099059 0.013056 5.971 0.081492 0.00010066 0.80861 0.0065689 0.007362 0.0016957 0.98277 0.98402 3.7027e-006 1.4811e-005 0.14249 0.66675 0.74758 0.0015531 0.73849 0.45786 0.0020862 0.42235 1.2882 1.2839 16.0034 144.9653 0.00041993 -84.4423 0.14395
3.248 0.98806 5.5047e-005 3.8182 0.012005 4.2601e-005 0.0011563 0.21981 0.00065919 0.22046 0.20307 0 0.032965 0.0389 0 1.0949 0.33954 0.099075 0.013058 5.9723 0.081503 0.00010067 0.8086 0.0065696 0.0073627 0.0016931 0.98281 0.98433 3.6967e-006 1.4787e-005 0.14249 0.66773 0.74848 0.0015518 0.73998 0.45804 0.0020846 0.42235 1.2902 1.2859 16.0035 144.9653 0.0004187 -84.4515 0.14495
3.249 0.98806 5.5047e-005 3.8182 0.012005 4.2614e-005 0.0011564 0.21982 0.00065919 0.22047 0.20308 0 0.032964 0.0389 0 1.095 0.33958 0.099091 0.01306 5.9736 0.081514 0.00010069 0.80859 0.0065703 0.0073635 0.0016906 0.98284 0.98463 3.6908e-006 1.4764e-005 0.1425 0.66871 0.74936 0.0015506 0.74145 0.45822 0.0020829 0.42236 1.2922 1.2879 16.0035 144.9653 0.00041747 -84.4605 0.14595
3.25 0.98806 5.5047e-005 3.8182 0.012005 4.2627e-005 0.0011564 0.21983 0.00065919 0.22049 0.20309 0 0.032963 0.0389 0 1.0951 0.33963 0.099107 0.013061 5.9748 0.081525 0.0001007 0.80858 0.0065711 0.0073643 0.001688 0.98288 0.98491 3.6849e-006 1.474e-005 0.1425 0.66969 0.75024 0.0015494 0.74292 0.4584 0.0020814 0.42236 1.2942 1.2899 16.0036 144.9653 0.00041626 -84.4695 0.14695
3.251 0.98806 5.5047e-005 3.8182 0.012005 4.264e-005 0.0011564 0.21984 0.00065919 0.2205 0.20311 0 0.032963 0.0389 0 1.0952 0.33968 0.099123 0.013063 5.9761 0.081535 0.00010072 0.80857 0.0065718 0.007365 0.0016855 0.98291 0.98518 3.6791e-006 1.4717e-005 0.14251 0.67066 0.75112 0.0015482 0.74438 0.45858 0.0020798 0.42236 1.2962 1.2919 16.0036 144.9654 0.00041505 -84.4784 0.14795
3.252 0.98806 5.5047e-005 3.8182 0.012005 4.2653e-005 0.0011564 0.21986 0.00065919 0.22051 0.20312 0 0.032962 0.0389 0 1.0953 0.33972 0.099139 0.013065 5.9773 0.081546 0.00010073 0.80855 0.0065725 0.0073658 0.0016831 0.98295 0.98543 3.6734e-006 1.4694e-005 0.14252 0.67163 0.75199 0.001547 0.74584 0.45876 0.0020782 0.42236 1.2982 1.294 16.0037 144.9654 0.00041384 -84.4872 0.14895
3.253 0.98806 5.5047e-005 3.8182 0.012005 4.2666e-005 0.0011564 0.21987 0.00065919 0.22052 0.20313 0 0.032961 0.0389 0 1.0954 0.33977 0.099155 0.013067 5.9786 0.081557 0.00010074 0.80854 0.0065732 0.0073666 0.0016807 0.98298 0.98566 3.6677e-006 1.4671e-005 0.14252 0.6726 0.75285 0.0015458 0.74729 0.45894 0.0020767 0.42236 1.3002 1.296 16.0038 144.9654 0.00041264 -84.4959 0.14995
3.254 0.98806 5.5046e-005 3.8182 0.012005 4.268e-005 0.0011564 0.21988 0.00065919 0.22054 0.20314 0 0.032961 0.0389 0 1.0955 0.33981 0.099171 0.013068 5.9798 0.081568 0.00010076 0.80853 0.006574 0.0073674 0.0016784 0.98302 0.98589 3.6621e-006 1.4649e-005 0.14253 0.67357 0.75371 0.0015446 0.74873 0.45913 0.0020751 0.42237 1.3022 1.298 16.0038 144.9654 0.00041145 -84.5046 0.15095
3.255 0.98806 5.5046e-005 3.8182 0.012005 4.2693e-005 0.0011564 0.21989 0.00065919 0.22055 0.20315 0 0.03296 0.0389 0 1.0956 0.33986 0.099188 0.01307 5.9811 0.081579 0.00010077 0.80852 0.0065747 0.0073681 0.001676 0.98305 0.9861 3.6565e-006 1.4627e-005 0.14253 0.67453 0.75456 0.0015434 0.75017 0.45931 0.0020736 0.42237 1.3042 1.3 16.0039 144.9654 0.00041027 -84.5132 0.15195
3.256 0.98806 5.5046e-005 3.8182 0.012005 4.2706e-005 0.0011564 0.2199 0.00065919 0.22056 0.20316 0 0.03296 0.0389 0 1.0957 0.33991 0.099204 0.013072 5.9824 0.08159 0.00010079 0.80851 0.0065754 0.0073689 0.0016737 0.98308 0.9863 3.651e-006 1.4605e-005 0.14254 0.67549 0.7554 0.0015423 0.75159 0.45949 0.0020721 0.42237 1.3062 1.302 16.0039 144.9654 0.00040909 -84.5218 0.15295
3.257 0.98806 5.5046e-005 3.8182 0.012005 4.2719e-005 0.0011564 0.21992 0.00065919 0.22057 0.20318 0 0.032959 0.0389 0 1.0958 0.33995 0.09922 0.013074 5.9836 0.081601 0.0001008 0.8085 0.0065761 0.0073697 0.0016714 0.98312 0.98649 3.6455e-006 1.4583e-005 0.14254 0.67644 0.75624 0.0015411 0.75301 0.45967 0.0020706 0.42237 1.3081 1.3039 16.004 144.9654 0.00040791 -84.5303 0.15395
3.258 0.98806 5.5046e-005 3.8182 0.012005 4.2732e-005 0.0011564 0.21993 0.00065919 0.22058 0.20319 0 0.032958 0.0389 0 1.0959 0.34 0.099236 0.013075 5.9849 0.081612 0.00010082 0.80849 0.0065769 0.0073704 0.0016691 0.98315 0.98667 3.6401e-006 1.4561e-005 0.14255 0.67739 0.75708 0.00154 0.75443 0.45985 0.0020691 0.42238 1.3101 1.3059 16.0041 144.9654 0.00040674 -84.5387 0.15495
3.259 0.98806 5.5046e-005 3.8182 0.012005 4.2745e-005 0.0011564 0.21994 0.00065919 0.2206 0.2032 0 0.032958 0.0389 0 1.096 0.34004 0.099252 0.013077 5.9862 0.081623 0.00010083 0.80848 0.0065776 0.0073712 0.0016667 0.98318 0.98684 3.6347e-006 1.4539e-005 0.14256 0.67834 0.75791 0.0015389 0.75583 0.46003 0.0020677 0.42238 1.3121 1.3079 16.0041 144.9654 0.00040558 -84.547 0.15595
3.26 0.98806 5.5046e-005 3.8182 0.012005 4.2758e-005 0.0011564 0.21995 0.00065919 0.22061 0.20321 0 0.032957 0.0389 0 1.0961 0.34009 0.099268 0.013079 5.9874 0.081633 0.00010085 0.80847 0.0065783 0.007372 0.0016644 0.98321 0.987 3.6294e-006 1.4518e-005 0.14256 0.67929 0.75873 0.0015378 0.75723 0.46021 0.0020662 0.42238 1.314 1.3099 16.0042 144.9655 0.00040443 -84.5553 0.15695
3.261 0.98806 5.5046e-005 3.8182 0.012005 4.2771e-005 0.0011564 0.21997 0.00065919 0.22062 0.20322 0 0.032956 0.0389 0 1.0962 0.34013 0.099284 0.01308 5.9887 0.081644 0.00010086 0.80846 0.006579 0.0073728 0.0016621 0.98325 0.98716 3.6241e-006 1.4497e-005 0.14257 0.68024 0.75955 0.0015367 0.75863 0.46039 0.0020648 0.42239 1.316 1.3119 16.0042 144.9655 0.00040328 -84.5635 0.15795
3.262 0.98806 5.5046e-005 3.8182 0.012005 4.2784e-005 0.0011564 0.21998 0.0006592 0.22063 0.20323 0 0.032956 0.0389 0 1.0963 0.34018 0.0993 0.013082 5.9899 0.081655 0.00010088 0.80845 0.0065797 0.0073735 0.0016598 0.98328 0.9873 3.6189e-006 1.4476e-005 0.14257 0.68118 0.76036 0.0015356 0.76001 0.46058 0.0020633 0.42239 1.318 1.3138 16.0043 144.9655 0.00040213 -84.5717 0.15895
3.263 0.98806 5.5046e-005 3.8182 0.012005 4.2797e-005 0.0011564 0.21999 0.0006592 0.22064 0.20325 0 0.032955 0.0389 0 1.0964 0.34023 0.099316 0.013084 5.9912 0.081666 0.00010089 0.80843 0.0065805 0.0073743 0.0016575 0.98331 0.98744 3.6137e-006 1.4455e-005 0.14258 0.68211 0.76117 0.0015345 0.76139 0.46076 0.0020619 0.42239 1.3199 1.3158 16.0044 144.9655 0.000401 -84.5797 0.15995
3.264 0.98806 5.5046e-005 3.8182 0.012005 4.281e-005 0.0011564 0.22 0.0006592 0.22066 0.20326 0 0.032954 0.0389 0 1.0965 0.34027 0.099333 0.013086 5.9925 0.081677 0.00010091 0.80842 0.0065812 0.0073751 0.0016551 0.98334 0.98757 3.6086e-006 1.4435e-005 0.14259 0.68305 0.76197 0.0015335 0.76276 0.46094 0.0020605 0.4224 1.3219 1.3178 16.0044 144.9655 0.00039986 -84.5878 0.16095
3.265 0.98806 5.5046e-005 3.8182 0.012005 4.2823e-005 0.0011564 0.22001 0.0006592 0.22067 0.20327 0 0.032954 0.0389 0 1.0966 0.34032 0.099349 0.013087 5.9937 0.081688 0.00010092 0.80841 0.0065819 0.0073758 0.0016528 0.98337 0.98769 3.6035e-006 1.4415e-005 0.14259 0.68398 0.76277 0.0015324 0.76413 0.46112 0.0020591 0.4224 1.3238 1.3197 16.0045 144.9655 0.00039874 -84.5957 0.16195
3.266 0.98806 5.5046e-005 3.8182 0.012005 4.2836e-005 0.0011564 0.22003 0.0006592 0.22068 0.20328 0 0.032953 0.0389 0 1.0967 0.34036 0.099365 0.013089 5.995 0.081699 0.00010094 0.8084 0.0065826 0.0073766 0.0016506 0.9834 0.98781 3.5985e-006 1.4394e-005 0.1426 0.68491 0.76356 0.0015313 0.76549 0.4613 0.0020577 0.4224 1.3257 1.3217 16.0045 144.9655 0.00039762 -84.6036 0.16295
3.267 0.98806 5.5046e-005 3.8182 0.012005 4.2849e-005 0.0011564 0.22004 0.0006592 0.22069 0.20329 0 0.032953 0.0389 0 1.0968 0.34041 0.099381 0.013091 5.9963 0.08171 0.00010095 0.80839 0.0065834 0.0073774 0.0016484 0.98343 0.98792 3.5935e-006 1.4374e-005 0.1426 0.68584 0.76435 0.0015303 0.76684 0.46148 0.0020563 0.42241 1.3277 1.3236 16.0046 144.9655 0.0003965 -84.6115 0.16395
3.268 0.98806 5.5045e-005 3.8182 0.012005 4.2862e-005 0.0011564 0.22005 0.0006592 0.22071 0.2033 0 0.032952 0.0389 0 1.0969 0.34046 0.099397 0.013093 5.9975 0.081721 0.00010097 0.80838 0.0065841 0.0073781 0.0016463 0.98346 0.98803 3.5885e-006 1.4355e-005 0.14261 0.68676 0.76513 0.0015292 0.76818 0.46166 0.002055 0.42241 1.3296 1.3255 16.0046 144.9656 0.00039539 -84.6192 0.16495
3.269 0.98806 5.5045e-005 3.8182 0.012005 4.2875e-005 0.0011564 0.22006 0.0006592 0.22072 0.20331 0 0.032951 0.0389 0 1.097 0.3405 0.099413 0.013094 5.9988 0.081731 0.00010098 0.80837 0.0065848 0.0073789 0.0016443 0.98349 0.98813 3.5837e-006 1.4335e-005 0.14262 0.68768 0.7659 0.0015282 0.76952 0.46184 0.0020536 0.42242 1.3315 1.3275 16.0047 144.9656 0.00039429 -84.6269 0.16595
3.27 0.98806 5.5045e-005 3.8182 0.012005 4.2888e-005 0.0011564 0.22008 0.0006592 0.22073 0.20333 0 0.032951 0.0389 0 1.0971 0.34055 0.099429 0.013096 6.0001 0.081742 0.000101 0.80836 0.0065855 0.0073797 0.0016422 0.98352 0.98822 3.5788e-006 1.4316e-005 0.14262 0.6886 0.76668 0.0015271 0.77085 0.46203 0.0020523 0.42242 1.3334 1.3294 16.0047 144.9656 0.00039319 -84.6346 0.16695
3.271 0.98806 5.5045e-005 3.8182 0.012005 4.2901e-005 0.0011564 0.22009 0.0006592 0.22074 0.20334 0 0.03295 0.0389 0 1.0972 0.34059 0.099445 0.013098 6.0013 0.081753 0.00010101 0.80835 0.0065863 0.0073805 0.0016402 0.98355 0.98831 3.574e-006 1.4296e-005 0.14263 0.68952 0.76744 0.0015261 0.77218 0.46221 0.002051 0.42242 1.3353 1.3313 16.0048 144.9656 0.0003921 -84.6422 0.16795
3.272 0.98806 5.5045e-005 3.8182 0.012005 4.2914e-005 0.0011564 0.2201 0.0006592 0.22075 0.20335 0 0.032949 0.0389 0 1.0973 0.34064 0.099462 0.0131 6.0026 0.081764 0.00010103 0.80834 0.006587 0.0073812 0.0016381 0.98357 0.9884 3.5692e-006 1.4277e-005 0.14263 0.69043 0.7682 0.0015251 0.77349 0.46239 0.0020497 0.42243 1.3373 1.3333 16.0048 144.9656 0.00039101 -84.6497 0.16895
3.273 0.98806 5.5045e-005 3.8182 0.012005 4.2927e-005 0.0011564 0.22011 0.0006592 0.22077 0.20336 0 0.032949 0.0389 0 1.0974 0.34069 0.099478 0.013101 6.0039 0.081775 0.00010104 0.80833 0.0065877 0.007382 0.0016361 0.9836 0.98848 3.5645e-006 1.4259e-005 0.14264 0.69134 0.76896 0.0015241 0.7748 0.46257 0.0020484 0.42243 1.3392 1.3352 16.0049 144.9656 0.00038993 -84.6572 0.16995
3.274 0.98806 5.5045e-005 3.8182 0.012005 4.294e-005 0.0011564 0.22012 0.0006592 0.22078 0.20337 0 0.032948 0.0389 0 1.0975 0.34073 0.099494 0.013103 6.0051 0.081786 0.00010106 0.80832 0.0065884 0.0073828 0.0016341 0.98363 0.98856 3.5598e-006 1.424e-005 0.14264 0.69225 0.76971 0.0015232 0.77611 0.46275 0.0020471 0.42244 1.3411 1.3371 16.005 144.9656 0.00038886 -84.6646 0.17095
3.275 0.98806 5.5045e-005 3.8182 0.012005 4.2953e-005 0.0011564 0.22014 0.0006592 0.22079 0.20338 0 0.032948 0.0389 0 1.0976 0.34078 0.09951 0.013105 6.0064 0.081797 0.00010107 0.8083 0.0065892 0.0073835 0.0016321 0.98366 0.98863 3.5552e-006 1.4221e-005 0.14265 0.69315 0.77046 0.0015222 0.77741 0.46293 0.0020458 0.42244 1.343 1.339 16.005 144.9656 0.00038779 -84.672 0.17195
3.276 0.98806 5.5045e-005 3.8182 0.012005 4.2966e-005 0.0011564 0.22015 0.0006592 0.2208 0.20339 0 0.032947 0.0389 0 1.0977 0.34082 0.099526 0.013107 6.0077 0.081808 0.00010109 0.80829 0.0065899 0.0073843 0.0016301 0.98369 0.98871 3.5506e-006 1.4203e-005 0.14266 0.69405 0.77121 0.0015212 0.7787 0.46311 0.0020445 0.42245 1.3449 1.3409 16.0051 144.9657 0.00038672 -84.6793 0.17295
3.277 0.98806 5.5045e-005 3.8182 0.012005 4.298e-005 0.0011564 0.22016 0.0006592 0.22081 0.20341 0 0.032946 0.0389 0 1.0978 0.34087 0.099542 0.013108 6.0089 0.081819 0.0001011 0.80828 0.0065906 0.0073851 0.0016282 0.98371 0.98877 3.5461e-006 1.4185e-005 0.14266 0.69495 0.77194 0.0015203 0.77998 0.46329 0.0020432 0.42245 1.3467 1.3428 16.0051 144.9657 0.00038566 -84.6865 0.17395
3.278 0.98806 5.5045e-005 3.8182 0.012005 4.2993e-005 0.0011564 0.22017 0.0006592 0.22083 0.20342 0 0.032946 0.0389 0 1.0979 0.34092 0.099558 0.01311 6.0102 0.081829 0.00010111 0.80827 0.0065913 0.0073859 0.0016262 0.98374 0.98884 3.5416e-006 1.4167e-005 0.14267 0.69585 0.77268 0.0015193 0.78126 0.46347 0.002042 0.42245 1.3486 1.3447 16.0052 144.9657 0.00038461 -84.6937 0.17495
3.279 0.98806 5.5045e-005 3.8182 0.012005 4.3006e-005 0.0011564 0.22018 0.0006592 0.22084 0.20343 0 0.032945 0.0389 0 1.098 0.34096 0.099574 0.013112 6.0115 0.08184 0.00010113 0.80826 0.006592 0.0073866 0.0016243 0.98377 0.9889 3.5371e-006 1.4149e-005 0.14267 0.69674 0.77341 0.0015184 0.78253 0.46366 0.0020408 0.42246 1.3505 1.3466 16.0052 144.9657 0.00038356 -84.7008 0.17595
3.28 0.98806 5.5045e-005 3.8182 0.012005 4.3019e-005 0.0011564 0.2202 0.0006592 0.22085 0.20344 0 0.032944 0.0389 0 1.0981 0.34101 0.099591 0.013114 6.0127 0.081851 0.00010114 0.80825 0.0065928 0.0073874 0.0016223 0.98379 0.98896 3.5327e-006 1.4131e-005 0.14268 0.69763 0.77413 0.0015175 0.78379 0.46384 0.0020395 0.42246 1.3524 1.3485 16.0053 144.9657 0.00038252 -84.7079 0.17695
3.281 0.98806 5.5045e-005 3.8182 0.012005 4.3032e-005 0.0011564 0.22021 0.0006592 0.22086 0.20345 0 0.032944 0.0389 0 1.0982 0.34105 0.099607 0.013115 6.014 0.081862 0.00010116 0.80824 0.0065935 0.0073882 0.0016204 0.98382 0.98902 3.5283e-006 1.4114e-005 0.14269 0.69852 0.77485 0.0015165 0.78505 0.46402 0.0020383 0.42247 1.3543 1.3504 16.0053 144.9657 0.00038148 -84.7149 0.17795
3.282 0.98806 5.5045e-005 3.8182 0.012005 4.3045e-005 0.0011564 0.22022 0.0006592 0.22087 0.20346 0 0.032943 0.0389 0 1.0983 0.3411 0.099623 0.013117 6.0153 0.081873 0.00010117 0.80823 0.0065942 0.0073889 0.0016186 0.98385 0.98907 3.5239e-006 1.4096e-005 0.14269 0.6994 0.77557 0.0015156 0.7863 0.4642 0.0020371 0.42247 1.3561 1.3523 16.0054 144.9657 0.00038045 -84.7219 0.17895
3.283 0.98806 5.5044e-005 3.8182 0.012005 4.3058e-005 0.0011564 0.22023 0.0006592 0.22089 0.20347 0 0.032943 0.0389 0 1.0984 0.34115 0.099639 0.013119 6.0165 0.081884 0.00010119 0.80822 0.0065949 0.0073897 0.0016167 0.98387 0.98912 3.5196e-006 1.4079e-005 0.1427 0.70029 0.77628 0.0015147 0.78755 0.46438 0.0020359 0.42248 1.358 1.3542 16.0054 144.9658 0.00037942 -84.7288 0.17995
3.284 0.98806 5.5044e-005 3.8182 0.012005 4.3071e-005 0.0011564 0.22024 0.0006592 0.2209 0.20349 0 0.032942 0.0389 0 1.0985 0.34119 0.099655 0.013121 6.0178 0.081895 0.0001012 0.80821 0.0065957 0.0073905 0.0016149 0.9839 0.98917 3.5153e-006 1.4062e-005 0.1427 0.70117 0.77699 0.0015137 0.78879 0.46456 0.0020347 0.42248 1.3598 1.356 16.0055 144.9658 0.0003784 -84.7357 0.18095
3.285 0.98806 5.5044e-005 3.8182 0.012005 4.3084e-005 0.0011564 0.22026 0.0006592 0.22091 0.2035 0 0.032941 0.0389 0 1.0986 0.34124 0.099671 0.013122 6.0191 0.081906 0.00010122 0.8082 0.0065964 0.0073912 0.0016131 0.98392 0.98922 3.5111e-006 1.4045e-005 0.14271 0.70204 0.77769 0.0015128 0.79002 0.46474 0.0020335 0.42249 1.3617 1.3579 16.0055 144.9658 0.00037738 -84.7425 0.18195
3.286 0.98806 5.5044e-005 3.8182 0.012004 4.3097e-005 0.0011564 0.22027 0.0006592 0.22092 0.20351 0 0.032941 0.0389 0 1.0987 0.34128 0.099687 0.013124 6.0204 0.081916 0.00010123 0.80818 0.0065971 0.007392 0.0016113 0.98395 0.98926 3.5069e-006 1.4028e-005 0.14271 0.70292 0.77839 0.0015119 0.79125 0.46492 0.0020324 0.42249 1.3636 1.3598 16.0056 144.9658 0.00037637 -84.7493 0.18295
3.287 0.98806 5.5044e-005 3.8182 0.012004 4.311e-005 0.0011564 0.22028 0.0006592 0.22093 0.20352 0 0.03294 0.0389 0 1.0988 0.34133 0.099703 0.013126 6.0216 0.081927 0.00010125 0.80817 0.0065978 0.0073928 0.0016095 0.98397 0.98931 3.5028e-006 1.4011e-005 0.14272 0.70379 0.77908 0.0015109 0.79247 0.4651 0.0020312 0.4225 1.3654 1.3616 16.0056 144.9658 0.00037536 -84.756 0.18395
3.288 0.98806 5.5044e-005 3.8182 0.012004 4.3123e-005 0.0011564 0.22029 0.0006592 0.22095 0.20353 0 0.03294 0.0389 0 1.0989 0.34137 0.09972 0.013128 6.0229 0.081938 0.00010126 0.80816 0.0065986 0.0073936 0.0016078 0.984 0.98935 3.4986e-006 1.3995e-005 0.14273 0.70466 0.77977 0.00151 0.79368 0.46528 0.0020301 0.42251 1.3672 1.3635 16.0057 144.9658 0.00037436 -84.7626 0.18495
3.289 0.98806 5.5044e-005 3.8182 0.012004 4.3136e-005 0.0011564 0.2203 0.0006592 0.22096 0.20354 0 0.032939 0.0389 0 1.099 0.34142 0.099736 0.013129 6.0242 0.081949 0.00010128 0.80815 0.0065993 0.0073943 0.0016061 0.98402 0.98939 3.4946e-006 1.3979e-005 0.14273 0.70552 0.78046 0.0015092 0.79489 0.46546 0.0020289 0.42251 1.3691 1.3653 16.0057 144.9658 0.00037337 -84.7692 0.18595
3.29 0.98806 5.5044e-005 3.8182 0.012004 4.3149e-005 0.0011564 0.22031 0.0006592 0.22097 0.20355 0 0.032938 0.0389 0 1.0991 0.34147 0.099752 0.013131 6.0255 0.08196 0.00010129 0.80814 0.0066 0.0073951 0.0016044 0.98404 0.98943 3.4905e-006 1.3962e-005 0.14274 0.70639 0.78114 0.0015083 0.79609 0.46565 0.0020278 0.42252 1.3709 1.3672 16.0057 144.9658 0.00037237 -84.7758 0.18695
3.291 0.98806 5.5044e-005 3.8182 0.012004 4.3162e-005 0.0011564 0.22033 0.0006592 0.22098 0.20356 0 0.032938 0.0389 0 1.0992 0.34151 0.099768 0.013133 6.0267 0.081971 0.00010131 0.80813 0.0066007 0.0073959 0.0016026 0.98407 0.98946 3.4865e-006 1.3946e-005 0.14274 0.70725 0.78182 0.0015074 0.79728 0.46583 0.0020267 0.42252 1.3727 1.369 16.0058 144.9659 0.00037139 -84.7823 0.18795
3.292 0.98806 5.5044e-005 3.8182 0.012004 4.3175e-005 0.0011564 0.22034 0.0006592 0.22099 0.20358 0 0.032937 0.0389 0 1.0993 0.34156 0.099784 0.013135 6.028 0.081982 0.00010132 0.80812 0.0066015 0.0073966 0.0016009 0.98409 0.9895 3.4825e-006 1.393e-005 0.14275 0.70811 0.78249 0.0015066 0.79847 0.46601 0.0020256 0.42253 1.3746 1.3709 16.0058 144.9659 0.00037041 -84.7887 0.18895
3.293 0.98806 5.5044e-005 3.8182 0.012004 4.3188e-005 0.0011564 0.22035 0.0006592 0.221 0.20359 0 0.032936 0.0389 0 1.0994 0.3416 0.0998 0.013136 6.0293 0.081992 0.00010134 0.80811 0.0066022 0.0073974 0.0015992 0.98411 0.98953 3.4786e-006 1.3915e-005 0.14276 0.70896 0.78316 0.0015058 0.79965 0.46619 0.0020245 0.42253 1.3764 1.3727 16.0059 144.9659 0.00036943 -84.7951 0.18995
3.294 0.98806 5.5044e-005 3.8182 0.012004 4.3201e-005 0.0011564 0.22036 0.0006592 0.22102 0.2036 0 0.032936 0.0389 0 1.0995 0.34165 0.099816 0.013138 6.0306 0.082003 0.00010135 0.8081 0.0066029 0.0073982 0.0015975 0.98414 0.98957 3.4747e-006 1.3899e-005 0.14276 0.70982 0.78382 0.001505 0.80082 0.46637 0.0020234 0.42254 1.3782 1.3745 16.0059 144.9659 0.00036846 -84.8015 0.19095
3.295 0.98806 5.5044e-005 3.8182 0.012004 4.3214e-005 0.0011564 0.22037 0.0006592 0.22103 0.20361 0 0.032935 0.0389 0 1.0996 0.3417 0.099832 0.01314 6.0318 0.082014 0.00010137 0.80809 0.0066036 0.007399 0.0015958 0.98416 0.9896 3.4708e-006 1.3884e-005 0.14277 0.71067 0.78449 0.0015042 0.80199 0.46655 0.0020223 0.42255 1.38 1.3763 16.006 144.9659 0.00036749 -84.8078 0.19195
3.296 0.98806 5.5044e-005 3.8182 0.012004 4.3227e-005 0.0011564 0.22039 0.0006592 0.22104 0.20362 0 0.032935 0.0389 0 1.0997 0.34174 0.099848 0.013142 6.0331 0.082025 0.00010138 0.80808 0.0066043 0.0073997 0.0015941 0.98418 0.98963 3.467e-006 1.3868e-005 0.14277 0.71151 0.78514 0.0015034 0.80316 0.46673 0.0020212 0.42255 1.3818 1.3782 16.006 144.9659 0.00036653 -84.814 0.19295
3.297 0.98806 5.5043e-005 3.8182 0.012004 4.324e-005 0.0011564 0.2204 0.0006592 0.22105 0.20363 0 0.032934 0.0389 0 1.0998 0.34179 0.099865 0.013143 6.0344 0.082036 0.0001014 0.80807 0.0066051 0.0074005 0.0015924 0.98421 0.98966 3.4631e-006 1.3853e-005 0.14278 0.71236 0.7858 0.0015026 0.80431 0.46691 0.0020201 0.42256 1.3836 1.38 16.0061 144.9659 0.00036557 -84.8202 0.19395
3.298 0.98806 5.5043e-005 3.8182 0.012004 4.3253e-005 0.0011564 0.22041 0.0006592 0.22106 0.20364 0 0.032933 0.0389 0 1.0999 0.34183 0.099881 0.013145 6.0357 0.082047 0.00010141 0.80805 0.0066058 0.0074013 0.0015908 0.98423 0.98969 3.4594e-006 1.3838e-005 0.14279 0.7132 0.78645 0.0015018 0.80546 0.46709 0.0020191 0.42256 1.3854 1.3818 16.0061 144.966 0.00036462 -84.8264 0.19495
3.299 0.98806 5.5043e-005 3.8182 0.012004 4.3266e-005 0.0011564 0.22042 0.0006592 0.22108 0.20365 0 0.032933 0.0389 0 1.1 0.34188 0.099897 0.013147 6.0369 0.082058 0.00010143 0.80804 0.0066065 0.007402 0.0015891 0.98425 0.98971 3.4556e-006 1.3823e-005 0.14279 0.71404 0.78709 0.001501 0.80661 0.46727 0.002018 0.42257 1.3872 1.3836 16.0061 144.966 0.00036367 -84.8325 0.19595
3.3 0.98806 5.5043e-005 3.8182 0.012004 4.3279e-005 0.0011564 0.22043 0.0006592 0.22109 0.20367 0 0.032932 0.0389 0 1.1001 0.34193 0.099913 0.013148 6.0382 0.082069 0.00010144 0.80803 0.0066072 0.0074028 0.0015875 0.98427 0.98974 3.4519e-006 1.3808e-005 0.1428 0.71488 0.78774 0.0015002 0.80775 0.46745 0.002017 0.42258 1.389 1.3854 16.0062 144.966 0.00036273 -84.8386 0.19695
3.301 0.98806 5.5043e-005 3.8182 0.012004 4.3293e-005 0.0011564 0.22044 0.0006592 0.2211 0.20368 0 0.032932 0.0389 0 1.1002 0.34197 0.099929 0.01315 6.0395 0.082079 0.00010146 0.80802 0.006608 0.0074036 0.0015859 0.98429 0.98977 3.4483e-006 1.3793e-005 0.1428 0.71571 0.78837 0.0014994 0.80888 0.46763 0.0020159 0.42258 1.3908 1.3872 16.0062 144.966 0.00036179 -84.8446 0.19795
3.302 0.98806 5.5043e-005 3.8182 0.012004 4.3306e-005 0.0011564 0.22046 0.0006592 0.22111 0.20369 0 0.032931 0.0389 0 1.1003 0.34202 0.099945 0.013152 6.0408 0.08209 0.00010147 0.80801 0.0066087 0.0074044 0.0015843 0.98432 0.98979 3.4446e-006 1.3779e-005 0.14281 0.71654 0.78901 0.0014986 0.81 0.46781 0.0020149 0.42259 1.3926 1.389 16.0063 144.966 0.00036086 -84.8505 0.19895
3.303 0.98806 5.5043e-005 3.8182 0.012004 4.3319e-005 0.0011564 0.22047 0.0006592 0.22112 0.2037 0 0.03293 0.0389 0 1.1004 0.34206 0.099961 0.013154 6.042 0.082101 0.00010148 0.808 0.0066094 0.0074051 0.0015827 0.98434 0.98982 3.441e-006 1.3764e-005 0.14281 0.71737 0.78964 0.0014978 0.81112 0.46799 0.0020139 0.4226 1.3944 1.3908 16.0063 144.966 0.00035993 -84.8565 0.19995
3.304 0.98806 5.5043e-005 3.8182 0.012004 4.3332e-005 0.0011564 0.22048 0.0006592 0.22113 0.20371 0 0.03293 0.0389 0 1.1005 0.34211 0.099977 0.013155 6.0433 0.082112 0.0001015 0.80799 0.0066101 0.0074059 0.0015812 0.98436 0.98984 3.4374e-006 1.375e-005 0.14282 0.7182 0.79027 0.001497 0.81224 0.46817 0.0020129 0.4226 1.3961 1.3926 16.0064 144.966 0.000359 -84.8624 0.20095
3.305 0.98806 5.5043e-005 3.8182 0.012004 4.3345e-005 0.0011564 0.22049 0.0006592 0.22115 0.20372 0 0.032929 0.0389 0 1.1006 0.34216 0.099994 0.013157 6.0446 0.082123 0.00010151 0.80798 0.0066109 0.0074067 0.0015797 0.98438 0.98986 3.4339e-006 1.3736e-005 0.14283 0.71903 0.79089 0.0014963 0.81335 0.46835 0.0020119 0.42261 1.3979 1.3944 16.0064 144.9661 0.00035808 -84.8682 0.20195
3.306 0.98806 5.5043e-005 3.8182 0.012004 4.3358e-005 0.0011565 0.2205 0.0006592 0.22116 0.20373 0 0.032929 0.0389 0 1.1007 0.3422 0.10001 0.013159 6.0459 0.082134 0.00010153 0.80797 0.0066116 0.0074074 0.0015782 0.9844 0.98988 3.4304e-006 1.3722e-005 0.14283 0.71985 0.79151 0.0014955 0.81445 0.46853 0.0020109 0.42261 1.3997 1.3961 16.0064 144.9661 0.00035717 -84.874 0.20295
3.307 0.98806 5.5043e-005 3.8182 0.012004 4.3371e-005 0.0011565 0.22052 0.0006592 0.22117 0.20374 0 0.032928 0.0389 0 1.1008 0.34225 0.10003 0.013161 6.0472 0.082145 0.00010154 0.80796 0.0066123 0.0074082 0.0015767 0.98442 0.98991 3.4269e-006 1.3708e-005 0.14284 0.72067 0.79213 0.0014947 0.81554 0.46872 0.0020099 0.42262 1.4014 1.3979 16.0065 144.9661 0.00035626 -84.8797 0.20395
3.308 0.98806 5.5043e-005 3.8182 0.012004 4.3384e-005 0.0011565 0.22053 0.0006592 0.22118 0.20375 0 0.032927 0.0389 0 1.1009 0.34229 0.10004 0.013162 6.0484 0.082155 0.00010156 0.80795 0.006613 0.007409 0.0015753 0.98444 0.98993 3.4234e-006 1.3694e-005 0.14284 0.72148 0.79274 0.0014939 0.81663 0.4689 0.002009 0.42263 1.4032 1.3997 16.0065 144.9661 0.00035535 -84.8854 0.20495
3.309 0.98806 5.5043e-005 3.8182 0.012004 4.3397e-005 0.0011565 0.22054 0.0006592 0.22119 0.20377 0 0.032927 0.0389 0 1.101 0.34234 0.10006 0.013164 6.0497 0.082166 0.00010157 0.80794 0.0066137 0.0074097 0.0015738 0.98446 0.98995 3.42e-006 1.368e-005 0.14285 0.7223 0.79335 0.0014932 0.81772 0.46908 0.002008 0.42264 1.4049 1.4014 16.0066 144.9661 0.00035445 -84.8911 0.20595
3.31 0.98806 5.5043e-005 3.8182 0.012004 4.341e-005 0.0011565 0.22055 0.0006592 0.22121 0.20378 0 0.032926 0.0389 0 1.1011 0.34239 0.10007 0.013166 6.051 0.082177 0.00010159 0.80792 0.0066145 0.0074105 0.0015724 0.98448 0.98997 3.4166e-006 1.3667e-005 0.14286 0.72311 0.79396 0.0014924 0.8188 0.46926 0.002007 0.42264 1.4067 1.4032 16.0066 144.9661 0.00035355 -84.8967 0.20695
3.311 0.98806 5.5043e-005 3.8182 0.012004 4.3423e-005 0.0011565 0.22056 0.0006592 0.22122 0.20379 0 0.032925 0.0389 0 1.1012 0.34243 0.10009 0.013168 6.0523 0.082188 0.0001016 0.80791 0.0066152 0.0074113 0.0015709 0.9845 0.98999 3.4132e-006 1.3653e-005 0.14286 0.72392 0.79456 0.0014917 0.81987 0.46944 0.0020061 0.42265 1.4084 1.405 16.0066 144.9661 0.00035266 -84.9023 0.20795
3.312 0.98806 5.5042e-005 3.8182 0.012004 4.3436e-005 0.0011565 0.22057 0.0006592 0.22123 0.2038 0 0.032925 0.0389 0 1.1013 0.34248 0.10011 0.013169 6.0536 0.082199 0.00010162 0.8079 0.0066159 0.0074121 0.0015695 0.98452 0.99001 3.4099e-006 1.364e-005 0.14287 0.72473 0.79516 0.001491 0.82094 0.46962 0.0020051 0.42266 1.4102 1.4067 16.0067 144.9662 0.00035177 -84.9078 0.20895
3.313 0.98806 5.5042e-005 3.8182 0.012004 4.3449e-005 0.0011565 0.22059 0.0006592 0.22124 0.20381 0 0.032924 0.0389 0 1.1014 0.34252 0.10012 0.013171 6.0549 0.08221 0.00010163 0.80789 0.0066166 0.0074128 0.001568 0.98454 0.99002 3.4066e-006 1.3627e-005 0.14287 0.72553 0.79575 0.0014903 0.822 0.4698 0.0020042 0.42266 1.4119 1.4085 16.0067 144.9662 0.00035088 -84.9133 0.20995
3.314 0.98806 5.5042e-005 3.8182 0.012004 4.3462e-005 0.0011565 0.2206 0.0006592 0.22125 0.20382 0 0.032924 0.0389 0 1.1015 0.34257 0.10014 0.013173 6.0561 0.082221 0.00010165 0.80788 0.0066174 0.0074136 0.0015666 0.98456 0.99004 3.4033e-006 1.3613e-005 0.14288 0.72633 0.79634 0.0014896 0.82305 0.46998 0.0020033 0.42267 1.4136 1.4102 16.0068 144.9662 0.00035 -84.9188 0.21095
3.315 0.98806 5.5042e-005 3.8182 0.012004 4.3475e-005 0.0011565 0.22061 0.0006592 0.22126 0.20383 0 0.032923 0.0389 0 1.1016 0.34262 0.10015 0.013175 6.0574 0.082231 0.00010166 0.80787 0.0066181 0.0074144 0.0015651 0.98458 0.99006 3.4e-006 1.36e-005 0.14288 0.72713 0.79693 0.0014889 0.8241 0.47016 0.0020023 0.42268 1.4154 1.4119 16.0068 144.9662 0.00034913 -84.9242 0.21195
3.316 0.98806 5.5042e-005 3.8182 0.012004 4.3488e-005 0.0011565 0.22062 0.0006592 0.22128 0.20384 0 0.032922 0.0389 0 1.1017 0.34266 0.10017 0.013176 6.0587 0.082242 0.00010168 0.80786 0.0066188 0.0074151 0.0015637 0.9846 0.99008 3.3968e-006 1.3587e-005 0.14289 0.72793 0.79752 0.0014883 0.82515 0.47034 0.0020014 0.42268 1.4171 1.4137 16.0068 144.9662 0.00034826 -84.9295 0.21295
3.317 0.98806 5.5042e-005 3.8182 0.012004 4.3501e-005 0.0011565 0.22063 0.0006592 0.22129 0.20385 0 0.032922 0.0389 0 1.1018 0.34271 0.10019 0.013178 6.06 0.082253 0.00010169 0.80785 0.0066195 0.0074159 0.0015623 0.98462 0.99009 3.3936e-006 1.3575e-005 0.1429 0.72872 0.7981 0.0014876 0.82618 0.47052 0.0020005 0.42269 1.4188 1.4154 16.0069 144.9662 0.00034739 -84.9349 0.21395
3.318 0.98806 5.5042e-005 3.8182 0.012004 4.3514e-005 0.0011565 0.22064 0.0006592 0.2213 0.20387 0 0.032921 0.0389 0 1.1019 0.34275 0.1002 0.01318 6.0613 0.082264 0.00010171 0.80784 0.0066203 0.0074167 0.0015609 0.98463 0.99011 3.3904e-006 1.3562e-005 0.1429 0.72952 0.79868 0.0014869 0.82722 0.4707 0.0019996 0.4227 1.4205 1.4171 16.0069 144.9662 0.00034653 -84.9401 0.21495
3.319 0.98806 5.5042e-005 3.8182 0.012004 4.3527e-005 0.0011565 0.22066 0.0006592 0.22131 0.20388 0 0.032921 0.0389 0 1.102 0.3428 0.10022 0.013182 6.0626 0.082275 0.00010172 0.80783 0.006621 0.0074175 0.0015595 0.98465 0.99013 3.3873e-006 1.3549e-005 0.14291 0.73031 0.79926 0.0014863 0.82824 0.47088 0.0019987 0.42271 1.4222 1.4189 16.007 144.9663 0.00034567 -84.9454 0.21595
3.32 0.98806 5.5042e-005 3.8182 0.012004 4.354e-005 0.0011565 0.22067 0.0006592 0.22132 0.20389 0 0.03292 0.0389 0 1.1021 0.34285 0.10024 0.013183 6.0638 0.082286 0.00010174 0.80782 0.0066217 0.0074182 0.0015581 0.98467 0.99014 3.3842e-006 1.3537e-005 0.14291 0.73109 0.79983 0.0014856 0.82926 0.47106 0.0019978 0.42271 1.4239 1.4206 16.007 144.9663 0.00034481 -84.9506 0.21695
3.321 0.98806 5.5042e-005 3.8182 0.012004 4.3553e-005 0.0011565 0.22068 0.0006592 0.22133 0.2039 0 0.032919 0.0389 0 1.1022 0.34289 0.10025 0.013185 6.0651 0.082296 0.00010175 0.80781 0.0066224 0.007419 0.0015568 0.98469 0.99016 3.3811e-006 1.3525e-005 0.14292 0.73188 0.8004 0.0014849 0.83028 0.47124 0.001997 0.42272 1.4256 1.4223 16.007 144.9663 0.00034396 -84.9558 0.21795
3.322 0.98806 5.5042e-005 3.8182 0.012004 4.3566e-005 0.0011565 0.22069 0.0006592 0.22134 0.20391 0 0.032919 0.0389 0 1.1023 0.34294 0.10027 0.013187 6.0664 0.082307 0.00010177 0.80779 0.0066232 0.0074198 0.0015555 0.98471 0.99017 3.378e-006 1.3512e-005 0.14293 0.73266 0.80096 0.0014843 0.83129 0.47142 0.0019961 0.42273 1.4273 1.424 16.0071 144.9663 0.00034312 -84.9609 0.21895
3.323 0.98806 5.5042e-005 3.8182 0.012004 4.3579e-005 0.0011565 0.2207 0.0006592 0.22136 0.20392 0 0.032918 0.0389 0 1.1024 0.34298 0.10028 0.013188 6.0677 0.082318 0.00010178 0.80778 0.0066239 0.0074205 0.0015542 0.98473 0.99019 3.375e-006 1.35e-005 0.14293 0.73344 0.80153 0.0014836 0.83229 0.4716 0.0019952 0.42274 1.429 1.4257 16.0071 144.9663 0.00034228 -84.966 0.21995
3.324 0.98806 5.5042e-005 3.8182 0.012004 4.3592e-005 0.0011565 0.22071 0.0006592 0.22137 0.20393 0 0.032918 0.0389 0 1.1025 0.34303 0.1003 0.01319 6.069 0.082329 0.0001018 0.80777 0.0066246 0.0074213 0.0015529 0.98474 0.9902 3.3719e-006 1.3488e-005 0.14294 0.73422 0.80209 0.0014829 0.83329 0.47178 0.0019944 0.42274 1.4307 1.4274 16.0071 144.9663 0.00034144 -84.971 0.22095
3.325 0.98806 5.5042e-005 3.8182 0.012004 4.3606e-005 0.0011565 0.22072 0.0006592 0.22138 0.20394 0 0.032917 0.0389 0 1.1026 0.34308 0.10032 0.013192 6.0703 0.08234 0.00010181 0.80776 0.0066253 0.0074221 0.0015516 0.98476 0.99022 3.369e-006 1.3476e-005 0.14294 0.73499 0.80264 0.0014822 0.83428 0.47196 0.0019935 0.42275 1.4324 1.4291 16.0072 144.9664 0.0003406 -84.976 0.22195
3.326 0.98806 5.5041e-005 3.8182 0.012004 4.3619e-005 0.0011565 0.22074 0.0006592 0.22139 0.20395 0 0.032916 0.0389 0 1.1027 0.34312 0.10033 0.013194 6.0716 0.082351 0.00010182 0.80775 0.006626 0.0074229 0.0015503 0.98478 0.99023 3.366e-006 1.3464e-005 0.14295 0.73577 0.8032 0.0014815 0.83527 0.47214 0.0019927 0.42276 1.4341 1.4308 16.0072 144.9664 0.00033977 -84.981 0.22295
3.327 0.98806 5.5041e-005 3.8182 0.012004 4.3632e-005 0.0011565 0.22075 0.0006592 0.2214 0.20396 0 0.032916 0.0389 0 1.1028 0.34317 0.10035 0.013195 6.0729 0.082362 0.00010184 0.80774 0.0066268 0.0074236 0.0015491 0.9848 0.99025 3.3631e-006 1.3452e-005 0.14296 0.73654 0.80375 0.0014809 0.83625 0.47232 0.0019918 0.42277 1.4358 1.4325 16.0072 144.9664 0.00033895 -84.9859 0.22395
3.328 0.98806 5.5041e-005 3.8182 0.012004 4.3645e-005 0.0011565 0.22076 0.0006592 0.22141 0.20397 0 0.032915 0.0389 0 1.1029 0.34321 0.10036 0.013197 6.0741 0.082372 0.00010185 0.80773 0.0066275 0.0074244 0.0015478 0.98481 0.99026 3.3601e-006 1.3441e-005 0.14296 0.7373 0.8043 0.0014802 0.83723 0.4725 0.001991 0.42278 1.4374 1.4342 16.0073 144.9664 0.00033813 -84.9908 0.22495
3.329 0.98806 5.5041e-005 3.8182 0.012004 4.3658e-005 0.0011565 0.22077 0.0006592 0.22143 0.20399 0 0.032915 0.0389 0 1.103 0.34326 0.10038 0.013199 6.0754 0.082383 0.00010187 0.80772 0.0066282 0.0074252 0.0015466 0.98483 0.99027 3.3572e-006 1.3429e-005 0.14297 0.73807 0.80484 0.0014796 0.8382 0.47268 0.0019902 0.42278 1.4391 1.4358 16.0073 144.9664 0.00033731 -84.9957 0.22595
3.33 0.98806 5.5041e-005 3.8182 0.012004 4.3671e-005 0.0011565 0.22078 0.0006592 0.22144 0.204 0 0.032914 0.0389 0 1.1031 0.34331 0.1004 0.013201 6.0767 0.082394 0.00010188 0.80771 0.0066289 0.0074259 0.0015454 0.98485 0.99029 3.3544e-006 1.3418e-005 0.14297 0.73883 0.80538 0.0014789 0.83917 0.47286 0.0019894 0.42279 1.4408 1.4375 16.0073 144.9664 0.00033649 -85.0005 0.22695
3.331 0.98806 5.5041e-005 3.8182 0.012004 4.3684e-005 0.0011565 0.22079 0.0006592 0.22145 0.20401 0 0.032914 0.0389 0 1.1032 0.34335 0.10041 0.013202 6.078 0.082405 0.0001019 0.8077 0.0066297 0.0074267 0.0015442 0.98486 0.9903 3.3515e-006 1.3406e-005 0.14298 0.73959 0.80592 0.0014783 0.84013 0.47304 0.0019886 0.4228 1.4424 1.4392 16.0074 144.9664 0.00033568 -85.0053 0.22795
3.332 0.98806 5.5041e-005 3.8182 0.012004 4.3697e-005 0.0011565 0.22081 0.0006592 0.22146 0.20402 0 0.032913 0.0389 0 1.1033 0.3434 0.10043 0.013204 6.0793 0.082416 0.00010191 0.80769 0.0066304 0.0074275 0.0015429 0.98488 0.99031 3.3487e-006 1.3395e-005 0.14298 0.74035 0.80646 0.0014777 0.84108 0.47322 0.0019878 0.42281 1.4441 1.4409 16.0074 144.9665 0.00033488 -85.0101 0.22895
3.333 0.98806 5.5041e-005 3.8182 0.012004 4.371e-005 0.0011565 0.22082 0.0006592 0.22147 0.20403 0 0.032912 0.0389 0 1.1034 0.34344 0.10045 0.013206 6.0806 0.082427 0.00010193 0.80768 0.0066311 0.0074282 0.0015417 0.9849 0.99032 3.3459e-006 1.3384e-005 0.14299 0.74111 0.80699 0.0014771 0.84203 0.47339 0.001987 0.42282 1.4457 1.4425 16.0074 144.9665 0.00033408 -85.0148 0.22995
3.334 0.98806 5.5041e-005 3.8182 0.012004 4.3723e-005 0.0011565 0.22083 0.0006592 0.22148 0.20404 0 0.032912 0.0389 0 1.1035 0.34349 0.10046 0.013208 6.0819 0.082437 0.00010194 0.80766 0.0066318 0.007429 0.0015405 0.98491 0.99034 3.3432e-006 1.3373e-005 0.143 0.74186 0.80752 0.0014765 0.84298 0.47357 0.0019862 0.42282 1.4474 1.4442 16.0075 144.9665 0.00033328 -85.0195 0.23095
3.335 0.98806 5.5041e-005 3.8182 0.012004 4.3736e-005 0.0011565 0.22084 0.0006592 0.22149 0.20405 0 0.032911 0.0389 0 1.1036 0.34354 0.10048 0.013209 6.0832 0.082448 0.00010196 0.80765 0.0066326 0.0074298 0.0015393 0.98493 0.99035 3.3404e-006 1.3362e-005 0.143 0.74261 0.80805 0.0014759 0.84392 0.47375 0.0019854 0.42283 1.449 1.4458 16.0075 144.9665 0.00033248 -85.0241 0.23195
3.336 0.98806 5.5041e-005 3.8182 0.012004 4.3749e-005 0.0011565 0.22085 0.0006592 0.22151 0.20406 0 0.032911 0.0389 0 1.1037 0.34358 0.10049 0.013211 6.0845 0.082459 0.00010197 0.80764 0.0066333 0.0074306 0.0015381 0.98494 0.99036 3.3377e-006 1.3351e-005 0.14301 0.74336 0.80857 0.0014754 0.84485 0.47393 0.0019846 0.42284 1.4507 1.4475 16.0075 144.9665 0.00033169 -85.0287 0.23295
3.337 0.98806 5.5041e-005 3.8182 0.012004 4.3762e-005 0.0011565 0.22086 0.0006592 0.22152 0.20407 0 0.03291 0.0389 0 1.1038 0.34363 0.10051 0.013213 6.0858 0.08247 0.00010199 0.80763 0.006634 0.0074313 0.0015369 0.98496 0.99037 3.335e-006 1.334e-005 0.14301 0.74411 0.80909 0.0014748 0.84578 0.47411 0.0019838 0.42285 1.4523 1.4491 16.0076 144.9665 0.00033091 -85.0333 0.23395
3.338 0.98806 5.5041e-005 3.8182 0.012004 4.3775e-005 0.0011565 0.22087 0.0006592 0.22153 0.20408 0 0.032909 0.0389 0 1.1039 0.34367 0.10053 0.013215 6.0871 0.082481 0.000102 0.80762 0.0066347 0.0074321 0.0015357 0.98498 0.99038 3.3323e-006 1.3329e-005 0.14302 0.74486 0.80961 0.0014743 0.8467 0.47429 0.0019831 0.42286 1.4539 1.4508 16.0076 144.9666 0.00033012 -85.0379 0.23495
3.339 0.98806 5.5041e-005 3.8182 0.012004 4.3788e-005 0.0011565 0.22089 0.0006592 0.22154 0.20409 0 0.032909 0.0389 0 1.104 0.34372 0.10054 0.013216 6.0883 0.082492 0.00010202 0.80761 0.0066354 0.0074329 0.0015345 0.98499 0.9904 3.3296e-006 1.3319e-005 0.14303 0.7456 0.81013 0.0014737 0.84762 0.47447 0.0019823 0.42287 1.4555 1.4524 16.0076 144.9666 0.00032935 -85.0424 0.23595
3.34 0.98806 5.5041e-005 3.8182 0.012004 4.3801e-005 0.0011565 0.2209 0.0006592 0.22155 0.20411 0 0.032908 0.0389 0 1.1041 0.34377 0.10056 0.013218 6.0896 0.082502 0.00010203 0.8076 0.0066362 0.0074336 0.0015334 0.98501 0.99041 3.327e-006 1.3308e-005 0.14303 0.74634 0.81064 0.0014731 0.84853 0.47465 0.0019816 0.42287 1.4572 1.454 16.0077 144.9666 0.00032857 -85.0468 0.23695
3.341 0.98806 5.504e-005 3.8182 0.012004 4.3814e-005 0.0011565 0.22091 0.0006592 0.22156 0.20412 0 0.032908 0.0389 0 1.1042 0.34381 0.10057 0.01322 6.0909 0.082513 0.00010205 0.80759 0.0066369 0.0074344 0.0015322 0.98502 0.99042 3.3244e-006 1.3298e-005 0.14304 0.74708 0.81115 0.0014726 0.84944 0.47483 0.0019808 0.42288 1.4588 1.4557 16.0077 144.9666 0.0003278 -85.0513 0.23795
3.342 0.98806 5.504e-005 3.8182 0.012004 4.3827e-005 0.0011565 0.22092 0.0006592 0.22157 0.20413 0 0.032907 0.0389 0 1.1043 0.34386 0.10059 0.013222 6.0922 0.082524 0.00010206 0.80758 0.0066376 0.0074352 0.0015311 0.98504 0.99043 3.3218e-006 1.3287e-005 0.14304 0.74781 0.81166 0.001472 0.85035 0.47501 0.0019801 0.42289 1.4604 1.4573 16.0077 144.9666 0.00032703 -85.0557 0.23895
3.343 0.98806 5.504e-005 3.8182 0.012004 4.384e-005 0.0011565 0.22093 0.0006592 0.22159 0.20414 0 0.032906 0.0389 0 1.1044 0.3439 0.10061 0.013223 6.0935 0.082535 0.00010208 0.80757 0.0066383 0.007436 0.00153 0.98505 0.99044 3.3192e-006 1.3277e-005 0.14305 0.74854 0.81216 0.0014714 0.85124 0.47519 0.0019793 0.4229 1.462 1.4589 16.0078 144.9666 0.00032627 -85.0601 0.23995
3.344 0.98806 5.504e-005 3.8182 0.012004 4.3853e-005 0.0011565 0.22094 0.0006592 0.2216 0.20415 0 0.032906 0.0389 0 1.1045 0.34395 0.10062 0.013225 6.0948 0.082546 0.00010209 0.80756 0.0066391 0.0074367 0.0015289 0.98507 0.99045 3.3167e-006 1.3267e-005 0.14305 0.74928 0.81267 0.0014708 0.85214 0.47537 0.0019786 0.42291 1.4636 1.4605 16.0078 144.9666 0.00032551 -85.0644 0.24095
3.345 0.98806 5.504e-005 3.8182 0.012004 4.3866e-005 0.0011565 0.22095 0.0006592 0.22161 0.20416 0 0.032905 0.0389 0 1.1046 0.344 0.10064 0.013227 6.0961 0.082557 0.00010211 0.80755 0.0066398 0.0074375 0.0015278 0.98508 0.99046 3.3141e-006 1.3257e-005 0.14306 0.75 0.81317 0.0014703 0.85302 0.47555 0.0019779 0.42292 1.4652 1.4621 16.0078 144.9667 0.00032475 -85.0687 0.24195
3.346 0.98806 5.504e-005 3.8182 0.012004 4.3879e-005 0.0011565 0.22097 0.0006592 0.22162 0.20417 0 0.032905 0.0389 0 1.1047 0.34404 0.10065 0.013228 6.0974 0.082567 0.00010212 0.80753 0.0066405 0.0074383 0.0015268 0.9851 0.99047 3.3116e-006 1.3247e-005 0.14307 0.75073 0.81366 0.0014697 0.85391 0.47573 0.0019772 0.42293 1.4668 1.4638 16.0079 144.9667 0.00032399 -85.073 0.24295
3.347 0.98806 5.504e-005 3.8182 0.012004 4.3892e-005 0.0011565 0.22098 0.0006592 0.22163 0.20418 0 0.032904 0.0389 0 1.1047 0.34409 0.10067 0.01323 6.0987 0.082578 0.00010213 0.80752 0.0066412 0.007439 0.0015257 0.98511 0.99048 3.3091e-006 1.3237e-005 0.14307 0.75146 0.81416 0.0014691 0.85478 0.47591 0.0019764 0.42294 1.4684 1.4654 16.0079 144.9667 0.00032325 -85.0773 0.24395
3.348 0.98806 5.504e-005 3.8182 0.012004 4.3905e-005 0.0011565 0.22099 0.0006592 0.22164 0.20419 0 0.032903 0.0389 0 1.1048 0.34413 0.10069 0.013232 6.1 0.082589 0.00010215 0.80751 0.006642 0.0074398 0.0015247 0.98512 0.99049 3.3067e-006 1.3227e-005 0.14308 0.75218 0.81465 0.0014685 0.85566 0.47608 0.0019757 0.42294 1.47 1.467 16.0079 144.9667 0.0003225 -85.0815 0.24495
3.349 0.98806 5.504e-005 3.8182 0.012004 4.3918e-005 0.0011565 0.221 0.0006592 0.22165 0.2042 0 0.032903 0.0389 0 1.1049 0.34418 0.1007 0.013234 6.1013 0.0826 0.00010216 0.8075 0.0066427 0.0074406 0.0015236 0.98514 0.9905 3.3042e-006 1.3217e-005 0.14308 0.7529 0.81514 0.001468 0.85652 0.47626 0.001975 0.42295 1.4716 1.4686 16.0079 144.9667 0.00032176 -85.0857 0.24595
3.35 0.98806 5.504e-005 3.8182 0.012004 4.3932e-005 0.0011565 0.22101 0.0006592 0.22167 0.20421 0 0.032902 0.0389 0 1.105 0.34423 0.10072 0.013235 6.1026 0.082611 0.00010218 0.80749 0.0066434 0.0074414 0.0015226 0.98515 0.99051 3.3018e-006 1.3207e-005 0.14309 0.75361 0.81563 0.0014674 0.85739 0.47644 0.0019743 0.42296 1.4732 1.4701 16.008 144.9667 0.00032102 -85.0898 0.24695
3.351 0.98806 5.504e-005 3.8182 0.012004 4.3945e-005 0.0011565 0.22102 0.0006592 0.22168 0.20422 0 0.032902 0.0389 0 1.1051 0.34427 0.10074 0.013237 6.1039 0.082622 0.00010219 0.80748 0.0066441 0.0074421 0.0015215 0.98517 0.99052 3.2994e-006 1.3198e-005 0.1431 0.75433 0.81611 0.0014669 0.85824 0.47662 0.0019736 0.42297 1.4747 1.4717 16.008 144.9668 0.00032028 -85.0939 0.24795
3.352 0.98806 5.504e-005 3.8182 0.012004 4.3958e-005 0.0011565 0.22103 0.0006592 0.22169 0.20423 0 0.032901 0.0389 0 1.1052 0.34432 0.10075 0.013239 6.1052 0.082632 0.00010221 0.80747 0.0066448 0.0074429 0.0015205 0.98518 0.99053 3.297e-006 1.3188e-005 0.1431 0.75504 0.81659 0.0014664 0.8591 0.4768 0.0019729 0.42298 1.4763 1.4733 16.008 144.9668 0.00031955 -85.098 0.24895
3.353 0.98806 5.504e-005 3.8182 0.012003 4.3971e-005 0.0011565 0.22104 0.0006592 0.2217 0.20425 0 0.032901 0.0389 0 1.1053 0.34436 0.10077 0.013241 6.1065 0.082643 0.00010222 0.80746 0.0066456 0.0074437 0.0015195 0.98519 0.99054 3.2946e-006 1.3179e-005 0.14311 0.75575 0.81707 0.0014658 0.85994 0.47698 0.0019723 0.42299 1.4779 1.4749 16.008 144.9668 0.00031882 -85.1021 0.24995
3.354 0.98806 5.504e-005 3.8182 0.012003 4.3984e-005 0.0011565 0.22106 0.0006592 0.22171 0.20426 0 0.0329 0.0389 0 1.1054 0.34441 0.10078 0.013242 6.1078 0.082654 0.00010224 0.80745 0.0066463 0.0074444 0.0015184 0.98521 0.99055 3.2923e-006 1.3169e-005 0.14311 0.75646 0.81755 0.0014654 0.86079 0.47716 0.0019716 0.423 1.4795 1.4765 16.0081 144.9668 0.0003181 -85.1061 0.25095
3.355 0.98806 5.5039e-005 3.8182 0.012003 4.3997e-005 0.0011565 0.22107 0.0006592 0.22172 0.20427 0 0.032899 0.0389 0 1.1055 0.34446 0.1008 0.013244 6.1091 0.082665 0.00010225 0.80744 0.006647 0.0074452 0.0015174 0.98522 0.99056 3.29e-006 1.316e-005 0.14312 0.75717 0.81802 0.0014649 0.86163 0.47734 0.0019709 0.42301 1.481 1.478 16.0081 144.9668 0.00031737 -85.1101 0.25195
3.356 0.98806 5.5039e-005 3.8182 0.012003 4.401e-005 0.0011565 0.22108 0.0006592 0.22173 0.20428 0 0.032899 0.0389 0 1.1056 0.3445 0.10082 0.013246 6.1104 0.082676 0.00010227 0.80743 0.0066477 0.007446 0.0015164 0.98524 0.99057 3.2877e-006 1.3151e-005 0.14312 0.75787 0.81849 0.0014644 0.86246 0.47752 0.0019703 0.42302 1.4826 1.4796 16.0081 144.9668 0.00031666 -85.1141 0.25295
3.357 0.98806 5.5039e-005 3.8182 0.012003 4.4023e-005 0.0011565 0.22109 0.0006592 0.22174 0.20429 0 0.032898 0.0389 0 1.1057 0.34455 0.10083 0.013248 6.1117 0.082687 0.00010228 0.80742 0.0066485 0.0074467 0.0015154 0.98525 0.99058 3.2854e-006 1.3142e-005 0.14313 0.75858 0.81896 0.0014639 0.86329 0.47769 0.0019696 0.42303 1.4841 1.4812 16.0082 144.9669 0.00031594 -85.118 0.25395
3.358 0.98806 5.5039e-005 3.8182 0.012003 4.4036e-005 0.0011565 0.2211 0.0006592 0.22176 0.2043 0 0.032898 0.0389 0 1.1058 0.34459 0.10085 0.013249 6.113 0.082697 0.0001023 0.8074 0.0066492 0.0074475 0.0015143 0.98526 0.99059 3.2831e-006 1.3133e-005 0.14314 0.75928 0.81943 0.0014634 0.86411 0.47787 0.0019689 0.42303 1.4857 1.4827 16.0082 144.9669 0.00031523 -85.1219 0.25495
3.359 0.98806 5.5039e-005 3.8182 0.012003 4.4049e-005 0.0011565 0.22111 0.00065921 0.22177 0.20431 0 0.032897 0.0389 0 1.1059 0.34464 0.10086 0.013251 6.1143 0.082708 0.00010231 0.80739 0.0066499 0.0074483 0.0015133 0.98528 0.9906 3.2808e-006 1.3123e-005 0.14314 0.75997 0.81989 0.001463 0.86493 0.47805 0.0019683 0.42304 1.4872 1.4843 16.0082 144.9669 0.00031452 -85.1258 0.25595
3.36 0.98806 5.5039e-005 3.8182 0.012003 4.4062e-005 0.0011565 0.22112 0.00065921 0.22178 0.20432 0 0.032896 0.0389 0 1.106 0.34469 0.10088 0.013253 6.1156 0.082719 0.00010233 0.80738 0.0066506 0.0074491 0.0015123 0.98529 0.99061 3.2786e-006 1.3115e-005 0.14315 0.76067 0.82036 0.0014625 0.86575 0.47823 0.0019676 0.42305 1.4888 1.4858 16.0082 144.9669 0.00031382 -85.1297 0.25695
3.361 0.98806 5.5039e-005 3.8182 0.012003 4.4075e-005 0.0011566 0.22113 0.00065921 0.22179 0.20433 0 0.032896 0.0389 0 1.1061 0.34473 0.1009 0.013254 6.1169 0.08273 0.00010234 0.80737 0.0066514 0.0074498 0.0015114 0.9853 0.99062 3.2764e-006 1.3106e-005 0.14315 0.76136 0.82082 0.001462 0.86656 0.47841 0.001967 0.42306 1.4903 1.4874 16.0083 144.9669 0.00031311 -85.1335 0.25795
3.362 0.98806 5.5039e-005 3.8182 0.012003 4.4088e-005 0.0011566 0.22115 0.00065921 0.2218 0.20434 0 0.032895 0.0389 0 1.1062 0.34478 0.10091 0.013256 6.1182 0.082741 0.00010236 0.80736 0.0066521 0.0074506 0.0015104 0.98531 0.99063 3.2742e-006 1.3097e-005 0.14316 0.76205 0.82127 0.0014615 0.86736 0.47859 0.0019664 0.42307 1.4918 1.4889 16.0083 144.9669 0.00031242 -85.1373 0.25895
3.363 0.98806 5.5039e-005 3.8182 0.012003 4.4101e-005 0.0011566 0.22116 0.00065921 0.22181 0.20435 0 0.032895 0.0389 0 1.1063 0.34482 0.10093 0.013258 6.1195 0.082751 0.00010237 0.80735 0.0066528 0.0074514 0.0015095 0.98533 0.99063 3.272e-006 1.3088e-005 0.14317 0.76274 0.82173 0.0014611 0.86816 0.47877 0.0019657 0.42308 1.4934 1.4905 16.0083 144.967 0.00031172 -85.1411 0.25995
3.364 0.98806 5.5039e-005 3.8182 0.012003 4.4114e-005 0.0011566 0.22117 0.00065921 0.22182 0.20436 0 0.032894 0.0389 0 1.1064 0.34487 0.10094 0.01326 6.1208 0.082762 0.00010239 0.80734 0.0066535 0.0074521 0.0015086 0.98534 0.99064 3.2698e-006 1.3079e-005 0.14317 0.76343 0.82218 0.0014606 0.86896 0.47894 0.0019651 0.42309 1.4949 1.492 16.0083 144.967 0.00031103 -85.1448 0.26095
3.365 0.98806 5.5039e-005 3.8182 0.012003 4.4127e-005 0.0011566 0.22118 0.00065921 0.22183 0.20437 0 0.032894 0.0389 0 1.1065 0.34492 0.10096 0.013261 6.1221 0.082773 0.0001024 0.80733 0.0066542 0.0074529 0.0015077 0.98535 0.99065 3.2677e-006 1.3071e-005 0.14318 0.76412 0.82263 0.0014601 0.86975 0.47912 0.0019645 0.4231 1.4964 1.4935 16.0084 144.967 0.00031034 -85.1485 0.26195
3.366 0.98806 5.5039e-005 3.8182 0.012003 4.414e-005 0.0011566 0.22119 0.00065921 0.22185 0.20438 0 0.032893 0.0389 0 1.1066 0.34496 0.10098 0.013263 6.1234 0.082784 0.00010242 0.80732 0.006655 0.0074537 0.0015067 0.98536 0.99066 3.2655e-006 1.3062e-005 0.14318 0.7648 0.82308 0.0014596 0.87053 0.4793 0.0019639 0.42311 1.4979 1.4951 16.0084 144.967 0.00030966 -85.1522 0.26295
3.367 0.98806 5.5039e-005 3.8182 0.012003 4.4153e-005 0.0011566 0.2212 0.00065921 0.22186 0.20439 0 0.032892 0.0389 0 1.1067 0.34501 0.10099 0.013265 6.1247 0.082795 0.00010243 0.80731 0.0066557 0.0074545 0.0015059 0.98538 0.99067 3.2634e-006 1.3054e-005 0.14319 0.76548 0.82353 0.0014591 0.87132 0.47948 0.0019633 0.42312 1.4994 1.4966 16.0084 144.967 0.00030897 -85.1559 0.26395
3.368 0.98806 5.5039e-005 3.8182 0.012003 4.4166e-005 0.0011566 0.22121 0.00065921 0.22187 0.2044 0 0.032892 0.0389 0 1.1068 0.34505 0.10101 0.013267 6.126 0.082806 0.00010244 0.8073 0.0066564 0.0074552 0.001505 0.98539 0.99068 3.2613e-006 1.3045e-005 0.1432 0.76616 0.82397 0.0014586 0.87209 0.47966 0.0019627 0.42313 1.5009 1.4981 16.0084 144.967 0.00030829 -85.1595 0.26495
3.369 0.98806 5.5039e-005 3.8182 0.012003 4.4179e-005 0.0011566 0.22122 0.00065921 0.22188 0.20442 0 0.032891 0.0389 0 1.1069 0.3451 0.10103 0.013268 6.1273 0.082816 0.00010246 0.80729 0.0066571 0.007456 0.0015041 0.9854 0.99068 3.2593e-006 1.3037e-005 0.1432 0.76683 0.82441 0.0014581 0.87287 0.47984 0.0019621 0.42314 1.5024 1.4996 16.0085 144.967 0.00030762 -85.1631 0.26595
3.37 0.98806 5.5038e-005 3.8182 0.012003 4.4192e-005 0.0011566 0.22124 0.00065921 0.22189 0.20443 0 0.032891 0.0389 0 1.107 0.34515 0.10104 0.01327 6.1286 0.082827 0.00010247 0.80728 0.0066579 0.0074568 0.0015032 0.98541 0.99069 3.2572e-006 1.3029e-005 0.14321 0.76751 0.82485 0.0014576 0.87364 0.48001 0.0019615 0.42315 1.504 1.5011 16.0085 144.9671 0.00030695 -85.1667 0.26695
3.371 0.98806 5.5038e-005 3.8182 0.012003 4.4205e-005 0.0011566 0.22125 0.00065921 0.2219 0.20444 0 0.03289 0.0389 0 1.1071 0.34519 0.10106 0.013272 6.1299 0.082838 0.00010249 0.80726 0.0066586 0.0074575 0.0015023 0.98542 0.9907 3.2552e-006 1.3021e-005 0.14321 0.76818 0.82529 0.0014571 0.8744 0.48019 0.0019609 0.42316 1.5054 1.5026 16.0085 144.9671 0.00030628 -85.1702 0.26795
3.372 0.98806 5.5038e-005 3.8182 0.012003 4.4218e-005 0.0011566 0.22126 0.00065921 0.22191 0.20445 0 0.03289 0.0389 0 1.1072 0.34524 0.10107 0.013274 6.1312 0.082849 0.0001025 0.80725 0.0066593 0.0074583 0.0015014 0.98544 0.99071 3.2531e-006 1.3013e-005 0.14322 0.76885 0.82572 0.0014566 0.87516 0.48037 0.0019603 0.42317 1.5069 1.5042 16.0085 144.9671 0.00030561 -85.1737 0.26895
3.373 0.98806 5.5038e-005 3.8182 0.012003 4.4231e-005 0.0011566 0.22127 0.00065921 0.22192 0.20446 0 0.032889 0.0389 0 1.1073 0.34528 0.10109 0.013275 6.1325 0.08286 0.00010252 0.80724 0.00666 0.0074591 0.0015006 0.98545 0.99072 3.2511e-006 1.3005e-005 0.14322 0.76952 0.82615 0.0014562 0.87592 0.48055 0.0019597 0.42318 1.5084 1.5057 16.0085 144.9671 0.00030495 -85.1772 0.26995
3.374 0.98806 5.5038e-005 3.8182 0.012003 4.4244e-005 0.0011566 0.22128 0.00065921 0.22193 0.20447 0 0.032888 0.0389 0 1.1074 0.34533 0.10111 0.013277 6.1338 0.08287 0.00010253 0.80723 0.0066607 0.0074599 0.0014997 0.98546 0.99073 3.2491e-006 1.2997e-005 0.14323 0.77019 0.82658 0.0014558 0.87667 0.48073 0.0019591 0.42319 1.5099 1.5071 16.0086 144.9671 0.00030429 -85.1807 0.27095
3.375 0.98806 5.5038e-005 3.8182 0.012003 4.4258e-005 0.0011566 0.22129 0.00065921 0.22195 0.20448 0 0.032888 0.0389 0 1.1075 0.34538 0.10112 0.013279 6.1351 0.082881 0.00010255 0.80722 0.0066615 0.0074606 0.0014988 0.98547 0.99073 3.2471e-006 1.2989e-005 0.14324 0.77085 0.82701 0.0014554 0.87741 0.48091 0.0019585 0.4232 1.5114 1.5086 16.0086 144.9671 0.00030363 -85.1842 0.27195
3.376 0.98806 5.5038e-005 3.8182 0.012003 4.4271e-005 0.0011566 0.2213 0.00065921 0.22196 0.20449 0 0.032887 0.0389 0 1.1076 0.34542 0.10114 0.013281 6.1365 0.082892 0.00010256 0.80721 0.0066622 0.0074614 0.0014979 0.98548 0.99074 3.2452e-006 1.2981e-005 0.14324 0.77151 0.82744 0.0014549 0.87815 0.48108 0.001958 0.42321 1.5129 1.5101 16.0086 144.9672 0.00030298 -85.1876 0.27295
3.377 0.98806 5.5038e-005 3.8182 0.012003 4.4284e-005 0.0011566 0.22131 0.00065921 0.22197 0.2045 0 0.032887 0.0389 0 1.1077 0.34547 0.10115 0.013282 6.1378 0.082903 0.00010258 0.8072 0.0066629 0.0074622 0.0014971 0.98549 0.99075 3.2432e-006 1.2973e-005 0.14325 0.77217 0.82786 0.0014545 0.87889 0.48126 0.0019574 0.42322 1.5144 1.5116 16.0086 144.9672 0.00030233 -85.191 0.27395
3.378 0.98806 5.5038e-005 3.8182 0.012003 4.4297e-005 0.0011566 0.22132 0.00065921 0.22198 0.20451 0 0.032886 0.0389 0 1.1078 0.34551 0.10117 0.013284 6.1391 0.082914 0.00010259 0.80719 0.0066636 0.0074629 0.0014962 0.9855 0.99076 3.2413e-006 1.2965e-005 0.14325 0.77283 0.82828 0.0014541 0.87963 0.48144 0.0019569 0.42323 1.5158 1.5131 16.0087 144.9672 0.00030168 -85.1944 0.27495
3.379 0.98806 5.5038e-005 3.8182 0.012003 4.431e-005 0.0011566 0.22133 0.00065921 0.22199 0.20452 0 0.032886 0.0389 0 1.1079 0.34556 0.10119 0.013286 6.1404 0.082925 0.00010261 0.80718 0.0066644 0.0074637 0.0014954 0.98552 0.99076 3.2394e-006 1.2958e-005 0.14326 0.77349 0.8287 0.0014537 0.88036 0.48162 0.0019563 0.42324 1.5173 1.5146 16.0087 144.9672 0.00030103 -85.1977 0.27595
3.38 0.98806 5.5038e-005 3.8182 0.012003 4.4323e-005 0.0011566 0.22135 0.00065921 0.222 0.20453 0 0.032885 0.0389 0 1.108 0.34561 0.1012 0.013287 6.1417 0.082935 0.00010262 0.80717 0.0066651 0.0074645 0.0014945 0.98553 0.99077 3.2375e-006 1.295e-005 0.14327 0.77414 0.82912 0.0014533 0.88108 0.4818 0.0019557 0.42325 1.5187 1.516 16.0087 144.9672 0.00030039 -85.201 0.27695
3.381 0.98806 5.5038e-005 3.8182 0.012003 4.4336e-005 0.0011566 0.22136 0.00065921 0.22201 0.20454 0 0.032884 0.0389 0 1.1081 0.34565 0.10122 0.013289 6.143 0.082946 0.00010264 0.80716 0.0066658 0.0074652 0.0014937 0.98554 0.99078 3.2356e-006 1.2942e-005 0.14327 0.77479 0.82954 0.0014529 0.8818 0.48197 0.0019552 0.42326 1.5202 1.5175 16.0087 144.9673 0.00029975 -85.2043 0.27795
3.382 0.98806 5.5038e-005 3.8182 0.012003 4.4349e-005 0.0011566 0.22137 0.00065921 0.22202 0.20455 0 0.032884 0.0389 0 1.1082 0.3457 0.10124 0.013291 6.1443 0.082957 0.00010265 0.80715 0.0066665 0.007466 0.0014929 0.98555 0.99079 3.2337e-006 1.2935e-005 0.14328 0.77544 0.82995 0.0014525 0.88252 0.48215 0.0019546 0.42327 1.5217 1.519 16.0087 144.9673 0.00029912 -85.2076 0.27895
3.383 0.98806 5.5038e-005 3.8182 0.012003 4.4362e-005 0.0011566 0.22138 0.00065921 0.22203 0.20456 0 0.032883 0.0389 0 1.1083 0.34575 0.10125 0.013293 6.1456 0.082968 0.00010267 0.80713 0.0066672 0.0074668 0.0014921 0.98556 0.99079 3.2318e-006 1.2927e-005 0.14328 0.77609 0.83036 0.0014521 0.88323 0.48233 0.0019541 0.42328 1.5231 1.5204 16.0088 144.9673 0.00029848 -85.2109 0.27995
3.384 0.98806 5.5037e-005 3.8182 0.012003 4.4375e-005 0.0011566 0.22139 0.00065921 0.22204 0.20457 0 0.032883 0.0389 0 1.1084 0.34579 0.10127 0.013294 6.1469 0.082979 0.00010268 0.80712 0.006668 0.0074676 0.0014913 0.98557 0.9908 3.23e-006 1.292e-005 0.14329 0.77674 0.83077 0.0014517 0.88394 0.48251 0.0019536 0.42329 1.5246 1.5219 16.0088 144.9673 0.00029785 -85.2141 0.28095
3.385 0.98806 5.5037e-005 3.8182 0.012003 4.4388e-005 0.0011566 0.2214 0.00065921 0.22206 0.20458 0 0.032882 0.0389 0 1.1085 0.34584 0.10128 0.013296 6.1482 0.082989 0.0001027 0.80711 0.0066687 0.0074683 0.0014905 0.98558 0.99081 3.2282e-006 1.2913e-005 0.14329 0.77738 0.83118 0.0014513 0.88464 0.48268 0.001953 0.4233 1.526 1.5233 16.0088 144.9673 0.00029723 -85.2173 0.28195
3.386 0.98806 5.5037e-005 3.8182 0.012003 4.4401e-005 0.0011566 0.22141 0.00065921 0.22207 0.20459 0 0.032882 0.0389 0 1.1086 0.34588 0.1013 0.013298 6.1495 0.083 0.00010271 0.8071 0.0066694 0.0074691 0.0014897 0.98559 0.99081 3.2263e-006 1.2905e-005 0.1433 0.77802 0.83159 0.0014509 0.88534 0.48286 0.0019525 0.42331 1.5274 1.5248 16.0088 144.9673 0.0002966 -85.2205 0.28295
3.387 0.98806 5.5037e-005 3.8182 0.012003 4.4414e-005 0.0011566 0.22142 0.00065921 0.22208 0.2046 0 0.032881 0.0389 0 1.1087 0.34593 0.10132 0.0133 6.1509 0.083011 0.00010272 0.80709 0.0066701 0.0074699 0.0014889 0.9856 0.99082 3.2245e-006 1.2898e-005 0.14331 0.77866 0.83199 0.0014505 0.88604 0.48304 0.001952 0.42332 1.5289 1.5262 16.0088 144.9674 0.00029598 -85.2236 0.28395
3.388 0.98806 5.5037e-005 3.8182 0.012003 4.4427e-005 0.0011566 0.22143 0.00065921 0.22209 0.20461 0 0.03288 0.0389 0 1.1088 0.34598 0.10133 0.013301 6.1522 0.083022 0.00010274 0.80708 0.0066709 0.0074706 0.0014882 0.98561 0.99083 3.2228e-006 1.2891e-005 0.14331 0.7793 0.83239 0.0014501 0.88673 0.48322 0.0019515 0.42333 1.5303 1.5277 16.0089 144.9674 0.00029536 -85.2268 0.28495
3.389 0.98806 5.5037e-005 3.8182 0.012003 4.444e-005 0.0011566 0.22144 0.00065921 0.2221 0.20462 0 0.03288 0.0389 0 1.1089 0.34602 0.10135 0.013303 6.1535 0.083033 0.00010275 0.80707 0.0066716 0.0074714 0.0014874 0.98562 0.99083 3.221e-006 1.2884e-005 0.14332 0.77994 0.83279 0.0014497 0.88742 0.48339 0.001951 0.42334 1.5317 1.5291 16.0089 144.9674 0.00029475 -85.2299 0.28595
3.39 0.98806 5.5037e-005 3.8182 0.012003 4.4453e-005 0.0011566 0.22146 0.00065921 0.22211 0.20464 0 0.032879 0.0389 0 1.109 0.34607 0.10136 0.013305 6.1548 0.083043 0.00010277 0.80706 0.0066723 0.0074722 0.0014866 0.98563 0.99084 3.2192e-006 1.2877e-005 0.14332 0.78057 0.83319 0.0014493 0.8881 0.48357 0.0019504 0.42335 1.5332 1.5305 16.0089 144.9674 0.00029413 -85.233 0.28695
3.391 0.98806 5.5037e-005 3.8182 0.012003 4.4466e-005 0.0011566 0.22147 0.00065921 0.22212 0.20465 0 0.032879 0.0389 0 1.1091 0.34611 0.10138 0.013307 6.1561 0.083054 0.00010278 0.80705 0.006673 0.007473 0.0014859 0.98564 0.99085 3.2175e-006 1.287e-005 0.14333 0.7812 0.83358 0.0014489 0.88878 0.48375 0.0019499 0.42336 1.5346 1.532 16.0089 144.9674 0.00029352 -85.236 0.28795
3.392 0.98806 5.5037e-005 3.8182 0.012003 4.4479e-005 0.0011566 0.22148 0.00065921 0.22213 0.20466 0 0.032878 0.0389 0 1.1092 0.34616 0.1014 0.013308 6.1574 0.083065 0.0001028 0.80704 0.0066738 0.0074737 0.0014851 0.98565 0.99086 3.2157e-006 1.2863e-005 0.14334 0.78183 0.83398 0.0014485 0.88946 0.48393 0.0019494 0.42337 1.536 1.5334 16.0089 144.9674 0.00029292 -85.2391 0.28895
3.393 0.98806 5.5037e-005 3.8182 0.012003 4.4492e-005 0.0011566 0.22149 0.00065921 0.22214 0.20467 0 0.032878 0.0389 0 1.1093 0.34621 0.10141 0.01331 6.1587 0.083076 0.00010281 0.80703 0.0066745 0.0074745 0.0014844 0.98566 0.99086 3.214e-006 1.2856e-005 0.14334 0.78246 0.83437 0.0014481 0.89013 0.4841 0.0019489 0.42338 1.5374 1.5348 16.009 144.9675 0.00029231 -85.2421 0.28995
3.394 0.98806 5.5037e-005 3.8182 0.012003 4.4505e-005 0.0011566 0.2215 0.00065921 0.22215 0.20468 0 0.032877 0.0389 0 1.1094 0.34625 0.10143 0.013312 6.16 0.083087 0.00010283 0.80702 0.0066752 0.0074753 0.0014836 0.98567 0.99087 3.2123e-006 1.2849e-005 0.14335 0.78309 0.83476 0.0014477 0.89079 0.48428 0.0019484 0.42339 1.5388 1.5362 16.009 144.9675 0.00029171 -85.2451 0.29095
3.395 0.98806 5.5037e-005 3.8182 0.012003 4.4518e-005 0.0011566 0.22151 0.00065921 0.22217 0.20469 0 0.032877 0.0389 0 1.1095 0.3463 0.10144 0.013313 6.1614 0.083097 0.00010284 0.80701 0.0066759 0.007476 0.0014829 0.98568 0.99087 3.2106e-006 1.2843e-005 0.14335 0.78371 0.83515 0.0014473 0.89146 0.48446 0.0019479 0.4234 1.5402 1.5377 16.009 144.9675 0.00029111 -85.2481 0.29195
3.396 0.98806 5.5037e-005 3.8182 0.012003 4.4531e-005 0.0011566 0.22152 0.00065921 0.22218 0.2047 0 0.032876 0.0389 0 1.1096 0.34634 0.10146 0.013315 6.1627 0.083108 0.00010286 0.80699 0.0066766 0.0074768 0.0014822 0.98569 0.99088 3.2089e-006 1.2836e-005 0.14336 0.78433 0.83554 0.0014469 0.89212 0.48463 0.0019474 0.42341 1.5416 1.5391 16.009 144.9675 0.00029052 -85.251 0.29295
3.397 0.98806 5.5037e-005 3.8182 0.012003 4.4544e-005 0.0011566 0.22153 0.00065921 0.22219 0.20471 0 0.032875 0.0389 0 1.1097 0.34639 0.10148 0.013317 6.164 0.083119 0.00010287 0.80698 0.0066774 0.0074776 0.0014814 0.9857 0.99089 3.2073e-006 1.2829e-005 0.14336 0.78495 0.83592 0.0014466 0.89277 0.48481 0.001947 0.42342 1.543 1.5405 16.009 144.9675 0.00028992 -85.2539 0.29395
3.398 0.98806 5.5037e-005 3.8182 0.012003 4.4557e-005 0.0011566 0.22154 0.00065921 0.2222 0.20472 0 0.032875 0.0389 0 1.1098 0.34644 0.10149 0.013319 6.1653 0.08313 0.00010289 0.80697 0.0066781 0.0074784 0.0014807 0.98571 0.99089 3.2056e-006 1.2823e-005 0.14337 0.78557 0.8363 0.0014462 0.89343 0.48499 0.0019465 0.42343 1.5444 1.5419 16.009 144.9675 0.00028933 -85.2569 0.29495
3.399 0.98806 5.5036e-005 3.8182 0.012003 4.457e-005 0.0011566 0.22155 0.00065921 0.22221 0.20473 0 0.032874 0.0389 0 1.1099 0.34648 0.10151 0.01332 6.1666 0.08314 0.0001029 0.80696 0.0066788 0.0074791 0.00148 0.98572 0.9909 3.204e-006 1.2816e-005 0.14338 0.78619 0.83668 0.0014458 0.89407 0.48517 0.001946 0.42345 1.5458 1.5433 16.0091 144.9676 0.00028874 -85.2597 0.29595
3.4 0.98806 5.5036e-005 3.8182 0.012003 4.4583e-005 0.0011566 0.22156 0.00065921 0.22222 0.20474 0 0.032874 0.0389 0 1.11 0.34653 0.10153 0.013322 6.1679 0.083151 0.00010292 0.80695 0.0066795 0.0074799 0.0014793 0.98573 0.99091 3.2024e-006 1.281e-005 0.14338 0.7868 0.83706 0.0014455 0.89472 0.48534 0.0019455 0.42346 1.5472 1.5447 16.0091 144.9676 0.00028816 -85.2626 0.29695
3.401 0.98806 5.5036e-005 3.8182 0.012003 4.4596e-005 0.0011566 0.22158 0.00065921 0.22223 0.20475 0 0.032873 0.0389 0 1.1101 0.34657 0.10154 0.013324 6.1693 0.083162 0.00010293 0.80694 0.0066803 0.0074807 0.0014786 0.98574 0.99091 3.2008e-006 1.2803e-005 0.14339 0.78741 0.83744 0.0014451 0.89536 0.48552 0.0019451 0.42347 1.5486 1.5461 16.0091 144.9676 0.00028758 -85.2655 0.29795
3.402 0.98806 5.5036e-005 3.8182 0.012003 4.461e-005 0.0011566 0.22159 0.00065921 0.22224 0.20476 0 0.032873 0.0389 0 1.1102 0.34662 0.10156 0.013326 6.1706 0.083173 0.00010295 0.80693 0.006681 0.0074814 0.0014779 0.98575 0.99092 3.1991e-006 1.2797e-005 0.14339 0.78803 0.83781 0.0014448 0.89599 0.4857 0.0019446 0.42348 1.55 1.5474 16.0091 144.9676 0.000287 -85.2683 0.29895
3.403 0.98806 5.5036e-005 3.8182 0.012003 4.4623e-005 0.0011566 0.2216 0.00065921 0.22225 0.20477 0 0.032872 0.0389 0 1.1103 0.34667 0.10157 0.013327 6.1719 0.083184 0.00010296 0.80692 0.0066817 0.0074822 0.0014772 0.98576 0.99093 3.1976e-006 1.279e-005 0.1434 0.78863 0.83819 0.0014444 0.89663 0.48587 0.0019441 0.42349 1.5513 1.5488 16.0091 144.9676 0.00028642 -85.2711 0.29995
3.404 0.98806 5.5036e-005 3.8182 0.012003 4.4636e-005 0.0011566 0.22161 0.00065921 0.22226 0.20478 0 0.032871 0.0389 0 1.1104 0.34671 0.10159 0.013329 6.1732 0.083194 0.00010298 0.80691 0.0066824 0.007483 0.0014765 0.98577 0.99093 3.196e-006 1.2784e-005 0.14341 0.78924 0.83856 0.0014441 0.89726 0.48605 0.0019437 0.4235 1.5527 1.5502 16.0091 144.9676 0.00028584 -85.2739 0.30095
3.405 0.98806 5.5036e-005 3.8182 0.012003 4.4649e-005 0.0011566 0.22162 0.00065921 0.22227 0.20479 0 0.032871 0.0389 0 1.1105 0.34676 0.10161 0.013331 6.1745 0.083205 0.00010299 0.8069 0.0066831 0.0074837 0.0014758 0.98577 0.99094 3.1944e-006 1.2778e-005 0.14341 0.78985 0.83893 0.0014437 0.89788 0.48623 0.0019432 0.42351 1.5541 1.5516 16.0092 144.9677 0.00028527 -85.2767 0.30195
3.406 0.98806 5.5036e-005 3.8182 0.012003 4.4662e-005 0.0011566 0.22163 0.00065921 0.22228 0.2048 0 0.03287 0.0389 0 1.1106 0.3468 0.10162 0.013332 6.1758 0.083216 0.000103 0.80689 0.0066839 0.0074845 0.0014751 0.98578 0.99094 3.1929e-006 1.2772e-005 0.14342 0.79045 0.8393 0.0014434 0.8985 0.4864 0.0019428 0.42352 1.5554 1.553 16.0092 144.9677 0.0002847 -85.2794 0.30295
3.407 0.98806 5.5036e-005 3.8182 0.012003 4.4675e-005 0.0011566 0.22164 0.00065921 0.2223 0.20481 0 0.03287 0.0389 0 1.1107 0.34685 0.10164 0.013334 6.1772 0.083227 0.00010302 0.80688 0.0066846 0.0074853 0.0014745 0.98579 0.99095 3.1913e-006 1.2765e-005 0.14342 0.79105 0.83966 0.0014431 0.89912 0.48658 0.0019423 0.42353 1.5568 1.5543 16.0092 144.9677 0.00028414 -85.2821 0.30395
3.408 0.98806 5.5036e-005 3.8182 0.012003 4.4688e-005 0.0011566 0.22165 0.00065921 0.22231 0.20482 0 0.032869 0.0389 0 1.1108 0.3469 0.10165 0.013336 6.1785 0.083238 0.00010303 0.80687 0.0066853 0.0074861 0.0014738 0.9858 0.99096 3.1898e-006 1.2759e-005 0.14343 0.79165 0.84003 0.0014427 0.89973 0.48676 0.0019419 0.42354 1.5582 1.5557 16.0092 144.9677 0.00028357 -85.2848 0.30495
3.409 0.98806 5.5036e-005 3.8182 0.012003 4.4701e-005 0.0011566 0.22166 0.00065921 0.22232 0.20483 0 0.032869 0.0389 0 1.1109 0.34694 0.10167 0.013338 6.1798 0.083248 0.00010305 0.80685 0.006686 0.0074868 0.0014732 0.98581 0.99096 3.1883e-006 1.2753e-005 0.14343 0.79225 0.84039 0.0014424 0.90034 0.48693 0.0019414 0.42355 1.5595 1.5571 16.0092 144.9677 0.00028301 -85.2875 0.30595
3.41 0.98806 5.5036e-005 3.8182 0.012003 4.4714e-005 0.0011566 0.22167 0.00065921 0.22233 0.20484 0 0.032868 0.0389 0 1.111 0.34699 0.10169 0.013339 6.1811 0.083259 0.00010306 0.80684 0.0066868 0.0074876 0.0014725 0.98582 0.99097 3.1868e-006 1.2747e-005 0.14344 0.79284 0.84075 0.001442 0.90095 0.48711 0.001941 0.42356 1.5609 1.5584 16.0092 144.9678 0.00028245 -85.2902 0.30695
3.411 0.98806 5.5036e-005 3.8182 0.012003 4.4727e-005 0.0011566 0.22168 0.00065921 0.22234 0.20485 0 0.032868 0.0389 0 1.1111 0.34704 0.1017 0.013341 6.1825 0.08327 0.00010308 0.80683 0.0066875 0.0074884 0.0014719 0.98583 0.99097 3.1853e-006 1.2741e-005 0.14345 0.79344 0.84111 0.0014417 0.90155 0.48729 0.0019405 0.42358 1.5622 1.5598 16.0092 144.9678 0.00028189 -85.2928 0.30795
3.412 0.98806 5.5036e-005 3.8182 0.012003 4.474e-005 0.0011566 0.22169 0.00065921 0.22235 0.20486 0 0.032867 0.0389 0 1.1112 0.34708 0.10172 0.013343 6.1838 0.083281 0.00010309 0.80682 0.0066882 0.0074891 0.0014712 0.98584 0.99098 3.1838e-006 1.2735e-005 0.14345 0.79403 0.84147 0.0014413 0.90215 0.48746 0.0019401 0.42359 1.5635 1.5611 16.0093 144.9678 0.00028134 -85.2955 0.30895
3.413 0.98806 5.5035e-005 3.8182 0.012003 4.4753e-005 0.0011566 0.22171 0.00065921 0.22236 0.20487 0 0.032866 0.0389 0 1.1113 0.34713 0.10174 0.013345 6.1851 0.083292 0.00010311 0.80681 0.0066889 0.0074899 0.0014706 0.98584 0.99098 3.1823e-006 1.2729e-005 0.14346 0.79462 0.84183 0.001441 0.90275 0.48764 0.0019397 0.4236 1.5649 1.5625 16.0093 144.9678 0.00028079 -85.2981 0.30995
3.414 0.98806 5.5035e-005 3.8182 0.012003 4.4766e-005 0.0011566 0.22172 0.00065921 0.22237 0.20488 0 0.032866 0.0389 0 1.1114 0.34717 0.10175 0.013346 6.1864 0.083302 0.00010312 0.8068 0.0066896 0.0074907 0.0014699 0.98585 0.99099 3.1809e-006 1.2724e-005 0.14346 0.79521 0.84218 0.0014407 0.90334 0.48782 0.0019392 0.42361 1.5662 1.5638 16.0093 144.9678 0.00028024 -85.3007 0.31095
3.415 0.98806 5.5035e-005 3.8182 0.012003 4.4779e-005 0.0011566 0.22173 0.00065921 0.22238 0.20489 0 0.032865 0.0389 0 1.1115 0.34722 0.10177 0.013348 6.1877 0.083313 0.00010314 0.80679 0.0066904 0.0074915 0.0014693 0.98586 0.99099 3.1794e-006 1.2718e-005 0.14347 0.7958 0.84254 0.0014403 0.90393 0.48799 0.0019388 0.42362 1.5676 1.5652 16.0093 144.9678 0.00027969 -85.3032 0.31195
3.416 0.98806 5.5035e-005 3.8182 0.012003 4.4792e-005 0.0011567 0.22174 0.00065921 0.22239 0.2049 0 0.032865 0.0389 0 1.1116 0.34727 0.10178 0.01335 6.1891 0.083324 0.00010315 0.80678 0.0066911 0.0074922 0.0014687 0.98587 0.991 3.178e-006 1.2712e-005 0.14348 0.79638 0.84289 0.00144 0.90451 0.48817 0.0019384 0.42363 1.5689 1.5665 16.0093 144.9679 0.00027915 -85.3058 0.31295
3.417 0.98806 5.5035e-005 3.8182 0.012003 4.4805e-005 0.0011567 0.22175 0.00065921 0.2224 0.20491 0 0.032864 0.0389 0 1.1117 0.34731 0.1018 0.013351 6.1904 0.083335 0.00010317 0.80677 0.0066918 0.007493 0.0014681 0.98588 0.99101 3.1766e-006 1.2706e-005 0.14348 0.79696 0.84324 0.0014397 0.9051 0.48835 0.001938 0.42364 1.5702 1.5678 16.0093 144.9679 0.00027861 -85.3083 0.31395
3.418 0.98806 5.5035e-005 3.8182 0.012003 4.4818e-005 0.0011567 0.22176 0.00065921 0.22241 0.20492 0 0.032864 0.0389 0 1.1118 0.34736 0.10182 0.013353 6.1917 0.083345 0.00010318 0.80676 0.0066925 0.0074938 0.0014674 0.98589 0.99101 3.1752e-006 1.2701e-005 0.14349 0.79754 0.84358 0.0014394 0.90567 0.48852 0.0019376 0.42365 1.5715 1.5692 16.0093 144.9679 0.00027807 -85.3108 0.31495
3.419 0.98806 5.5035e-005 3.8182 0.012003 4.4831e-005 0.0011567 0.22177 0.00065921 0.22242 0.20493 0 0.032863 0.0389 0 1.1119 0.3474 0.10183 0.013355 6.193 0.083356 0.0001032 0.80675 0.0066932 0.0074945 0.0014668 0.98589 0.99102 3.1737e-006 1.2695e-005 0.14349 0.79812 0.84393 0.0014391 0.90625 0.4887 0.0019372 0.42366 1.5728 1.5705 16.0093 144.9679 0.00027753 -85.3133 0.31595
3.42 0.98806 5.5035e-005 3.8182 0.012002 4.4844e-005 0.0011567 0.22178 0.00065921 0.22243 0.20494 0 0.032863 0.0389 0 1.112 0.34745 0.10185 0.013357 6.1944 0.083367 0.00010321 0.80674 0.006694 0.0074953 0.0014662 0.9859 0.99102 3.1724e-006 1.2689e-005 0.1435 0.7987 0.84428 0.0014388 0.90682 0.48887 0.0019368 0.42367 1.5742 1.5718 16.0094 144.9679 0.00027699 -85.3158 0.31695
3.421 0.98806 5.5035e-005 3.8182 0.012002 4.4857e-005 0.0011567 0.22179 0.00065921 0.22245 0.20495 0 0.032862 0.0389 0 1.1121 0.3475 0.10186 0.013358 6.1957 0.083378 0.00010323 0.80673 0.0066947 0.0074961 0.0014656 0.98591 0.99103 3.171e-006 1.2684e-005 0.1435 0.79928 0.84462 0.0014384 0.90739 0.48905 0.0019363 0.42369 1.5755 1.5731 16.0094 144.9679 0.00027646 -85.3183 0.31795
3.422 0.98806 5.5035e-005 3.8182 0.012002 4.487e-005 0.0011567 0.2218 0.00065921 0.22246 0.20496 0 0.032862 0.0389 0 1.1122 0.34754 0.10188 0.01336 6.197 0.083389 0.00010324 0.80671 0.0066954 0.0074968 0.001465 0.98592 0.99103 3.1696e-006 1.2678e-005 0.14351 0.79985 0.84496 0.0014382 0.90795 0.48923 0.0019359 0.4237 1.5768 1.5744 16.0094 144.968 0.00027593 -85.3207 0.31895
3.423 0.98806 5.5035e-005 3.8182 0.012002 4.4883e-005 0.0011567 0.22181 0.00065921 0.22247 0.20497 0 0.032861 0.0389 0 1.1123 0.34759 0.1019 0.013362 6.1983 0.083399 0.00010325 0.8067 0.0066961 0.0074976 0.0014644 0.98593 0.99104 3.1682e-006 1.2673e-005 0.14352 0.80042 0.8453 0.0014379 0.90851 0.4894 0.0019355 0.42371 1.5781 1.5757 16.0094 144.968 0.00027541 -85.3231 0.31995
3.424 0.98806 5.5035e-005 3.8182 0.012002 4.4896e-005 0.0011567 0.22182 0.00065921 0.22248 0.20498 0 0.03286 0.0389 0 1.1124 0.34763 0.10191 0.013364 6.1997 0.08341 0.00010327 0.80669 0.0066969 0.0074984 0.0014638 0.98593 0.99104 3.1669e-006 1.2668e-005 0.14352 0.80099 0.84564 0.0014376 0.90907 0.48958 0.0019351 0.42372 1.5794 1.5771 16.0094 144.968 0.00027488 -85.3256 0.32095
3.425 0.98806 5.5035e-005 3.8182 0.012002 4.4909e-005 0.0011567 0.22183 0.00065921 0.22249 0.20499 0 0.03286 0.0389 0 1.1125 0.34768 0.10193 0.013365 6.201 0.083421 0.00010328 0.80668 0.0066976 0.0074992 0.0014632 0.98594 0.99105 3.1655e-006 1.2662e-005 0.14353 0.80156 0.84598 0.0014373 0.90962 0.48975 0.0019348 0.42373 1.5807 1.5784 16.0094 144.968 0.00027436 -85.3279 0.32195
3.426 0.98806 5.5035e-005 3.8182 0.012002 4.4922e-005 0.0011567 0.22184 0.00065921 0.2225 0.205 0 0.032859 0.0389 0 1.1126 0.34773 0.10194 0.013367 6.2023 0.083432 0.0001033 0.80667 0.0066983 0.0074999 0.0014627 0.98595 0.99105 3.1642e-006 1.2657e-005 0.14353 0.80213 0.84631 0.001437 0.91018 0.48993 0.0019344 0.42374 1.582 1.5797 16.0094 144.968 0.00027384 -85.3303 0.32295
3.427 0.98806 5.5035e-005 3.8182 0.012002 4.4935e-005 0.0011567 0.22185 0.00065921 0.22251 0.20501 0 0.032859 0.0389 0 1.1127 0.34777 0.10196 0.013369 6.2036 0.083442 0.00010331 0.80666 0.006699 0.0075007 0.0014621 0.98596 0.99106 3.1629e-006 1.2652e-005 0.14354 0.8027 0.84665 0.0014367 0.91072 0.4901 0.001934 0.42375 1.5833 1.581 16.0094 144.9681 0.00027332 -85.3327 0.32395
3.428 0.98806 5.5034e-005 3.8182 0.012002 4.4948e-005 0.0011567 0.22187 0.00065921 0.22252 0.20502 0 0.032858 0.0389 0 1.1128 0.34782 0.10198 0.013371 6.205 0.083453 0.00010333 0.80665 0.0066997 0.0075015 0.0014615 0.98596 0.99106 3.1616e-006 1.2646e-005 0.14355 0.80326 0.84698 0.0014364 0.91127 0.49028 0.0019336 0.42377 1.5845 1.5822 16.0095 144.9681 0.0002728 -85.335 0.32495
3.429 0.98806 5.5034e-005 3.8182 0.012002 4.4962e-005 0.0011567 0.22188 0.00065921 0.22253 0.20503 0 0.032858 0.0389 0 1.1129 0.34787 0.10199 0.013372 6.2063 0.083464 0.00010334 0.80664 0.0067005 0.0075022 0.001461 0.98597 0.99107 3.1603e-006 1.2641e-005 0.14355 0.80382 0.84731 0.0014361 0.91181 0.49046 0.0019332 0.42378 1.5858 1.5835 16.0095 144.9681 0.00027229 -85.3373 0.32595
3.43 0.98806 5.5034e-005 3.8182 0.012002 4.4975e-005 0.0011567 0.22189 0.00065921 0.22254 0.20504 0 0.032857 0.0389 0 1.113 0.34791 0.10201 0.013374 6.2076 0.083475 0.00010336 0.80663 0.0067012 0.007503 0.0014604 0.98598 0.99107 3.159e-006 1.2636e-005 0.14356 0.80438 0.84764 0.0014358 0.91235 0.49063 0.0019328 0.42379 1.5871 1.5848 16.0095 144.9681 0.00027178 -85.3397 0.32695
3.431 0.98806 5.5034e-005 3.8182 0.012002 4.4988e-005 0.0011567 0.2219 0.00065921 0.22255 0.20505 0 0.032857 0.0389 0 1.1131 0.34796 0.10203 0.013376 6.2089 0.083485 0.00010337 0.80662 0.0067019 0.0075038 0.0014599 0.98599 0.99108 3.1577e-006 1.2631e-005 0.14356 0.80494 0.84797 0.0014355 0.91288 0.49081 0.0019325 0.4238 1.5884 1.5861 16.0095 144.9681 0.00027127 -85.3419 0.32795
3.432 0.98806 5.5034e-005 3.8182 0.012002 4.5001e-005 0.0011567 0.22191 0.00065921 0.22256 0.20506 0 0.032856 0.0389 0 1.1132 0.348 0.10204 0.013377 6.2103 0.083496 0.00010339 0.80661 0.0067026 0.0075045 0.0014593 0.98599 0.99108 3.1564e-006 1.2626e-005 0.14357 0.8055 0.84829 0.0014352 0.91341 0.49098 0.0019321 0.42381 1.5896 1.5874 16.0095 144.9681 0.00027076 -85.3442 0.32895
3.433 0.98806 5.5034e-005 3.8182 0.012002 4.5014e-005 0.0011567 0.22192 0.00065921 0.22257 0.20507 0 0.032855 0.0389 0 1.1133 0.34805 0.10206 0.013379 6.2116 0.083507 0.0001034 0.8066 0.0067034 0.0075053 0.0014588 0.986 0.99109 3.1552e-006 1.2621e-005 0.14357 0.80605 0.84862 0.0014349 0.91394 0.49116 0.0019317 0.42382 1.5909 1.5887 16.0095 144.9682 0.00027026 -85.3465 0.32995
3.434 0.98806 5.5034e-005 3.8182 0.012002 4.5027e-005 0.0011567 0.22193 0.00065921 0.22258 0.20508 0 0.032855 0.0389 0 1.1134 0.3481 0.10207 0.013381 6.2129 0.083518 0.00010342 0.80659 0.0067041 0.0075061 0.0014582 0.98601 0.99109 3.1539e-006 1.2616e-005 0.14358 0.8066 0.84894 0.0014346 0.91446 0.49133 0.0019313 0.42383 1.5922 1.5899 16.0095 144.9682 0.00026976 -85.3487 0.33095
3.435 0.98806 5.5034e-005 3.8182 0.012002 4.504e-005 0.0011567 0.22194 0.00065921 0.22259 0.20509 0 0.032854 0.0389 0 1.1135 0.34814 0.10209 0.013383 6.2143 0.083529 0.00010343 0.80657 0.0067048 0.0075069 0.0014577 0.98601 0.9911 3.1527e-006 1.2611e-005 0.14359 0.80715 0.84926 0.0014343 0.91499 0.49151 0.001931 0.42385 1.5934 1.5912 16.0095 144.9682 0.00026926 -85.3509 0.33195
3.436 0.98806 5.5034e-005 3.8182 0.012002 4.5053e-005 0.0011567 0.22195 0.00065921 0.2226 0.2051 0 0.032854 0.0389 0 1.1136 0.34819 0.10211 0.013384 6.2156 0.083539 0.00010345 0.80656 0.0067055 0.0075076 0.0014571 0.98602 0.9911 3.1515e-006 1.2606e-005 0.14359 0.8077 0.84958 0.001434 0.9155 0.49168 0.0019306 0.42386 1.5947 1.5925 16.0095 144.9682 0.00026876 -85.3531 0.33295
3.437 0.98806 5.5034e-005 3.8182 0.012002 4.5066e-005 0.0011567 0.22196 0.00065921 0.22262 0.20511 0 0.032853 0.0389 0 1.1137 0.34823 0.10212 0.013386 6.2169 0.08355 0.00010346 0.80655 0.0067062 0.0075084 0.0014566 0.98603 0.99111 3.1502e-006 1.2601e-005 0.1436 0.80825 0.8499 0.0014338 0.91602 0.49186 0.0019303 0.42387 1.596 1.5937 16.0095 144.9682 0.00026826 -85.3553 0.33395
3.438 0.98806 5.5034e-005 3.8182 0.012002 4.5079e-005 0.0011567 0.22197 0.00065921 0.22263 0.20512 0 0.032853 0.0389 0 1.1138 0.34828 0.10214 0.013388 6.2183 0.083561 0.00010348 0.80654 0.006707 0.0075092 0.0014561 0.98604 0.99111 3.149e-006 1.2596e-005 0.1436 0.8088 0.85022 0.0014335 0.91653 0.49204 0.0019299 0.42388 1.5972 1.595 16.0096 144.9683 0.00026777 -85.3575 0.33495
3.439 0.98806 5.5034e-005 3.8182 0.012002 4.5092e-005 0.0011567 0.22198 0.00065921 0.22264 0.20513 0 0.032852 0.0389 0 1.1139 0.34833 0.10215 0.01339 6.2196 0.083572 0.00010349 0.80653 0.0067077 0.0075099 0.0014555 0.98604 0.99112 3.1478e-006 1.2591e-005 0.14361 0.80934 0.85053 0.0014332 0.91704 0.49221 0.0019295 0.42389 1.5985 1.5962 16.0096 144.9683 0.00026728 -85.3597 0.33595
3.44 0.98806 5.5034e-005 3.8182 0.012002 4.5105e-005 0.0011567 0.22199 0.00065921 0.22265 0.20514 0 0.032852 0.0389 0 1.114 0.34837 0.10217 0.013391 6.2209 0.083582 0.0001035 0.80652 0.0067084 0.0075107 0.001455 0.98605 0.99112 3.1466e-006 1.2587e-005 0.14362 0.80989 0.85085 0.0014329 0.91755 0.49239 0.0019292 0.4239 1.5997 1.5975 16.0096 144.9683 0.00026679 -85.3618 0.33695
3.441 0.98806 5.5034e-005 3.8182 0.012002 4.5118e-005 0.0011567 0.222 0.00065921 0.22266 0.20515 0 0.032851 0.0389 0 1.1141 0.34842 0.10219 0.013393 6.2223 0.083593 0.00010352 0.80651 0.0067091 0.0075115 0.0014545 0.98606 0.99112 3.1454e-006 1.2582e-005 0.14362 0.81043 0.85116 0.0014327 0.91805 0.49256 0.0019288 0.42391 1.6009 1.5987 16.0096 144.9683 0.0002663 -85.364 0.33795
3.442 0.98806 5.5033e-005 3.8182 0.012002 4.5131e-005 0.0011567 0.22201 0.00065921 0.22267 0.20516 0 0.032851 0.0389 0 1.1142 0.34846 0.1022 0.013395 6.2236 0.083604 0.00010353 0.8065 0.0067098 0.0075123 0.001454 0.98606 0.99113 3.1443e-006 1.2577e-005 0.14363 0.81097 0.85147 0.0014324 0.91855 0.49274 0.0019285 0.42393 1.6022 1.6 16.0096 144.9683 0.00026582 -85.3661 0.33895
3.443 0.98806 5.5033e-005 3.8182 0.012002 4.5144e-005 0.0011567 0.22202 0.00065921 0.22268 0.20517 0 0.03285 0.0389 0 1.1143 0.34851 0.10222 0.013396 6.2249 0.083615 0.00010355 0.80649 0.0067106 0.007513 0.0014535 0.98607 0.99113 3.1431e-006 1.2572e-005 0.14363 0.8115 0.85178 0.0014322 0.91905 0.49291 0.0019281 0.42394 1.6034 1.6012 16.0096 144.9683 0.00026534 -85.3682 0.33995
3.444 0.98806 5.5033e-005 3.8182 0.012002 4.5157e-005 0.0011567 0.22203 0.00065921 0.22269 0.20518 0 0.03285 0.0389 0 1.1144 0.34856 0.10224 0.013398 6.2263 0.083625 0.00010356 0.80648 0.0067113 0.0075138 0.001453 0.98608 0.99114 3.1419e-006 1.2568e-005 0.14364 0.81204 0.85209 0.0014319 0.91954 0.49309 0.0019278 0.42395 1.6046 1.6025 16.0096 144.9684 0.00026486 -85.3703 0.34095
3.445 0.98806 5.5033e-005 3.8182 0.012002 4.517e-005 0.0011567 0.22204 0.00065921 0.2227 0.20519 0 0.032849 0.0389 0 1.1145 0.3486 0.10225 0.0134 6.2276 0.083636 0.00010358 0.80647 0.006712 0.0075146 0.0014525 0.98608 0.99114 3.1408e-006 1.2563e-005 0.14364 0.81257 0.8524 0.0014317 0.92003 0.49326 0.0019275 0.42396 1.6059 1.6037 16.0096 144.9684 0.00026438 -85.3723 0.34195
3.446 0.98806 5.5033e-005 3.8182 0.012002 4.5183e-005 0.0011567 0.22206 0.00065921 0.22271 0.2052 0 0.032848 0.0389 0 1.1146 0.34865 0.10227 0.013402 6.2289 0.083647 0.00010359 0.80646 0.0067127 0.0075153 0.001452 0.98609 0.99115 3.1396e-006 1.2559e-005 0.14365 0.81311 0.85271 0.0014315 0.92052 0.49344 0.0019271 0.42397 1.6071 1.6049 16.0096 144.9684 0.0002639 -85.3744 0.34295
3.447 0.98806 5.5033e-005 3.8182 0.012002 4.5196e-005 0.0011567 0.22207 0.00065921 0.22272 0.20521 0 0.032848 0.0389 0 1.1147 0.3487 0.10228 0.013403 6.2303 0.083658 0.00010361 0.80645 0.0067135 0.0075161 0.0014515 0.9861 0.99115 3.1385e-006 1.2554e-005 0.14366 0.81364 0.85301 0.0014312 0.921 0.49361 0.0019268 0.42398 1.6083 1.6062 16.0096 144.9684 0.00026343 -85.3764 0.34395
3.448 0.98806 5.5033e-005 3.8182 0.012002 4.5209e-005 0.0011567 0.22208 0.00065921 0.22273 0.20522 0 0.032847 0.0389 0 1.1148 0.34874 0.1023 0.013405 6.2316 0.083668 0.00010362 0.80644 0.0067142 0.0075169 0.001451 0.9861 0.99115 3.1374e-006 1.255e-005 0.14366 0.81417 0.85332 0.001431 0.92148 0.49379 0.0019265 0.424 1.6095 1.6074 16.0096 144.9684 0.00026296 -85.3785 0.34495
3.449 0.98806 5.5033e-005 3.8182 0.012002 4.5222e-005 0.0011567 0.22209 0.00065921 0.22274 0.20523 0 0.032847 0.0389 0 1.1149 0.34879 0.10232 0.013407 6.2329 0.083679 0.00010364 0.80642 0.0067149 0.0075176 0.0014505 0.98611 0.99116 3.1363e-006 1.2545e-005 0.14367 0.8147 0.85362 0.0014307 0.92196 0.49396 0.0019261 0.42401 1.6108 1.6086 16.0096 144.9685 0.00026249 -85.3805 0.34595
3.45 0.98806 5.5033e-005 3.8182 0.012002 4.5235e-005 0.0011567 0.2221 0.00065921 0.22275 0.20524 0 0.032846 0.0389 0 1.115 0.34883 0.10233 0.013409 6.2343 0.08369 0.00010365 0.80641 0.0067156 0.0075184 0.00145 0.98612 0.99116 3.1352e-006 1.2541e-005 0.14367 0.81522 0.85392 0.0014305 0.92244 0.49413 0.0019258 0.42402 1.612 1.6098 16.0096 144.9685 0.00026202 -85.3825 0.34695
3.451 0.98806 5.5033e-005 3.8182 0.012002 4.5248e-005 0.0011567 0.22211 0.00065921 0.22276 0.20525 0 0.032846 0.0389 0 1.1151 0.34888 0.10235 0.01341 6.2356 0.083701 0.00010367 0.8064 0.0067163 0.0075192 0.0014495 0.98612 0.99117 3.1341e-006 1.2536e-005 0.14368 0.81575 0.85422 0.0014302 0.92291 0.49431 0.0019255 0.42403 1.6132 1.6111 16.0097 144.9685 0.00026155 -85.3844 0.34795
3.452 0.98806 5.5033e-005 3.8182 0.012002 4.5261e-005 0.0011567 0.22212 0.00065921 0.22277 0.20526 0 0.032845 0.0389 0 1.1152 0.34893 0.10236 0.013412 6.2369 0.083711 0.00010368 0.80639 0.0067171 0.00752 0.0014491 0.98613 0.99117 3.133e-006 1.2532e-005 0.14369 0.81627 0.85452 0.00143 0.92338 0.49448 0.0019252 0.42404 1.6144 1.6123 16.0097 144.9685 0.00026109 -85.3864 0.34895
3.453 0.98806 5.5033e-005 3.8182 0.012002 4.5274e-005 0.0011567 0.22213 0.00065921 0.22278 0.20527 0 0.032845 0.0389 0 1.1153 0.34897 0.10238 0.013414 6.2383 0.083722 0.0001037 0.80638 0.0067178 0.0075207 0.0014486 0.98613 0.99118 3.1319e-006 1.2528e-005 0.14369 0.81679 0.85481 0.0014297 0.92385 0.49466 0.0019248 0.42406 1.6156 1.6135 16.0097 144.9685 0.00026063 -85.3884 0.34995
3.454 0.98806 5.5033e-005 3.8182 0.012002 4.5287e-005 0.0011567 0.22214 0.00065921 0.22279 0.20528 0 0.032844 0.0389 0 1.1153 0.34902 0.1024 0.013415 6.2396 0.083733 0.00010371 0.80637 0.0067185 0.0075215 0.0014481 0.98614 0.99118 3.1308e-006 1.2523e-005 0.1437 0.81731 0.85511 0.0014294 0.92431 0.49483 0.0019245 0.42407 1.6168 1.6147 16.0097 144.9685 0.00026017 -85.3903 0.35095
3.455 0.98806 5.5033e-005 3.8182 0.012002 4.53e-005 0.0011567 0.22215 0.00065921 0.2228 0.20529 0 0.032844 0.0389 0 1.1154 0.34906 0.10241 0.013417 6.2409 0.083744 0.00010373 0.80636 0.0067192 0.0075223 0.0014477 0.98615 0.99118 3.1297e-006 1.2519e-005 0.1437 0.81783 0.8554 0.0014292 0.92477 0.49501 0.0019242 0.42408 1.618 1.6159 16.0097 144.9686 0.00025971 -85.3922 0.35195
3.456 0.98806 5.5032e-005 3.8182 0.012002 4.5313e-005 0.0011567 0.22216 0.00065921 0.22281 0.2053 0 0.032843 0.0389 0 1.1155 0.34911 0.10243 0.013419 6.2423 0.083754 0.00010374 0.80635 0.0067199 0.007523 0.0014472 0.98615 0.99119 3.1287e-006 1.2515e-005 0.14371 0.81835 0.8557 0.0014289 0.92523 0.49518 0.0019239 0.42409 1.6192 1.6171 16.0097 144.9686 0.00025925 -85.3941 0.35295
3.457 0.98806 5.5032e-005 3.8182 0.012002 4.5327e-005 0.0011567 0.22217 0.00065921 0.22282 0.20531 0 0.032843 0.0389 0 1.1156 0.34916 0.10244 0.013421 6.2436 0.083765 0.00010375 0.80634 0.0067207 0.0075238 0.0014467 0.98616 0.99119 3.1276e-006 1.2511e-005 0.14371 0.81886 0.85599 0.0014287 0.92569 0.49536 0.0019236 0.4241 1.6203 1.6183 16.0097 144.9686 0.0002588 -85.396 0.35395
3.458 0.98806 5.5032e-005 3.8182 0.012002 4.534e-005 0.0011567 0.22218 0.00065921 0.22283 0.20532 0 0.032842 0.0389 0 1.1157 0.3492 0.10246 0.013422 6.245 0.083776 0.00010377 0.80633 0.0067214 0.0075246 0.0014463 0.98616 0.9912 3.1266e-006 1.2506e-005 0.14372 0.81937 0.85628 0.0014284 0.92614 0.49553 0.0019233 0.42412 1.6215 1.6195 16.0097 144.9686 0.00025835 -85.3979 0.35495
3.459 0.98806 5.5032e-005 3.8182 0.012002 4.5353e-005 0.0011567 0.22219 0.00065921 0.22284 0.20533 0 0.032841 0.0389 0 1.1158 0.34925 0.10248 0.013424 6.2463 0.083787 0.00010378 0.80632 0.0067221 0.0075253 0.0014458 0.98617 0.9912 3.1255e-006 1.2502e-005 0.14373 0.81989 0.85657 0.0014282 0.92659 0.4957 0.001923 0.42413 1.6227 1.6207 16.0097 144.9686 0.0002579 -85.3998 0.35595
3.46 0.98806 5.5032e-005 3.8182 0.012002 4.5366e-005 0.0011567 0.2222 0.00065921 0.22286 0.20534 0 0.032841 0.0389 0 1.1159 0.3493 0.10249 0.013426 6.2476 0.083797 0.0001038 0.80631 0.0067228 0.0075261 0.0014454 0.98618 0.9912 3.1245e-006 1.2498e-005 0.14373 0.8204 0.85685 0.0014279 0.92704 0.49588 0.0019227 0.42414 1.6239 1.6218 16.0097 144.9687 0.00025745 -85.4017 0.35695
3.461 0.98806 5.5032e-005 3.8182 0.012002 4.5379e-005 0.0011567 0.22221 0.00065921 0.22287 0.20535 0 0.03284 0.0389 0 1.116 0.34934 0.10251 0.013427 6.249 0.083808 0.00010381 0.8063 0.0067236 0.0075269 0.0014449 0.98618 0.99121 3.1235e-006 1.2494e-005 0.14374 0.8209 0.85714 0.0014277 0.92748 0.49605 0.0019224 0.42415 1.6251 1.623 16.0097 144.9687 0.000257 -85.4035 0.35795
3.462 0.98806 5.5032e-005 3.8182 0.012002 4.5392e-005 0.0011567 0.22222 0.00065921 0.22288 0.20536 0 0.03284 0.0389 0 1.1161 0.34939 0.10253 0.013429 6.2503 0.083819 0.00010383 0.80628 0.0067243 0.0075277 0.0014445 0.98619 0.99121 3.1225e-006 1.249e-005 0.14374 0.82141 0.85743 0.0014275 0.92793 0.49623 0.0019221 0.42416 1.6262 1.6242 16.0097 144.9687 0.00025656 -85.4053 0.35895
3.463 0.98806 5.5032e-005 3.8182 0.012002 4.5405e-005 0.0011567 0.22223 0.00065921 0.22289 0.20537 0 0.032839 0.0389 0 1.1162 0.34943 0.10254 0.013431 6.2517 0.08383 0.00010384 0.80627 0.006725 0.0075284 0.0014441 0.98619 0.99121 3.1215e-006 1.2486e-005 0.14375 0.82192 0.85771 0.0014273 0.92837 0.4964 0.0019218 0.42417 1.6274 1.6254 16.0097 144.9687 0.00025612 -85.4072 0.35995
3.464 0.98806 5.5032e-005 3.8182 0.012002 4.5418e-005 0.0011567 0.22224 0.00065921 0.2229 0.20538 0 0.032839 0.0389 0 1.1163 0.34948 0.10256 0.013433 6.253 0.08384 0.00010386 0.80626 0.0067257 0.0075292 0.0014436 0.9862 0.99122 3.1205e-006 1.2482e-005 0.14376 0.82242 0.85799 0.001427 0.9288 0.49657 0.0019215 0.42419 1.6286 1.6266 16.0097 144.9687 0.00025568 -85.409 0.36095
3.465 0.98806 5.5032e-005 3.8182 0.012002 4.5431e-005 0.0011567 0.22225 0.00065922 0.22291 0.20539 0 0.032838 0.0389 0 1.1164 0.34953 0.10257 0.013434 6.2543 0.083851 0.00010387 0.80625 0.0067264 0.00753 0.0014432 0.9862 0.99122 3.1195e-006 1.2478e-005 0.14376 0.82292 0.85827 0.0014268 0.92924 0.49675 0.0019212 0.4242 1.6297 1.6277 16.0097 144.9687 0.00025524 -85.4108 0.36195
3.466 0.98806 5.5032e-005 3.8182 0.012002 4.5444e-005 0.0011567 0.22226 0.00065922 0.22292 0.2054 0 0.032838 0.0389 0 1.1165 0.34957 0.10259 0.013436 6.2557 0.083862 0.00010389 0.80624 0.0067272 0.0075307 0.0014428 0.98621 0.99123 3.1185e-006 1.2474e-005 0.14377 0.82342 0.85855 0.0014266 0.92967 0.49692 0.0019209 0.42421 1.6309 1.6289 16.0097 144.9688 0.0002548 -85.4126 0.36295
3.467 0.98806 5.5032e-005 3.8182 0.012002 4.5457e-005 0.0011567 0.22227 0.00065922 0.22293 0.20541 0 0.032837 0.0389 0 1.1166 0.34962 0.10261 0.013438 6.257 0.083873 0.0001039 0.80623 0.0067279 0.0075315 0.0014423 0.98622 0.99123 3.1175e-006 1.247e-005 0.14377 0.82392 0.85883 0.0014264 0.9301 0.4971 0.0019206 0.42422 1.6321 1.63 16.0097 144.9688 0.00025437 -85.4143 0.36395
3.468 0.98806 5.5032e-005 3.8182 0.012002 4.547e-005 0.0011567 0.22228 0.00065922 0.22294 0.20542 0 0.032837 0.0389 0 1.1167 0.34966 0.10262 0.01344 6.2584 0.083883 0.00010392 0.80622 0.0067286 0.0075323 0.0014419 0.98622 0.99123 3.1166e-006 1.2466e-005 0.14378 0.82442 0.85911 0.0014262 0.93052 0.49727 0.0019203 0.42424 1.6332 1.6312 16.0097 144.9688 0.00025393 -85.4161 0.36495
3.469 0.98806 5.5032e-005 3.8182 0.012002 4.5483e-005 0.0011568 0.22229 0.00065922 0.22295 0.20543 0 0.032836 0.0389 0 1.1168 0.34971 0.10264 0.013441 6.2597 0.083894 0.00010393 0.80621 0.0067293 0.007533 0.0014415 0.98623 0.99124 3.1156e-006 1.2462e-005 0.14378 0.82492 0.85939 0.001426 0.93095 0.49744 0.00192 0.42425 1.6344 1.6324 16.0097 144.9688 0.0002535 -85.4178 0.36595
3.47 0.98806 5.5032e-005 3.8182 0.012002 4.5496e-005 0.0011568 0.2223 0.00065922 0.22296 0.20544 0 0.032836 0.0389 0 1.1169 0.34976 0.10265 0.013443 6.2611 0.083905 0.00010395 0.8062 0.00673 0.0075338 0.0014411 0.98623 0.99124 3.1147e-006 1.2459e-005 0.14379 0.82541 0.85966 0.0014258 0.93137 0.49762 0.0019197 0.42426 1.6355 1.6335 16.0098 144.9688 0.00025307 -85.4196 0.36695
3.471 0.98806 5.5031e-005 3.8182 0.012002 4.5509e-005 0.0011568 0.22231 0.00065922 0.22297 0.20545 0 0.032835 0.0389 0 1.117 0.3498 0.10267 0.013445 6.2624 0.083916 0.00010396 0.80619 0.0067308 0.0075346 0.0014407 0.98624 0.99124 3.1137e-006 1.2455e-005 0.1438 0.8259 0.85994 0.0014256 0.93178 0.49779 0.0019195 0.42427 1.6367 1.6347 16.0098 144.9689 0.00025265 -85.4213 0.36795
3.472 0.98806 5.5031e-005 3.8182 0.012002 4.5522e-005 0.0011568 0.22232 0.00065922 0.22298 0.20546 0 0.032835 0.0389 0 1.1171 0.34985 0.10269 0.013446 6.2637 0.083926 0.00010398 0.80618 0.0067315 0.0075354 0.0014403 0.98624 0.99125 3.1128e-006 1.2451e-005 0.1438 0.8264 0.86021 0.0014254 0.9322 0.49796 0.0019192 0.42428 1.6378 1.6358 16.0098 144.9689 0.00025222 -85.423 0.36895
3.473 0.98806 5.5031e-005 3.8182 0.012002 4.5535e-005 0.0011568 0.22233 0.00065922 0.22299 0.20547 0 0.032834 0.0389 0 1.1172 0.3499 0.1027 0.013448 6.2651 0.083937 0.00010399 0.80617 0.0067322 0.0075361 0.0014398 0.98625 0.99125 3.1118e-006 1.2447e-005 0.14381 0.82688 0.86048 0.0014252 0.93261 0.49814 0.0019189 0.4243 1.6389 1.637 16.0098 144.9689 0.0002518 -85.4247 0.36995
3.474 0.98806 5.5031e-005 3.8182 0.012002 4.5548e-005 0.0011568 0.22234 0.00065922 0.223 0.20548 0 0.032834 0.0389 0 1.1173 0.34994 0.10272 0.01345 6.2664 0.083948 0.000104 0.80616 0.0067329 0.0075369 0.0014394 0.98625 0.99125 3.1109e-006 1.2444e-005 0.14381 0.82737 0.86075 0.001425 0.93302 0.49831 0.0019186 0.42431 1.6401 1.6381 16.0098 144.9689 0.00025138 -85.4264 0.37095
3.475 0.98806 5.5031e-005 3.8182 0.012002 4.5561e-005 0.0011568 0.22235 0.00065922 0.22301 0.20549 0 0.032833 0.0389 0 1.1174 0.34999 0.10274 0.013452 6.2678 0.083959 0.00010402 0.80615 0.0067336 0.0075377 0.001439 0.98626 0.99126 3.11e-006 1.244e-005 0.14382 0.82786 0.86102 0.0014248 0.93343 0.49849 0.0019184 0.42432 1.6412 1.6392 16.0098 144.9689 0.00025096 -85.428 0.37195
3.476 0.98806 5.5031e-005 3.8182 0.012002 4.5574e-005 0.0011568 0.22236 0.00065922 0.22302 0.2055 0 0.032833 0.0389 0 1.1175 0.35003 0.10275 0.013453 6.2691 0.083969 0.00010403 0.80613 0.0067344 0.0075384 0.0014386 0.98626 0.99126 3.1091e-006 1.2436e-005 0.14383 0.82835 0.86129 0.0014245 0.93384 0.49866 0.0019181 0.42433 1.6423 1.6404 16.0098 144.969 0.00025054 -85.4297 0.37295
3.477 0.98806 5.5031e-005 3.8182 0.012002 4.5587e-005 0.0011568 0.22238 0.00065922 0.22303 0.20551 0 0.032832 0.0389 0 1.1176 0.35008 0.10277 0.013455 6.2705 0.08398 0.00010405 0.80612 0.0067351 0.0075392 0.0014383 0.98627 0.99126 3.1082e-006 1.2433e-005 0.14383 0.82883 0.86156 0.0014243 0.93424 0.49883 0.0019178 0.42434 1.6435 1.6415 16.0098 144.969 0.00025012 -85.4313 0.37395
3.478 0.98806 5.5031e-005 3.8182 0.012002 4.56e-005 0.0011568 0.22239 0.00065922 0.22304 0.20552 0 0.032831 0.0389 0 1.1177 0.35013 0.10278 0.013457 6.2718 0.083991 0.00010406 0.80611 0.0067358 0.00754 0.0014379 0.98627 0.99127 3.1073e-006 1.2429e-005 0.14384 0.82931 0.86182 0.0014241 0.93464 0.49901 0.0019176 0.42436 1.6446 1.6426 16.0098 144.969 0.00024971 -85.433 0.37495
3.479 0.98806 5.5031e-005 3.8182 0.012002 4.5613e-005 0.0011568 0.2224 0.00065922 0.22305 0.20553 0 0.032831 0.0389 0 1.1178 0.35017 0.1028 0.013458 6.2732 0.084002 0.00010408 0.8061 0.0067365 0.0075407 0.0014375 0.98628 0.99127 3.1064e-006 1.2425e-005 0.14384 0.82979 0.86209 0.0014239 0.93504 0.49918 0.0019173 0.42437 1.6457 1.6438 16.0098 144.969 0.0002493 -85.4346 0.37595
3.48 0.98806 5.5031e-005 3.8182 0.012002 4.5626e-005 0.0011568 0.22241 0.00065922 0.22306 0.20554 0 0.03283 0.0389 0 1.1179 0.35022 0.10282 0.01346 6.2745 0.084012 0.00010409 0.80609 0.0067372 0.0075415 0.0014371 0.98628 0.99127 3.1055e-006 1.2422e-005 0.14385 0.83027 0.86235 0.0014237 0.93543 0.49935 0.001917 0.42438 1.6468 1.6449 16.0098 144.969 0.00024889 -85.4362 0.37695
3.481 0.98806 5.5031e-005 3.8182 0.012002 4.5639e-005 0.0011568 0.22242 0.00065922 0.22307 0.20555 0 0.03283 0.0389 0 1.118 0.35026 0.10283 0.013462 6.2759 0.084023 0.00010411 0.80608 0.006738 0.0075423 0.0014367 0.98629 0.99128 3.1046e-006 1.2418e-005 0.14385 0.83075 0.86261 0.0014235 0.93583 0.49952 0.0019168 0.42439 1.6479 1.646 16.0098 144.969 0.00024848 -85.4378 0.37795
3.482 0.98806 5.5031e-005 3.8182 0.012002 4.5652e-005 0.0011568 0.22243 0.00065922 0.22308 0.20556 0 0.032829 0.0389 0 1.1181 0.35031 0.10285 0.013464 6.2772 0.084034 0.00010412 0.80607 0.0067387 0.0075431 0.0014363 0.98629 0.99128 3.1037e-006 1.2415e-005 0.14386 0.83123 0.86288 0.0014233 0.93622 0.4997 0.0019165 0.42441 1.649 1.6471 16.0098 144.9691 0.00024807 -85.4394 0.37895
3.483 0.98806 5.5031e-005 3.8182 0.012002 4.5665e-005 0.0011568 0.22244 0.00065922 0.22309 0.20556 0 0.032829 0.0389 0 1.1182 0.35036 0.10286 0.013465 6.2786 0.084044 0.00010414 0.80606 0.0067394 0.0075438 0.0014359 0.9863 0.99128 3.1029e-006 1.2411e-005 0.14387 0.8317 0.86314 0.0014231 0.9366 0.49987 0.0019163 0.42442 1.6501 1.6482 16.0098 144.9691 0.00024766 -85.441 0.37995
3.484 0.98806 5.5031e-005 3.8182 0.012002 4.5678e-005 0.0011568 0.22245 0.00065922 0.2231 0.20557 0 0.032828 0.0389 0 1.1183 0.3504 0.10288 0.013467 6.2799 0.084055 0.00010415 0.80605 0.0067401 0.0075446 0.0014356 0.9863 0.99129 3.102e-006 1.2408e-005 0.14387 0.83217 0.86339 0.0014229 0.93699 0.50004 0.001916 0.42443 1.6512 1.6493 16.0098 144.9691 0.00024726 -85.4425 0.38095
3.485 0.98806 5.503e-005 3.8182 0.012002 4.5691e-005 0.0011568 0.22246 0.00065922 0.22311 0.20558 0 0.032828 0.0389 0 1.1184 0.35045 0.1029 0.013469 6.2813 0.084066 0.00010417 0.80604 0.0067409 0.0075454 0.0014352 0.98631 0.99129 3.1011e-006 1.2405e-005 0.14388 0.83265 0.86365 0.0014227 0.93737 0.50022 0.0019157 0.42444 1.6523 1.6505 16.0098 144.9691 0.00024686 -85.4441 0.38195
3.486 0.98806 5.503e-005 3.8182 0.012002 4.5705e-005 0.0011568 0.22247 0.00065922 0.22312 0.20559 0 0.032827 0.0389 0 1.1185 0.3505 0.10291 0.013471 6.2826 0.084077 0.00010418 0.80603 0.0067416 0.0075461 0.0014348 0.98631 0.99129 3.1003e-006 1.2401e-005 0.14388 0.83312 0.86391 0.0014225 0.93775 0.50039 0.0019155 0.42445 1.6534 1.6516 16.0098 144.9691 0.00024646 -85.4457 0.38295
3.487 0.98806 5.503e-005 3.8182 0.012001 4.5718e-005 0.0011568 0.22248 0.00065922 0.22313 0.2056 0 0.032827 0.0389 0 1.1186 0.35054 0.10293 0.013472 6.284 0.084087 0.0001042 0.80602 0.0067423 0.0075469 0.0014344 0.98632 0.9913 3.0995e-006 1.2398e-005 0.14389 0.83359 0.86417 0.0014223 0.93813 0.50056 0.0019152 0.42447 1.6545 1.6527 16.0098 144.9692 0.00024606 -85.4472 0.38395
3.488 0.98806 5.503e-005 3.8182 0.012001 4.5731e-005 0.0011568 0.22249 0.00065922 0.22314 0.20561 0 0.032826 0.0389 0 1.1187 0.35059 0.10294 0.013474 6.2853 0.084098 0.00010421 0.80601 0.006743 0.0075477 0.0014341 0.98632 0.9913 3.0986e-006 1.2394e-005 0.1439 0.83405 0.86442 0.0014221 0.93851 0.50074 0.001915 0.42448 1.6556 1.6538 16.0098 144.9692 0.00024566 -85.4487 0.38495
3.489 0.98806 5.503e-005 3.8182 0.012001 4.5744e-005 0.0011568 0.2225 0.00065922 0.22315 0.20562 0 0.032826 0.0389 0 1.1188 0.35063 0.10296 0.013476 6.2867 0.084109 0.00010422 0.806 0.0067437 0.0075484 0.0014337 0.98633 0.9913 3.0978e-006 1.2391e-005 0.1439 0.83452 0.86467 0.0014219 0.93888 0.50091 0.0019148 0.42449 1.6567 1.6549 16.0098 144.9692 0.00024526 -85.4502 0.38595
3.49 0.98806 5.503e-005 3.8182 0.012001 4.5757e-005 0.0011568 0.22251 0.00065922 0.22316 0.20563 0 0.032825 0.0389 0 1.1189 0.35068 0.10298 0.013477 6.288 0.08412 0.00010424 0.80598 0.0067445 0.0075492 0.0014334 0.98633 0.99131 3.097e-006 1.2388e-005 0.14391 0.83498 0.86493 0.0014218 0.93925 0.50108 0.0019145 0.4245 1.6578 1.6559 16.0098 144.9692 0.00024487 -85.4517 0.38695
3.491 0.98806 5.503e-005 3.8182 0.012001 4.577e-005 0.0011568 0.22252 0.00065922 0.22317 0.20564 0 0.032825 0.0389 0 1.119 0.35073 0.10299 0.013479 6.2894 0.08413 0.00010425 0.80597 0.0067452 0.00755 0.001433 0.98634 0.99131 3.0961e-006 1.2385e-005 0.14391 0.83545 0.86518 0.0014216 0.93962 0.50125 0.0019143 0.42452 1.6589 1.657 16.0098 144.9692 0.00024448 -85.4532 0.38795
3.492 0.98806 5.503e-005 3.8182 0.012001 4.5783e-005 0.0011568 0.22253 0.00065922 0.22318 0.20565 0 0.032824 0.0389 0 1.1191 0.35077 0.10301 0.013481 6.2907 0.084141 0.00010427 0.80596 0.0067459 0.0075507 0.0014327 0.98634 0.99131 3.0953e-006 1.2381e-005 0.14392 0.83591 0.86543 0.0014214 0.93999 0.50143 0.001914 0.42453 1.66 1.6581 16.0098 144.9693 0.00024409 -85.4547 0.38895
3.493 0.98806 5.503e-005 3.8182 0.012001 4.5796e-005 0.0011568 0.22254 0.00065922 0.22319 0.20566 0 0.032824 0.0389 0 1.1192 0.35082 0.10303 0.013483 6.2921 0.084152 0.00010428 0.80595 0.0067466 0.0075515 0.0014323 0.98635 0.99132 3.0945e-006 1.2378e-005 0.14392 0.83637 0.86568 0.0014212 0.94036 0.5016 0.0019138 0.42454 1.661 1.6592 16.0098 144.9693 0.0002437 -85.4562 0.38995
3.494 0.98806 5.503e-005 3.8182 0.012001 4.5809e-005 0.0011568 0.22255 0.00065922 0.2232 0.20567 0 0.032823 0.0389 0 1.1193 0.35087 0.10304 0.013484 6.2934 0.084162 0.0001043 0.80594 0.0067473 0.0075523 0.001432 0.98635 0.99132 3.0937e-006 1.2375e-005 0.14393 0.83683 0.86593 0.0014211 0.94072 0.50177 0.0019135 0.42455 1.6621 1.6603 16.0098 144.9693 0.00024331 -85.4576 0.39095
3.495 0.98806 5.503e-005 3.8182 0.012001 4.5822e-005 0.0011568 0.22256 0.00065922 0.22321 0.20568 0 0.032823 0.0389 0 1.1194 0.35091 0.10306 0.013486 6.2948 0.084173 0.00010431 0.80593 0.0067481 0.0075531 0.0014316 0.98636 0.99132 3.0929e-006 1.2372e-005 0.14394 0.83729 0.86617 0.0014209 0.94108 0.50194 0.0019133 0.42457 1.6632 1.6614 16.0098 144.9693 0.00024293 -85.4591 0.39195
3.496 0.98806 5.503e-005 3.8182 0.012001 4.5835e-005 0.0011568 0.22257 0.00065922 0.22322 0.20569 0 0.032822 0.0389 0 1.1195 0.35096 0.10307 0.013488 6.2961 0.084184 0.00010433 0.80592 0.0067488 0.0075538 0.0014313 0.98636 0.99132 3.0921e-006 1.2369e-005 0.14394 0.83774 0.86642 0.0014207 0.94144 0.50212 0.0019131 0.42458 1.6643 1.6624 16.0098 144.9693 0.00024254 -85.4605 0.39295
3.497 0.98806 5.503e-005 3.8182 0.012001 4.5848e-005 0.0011568 0.22258 0.00065922 0.22323 0.2057 0 0.032822 0.0389 0 1.1196 0.351 0.10309 0.013489 6.2975 0.084195 0.00010434 0.80591 0.0067495 0.0075546 0.0014309 0.98637 0.99133 3.0914e-006 1.2365e-005 0.14395 0.8382 0.86666 0.0014205 0.94179 0.50229 0.0019128 0.42459 1.6653 1.6635 16.0098 144.9693 0.00024216 -85.462 0.39395
3.498 0.98806 5.503e-005 3.8182 0.012001 4.5861e-005 0.0011568 0.22259 0.00065922 0.22324 0.20571 0 0.032821 0.0389 0 1.1197 0.35105 0.10311 0.013491 6.2988 0.084205 0.00010436 0.8059 0.0067502 0.0075554 0.0014306 0.98637 0.99133 3.0906e-006 1.2362e-005 0.14395 0.83865 0.86691 0.0014203 0.94215 0.50246 0.0019126 0.4246 1.6664 1.6646 16.0098 144.9694 0.00024178 -85.4634 0.39495
3.499 0.98806 5.503e-005 3.8182 0.012001 4.5874e-005 0.0011568 0.2226 0.00065922 0.22325 0.20572 0 0.032821 0.0389 0 1.1198 0.3511 0.10312 0.013493 6.3002 0.084216 0.00010437 0.80589 0.0067509 0.0075561 0.0014302 0.98637 0.99133 3.0898e-006 1.2359e-005 0.14396 0.8391 0.86715 0.0014202 0.9425 0.50263 0.0019124 0.42462 1.6675 1.6656 16.0098 144.9694 0.0002414 -85.4648 0.39595
3.5 0.98806 5.5029e-005 3.8182 0.012001 4.5887e-005 0.0011568 0.22261 0.00065922 0.22326 0.20573 0 0.03282 0.0389 0 1.1199 0.35114 0.10314 0.013495 6.3015 0.084227 0.00010439 0.80588 0.0067517 0.0075569 0.0014299 0.98638 0.99134 3.089e-006 1.2356e-005 0.14397 0.83955 0.86739 0.00142 0.94285 0.5028 0.0019122 0.42463 1.6685 1.6667 16.0098 144.9694 0.00024102 -85.4662 0.39695
3.501 0.98806 5.5029e-005 3.8182 0.012001 4.59e-005 0.0011568 0.22262 0.00065922 0.22327 0.20574 0 0.03282 0.0389 0 1.12 0.35119 0.10315 0.013496 6.3029 0.084237 0.0001044 0.80587 0.0067524 0.0075577 0.0014296 0.98638 0.99134 3.0883e-006 1.2353e-005 0.14397 0.84 0.86763 0.0014198 0.94319 0.50298 0.0019119 0.42464 1.6696 1.6678 16.0098 144.9694 0.00024065 -85.4676 0.39795
3.502 0.98806 5.5029e-005 3.8182 0.012001 4.5913e-005 0.0011568 0.22263 0.00065922 0.22328 0.20575 0 0.032819 0.0389 0 1.1201 0.35123 0.10317 0.013498 6.3043 0.084248 0.00010442 0.80586 0.0067531 0.0075584 0.0014292 0.98639 0.99134 3.0875e-006 1.235e-005 0.14398 0.84045 0.86787 0.0014196 0.94354 0.50315 0.0019117 0.42465 1.6706 1.6688 16.0098 144.9694 0.00024027 -85.469 0.39895
3.503 0.98806 5.5029e-005 3.8182 0.012001 4.5926e-005 0.0011568 0.22264 0.00065922 0.22329 0.20576 0 0.032819 0.0389 0 1.1202 0.35128 0.10319 0.0135 6.3056 0.084259 0.00010443 0.80585 0.0067538 0.0075592 0.0014289 0.98639 0.99134 3.0868e-006 1.2347e-005 0.14398 0.8409 0.86811 0.0014194 0.94388 0.50332 0.0019115 0.42467 1.6717 1.6699 16.0098 144.9695 0.0002399 -85.4703 0.39995
3.504 0.98806 5.5029e-005 3.8182 0.012001 4.5939e-005 0.0011568 0.22265 0.00065922 0.2233 0.20577 0 0.032818 0.0389 0 1.1203 0.35133 0.1032 0.013502 6.307 0.08427 0.00010444 0.80583 0.0067545 0.00756 0.0014286 0.9864 0.99135 3.086e-006 1.2344e-005 0.14399 0.84134 0.86835 0.0014193 0.94422 0.50349 0.0019113 0.42468 1.6727 1.6709 16.0098 144.9695 0.00023953 -85.4717 0.40095
3.505 0.98806 5.5029e-005 3.8182 0.012001 4.5952e-005 0.0011568 0.22266 0.00065922 0.22331 0.20577 0 0.032817 0.0389 0 1.1204 0.35137 0.10322 0.013503 6.3083 0.08428 0.00010446 0.80582 0.0067553 0.0075607 0.0014283 0.9864 0.99135 3.0853e-006 1.2341e-005 0.14399 0.84178 0.86859 0.0014191 0.94456 0.50366 0.001911 0.42469 1.6738 1.672 16.0098 144.9695 0.00023916 -85.473 0.40195
3.506 0.98806 5.5029e-005 3.8182 0.012001 4.5965e-005 0.0011568 0.22267 0.00065922 0.22332 0.20578 0 0.032817 0.0389 0 1.1205 0.35142 0.10324 0.013505 6.3097 0.084291 0.00010447 0.80581 0.006756 0.0075615 0.001428 0.9864 0.99135 3.0846e-006 1.2338e-005 0.144 0.84223 0.86882 0.0014189 0.94489 0.50384 0.0019108 0.4247 1.6748 1.673 16.0098 144.9695 0.00023879 -85.4744 0.40295
3.507 0.98806 5.5029e-005 3.8182 0.012001 4.5978e-005 0.0011568 0.22268 0.00065922 0.22333 0.20579 0 0.032816 0.0389 0 1.1206 0.35147 0.10325 0.013507 6.311 0.084302 0.00010449 0.8058 0.0067567 0.0075623 0.0014276 0.98641 0.99136 3.0838e-006 1.2335e-005 0.14401 0.84267 0.86906 0.0014188 0.94523 0.50401 0.0019106 0.42472 1.6758 1.6741 16.0098 144.9695 0.00023843 -85.4757 0.40395
3.508 0.98806 5.5029e-005 3.8182 0.012001 4.5991e-005 0.0011568 0.22269 0.00065922 0.22334 0.2058 0 0.032816 0.0389 0 1.1207 0.35151 0.10327 0.013508 6.3124 0.084312 0.0001045 0.80579 0.0067574 0.0075631 0.0014273 0.98641 0.99136 3.0831e-006 1.2332e-005 0.14401 0.84311 0.86929 0.0014186 0.94556 0.50418 0.0019104 0.42473 1.6769 1.6751 16.0098 144.9696 0.00023806 -85.477 0.40495
3.509 0.98806 5.5029e-005 3.8182 0.012001 4.6004e-005 0.0011568 0.2227 0.00065922 0.22335 0.20581 0 0.032815 0.0389 0 1.1208 0.35156 0.10328 0.01351 6.3138 0.084323 0.00010452 0.80578 0.0067581 0.0075638 0.001427 0.98642 0.99136 3.0824e-006 1.233e-005 0.14402 0.84354 0.86953 0.0014184 0.94589 0.50435 0.0019102 0.42474 1.6779 1.6762 16.0098 144.9696 0.0002377 -85.4783 0.40595
3.51 0.98806 5.5029e-005 3.8182 0.012001 4.6017e-005 0.0011568 0.22271 0.00065922 0.22336 0.20582 0 0.032815 0.0389 0 1.1209 0.3516 0.1033 0.013512 6.3151 0.084334 0.00010453 0.80577 0.0067589 0.0075646 0.0014267 0.98642 0.99136 3.0817e-006 1.2327e-005 0.14402 0.84398 0.86976 0.0014183 0.94622 0.50452 0.00191 0.42475 1.6789 1.6772 16.0098 144.9696 0.00023734 -85.4797 0.40695
3.511 0.98806 5.5029e-005 3.8182 0.012001 4.603e-005 0.0011568 0.22272 0.00065922 0.22337 0.20583 0 0.032814 0.0389 0 1.121 0.35165 0.10332 0.013514 6.3165 0.084345 0.00010455 0.80576 0.0067596 0.0075654 0.0014264 0.98642 0.99137 3.081e-006 1.2324e-005 0.14403 0.84442 0.86999 0.0014181 0.94654 0.50469 0.0019098 0.42477 1.68 1.6782 16.0098 144.9696 0.00023698 -85.4809 0.40795
3.512 0.98806 5.5029e-005 3.8182 0.012001 4.6043e-005 0.0011568 0.22273 0.00065922 0.22338 0.20584 0 0.032814 0.0389 0 1.1211 0.3517 0.10333 0.013515 6.3178 0.084355 0.00010456 0.80575 0.0067603 0.0075661 0.0014261 0.98643 0.99137 3.0803e-006 1.2321e-005 0.14404 0.84485 0.87022 0.001418 0.94687 0.50487 0.0019095 0.42478 1.681 1.6793 16.0098 144.9696 0.00023662 -85.4822 0.40895
3.513 0.98806 5.5029e-005 3.8182 0.012001 4.6056e-005 0.0011568 0.22274 0.00065922 0.22339 0.20585 0 0.032813 0.0389 0 1.1212 0.35174 0.10335 0.013517 6.3192 0.084366 0.00010458 0.80574 0.006761 0.0075669 0.0014258 0.98643 0.99137 3.0796e-006 1.2318e-005 0.14404 0.84528 0.87045 0.0014178 0.94719 0.50504 0.0019093 0.42479 1.682 1.6803 16.0098 144.9697 0.00023626 -85.4835 0.40995
3.514 0.98806 5.5028e-005 3.8182 0.012001 4.6069e-005 0.0011568 0.22275 0.00065922 0.2234 0.20586 0 0.032813 0.0389 0 1.1213 0.35179 0.10336 0.013519 6.3206 0.084377 0.00010459 0.80573 0.0067617 0.0075677 0.0014255 0.98644 0.99137 3.0789e-006 1.2316e-005 0.14405 0.84571 0.87068 0.0014177 0.94751 0.50521 0.0019091 0.4248 1.683 1.6813 16.0098 144.9697 0.0002359 -85.4848 0.41095
3.515 0.98806 5.5028e-005 3.8182 0.012001 4.6082e-005 0.0011568 0.22276 0.00065922 0.22341 0.20587 0 0.032812 0.0389 0 1.1214 0.35184 0.10338 0.01352 6.3219 0.084387 0.00010461 0.80572 0.0067625 0.0075684 0.0014252 0.98644 0.99138 3.0782e-006 1.2313e-005 0.14405 0.84614 0.8709 0.0014175 0.94783 0.50538 0.0019089 0.42482 1.684 1.6823 16.0098 144.9697 0.00023555 -85.486 0.41195
3.516 0.98806 5.5028e-005 3.8182 0.012001 4.6095e-005 0.0011568 0.22277 0.00065922 0.22342 0.20588 0 0.032812 0.0389 0 1.1215 0.35188 0.1034 0.013522 6.3233 0.084398 0.00010462 0.80571 0.0067632 0.0075692 0.0014249 0.98644 0.99138 3.0775e-006 1.231e-005 0.14406 0.84657 0.87113 0.0014174 0.94814 0.50555 0.0019087 0.42483 1.685 1.6833 16.0098 144.9697 0.0002352 -85.4873 0.41295
3.517 0.98806 5.5028e-005 3.8182 0.012001 4.6109e-005 0.0011568 0.22278 0.00065922 0.22343 0.20589 0 0.032811 0.0389 0 1.1216 0.35193 0.10341 0.013524 6.3246 0.084409 0.00010464 0.8057 0.0067639 0.00757 0.0014246 0.98645 0.99138 3.0768e-006 1.2307e-005 0.14406 0.847 0.87136 0.0014172 0.94846 0.50572 0.0019085 0.42484 1.6861 1.6844 16.0098 144.9697 0.00023484 -85.4885 0.41395
3.518 0.98806 5.5028e-005 3.8182 0.012001 4.6122e-005 0.0011568 0.22279 0.00065922 0.22344 0.2059 0 0.032811 0.0389 0 1.1217 0.35197 0.10343 0.013526 6.326 0.08442 0.00010465 0.80569 0.0067646 0.0075707 0.0014243 0.98645 0.99138 3.0762e-006 1.2305e-005 0.14407 0.84743 0.87158 0.0014171 0.94877 0.50589 0.0019083 0.42485 1.6871 1.6854 16.0098 144.9697 0.00023449 -85.4898 0.41495
3.519 0.98806 5.5028e-005 3.8182 0.012001 4.6135e-005 0.0011568 0.2228 0.00065922 0.22345 0.20591 0 0.03281 0.0389 0 1.1218 0.35202 0.10344 0.013527 6.3274 0.08443 0.00010466 0.80567 0.0067653 0.0075715 0.001424 0.98646 0.99139 3.0755e-006 1.2302e-005 0.14408 0.84785 0.8718 0.0014169 0.94908 0.50607 0.0019081 0.42487 1.6881 1.6864 16.0097 144.9698 0.00023415 -85.491 0.41595
3.52 0.98806 5.5028e-005 3.8182 0.012001 4.6148e-005 0.0011568 0.22281 0.00065922 0.22346 0.20592 0 0.03281 0.0389 0 1.1219 0.35207 0.10346 0.013529 6.3287 0.084441 0.00010468 0.80566 0.0067661 0.0075723 0.0014237 0.98646 0.99139 3.0748e-006 1.2299e-005 0.14408 0.84827 0.87203 0.0014168 0.94939 0.50624 0.0019079 0.42488 1.6891 1.6874 16.0097 144.9698 0.0002338 -85.4922 0.41695
3.521 0.98806 5.5028e-005 3.8182 0.012001 4.6161e-005 0.0011568 0.22282 0.00065922 0.22347 0.20592 0 0.032809 0.0389 0 1.122 0.35211 0.10348 0.013531 6.3301 0.084452 0.00010469 0.80565 0.0067668 0.0075731 0.0014234 0.98646 0.99139 3.0742e-006 1.2297e-005 0.14409 0.8487 0.87225 0.0014166 0.94969 0.50641 0.0019077 0.42489 1.6901 1.6884 16.0097 144.9698 0.00023345 -85.4934 0.41795
3.522 0.98806 5.5028e-005 3.8182 0.012001 4.6174e-005 0.0011569 0.22283 0.00065922 0.22348 0.20593 0 0.032809 0.0389 0 1.1221 0.35216 0.10349 0.013532 6.3315 0.084462 0.00010471 0.80564 0.0067675 0.0075738 0.0014231 0.98647 0.99139 3.0735e-006 1.2294e-005 0.14409 0.84912 0.87247 0.0014165 0.95 0.50658 0.0019075 0.4249 1.6911 1.6894 16.0097 144.9698 0.00023311 -85.4946 0.41895
3.523 0.98806 5.5028e-005 3.8182 0.012001 4.6187e-005 0.0011569 0.22284 0.00065922 0.22349 0.20594 0 0.032808 0.0389 0 1.1222 0.35221 0.10351 0.013534 6.3328 0.084473 0.00010472 0.80563 0.0067682 0.0075746 0.0014229 0.98647 0.9914 3.0729e-006 1.2292e-005 0.1441 0.84954 0.87269 0.0014163 0.9503 0.50675 0.0019073 0.42492 1.6921 1.6904 16.0097 144.9698 0.00023277 -85.4958 0.41995
3.524 0.98806 5.5028e-005 3.8182 0.012001 4.62e-005 0.0011569 0.22285 0.00065922 0.2235 0.20595 0 0.032808 0.0389 0 1.1223 0.35225 0.10353 0.013536 6.3342 0.084484 0.00010474 0.80562 0.0067689 0.0075754 0.0014226 0.98647 0.9914 3.0723e-006 1.2289e-005 0.1441 0.84995 0.87291 0.0014161 0.9506 0.50692 0.0019072 0.42493 1.6931 1.6914 16.0097 144.9699 0.00023242 -85.497 0.42095
3.525 0.98806 5.5028e-005 3.8182 0.012001 4.6213e-005 0.0011569 0.22285 0.00065922 0.22351 0.20596 0 0.032807 0.0389 0 1.1224 0.3523 0.10354 0.013538 6.3356 0.084494 0.00010475 0.80561 0.0067697 0.0075761 0.0014223 0.98648 0.9914 3.0716e-006 1.2286e-005 0.14411 0.85037 0.87312 0.001416 0.9509 0.50709 0.001907 0.42494 1.694 1.6924 16.0097 144.9699 0.00023208 -85.4982 0.42195
3.526 0.98806 5.5028e-005 3.8182 0.012001 4.6226e-005 0.0011569 0.22286 0.00065922 0.22352 0.20597 0 0.032807 0.0389 0 1.1225 0.35234 0.10356 0.013539 6.3369 0.084505 0.00010477 0.8056 0.0067704 0.0075769 0.001422 0.98648 0.9914 3.071e-006 1.2284e-005 0.14412 0.85079 0.87334 0.0014158 0.95119 0.50726 0.0019068 0.42496 1.695 1.6934 16.0097 144.9699 0.00023175 -85.4993 0.42295
3.527 0.98806 5.5028e-005 3.8182 0.012001 4.6239e-005 0.0011569 0.22287 0.00065922 0.22353 0.20598 0 0.032806 0.0389 0 1.1226 0.35239 0.10357 0.013541 6.3383 0.084516 0.00010478 0.80559 0.0067711 0.0075777 0.0014217 0.98648 0.99141 3.0704e-006 1.2281e-005 0.14412 0.8512 0.87356 0.0014157 0.95149 0.50743 0.0019066 0.42497 1.696 1.6944 16.0097 144.9699 0.00023141 -85.5005 0.42395
3.528 0.98806 5.5027e-005 3.8182 0.012001 4.6252e-005 0.0011569 0.22288 0.00065922 0.22354 0.20599 0 0.032806 0.0389 0 1.1227 0.35244 0.10359 0.013543 6.3396 0.084527 0.0001048 0.80558 0.0067718 0.0075784 0.0014215 0.98649 0.99141 3.0697e-006 1.2279e-005 0.14413 0.85161 0.87377 0.0014155 0.95178 0.5076 0.0019064 0.42498 1.697 1.6953 16.0097 144.9699 0.00023107 -85.5016 0.42495
3.529 0.98806 5.5027e-005 3.8182 0.012001 4.6265e-005 0.0011569 0.22289 0.00065922 0.22355 0.206 0 0.032805 0.0389 0 1.1228 0.35248 0.10361 0.013544 6.341 0.084537 0.00010481 0.80557 0.0067725 0.0075792 0.0014212 0.98649 0.99141 3.0691e-006 1.2276e-005 0.14413 0.85202 0.87399 0.0014154 0.95207 0.50777 0.0019062 0.42499 1.698 1.6963 16.0097 144.97 0.00023074 -85.5028 0.42595
3.53 0.98806 5.5027e-005 3.8182 0.012001 4.6278e-005 0.0011569 0.2229 0.00065922 0.22356 0.20601 0 0.032805 0.0389 0 1.1229 0.35253 0.10362 0.013546 6.3424 0.084548 0.00010483 0.80556 0.0067732 0.00758 0.0014209 0.9865 0.99141 3.0685e-006 1.2274e-005 0.14414 0.85243 0.8742 0.0014152 0.95236 0.50795 0.001906 0.42501 1.6989 1.6973 16.0097 144.97 0.0002304 -85.5039 0.42695
3.531 0.98806 5.5027e-005 3.8182 0.012001 4.6291e-005 0.0011569 0.22291 0.00065922 0.22357 0.20602 0 0.032804 0.0389 0 1.123 0.35257 0.10364 0.013548 6.3437 0.084559 0.00010484 0.80555 0.006774 0.0075807 0.0014207 0.9865 0.99141 3.0679e-006 1.2271e-005 0.14415 0.85284 0.87441 0.0014151 0.95265 0.50812 0.0019059 0.42502 1.6999 1.6983 16.0097 144.97 0.00023007 -85.505 0.42795
3.532 0.98806 5.5027e-005 3.8182 0.012001 4.6304e-005 0.0011569 0.22292 0.00065922 0.22358 0.20603 0 0.032804 0.0389 0 1.1231 0.35262 0.10365 0.01355 6.3451 0.084569 0.00010486 0.80554 0.0067747 0.0075815 0.0014204 0.9865 0.99142 3.0673e-006 1.2269e-005 0.14415 0.85325 0.87463 0.001415 0.95293 0.50829 0.0019057 0.42503 1.7009 1.6993 16.0097 144.97 0.00022974 -85.5062 0.42895
3.533 0.98806 5.5027e-005 3.8182 0.012001 4.6317e-005 0.0011569 0.22293 0.00065922 0.22359 0.20604 0 0.032803 0.0389 0 1.1232 0.35267 0.10367 0.013551 6.3465 0.08458 0.00010487 0.80552 0.0067754 0.0075823 0.0014201 0.98651 0.99142 3.0667e-006 1.2267e-005 0.14416 0.85366 0.87484 0.0014148 0.95322 0.50846 0.0019055 0.42504 1.7019 1.7002 16.0097 144.97 0.00022941 -85.5073 0.42995
3.534 0.98806 5.5027e-005 3.8182 0.012001 4.633e-005 0.0011569 0.22294 0.00065922 0.2236 0.20605 0 0.032803 0.0389 0 1.1233 0.35271 0.10369 0.013553 6.3479 0.084591 0.00010488 0.80551 0.0067761 0.0075831 0.0014199 0.98651 0.99142 3.0661e-006 1.2264e-005 0.14416 0.85406 0.87505 0.0014147 0.9535 0.50863 0.0019053 0.42506 1.7028 1.7012 16.0097 144.9701 0.00022909 -85.5084 0.43095
3.535 0.98806 5.5027e-005 3.8182 0.012001 4.6343e-005 0.0011569 0.22295 0.00065922 0.22361 0.20605 0 0.032802 0.0389 0 1.1234 0.35276 0.1037 0.013555 6.3492 0.084601 0.0001049 0.8055 0.0067768 0.0075838 0.0014196 0.98651 0.99142 3.0655e-006 1.2262e-005 0.14417 0.85447 0.87526 0.0014146 0.95378 0.5088 0.0019051 0.42507 1.7038 1.7022 16.0097 144.9701 0.00022876 -85.5095 0.43195
3.536 0.98806 5.5027e-005 3.8182 0.012001 4.6356e-005 0.0011569 0.22296 0.00065922 0.22362 0.20606 0 0.032802 0.0389 0 1.1235 0.35281 0.10372 0.013556 6.3506 0.084612 0.00010491 0.80549 0.0067776 0.0075846 0.0014194 0.98652 0.99143 3.0649e-006 1.2259e-005 0.14417 0.85487 0.87546 0.0014144 0.95406 0.50897 0.001905 0.42508 1.7047 1.7031 16.0097 144.9701 0.00022843 -85.5106 0.43295
3.537 0.98806 5.5027e-005 3.8182 0.012001 4.6369e-005 0.0011569 0.22297 0.00065922 0.22363 0.20607 0 0.032801 0.0389 0 1.1236 0.35285 0.10374 0.013558 6.352 0.084623 0.00010493 0.80548 0.0067783 0.0075854 0.0014191 0.98652 0.99143 3.0643e-006 1.2257e-005 0.14418 0.85527 0.87567 0.0014143 0.95433 0.50914 0.0019048 0.42509 1.7057 1.7041 16.0097 144.9701 0.00022811 -85.5116 0.43395
3.538 0.98806 5.5027e-005 3.8182 0.012001 4.6382e-005 0.0011569 0.22298 0.00065922 0.22364 0.20608 0 0.032801 0.0389 0 1.1237 0.3529 0.10375 0.01356 6.3533 0.084633 0.00010494 0.80547 0.006779 0.0075861 0.0014188 0.98652 0.99143 3.0637e-006 1.2255e-005 0.14419 0.85567 0.87588 0.0014142 0.95461 0.50931 0.0019046 0.42511 1.7067 1.7051 16.0097 144.9701 0.00022779 -85.5127 0.43495
3.539 0.98806 5.5027e-005 3.8182 0.012001 4.6395e-005 0.0011569 0.22299 0.00065922 0.22365 0.20609 0 0.0328 0.0389 0 1.1238 0.35294 0.10377 0.013562 6.3547 0.084644 0.00010496 0.80546 0.0067797 0.0075869 0.0014186 0.98653 0.99143 3.0631e-006 1.2252e-005 0.14419 0.85607 0.87608 0.001414 0.95488 0.50948 0.0019044 0.42512 1.7076 1.706 16.0097 144.9702 0.00022747 -85.5138 0.43595
3.54 0.98806 5.5027e-005 3.8182 0.012001 4.6408e-005 0.0011569 0.223 0.00065922 0.22366 0.2061 0 0.0328 0.0389 0 1.1239 0.35299 0.10378 0.013563 6.3561 0.084655 0.00010497 0.80545 0.0067804 0.0075877 0.0014183 0.98653 0.99143 3.0626e-006 1.225e-005 0.1442 0.85647 0.87629 0.0014139 0.95515 0.50965 0.0019043 0.42513 1.7086 1.707 16.0097 144.9702 0.00022715 -85.5148 0.43695
3.541 0.98806 5.5027e-005 3.8182 0.012001 4.6421e-005 0.0011569 0.22301 0.00065922 0.22367 0.20611 0 0.032799 0.0389 0 1.124 0.35304 0.1038 0.013565 6.3574 0.084666 0.00010499 0.80544 0.0067812 0.0075884 0.0014181 0.98653 0.99144 3.062e-006 1.2248e-005 0.1442 0.85686 0.87649 0.0014138 0.95542 0.50982 0.0019041 0.42515 1.7095 1.7079 16.0096 144.9702 0.00022683 -85.5159 0.43795
3.542 0.98806 5.5027e-005 3.8182 0.012001 4.6434e-005 0.0011569 0.22302 0.00065922 0.22367 0.20612 0 0.032799 0.0389 0 1.1241 0.35308 0.10382 0.013567 6.3588 0.084676 0.000105 0.80543 0.0067819 0.0075892 0.0014178 0.98654 0.99144 3.0614e-006 1.2246e-005 0.14421 0.85726 0.8767 0.0014136 0.95569 0.50999 0.0019039 0.42516 1.7104 1.7089 16.0096 144.9702 0.00022651 -85.5169 0.43895
3.543 0.98806 5.5026e-005 3.8182 0.012001 4.6447e-005 0.0011569 0.22303 0.00065922 0.22368 0.20613 0 0.032798 0.0389 0 1.1242 0.35313 0.10383 0.013569 6.3602 0.084687 0.00010502 0.80542 0.0067826 0.00759 0.0014176 0.98654 0.99144 3.0609e-006 1.2243e-005 0.14422 0.85765 0.8769 0.0014135 0.95596 0.51016 0.0019038 0.42517 1.7114 1.7098 16.0096 144.9702 0.0002262 -85.518 0.43995
3.544 0.98806 5.5026e-005 3.8182 0.012001 4.646e-005 0.0011569 0.22304 0.00065922 0.22369 0.20614 0 0.032798 0.0389 0 1.1243 0.35318 0.10385 0.01357 6.3616 0.084698 0.00010503 0.80541 0.0067833 0.0075907 0.0014174 0.98654 0.99144 3.0603e-006 1.2241e-005 0.14422 0.85805 0.8771 0.0014134 0.95622 0.51033 0.0019036 0.42518 1.7123 1.7108 16.0096 144.9702 0.00022588 -85.519 0.44095
3.545 0.98806 5.5026e-005 3.8182 0.012001 4.6473e-005 0.0011569 0.22305 0.00065922 0.2237 0.20615 0 0.032797 0.0389 0 1.1244 0.35322 0.10386 0.013572 6.3629 0.084708 0.00010505 0.8054 0.006784 0.0075915 0.0014171 0.98654 0.99145 3.0598e-006 1.2239e-005 0.14423 0.85844 0.8773 0.0014133 0.95649 0.5105 0.0019034 0.4252 1.7133 1.7117 16.0096 144.9703 0.00022557 -85.52 0.44195
3.546 0.98806 5.5026e-005 3.8182 0.012001 4.6486e-005 0.0011569 0.22306 0.00065922 0.22371 0.20616 0 0.032797 0.0389 0 1.1245 0.35327 0.10388 0.013574 6.3643 0.084719 0.00010506 0.80539 0.0067848 0.0075923 0.0014169 0.98655 0.99145 3.0592e-006 1.2237e-005 0.14423 0.85883 0.8775 0.0014131 0.95675 0.51067 0.0019033 0.42521 1.7142 1.7126 16.0096 144.9703 0.00022526 -85.521 0.44295
3.547 0.98806 5.5026e-005 3.8182 0.012001 4.6499e-005 0.0011569 0.22307 0.00065922 0.22372 0.20616 0 0.032796 0.0389 0 1.1246 0.35331 0.1039 0.013575 6.3657 0.08473 0.00010507 0.80538 0.0067855 0.007593 0.0014166 0.98655 0.99145 3.0587e-006 1.2235e-005 0.14424 0.85922 0.8777 0.001413 0.95701 0.51084 0.0019031 0.42522 1.7151 1.7136 16.0096 144.9703 0.00022494 -85.5221 0.44395
3.548 0.98806 5.5026e-005 3.8182 0.012001 4.6513e-005 0.0011569 0.22308 0.00065922 0.22373 0.20617 0 0.032796 0.0389 0 1.1247 0.35336 0.10391 0.013577 6.367 0.08474 0.00010509 0.80536 0.0067862 0.0075938 0.0014164 0.98655 0.99145 3.0581e-006 1.2232e-005 0.14424 0.85961 0.8779 0.0014129 0.95726 0.51101 0.0019029 0.42524 1.7161 1.7145 16.0096 144.9703 0.00022464 -85.5231 0.44495
3.549 0.98806 5.5026e-005 3.8182 0.012001 4.6526e-005 0.0011569 0.22309 0.00065922 0.22374 0.20618 0 0.032795 0.0389 0 1.1248 0.35341 0.10393 0.013579 6.3684 0.084751 0.0001051 0.80535 0.0067869 0.0075946 0.0014162 0.98656 0.99145 3.0576e-006 1.223e-005 0.14425 0.85999 0.8781 0.0014128 0.95752 0.51118 0.0019028 0.42525 1.717 1.7154 16.0096 144.9703 0.00022433 -85.524 0.44595
3.55 0.98806 5.5026e-005 3.8182 0.012001 4.6539e-005 0.0011569 0.2231 0.00065922 0.22375 0.20619 0 0.032795 0.0389 0 1.1249 0.35345 0.10394 0.013581 6.3698 0.084762 0.00010512 0.80534 0.0067876 0.0075953 0.0014159 0.98656 0.99146 3.0571e-006 1.2228e-005 0.14426 0.86038 0.87829 0.0014127 0.95778 0.51135 0.0019026 0.42526 1.7179 1.7164 16.0096 144.9704 0.00022402 -85.525 0.44695
3.551 0.98806 5.5026e-005 3.8182 0.012001 4.6552e-005 0.0011569 0.22311 0.00065922 0.22376 0.2062 0 0.032794 0.0389 0 1.125 0.3535 0.10396 0.013582 6.3712 0.084772 0.00010513 0.80533 0.0067883 0.0075961 0.0014157 0.98656 0.99146 3.0565e-006 1.2226e-005 0.14426 0.86076 0.87849 0.0014126 0.95803 0.51152 0.0019025 0.42527 1.7188 1.7173 16.0096 144.9704 0.00022371 -85.526 0.44795
3.552 0.98806 5.5026e-005 3.8182 0.012001 4.6565e-005 0.0011569 0.22312 0.00065922 0.22377 0.20621 0 0.032794 0.0389 0 1.1251 0.35355 0.10398 0.013584 6.3725 0.084783 0.00010515 0.80532 0.0067891 0.0075969 0.0014155 0.98657 0.99146 3.056e-006 1.2224e-005 0.14427 0.86114 0.87868 0.0014125 0.95828 0.51168 0.0019023 0.42529 1.7198 1.7182 16.0096 144.9704 0.00022341 -85.527 0.44895
3.553 0.98806 5.5026e-005 3.8182 0.012001 4.6578e-005 0.0011569 0.22313 0.00065922 0.22378 0.20622 0 0.032793 0.0389 0 1.1252 0.35359 0.10399 0.013586 6.3739 0.084794 0.00010516 0.80531 0.0067898 0.0075977 0.0014153 0.98657 0.99146 3.0555e-006 1.2222e-005 0.14427 0.86153 0.87888 0.0014123 0.95853 0.51185 0.0019021 0.4253 1.7207 1.7192 16.0096 144.9704 0.00022311 -85.528 0.44995
3.554 0.98806 5.5026e-005 3.8182 0.012 4.6591e-005 0.0011569 0.22314 0.00065922 0.22379 0.20623 0 0.032793 0.0389 0 1.1253 0.35364 0.10401 0.013587 6.3753 0.084804 0.00010518 0.8053 0.0067905 0.0075984 0.001415 0.98657 0.99146 3.055e-006 1.222e-005 0.14428 0.86191 0.87907 0.0014122 0.95878 0.51202 0.001902 0.42531 1.7216 1.7201 16.0096 144.9704 0.0002228 -85.5289 0.45095
3.555 0.98806 5.5026e-005 3.8182 0.012 4.6604e-005 0.0011569 0.22315 0.00065922 0.2238 0.20624 0 0.032792 0.0389 0 1.1254 0.35368 0.10403 0.013589 6.3767 0.084815 0.00010519 0.80529 0.0067912 0.0075992 0.0014148 0.98657 0.99146 3.0544e-006 1.2218e-005 0.14428 0.86229 0.87927 0.0014121 0.95903 0.51219 0.0019018 0.42533 1.7225 1.721 16.0095 144.9705 0.0002225 -85.5299 0.45195
3.556 0.98806 5.5026e-005 3.8182 0.012 4.6617e-005 0.0011569 0.22315 0.00065922 0.22381 0.20625 0 0.032792 0.0389 0 1.1255 0.35373 0.10404 0.013591 6.378 0.084826 0.00010521 0.80528 0.0067919 0.0076 0.0014146 0.98658 0.99147 3.0539e-006 1.2216e-005 0.14429 0.86267 0.87946 0.001412 0.95927 0.51236 0.0019017 0.42534 1.7234 1.7219 16.0095 144.9705 0.0002222 -85.5308 0.45295
3.557 0.98806 5.5025e-005 3.8182 0.012 4.663e-005 0.0011569 0.22316 0.00065922 0.22382 0.20626 0 0.032791 0.0389 0 1.1256 0.35378 0.10406 0.013593 6.3794 0.084836 0.00010522 0.80527 0.0067927 0.0076007 0.0014144 0.98658 0.99147 3.0534e-006 1.2214e-005 0.1443 0.86304 0.87965 0.0014119 0.95951 0.51253 0.0019015 0.42535 1.7243 1.7228 16.0095 144.9705 0.00022191 -85.5318 0.45395
3.558 0.98806 5.5025e-005 3.8182 0.012 4.6643e-005 0.0011569 0.22317 0.00065922 0.22383 0.20626 0 0.032791 0.0389 0 1.1257 0.35382 0.10407 0.013594 6.3808 0.084847 0.00010524 0.80526 0.0067934 0.0076015 0.0014141 0.98658 0.99147 3.0529e-006 1.2212e-005 0.1443 0.86342 0.87984 0.0014117 0.95976 0.5127 0.0019014 0.42536 1.7252 1.7237 16.0095 144.9705 0.00022161 -85.5327 0.45495
3.559 0.98806 5.5025e-005 3.8182 0.012 4.6656e-005 0.0011569 0.22318 0.00065922 0.22384 0.20627 0 0.03279 0.0389 0 1.1257 0.35387 0.10409 0.013596 6.3822 0.084858 0.00010525 0.80525 0.0067941 0.0076023 0.0014139 0.98659 0.99147 3.0524e-006 1.221e-005 0.14431 0.86379 0.88003 0.0014116 0.96 0.51287 0.0019012 0.42538 1.7261 1.7246 16.0095 144.9705 0.00022131 -85.5336 0.45595
3.56 0.98806 5.5025e-005 3.8182 0.012 4.6669e-005 0.0011569 0.22319 0.00065922 0.22385 0.20628 0 0.03279 0.0389 0 1.1258 0.35392 0.10411 0.013598 6.3836 0.084868 0.00010526 0.80524 0.0067948 0.007603 0.0014137 0.98659 0.99147 3.0519e-006 1.2208e-005 0.14431 0.86417 0.88022 0.0014115 0.96024 0.51304 0.0019011 0.42539 1.727 1.7255 16.0095 144.9706 0.00022102 -85.5345 0.45695
3.561 0.98806 5.5025e-005 3.8182 0.012 4.6682e-005 0.0011569 0.2232 0.00065922 0.22386 0.20629 0 0.032789 0.0389 0 1.1259 0.35396 0.10412 0.013599 6.3849 0.084879 0.00010528 0.80523 0.0067955 0.0076038 0.0014135 0.98659 0.99148 3.0514e-006 1.2206e-005 0.14432 0.86454 0.88041 0.0014114 0.96047 0.51321 0.0019009 0.4254 1.7279 1.7264 16.0095 144.9706 0.00022072 -85.5355 0.45795
3.562 0.98806 5.5025e-005 3.8182 0.012 4.6695e-005 0.0011569 0.22321 0.00065922 0.22387 0.2063 0 0.032789 0.0389 0 1.126 0.35401 0.10414 0.013601 6.3863 0.08489 0.00010529 0.80522 0.0067963 0.0076046 0.0014133 0.98659 0.99148 3.0509e-006 1.2204e-005 0.14433 0.86491 0.88059 0.0014113 0.96071 0.51338 0.0019008 0.42542 1.7288 1.7273 16.0095 144.9706 0.00022043 -85.5364 0.45895
3.563 0.98806 5.5025e-005 3.8182 0.012 4.6708e-005 0.0011569 0.22322 0.00065922 0.22388 0.20631 0 0.032789 0.0389 0 1.1261 0.35405 0.10415 0.013603 6.3877 0.0849 0.00010531 0.8052 0.006797 0.0076053 0.0014131 0.9866 0.99148 3.0504e-006 1.2202e-005 0.14433 0.86528 0.88078 0.0014112 0.96094 0.51355 0.0019006 0.42543 1.7297 1.7282 16.0095 144.9706 0.00022014 -85.5373 0.45995
3.564 0.98806 5.5025e-005 3.8182 0.012 4.6721e-005 0.0011569 0.22323 0.00065922 0.22389 0.20632 0 0.032788 0.0389 0 1.1262 0.3541 0.10417 0.013604 6.3891 0.084911 0.00010532 0.80519 0.0067977 0.0076061 0.0014128 0.9866 0.99148 3.05e-006 1.22e-005 0.14434 0.86565 0.88097 0.001411 0.96118 0.51371 0.0019005 0.42544 1.7306 1.7291 16.0095 144.9706 0.00021985 -85.5382 0.46095
3.565 0.98806 5.5025e-005 3.8182 0.012 4.6734e-005 0.0011569 0.22324 0.00065922 0.2239 0.20633 0 0.032788 0.0389 0 1.1263 0.35415 0.10419 0.013606 6.3905 0.084922 0.00010534 0.80518 0.0067984 0.0076069 0.0014126 0.9866 0.99148 3.0495e-006 1.2198e-005 0.14434 0.86602 0.88115 0.0014109 0.96141 0.51388 0.0019004 0.42545 1.7315 1.73 16.0095 144.9707 0.00021956 -85.539 0.46195
3.566 0.98806 5.5025e-005 3.8182 0.012 4.6747e-005 0.0011569 0.22325 0.00065922 0.2239 0.20634 0 0.032787 0.0389 0 1.1264 0.35419 0.1042 0.013608 6.3918 0.084932 0.00010535 0.80517 0.0067991 0.0076076 0.0014124 0.98661 0.99148 3.049e-006 1.2196e-005 0.14435 0.86638 0.88134 0.0014108 0.96164 0.51405 0.0019002 0.42547 1.7324 1.7309 16.0095 144.9707 0.00021927 -85.5399 0.46295
3.567 0.98806 5.5025e-005 3.8182 0.012 4.676e-005 0.0011569 0.22326 0.00065922 0.22391 0.20635 0 0.032787 0.0389 0 1.1265 0.35424 0.10422 0.01361 6.3932 0.084943 0.00010537 0.80516 0.0067998 0.0076084 0.0014122 0.98661 0.99149 3.0485e-006 1.2194e-005 0.14435 0.86675 0.88152 0.0014107 0.96187 0.51422 0.0019001 0.42548 1.7333 1.7318 16.0094 144.9707 0.00021899 -85.5408 0.46395
3.568 0.98806 5.5025e-005 3.8182 0.012 4.6773e-005 0.0011569 0.22327 0.00065922 0.22392 0.20635 0 0.032786 0.0389 0 1.1266 0.35429 0.10423 0.013611 6.3946 0.084954 0.00010538 0.80515 0.0068006 0.0076092 0.001412 0.98661 0.99149 3.0481e-006 1.2192e-005 0.14436 0.86712 0.8817 0.0014106 0.96209 0.51439 0.0018999 0.42549 1.7341 1.7327 16.0094 144.9707 0.0002187 -85.5417 0.46495
3.569 0.98806 5.5025e-005 3.8182 0.012 4.6786e-005 0.0011569 0.22328 0.00065922 0.22393 0.20636 0 0.032786 0.0389 0 1.1267 0.35433 0.10425 0.013613 6.396 0.084964 0.0001054 0.80514 0.0068013 0.0076099 0.0014118 0.98661 0.99149 3.0476e-006 1.219e-005 0.14437 0.86748 0.88188 0.0014105 0.96232 0.51456 0.0018998 0.42551 1.735 1.7336 16.0094 144.9707 0.00021842 -85.5425 0.46595
3.57 0.98806 5.5025e-005 3.8182 0.012 4.6799e-005 0.0011569 0.22329 0.00065922 0.22394 0.20637 0 0.032785 0.0389 0 1.1268 0.35438 0.10427 0.013615 6.3974 0.084975 0.00010541 0.80513 0.006802 0.0076107 0.0014116 0.98662 0.99149 3.0471e-006 1.2188e-005 0.14437 0.86784 0.88207 0.0014104 0.96254 0.51473 0.0018997 0.42552 1.7359 1.7345 16.0094 144.9708 0.00021813 -85.5434 0.46695
3.571 0.98806 5.5024e-005 3.8182 0.012 4.6812e-005 0.0011569 0.2233 0.00065922 0.22395 0.20638 0 0.032785 0.0389 0 1.1269 0.35442 0.10428 0.013616 6.3987 0.084986 0.00010543 0.80512 0.0068027 0.0076115 0.0014114 0.98662 0.99149 3.0467e-006 1.2187e-005 0.14438 0.8682 0.88225 0.0014103 0.96277 0.51489 0.0018995 0.42553 1.7368 1.7353 16.0094 144.9708 0.00021785 -85.5443 0.46795
3.572 0.98806 5.5024e-005 3.8182 0.012 4.6825e-005 0.0011569 0.22331 0.00065922 0.22396 0.20639 0 0.032784 0.0389 0 1.127 0.35447 0.1043 0.013618 6.4001 0.084996 0.00010544 0.80511 0.0068034 0.0076122 0.0014112 0.98662 0.9915 3.0462e-006 1.2185e-005 0.14438 0.86856 0.88243 0.0014102 0.96299 0.51506 0.0018994 0.42554 1.7376 1.7362 16.0094 144.9708 0.00021757 -85.5451 0.46895
3.573 0.98806 5.5024e-005 3.8182 0.012 4.6838e-005 0.001157 0.22332 0.00065922 0.22397 0.2064 0 0.032784 0.0389 0 1.1271 0.35452 0.10432 0.01362 6.4015 0.085007 0.00010545 0.8051 0.0068042 0.007613 0.001411 0.98662 0.9915 3.0457e-006 1.2183e-005 0.14439 0.86892 0.88261 0.0014101 0.96321 0.51523 0.0018992 0.42556 1.7385 1.7371 16.0094 144.9708 0.00021729 -85.5459 0.46995
3.574 0.98806 5.5024e-005 3.8182 0.012 4.6851e-005 0.001157 0.22333 0.00065922 0.22398 0.20641 0 0.032783 0.0389 0 1.1272 0.35456 0.10433 0.013622 6.4029 0.085018 0.00010547 0.80509 0.0068049 0.0076138 0.0014108 0.98663 0.9915 3.0453e-006 1.2181e-005 0.14439 0.86928 0.88279 0.00141 0.96343 0.5154 0.0018991 0.42557 1.7394 1.738 16.0094 144.9708 0.00021701 -85.5468 0.47095
3.575 0.98806 5.5024e-005 3.8182 0.012 4.6864e-005 0.001157 0.22333 0.00065922 0.22399 0.20642 0 0.032783 0.0389 0 1.1273 0.35461 0.10435 0.013623 6.4043 0.085028 0.00010548 0.80508 0.0068056 0.0076146 0.0014106 0.98663 0.9915 3.0449e-006 1.2179e-005 0.1444 0.86963 0.88296 0.0014099 0.96365 0.51557 0.001899 0.42558 1.7402 1.7388 16.0094 144.9709 0.00021673 -85.5476 0.47195
3.576 0.98806 5.5024e-005 3.8182 0.012 4.6877e-005 0.001157 0.22334 0.00065922 0.224 0.20643 0 0.032782 0.0389 0 1.1274 0.35466 0.10436 0.013625 6.4057 0.085039 0.0001055 0.80507 0.0068063 0.0076153 0.0014104 0.98663 0.9915 3.0444e-006 1.2178e-005 0.14441 0.86999 0.88314 0.0014098 0.96386 0.51574 0.0018988 0.4256 1.7411 1.7397 16.0094 144.9709 0.00021646 -85.5484 0.47295
3.577 0.98806 5.5024e-005 3.8182 0.012 4.689e-005 0.001157 0.22335 0.00065922 0.22401 0.20644 0 0.032782 0.0389 0 1.1275 0.3547 0.10438 0.013627 6.407 0.08505 0.00010551 0.80506 0.006807 0.0076161 0.0014102 0.98663 0.9915 3.044e-006 1.2176e-005 0.14441 0.87034 0.88332 0.0014097 0.96408 0.5159 0.0018987 0.42561 1.742 1.7406 16.0094 144.9709 0.00021618 -85.5493 0.47395
3.578 0.98806 5.5024e-005 3.8182 0.012 4.6903e-005 0.001157 0.22336 0.00065922 0.22402 0.20644 0 0.032781 0.0389 0 1.1276 0.35475 0.1044 0.013628 6.4084 0.08506 0.00010553 0.80505 0.0068077 0.0076169 0.00141 0.98664 0.9915 3.0435e-006 1.2174e-005 0.14442 0.8707 0.88349 0.0014096 0.96429 0.51607 0.0018986 0.42562 1.7428 1.7414 16.0093 144.9709 0.00021591 -85.5501 0.47495
3.579 0.98806 5.5024e-005 3.8182 0.012 4.6916e-005 0.001157 0.22337 0.00065922 0.22403 0.20645 0 0.032781 0.0389 0 1.1277 0.35479 0.10441 0.01363 6.4098 0.085071 0.00010554 0.80503 0.0068085 0.0076176 0.0014098 0.98664 0.99151 3.0431e-006 1.2172e-005 0.14442 0.87105 0.88367 0.0014095 0.9645 0.51624 0.0018984 0.42564 1.7437 1.7423 16.0093 144.9709 0.00021563 -85.5509 0.47595
3.58 0.98806 5.5024e-005 3.8182 0.012 4.6929e-005 0.001157 0.22338 0.00065922 0.22404 0.20646 0 0.03278 0.0389 0 1.1278 0.35484 0.10443 0.013632 6.4112 0.085082 0.00010556 0.80502 0.0068092 0.0076184 0.0014097 0.98664 0.99151 3.0427e-006 1.2171e-005 0.14443 0.8714 0.88384 0.0014094 0.96471 0.51641 0.0018983 0.42565 1.7445 1.7431 16.0093 144.971 0.00021536 -85.5517 0.47695
3.581 0.98806 5.5024e-005 3.8182 0.012 4.6942e-005 0.001157 0.22339 0.00065922 0.22405 0.20647 0 0.03278 0.0389 0 1.1279 0.35489 0.10444 0.013634 6.4126 0.085092 0.00010557 0.80501 0.0068099 0.0076192 0.0014095 0.98664 0.99151 3.0422e-006 1.2169e-005 0.14444 0.87175 0.88402 0.0014093 0.96492 0.51658 0.0018982 0.42566 1.7454 1.744 16.0093 144.971 0.00021509 -85.5525 0.47795
3.582 0.98806 5.5024e-005 3.8182 0.012 4.6956e-005 0.001157 0.2234 0.00065923 0.22406 0.20648 0 0.032779 0.0389 0 1.128 0.35493 0.10446 0.013635 6.414 0.085103 0.00010559 0.805 0.0068106 0.0076199 0.0014093 0.98665 0.99151 3.0418e-006 1.2167e-005 0.14444 0.8721 0.88419 0.0014092 0.96513 0.51674 0.0018981 0.42567 1.7462 1.7449 16.0093 144.971 0.00021482 -85.5533 0.47895
3.583 0.98806 5.5024e-005 3.8182 0.012 4.6969e-005 0.001157 0.22341 0.00065923 0.22406 0.20649 0 0.032779 0.0389 0 1.1281 0.35498 0.10448 0.013637 6.4154 0.085114 0.0001056 0.80499 0.0068113 0.0076207 0.0014091 0.98665 0.99151 3.0414e-006 1.2165e-005 0.14445 0.87245 0.88436 0.0014091 0.96533 0.51691 0.0018979 0.42569 1.7471 1.7457 16.0093 144.971 0.00021455 -85.5541 0.47995
3.584 0.98806 5.5024e-005 3.8182 0.012 4.6982e-005 0.001157 0.22342 0.00065923 0.22407 0.2065 0 0.032778 0.0389 0 1.1282 0.35503 0.10449 0.013639 6.4167 0.085124 0.00010562 0.80498 0.0068121 0.0076215 0.0014089 0.98665 0.99151 3.041e-006 1.2164e-005 0.14445 0.87279 0.88453 0.001409 0.96554 0.51708 0.0018978 0.4257 1.7479 1.7466 16.0093 144.971 0.00021428 -85.5548 0.48095
3.585 0.98806 5.5024e-005 3.8182 0.012 4.6995e-005 0.001157 0.22343 0.00065923 0.22408 0.20651 0 0.032778 0.0389 0 1.1283 0.35507 0.10451 0.01364 6.4181 0.085135 0.00010563 0.80497 0.0068128 0.0076222 0.0014087 0.98665 0.99152 3.0405e-006 1.2162e-005 0.14446 0.87314 0.8847 0.0014089 0.96574 0.51725 0.0018977 0.42571 1.7488 1.7474 16.0093 144.9711 0.00021402 -85.5556 0.48195
3.586 0.98806 5.5023e-005 3.8182 0.012 4.7008e-005 0.001157 0.22344 0.00065923 0.22409 0.20652 0 0.032777 0.0389 0 1.1284 0.35512 0.10453 0.013642 6.4195 0.085146 0.00010564 0.80496 0.0068135 0.007623 0.0014085 0.98666 0.99152 3.0401e-006 1.216e-005 0.14446 0.87348 0.88487 0.0014088 0.96595 0.51741 0.0018976 0.42573 1.7496 1.7482 16.0093 144.9711 0.00021375 -85.5564 0.48295
3.587 0.98806 5.5023e-005 3.8182 0.012 4.7021e-005 0.001157 0.22345 0.00065923 0.2241 0.20652 0 0.032777 0.0389 0 1.1285 0.35516 0.10454 0.013644 6.4209 0.085156 0.00010566 0.80495 0.0068142 0.0076238 0.0014084 0.98666 0.99152 3.0397e-006 1.2159e-005 0.14447 0.87383 0.88504 0.0014087 0.96615 0.51758 0.0018974 0.42574 1.7505 1.7491 16.0092 144.9711 0.00021349 -85.5571 0.48395
3.588 0.98806 5.5023e-005 3.8182 0.012 4.7034e-005 0.001157 0.22346 0.00065923 0.22411 0.20653 0 0.032776 0.0389 0 1.1286 0.35521 0.10456 0.013646 6.4223 0.085167 0.00010567 0.80494 0.0068149 0.0076245 0.0014082 0.98666 0.99152 3.0393e-006 1.2157e-005 0.14448 0.87417 0.88521 0.0014086 0.96635 0.51775 0.0018973 0.42575 1.7513 1.7499 16.0092 144.9711 0.00021322 -85.5579 0.48495
3.589 0.98806 5.5023e-005 3.8182 0.012 4.7047e-005 0.001157 0.22347 0.00065923 0.22412 0.20654 0 0.032776 0.0389 0 1.1287 0.35526 0.10457 0.013647 6.4237 0.085177 0.00010569 0.80493 0.0068156 0.0076253 0.001408 0.98666 0.99152 3.0389e-006 1.2156e-005 0.14448 0.87451 0.88538 0.0014085 0.96655 0.51792 0.0018972 0.42576 1.7521 1.7508 16.0092 144.9711 0.00021296 -85.5587 0.48595
3.59 0.98806 5.5023e-005 3.8182 0.012 4.706e-005 0.001157 0.22347 0.00065923 0.22413 0.20655 0 0.032776 0.0389 0 1.1288 0.3553 0.10459 0.013649 6.4251 0.085188 0.0001057 0.80492 0.0068164 0.0076261 0.0014078 0.98667 0.99152 3.0385e-006 1.2154e-005 0.14449 0.87485 0.88555 0.0014084 0.96674 0.51808 0.0018971 0.42578 1.753 1.7516 16.0092 144.9711 0.0002127 -85.5594 0.48695
3.591 0.98806 5.5023e-005 3.8182 0.012 4.7073e-005 0.001157 0.22348 0.00065923 0.22414 0.20656 0 0.032775 0.0389 0 1.1289 0.35535 0.10461 0.013651 6.4265 0.085199 0.00010572 0.80491 0.0068171 0.0076268 0.0014077 0.98667 0.99152 3.0381e-006 1.2152e-005 0.14449 0.87519 0.88572 0.0014083 0.96694 0.51825 0.0018969 0.42579 1.7538 1.7524 16.0092 144.9712 0.00021244 -85.5602 0.48795
3.592 0.98806 5.5023e-005 3.8182 0.012 4.7086e-005 0.001157 0.22349 0.00065923 0.22415 0.20657 0 0.032775 0.0389 0 1.129 0.3554 0.10462 0.013652 6.4279 0.085209 0.00010573 0.8049 0.0068178 0.0076276 0.0014075 0.98667 0.99153 3.0377e-006 1.2151e-005 0.1445 0.87553 0.88588 0.0014082 0.96714 0.51842 0.0018968 0.4258 1.7546 1.7533 16.0092 144.9712 0.00021218 -85.5609 0.48895
3.593 0.98806 5.5023e-005 3.8182 0.012 4.7099e-005 0.001157 0.2235 0.00065923 0.22416 0.20658 0 0.032774 0.0389 0 1.1291 0.35544 0.10464 0.013654 6.4293 0.08522 0.00010575 0.80489 0.0068185 0.0076284 0.0014073 0.98667 0.99153 3.0373e-006 1.2149e-005 0.14451 0.87587 0.88605 0.0014082 0.96733 0.51859 0.0018967 0.42582 1.7554 1.7541 16.0092 144.9712 0.00021192 -85.5616 0.48995
3.594 0.98806 5.5023e-005 3.8182 0.012 4.7112e-005 0.001157 0.22351 0.00065923 0.22417 0.20659 0 0.032774 0.0389 0 1.1292 0.35549 0.10465 0.013656 6.4306 0.085231 0.00010576 0.80488 0.0068192 0.0076291 0.0014072 0.98667 0.99153 3.0369e-006 1.2148e-005 0.14451 0.8762 0.88621 0.0014081 0.96752 0.51875 0.0018966 0.42583 1.7563 1.7549 16.0092 144.9712 0.00021166 -85.5624 0.49095
3.595 0.98806 5.5023e-005 3.8182 0.012 4.7125e-005 0.001157 0.22352 0.00065923 0.22418 0.20659 0 0.032773 0.0389 0 1.1293 0.35553 0.10467 0.013658 6.432 0.085241 0.00010578 0.80486 0.0068199 0.0076299 0.001407 0.98668 0.99153 3.0365e-006 1.2146e-005 0.14452 0.87654 0.88638 0.001408 0.96771 0.51892 0.0018965 0.42584 1.7571 1.7558 16.0092 144.9712 0.00021141 -85.5631 0.49195
3.596 0.98806 5.5023e-005 3.8182 0.012 4.7138e-005 0.001157 0.22353 0.00065923 0.22419 0.2066 0 0.032773 0.0389 0 1.1294 0.35558 0.10469 0.013659 6.4334 0.085252 0.00010579 0.80485 0.0068207 0.0076307 0.0014068 0.98668 0.99153 3.0362e-006 1.2145e-005 0.14452 0.87687 0.88654 0.0014079 0.9679 0.51909 0.0018964 0.42586 1.7579 1.7566 16.0091 144.9713 0.00021115 -85.5638 0.49295
3.597 0.98806 5.5023e-005 3.8182 0.012 4.7151e-005 0.001157 0.22354 0.00065923 0.22419 0.20661 0 0.032772 0.0389 0 1.1295 0.35563 0.1047 0.013661 6.4348 0.085263 0.00010581 0.80484 0.0068214 0.0076314 0.0014067 0.98668 0.99153 3.0358e-006 1.2143e-005 0.14453 0.87721 0.88671 0.0014078 0.96809 0.51925 0.0018962 0.42587 1.7587 1.7574 16.0091 144.9713 0.0002109 -85.5645 0.49395
3.598 0.98806 5.5023e-005 3.8182 0.012 4.7164e-005 0.001157 0.22355 0.00065923 0.2242 0.20662 0 0.032772 0.0389 0 1.1296 0.35567 0.10472 0.013663 6.4362 0.085273 0.00010582 0.80483 0.0068221 0.0076322 0.0014065 0.98668 0.99153 3.0354e-006 1.2141e-005 0.14453 0.87754 0.88687 0.0014077 0.96828 0.51942 0.0018961 0.42588 1.7595 1.7582 16.0091 144.9713 0.00021064 -85.5652 0.49495
3.599 0.98806 5.5023e-005 3.8182 0.012 4.7177e-005 0.001157 0.22356 0.00065923 0.22421 0.20663 0 0.032771 0.0389 0 1.1297 0.35572 0.10473 0.013664 6.4376 0.085284 0.00010583 0.80482 0.0068228 0.007633 0.0014063 0.98668 0.99154 3.035e-006 1.214e-005 0.14454 0.87787 0.88703 0.0014077 0.96847 0.51959 0.001896 0.42589 1.7604 1.759 16.0091 144.9713 0.00021039 -85.5659 0.49595
3.6 0.98806 5.5022e-005 3.8182 0.012 4.719e-005 0.001157 0.22357 0.00065923 0.22422 0.20664 0 0.032771 0.0389 0 1.1298 0.35577 0.10475 0.013666 6.439 0.085295 0.00010585 0.80481 0.0068235 0.0076337 0.0014062 0.98669 0.99154 3.0346e-006 1.2138e-005 0.14455 0.8782 0.88719 0.0014076 0.96865 0.51975 0.0018959 0.42591 1.7612 1.7599 16.0091 144.9713 0.00021014 -85.5666 0.49695
3.601 0.98806 5.5022e-005 3.8182 0.012 4.7203e-005 0.001157 0.22358 0.00065923 0.22423 0.20665 0 0.03277 0.0389 0 1.1299 0.35581 0.10477 0.013668 6.4404 0.085305 0.00010586 0.8048 0.0068242 0.0076345 0.001406 0.98669 0.99154 3.0343e-006 1.2137e-005 0.14455 0.87853 0.88735 0.0014075 0.96884 0.51992 0.0018958 0.42592 1.762 1.7607 16.0091 144.9714 0.00020989 -85.5673 0.49795
3.602 0.98806 5.5022e-005 3.8182 0.012 4.7216e-005 0.001157 0.22359 0.00065923 0.22424 0.20666 0 0.03277 0.0389 0 1.13 0.35586 0.10478 0.013669 6.4418 0.085316 0.00010588 0.80479 0.006825 0.0076353 0.0014058 0.98669 0.99154 3.0339e-006 1.2135e-005 0.14456 0.87885 0.88751 0.0014074 0.96902 0.52009 0.0018957 0.42593 1.7628 1.7615 16.0091 144.9714 0.00020964 -85.568 0.49895
3.603 0.98806 5.5022e-005 3.8182 0.012 4.7229e-005 0.001157 0.2236 0.00065923 0.22425 0.20666 0 0.032769 0.0389 0 1.1301 0.35591 0.1048 0.013671 6.4432 0.085326 0.00010589 0.80478 0.0068257 0.007636 0.0014057 0.98669 0.99154 3.0335e-006 1.2134e-005 0.14456 0.87918 0.88767 0.0014073 0.9692 0.52025 0.0018956 0.42595 1.7636 1.7623 16.0091 144.9714 0.00020939 -85.5687 0.49995
3.604 0.98806 5.5022e-005 3.8182 0.012 4.7242e-005 0.001157 0.2236 0.00065923 0.22426 0.20667 0 0.032769 0.0389 0 1.1302 0.35595 0.10482 0.013673 6.4446 0.085337 0.00010591 0.80477 0.0068264 0.0076368 0.0014055 0.9867 0.99154 3.0332e-006 1.2133e-005 0.14457 0.87951 0.88783 0.0014072 0.96938 0.52042 0.0018955 0.42596 1.7644 1.7631 16.009 144.9714 0.00020914 -85.5694 0.50095
3.605 0.98806 5.5022e-005 3.8182 0.012 4.7255e-005 0.001157 0.22361 0.00065923 0.22427 0.20668 0 0.032768 0.0389 0 1.1303 0.356 0.10483 0.013675 6.446 0.085348 0.00010592 0.80476 0.0068271 0.0076376 0.0014053 0.9867 0.99154 3.0328e-006 1.2131e-005 0.14457 0.87983 0.88799 0.0014071 0.96956 0.52059 0.0018954 0.42597 1.7652 1.7639 16.009 144.9714 0.0002089 -85.57 0.50195
3.606 0.98806 5.5022e-005 3.8182 0.012 4.7268e-005 0.001157 0.22362 0.00065923 0.22428 0.20669 0 0.032768 0.0389 0 1.1304 0.35604 0.10485 0.013676 6.4474 0.085358 0.00010594 0.80475 0.0068278 0.0076383 0.0014052 0.9867 0.99155 3.0324e-006 1.213e-005 0.14458 0.88016 0.88815 0.001407 0.96974 0.52075 0.0018952 0.42599 1.766 1.7647 16.009 144.9715 0.00020865 -85.5707 0.50295
3.607 0.98806 5.5022e-005 3.8182 0.012 4.7281e-005 0.001157 0.22363 0.00065923 0.22429 0.2067 0 0.032767 0.0389 0 1.1305 0.35609 0.10486 0.013678 6.4488 0.085369 0.00010595 0.80474 0.0068286 0.0076391 0.001405 0.9867 0.99155 3.0321e-006 1.2128e-005 0.14459 0.88048 0.8883 0.001407 0.96992 0.52092 0.0018951 0.426 1.7668 1.7655 16.009 144.9715 0.00020841 -85.5714 0.50395
3.608 0.98806 5.5022e-005 3.8182 0.012 4.7294e-005 0.001157 0.22364 0.00065923 0.2243 0.20671 0 0.032767 0.0389 0 1.1306 0.35614 0.10488 0.01368 6.4502 0.08538 0.00010597 0.80473 0.0068293 0.0076399 0.0014049 0.9867 0.99155 3.0317e-006 1.2127e-005 0.14459 0.8808 0.88846 0.0014069 0.97009 0.52109 0.001895 0.42601 1.7676 1.7663 16.009 144.9715 0.00020816 -85.572 0.50495
3.609 0.98806 5.5022e-005 3.8182 0.012 4.7307e-005 0.001157 0.22365 0.00065923 0.2243 0.20672 0 0.032767 0.0389 0 1.1307 0.35618 0.1049 0.013681 6.4516 0.08539 0.00010598 0.80472 0.00683 0.0076406 0.0014047 0.98671 0.99155 3.0314e-006 1.2125e-005 0.1446 0.88112 0.88861 0.0014068 0.97027 0.52125 0.0018949 0.42602 1.7684 1.7671 16.009 144.9715 0.00020792 -85.5727 0.50595
3.61 0.98806 5.5022e-005 3.8182 0.012 4.732e-005 0.001157 0.22366 0.00065923 0.22431 0.20673 0 0.032766 0.0389 0 1.1308 0.35623 0.10491 0.013683 6.453 0.085401 0.000106 0.80471 0.0068307 0.0076414 0.0014046 0.98671 0.99155 3.031e-006 1.2124e-005 0.1446 0.88144 0.88877 0.0014067 0.97044 0.52142 0.0018948 0.42604 1.7692 1.7679 16.009 144.9715 0.00020768 -85.5734 0.50695
3.611 0.98806 5.5022e-005 3.8182 0.012 4.7333e-005 0.001157 0.22367 0.00065923 0.22432 0.20673 0 0.032766 0.0389 0 1.1309 0.35628 0.10493 0.013685 6.4543 0.085412 0.00010601 0.80469 0.0068314 0.0076422 0.0014044 0.98671 0.99155 3.0307e-006 1.2123e-005 0.14461 0.88176 0.88892 0.0014066 0.97061 0.52159 0.0018947 0.42605 1.77 1.7687 16.009 144.9716 0.00020744 -85.574 0.50795
3.612 0.98806 5.5022e-005 3.8182 0.012 4.7346e-005 0.001157 0.22368 0.00065923 0.22433 0.20674 0 0.032765 0.0389 0 1.131 0.35632 0.10494 0.013687 6.4557 0.085422 0.00010602 0.80468 0.0068321 0.0076429 0.0014043 0.98671 0.99155 3.0303e-006 1.2121e-005 0.14461 0.88208 0.88908 0.0014065 0.97078 0.52175 0.0018946 0.42606 1.7707 1.7695 16.0089 144.9716 0.0002072 -85.5747 0.50895
3.613 0.98806 5.5022e-005 3.8182 0.012 4.7359e-005 0.001157 0.22369 0.00065923 0.22434 0.20675 0 0.032765 0.0389 0 1.1311 0.35637 0.10496 0.013688 6.4571 0.085433 0.00010604 0.80467 0.0068329 0.0076437 0.0014041 0.98671 0.99155 3.03e-006 1.212e-005 0.14462 0.88239 0.88923 0.0014065 0.97095 0.52192 0.0018945 0.42608 1.7715 1.7703 16.0089 144.9716 0.00020696 -85.5753 0.50995
3.614 0.98806 5.5021e-005 3.8182 0.012 4.7372e-005 0.001157 0.2237 0.00065923 0.22435 0.20676 0 0.032764 0.0389 0 1.1312 0.35641 0.10498 0.01369 6.4585 0.085443 0.00010605 0.80466 0.0068336 0.0076445 0.001404 0.98672 0.99156 3.0296e-006 1.2118e-005 0.14463 0.88271 0.88938 0.0014064 0.97112 0.52208 0.0018944 0.42609 1.7723 1.771 16.0089 144.9716 0.00020672 -85.5759 0.51095
3.615 0.98806 5.5021e-005 3.8182 0.012 4.7385e-005 0.001157 0.2237 0.00065923 0.22436 0.20677 0 0.032764 0.0389 0 1.1313 0.35646 0.10499 0.013692 6.4599 0.085454 0.00010607 0.80465 0.0068343 0.0076452 0.0014038 0.98672 0.99156 3.0293e-006 1.2117e-005 0.14463 0.88302 0.88954 0.0014063 0.97129 0.52225 0.0018943 0.4261 1.7731 1.7718 16.0089 144.9716 0.00020648 -85.5766 0.51195
3.616 0.98806 5.5021e-005 3.8182 0.012 4.7398e-005 0.001157 0.22371 0.00065923 0.22437 0.20678 0 0.032763 0.0389 0 1.1314 0.35651 0.10501 0.013693 6.4613 0.085465 0.00010608 0.80464 0.006835 0.007646 0.0014037 0.98672 0.99156 3.029e-006 1.2116e-005 0.14464 0.88334 0.88969 0.0014062 0.97146 0.52242 0.0018942 0.42612 1.7739 1.7726 16.0089 144.9717 0.00020624 -85.5772 0.51295
3.617 0.98806 5.5021e-005 3.8182 0.012 4.7412e-005 0.001157 0.22372 0.00065923 0.22438 0.20679 0 0.032763 0.0389 0 1.1315 0.35655 0.10502 0.013695 6.4627 0.085475 0.0001061 0.80463 0.0068357 0.0076468 0.0014035 0.98672 0.99156 3.0286e-006 1.2114e-005 0.14464 0.88365 0.88984 0.0014062 0.97163 0.52258 0.0018941 0.42613 1.7746 1.7734 16.0089 144.9717 0.00020601 -85.5778 0.51395
3.618 0.98806 5.5021e-005 3.8182 0.012 4.7425e-005 0.001157 0.22373 0.00065923 0.22439 0.20679 0 0.032762 0.0389 0 1.1316 0.3566 0.10504 0.013697 6.4641 0.085486 0.00010611 0.80462 0.0068364 0.0076475 0.0014034 0.98672 0.99156 3.0283e-006 1.2113e-005 0.14465 0.88396 0.88999 0.0014061 0.97179 0.52275 0.001894 0.42614 1.7754 1.7742 16.0089 144.9717 0.00020577 -85.5784 0.51495
3.619 0.98806 5.5021e-005 3.8182 0.012 4.7438e-005 0.001157 0.22374 0.00065923 0.2244 0.2068 0 0.032762 0.0389 0 1.1317 0.35665 0.10506 0.013699 6.4655 0.085497 0.00010613 0.80461 0.0068372 0.0076483 0.0014032 0.98672 0.99156 3.028e-006 1.2112e-005 0.14466 0.88427 0.89014 0.001406 0.97195 0.52291 0.0018939 0.42616 1.7762 1.7749 16.0088 144.9717 0.00020554 -85.579 0.51595
3.62 0.98806 5.5021e-005 3.8182 0.012 4.7451e-005 0.001157 0.22375 0.00065923 0.2244 0.20681 0 0.032761 0.0389 0 1.1318 0.35669 0.10507 0.0137 6.4669 0.085507 0.00010614 0.8046 0.0068379 0.0076491 0.0014031 0.98673 0.99156 3.0276e-006 1.211e-005 0.14466 0.88458 0.89029 0.001406 0.97212 0.52308 0.0018938 0.42617 1.777 1.7757 16.0088 144.9717 0.00020531 -85.5796 0.51695
3.621 0.98806 5.5021e-005 3.8182 0.011999 4.7464e-005 0.001157 0.22376 0.00065923 0.22441 0.20682 0 0.032761 0.0389 0 1.1319 0.35674 0.10509 0.013702 6.4683 0.085518 0.00010616 0.80459 0.0068386 0.0076498 0.001403 0.98673 0.99156 3.0273e-006 1.2109e-005 0.14467 0.88489 0.89044 0.0014059 0.97228 0.52325 0.0018937 0.42618 1.7777 1.7765 16.0088 144.9718 0.00020508 -85.5803 0.51795
3.622 0.98806 5.5021e-005 3.8182 0.011999 4.7477e-005 0.001157 0.22377 0.00065923 0.22442 0.20683 0 0.03276 0.0389 0 1.132 0.35678 0.10511 0.013704 6.4697 0.085528 0.00010617 0.80458 0.0068393 0.0076506 0.0014028 0.98673 0.99157 3.027e-006 1.2108e-005 0.14467 0.8852 0.89058 0.0014058 0.97244 0.52341 0.0018936 0.42619 1.7785 1.7773 16.0088 144.9718 0.00020485 -85.5809 0.51895
3.623 0.98806 5.5021e-005 3.8182 0.011999 4.749e-005 0.001157 0.22378 0.00065923 0.22443 0.20684 0 0.03276 0.0389 0 1.1321 0.35683 0.10512 0.013705 6.4711 0.085539 0.00010618 0.80457 0.00684 0.0076514 0.0014027 0.98673 0.99157 3.0267e-006 1.2107e-005 0.14468 0.88551 0.89073 0.0014057 0.9726 0.52358 0.0018935 0.42621 1.7793 1.778 16.0088 144.9718 0.00020462 -85.5815 0.51995
3.624 0.98806 5.5021e-005 3.8182 0.011999 4.7503e-005 0.0011571 0.22379 0.00065923 0.22444 0.20685 0 0.03276 0.0389 0 1.1322 0.35688 0.10514 0.013707 6.4726 0.08555 0.0001062 0.80456 0.0068407 0.0076521 0.0014025 0.98673 0.99157 3.0264e-006 1.2105e-005 0.14468 0.88581 0.89088 0.0014057 0.97276 0.52374 0.0018934 0.42622 1.78 1.7788 16.0088 144.9718 0.00020439 -85.582 0.52095
3.625 0.98806 5.5021e-005 3.8182 0.011999 4.7516e-005 0.0011571 0.2238 0.00065923 0.22445 0.20685 0 0.032759 0.0389 0 1.1323 0.35692 0.10515 0.013709 6.474 0.08556 0.00010621 0.80455 0.0068415 0.0076529 0.0014024 0.98674 0.99157 3.026e-006 1.2104e-005 0.14469 0.88612 0.89102 0.0014056 0.97292 0.52391 0.0018933 0.42623 1.7808 1.7796 16.0088 144.9718 0.00020416 -85.5826 0.52195
3.626 0.98806 5.5021e-005 3.8182 0.011999 4.7529e-005 0.0011571 0.2238 0.00065923 0.22446 0.20686 0 0.032759 0.0389 0 1.1324 0.35697 0.10517 0.01371 6.4754 0.085571 0.00010623 0.80454 0.0068422 0.0076537 0.0014023 0.98674 0.99157 3.0257e-006 1.2103e-005 0.1447 0.88642 0.89117 0.0014055 0.97307 0.52407 0.0018932 0.42625 1.7815 1.7803 16.0087 144.9719 0.00020393 -85.5832 0.52295
3.627 0.98806 5.5021e-005 3.8182 0.011999 4.7542e-005 0.0011571 0.22381 0.00065923 0.22447 0.20687 0 0.032758 0.0389 0 1.1325 0.35702 0.10519 0.013712 6.4768 0.085581 0.00010624 0.80452 0.0068429 0.0076544 0.0014021 0.98674 0.99157 3.0254e-006 1.2102e-005 0.1447 0.88673 0.89132 0.0014054 0.97323 0.52424 0.0018931 0.42626 1.7823 1.7811 16.0087 144.9719 0.0002037 -85.5838 0.52395
3.628 0.98806 5.5021e-005 3.8182 0.011999 4.7555e-005 0.0011571 0.22382 0.00065923 0.22448 0.20688 0 0.032758 0.0389 0 1.1326 0.35706 0.1052 0.013714 6.4782 0.085592 0.00010626 0.80451 0.0068436 0.0076552 0.001402 0.98674 0.99157 3.0251e-006 1.21e-005 0.14471 0.88703 0.89146 0.0014054 0.97338 0.5244 0.001893 0.42627 1.7831 1.7818 16.0087 144.9719 0.00020348 -85.5844 0.52495
3.629 0.98806 5.502e-005 3.8182 0.011999 4.7568e-005 0.0011571 0.22383 0.00065923 0.22449 0.20689 0 0.032757 0.0389 0 1.1327 0.35711 0.10522 0.013716 6.4796 0.085603 0.00010627 0.8045 0.0068443 0.007656 0.0014019 0.98674 0.99157 3.0248e-006 1.2099e-005 0.14471 0.88733 0.8916 0.0014053 0.97354 0.52457 0.001893 0.42629 1.7838 1.7826 16.0087 144.9719 0.00020325 -85.585 0.52595
3.63 0.98806 5.502e-005 3.8182 0.011999 4.7581e-005 0.0011571 0.22384 0.00065923 0.2245 0.2069 0 0.032757 0.0389 0 1.1328 0.35716 0.10523 0.013717 6.481 0.085613 0.00010629 0.80449 0.006845 0.0076567 0.0014017 0.98674 0.99157 3.0245e-006 1.2098e-005 0.14472 0.88763 0.89175 0.0014052 0.97369 0.52473 0.0018929 0.4263 1.7846 1.7834 16.0087 144.9719 0.00020303 -85.5855 0.52695
3.631 0.98806 5.502e-005 3.8182 0.011999 4.7594e-005 0.0011571 0.22385 0.00065923 0.2245 0.20691 0 0.032756 0.0389 0 1.1329 0.3572 0.10525 0.013719 6.4824 0.085624 0.0001063 0.80448 0.0068457 0.0076575 0.0014016 0.98675 0.99158 3.0242e-006 1.2097e-005 0.14472 0.88793 0.89189 0.0014051 0.97384 0.5249 0.0018928 0.42631 1.7853 1.7841 16.0087 144.972 0.00020281 -85.5861 0.52795
3.632 0.98806 5.502e-005 3.8182 0.011999 4.7607e-005 0.0011571 0.22386 0.00065923 0.22451 0.20691 0 0.032756 0.0389 0 1.133 0.35725 0.10527 0.013721 6.4838 0.085635 0.00010632 0.80447 0.0068465 0.0076583 0.0014015 0.98675 0.99158 3.0239e-006 1.2096e-005 0.14473 0.88823 0.89203 0.0014051 0.97399 0.52506 0.0018927 0.42632 1.7861 1.7849 16.0087 144.972 0.00020258 -85.5867 0.52895
3.633 0.98806 5.502e-005 3.8182 0.011999 4.762e-005 0.0011571 0.22387 0.00065923 0.22452 0.20692 0 0.032755 0.0389 0 1.1331 0.35729 0.10528 0.013722 6.4852 0.085645 0.00010633 0.80446 0.0068472 0.007659 0.0014013 0.98675 0.99158 3.0236e-006 1.2094e-005 0.14474 0.88853 0.89218 0.001405 0.97414 0.52523 0.0018926 0.42634 1.7868 1.7856 16.0086 144.972 0.00020236 -85.5872 0.52995
3.634 0.98806 5.502e-005 3.8182 0.011999 4.7633e-005 0.0011571 0.22388 0.00065923 0.22453 0.20693 0 0.032755 0.0389 0 1.1332 0.35734 0.1053 0.013724 6.4866 0.085656 0.00010635 0.80445 0.0068479 0.0076598 0.0014012 0.98675 0.99158 3.0233e-006 1.2093e-005 0.14474 0.88882 0.89232 0.0014049 0.97429 0.52539 0.0018925 0.42635 1.7875 1.7864 16.0086 144.972 0.00020214 -85.5878 0.53095
3.635 0.98806 5.502e-005 3.8182 0.011999 4.7646e-005 0.0011571 0.22389 0.00065923 0.22454 0.20694 0 0.032754 0.0389 0 1.1333 0.35739 0.10531 0.013726 6.488 0.085666 0.00010636 0.80444 0.0068486 0.0076606 0.0014011 0.98675 0.99158 3.023e-006 1.2092e-005 0.14475 0.88912 0.89246 0.0014049 0.97444 0.52556 0.0018924 0.42636 1.7883 1.7871 16.0086 144.972 0.00020192 -85.5883 0.53195
3.636 0.98806 5.502e-005 3.8182 0.011999 4.7659e-005 0.0011571 0.22389 0.00065923 0.22455 0.20695 0 0.032754 0.0389 0 1.1334 0.35743 0.10533 0.013728 6.4894 0.085677 0.00010637 0.80443 0.0068493 0.0076613 0.0014009 0.98675 0.99158 3.0227e-006 1.2091e-005 0.14475 0.88941 0.8926 0.0014048 0.97459 0.52572 0.0018923 0.42638 1.789 1.7878 16.0086 144.9721 0.0002017 -85.5889 0.53295
3.637 0.98806 5.502e-005 3.8182 0.011999 4.7672e-005 0.0011571 0.2239 0.00065923 0.22456 0.20696 0 0.032754 0.0389 0 1.1335 0.35748 0.10535 0.013729 6.4908 0.085688 0.00010639 0.80442 0.00685 0.0076621 0.0014008 0.98676 0.99158 3.0224e-006 1.209e-005 0.14476 0.88971 0.89274 0.0014047 0.97473 0.52589 0.0018922 0.42639 1.7898 1.7886 16.0086 144.9721 0.00020149 -85.5894 0.53395
3.638 0.98806 5.502e-005 3.8182 0.011999 4.7685e-005 0.0011571 0.22391 0.00065923 0.22457 0.20697 0 0.032753 0.0389 0 1.1336 0.35753 0.10536 0.013731 6.4922 0.085698 0.0001064 0.80441 0.0068508 0.0076629 0.0014007 0.98676 0.99158 3.0221e-006 1.2088e-005 0.14477 0.89 0.89288 0.0014047 0.97488 0.52605 0.0018922 0.4264 1.7905 1.7893 16.0086 144.9721 0.00020127 -85.5899 0.53495
3.639 0.98806 5.502e-005 3.8182 0.011999 4.7698e-005 0.0011571 0.22392 0.00065923 0.22458 0.20697 0 0.032753 0.0389 0 1.1337 0.35757 0.10538 0.013733 6.4936 0.085709 0.00010642 0.8044 0.0068515 0.0076636 0.0014006 0.98676 0.99158 3.0218e-006 1.2087e-005 0.14477 0.89029 0.89302 0.0014046 0.97502 0.52622 0.0018921 0.42642 1.7912 1.7901 16.0085 144.9721 0.00020105 -85.5905 0.53595
3.64 0.98806 5.502e-005 3.8182 0.011999 4.7711e-005 0.0011571 0.22393 0.00065923 0.22458 0.20698 0 0.032752 0.0389 0 1.1338 0.35762 0.1054 0.013734 6.495 0.085719 0.00010643 0.80439 0.0068522 0.0076644 0.0014004 0.98676 0.99159 3.0216e-006 1.2086e-005 0.14478 0.89058 0.89315 0.0014045 0.97517 0.52638 0.001892 0.42643 1.792 1.7908 16.0085 144.9721 0.00020084 -85.591 0.53695
3.641 0.98806 5.502e-005 3.8182 0.011999 4.7724e-005 0.0011571 0.22394 0.00065923 0.22459 0.20699 0 0.032752 0.0389 0 1.1339 0.35766 0.10541 0.013736 6.4965 0.08573 0.00010645 0.80438 0.0068529 0.0076652 0.0014003 0.98676 0.99159 3.0213e-006 1.2085e-005 0.14478 0.89087 0.89329 0.0014045 0.97531 0.52655 0.0018919 0.42644 1.7927 1.7915 16.0085 144.9722 0.00020062 -85.5915 0.53795
3.642 0.98806 5.502e-005 3.8182 0.011999 4.7737e-005 0.0011571 0.22395 0.00065923 0.2246 0.207 0 0.032751 0.0389 0 1.134 0.35771 0.10543 0.013738 6.4979 0.085741 0.00010646 0.80437 0.0068536 0.0076659 0.0014002 0.98676 0.99159 3.021e-006 1.2084e-005 0.14479 0.89116 0.89343 0.0014044 0.97545 0.52671 0.0018918 0.42645 1.7934 1.7923 16.0085 144.9722 0.00020041 -85.5921 0.53895
3.643 0.98806 5.5019e-005 3.8182 0.011999 4.775e-005 0.0011571 0.22396 0.00065923 0.22461 0.20701 0 0.032751 0.0389 0 1.1341 0.35776 0.10544 0.013739 6.4993 0.085751 0.00010648 0.80436 0.0068543 0.0076667 0.0014001 0.98677 0.99159 3.0207e-006 1.2083e-005 0.14479 0.89145 0.89357 0.0014044 0.97559 0.52688 0.0018917 0.42647 1.7942 1.793 16.0085 144.9722 0.00020019 -85.5926 0.53995
3.644 0.98806 5.5019e-005 3.8182 0.011999 4.7763e-005 0.0011571 0.22397 0.00065923 0.22462 0.20702 0 0.03275 0.0389 0 1.1342 0.3578 0.10546 0.013741 6.5007 0.085762 0.00010649 0.80434 0.0068551 0.0076675 0.0013999 0.98677 0.99159 3.0204e-006 1.2082e-005 0.1448 0.89174 0.8937 0.0014043 0.97573 0.52704 0.0018916 0.42648 1.7949 1.7937 16.0085 144.9722 0.00019998 -85.5931 0.54095
3.645 0.98806 5.5019e-005 3.8182 0.011999 4.7776e-005 0.0011571 0.22397 0.00065923 0.22463 0.20702 0 0.03275 0.0389 0 1.1343 0.35785 0.10548 0.013743 6.5021 0.085772 0.00010651 0.80433 0.0068558 0.0076682 0.0013998 0.98677 0.99159 3.0202e-006 1.2081e-005 0.14481 0.89202 0.89384 0.0014042 0.97587 0.52721 0.0018916 0.42649 1.7956 1.7945 16.0084 144.9722 0.00019977 -85.5936 0.54195
3.646 0.98806 5.5019e-005 3.8182 0.011999 4.7789e-005 0.0011571 0.22398 0.00065923 0.22464 0.20703 0 0.032749 0.0389 0 1.1344 0.3579 0.10549 0.013745 6.5035 0.085783 0.00010652 0.80432 0.0068565 0.007669 0.0013997 0.98677 0.99159 3.0199e-006 1.2079e-005 0.14481 0.89231 0.89397 0.0014042 0.97601 0.52737 0.0018915 0.42651 1.7963 1.7952 16.0084 144.9723 0.00019956 -85.5941 0.54295
3.647 0.98806 5.5019e-005 3.8182 0.011999 4.7802e-005 0.0011571 0.22399 0.00065923 0.22465 0.20704 0 0.032749 0.0389 0 1.1345 0.35794 0.10551 0.013746 6.5049 0.085794 0.00010653 0.80431 0.0068572 0.0076698 0.0013996 0.98677 0.99159 3.0196e-006 1.2078e-005 0.14482 0.8926 0.89411 0.0014041 0.97614 0.52753 0.0018914 0.42652 1.797 1.7959 16.0084 144.9723 0.00019935 -85.5946 0.54395
3.648 0.98806 5.5019e-005 3.8182 0.011999 4.7815e-005 0.0011571 0.224 0.00065923 0.22466 0.20705 0 0.032749 0.0389 0 1.1346 0.35799 0.10552 0.013748 6.5063 0.085804 0.00010655 0.8043 0.0068579 0.0076705 0.0013995 0.98677 0.99159 3.0194e-006 1.2077e-005 0.14482 0.89288 0.89424 0.001404 0.97628 0.5277 0.0018913 0.42653 1.7978 1.7966 16.0084 144.9723 0.00019914 -85.5951 0.54495
3.649 0.98806 5.5019e-005 3.8182 0.011999 4.7828e-005 0.0011571 0.22401 0.00065923 0.22466 0.20706 0 0.032748 0.0389 0 1.1347 0.35804 0.10554 0.01375 6.5077 0.085815 0.00010656 0.80429 0.0068586 0.0076713 0.0013994 0.98677 0.99159 3.0191e-006 1.2076e-005 0.14483 0.89316 0.89437 0.001404 0.97641 0.52786 0.0018912 0.42655 1.7985 1.7973 16.0084 144.9723 0.00019893 -85.5956 0.54595
3.65 0.98806 5.5019e-005 3.8182 0.011999 4.7841e-005 0.0011571 0.22402 0.00065923 0.22467 0.20707 0 0.032748 0.0389 0 1.1348 0.35808 0.10556 0.013751 6.5092 0.085825 0.00010658 0.80428 0.0068594 0.0076721 0.0013992 0.98678 0.9916 3.0188e-006 1.2075e-005 0.14483 0.89344 0.89451 0.0014039 0.97655 0.52803 0.0018912 0.42656 1.7992 1.7981 16.0084 144.9723 0.00019873 -85.5961 0.54695
3.651 0.98806 5.5019e-005 3.8182 0.011999 4.7854e-005 0.0011571 0.22403 0.00065923 0.22468 0.20707 0 0.032747 0.0389 0 1.1349 0.35813 0.10557 0.013753 6.5106 0.085836 0.00010659 0.80427 0.0068601 0.0076728 0.0013991 0.98678 0.9916 3.0186e-006 1.2074e-005 0.14484 0.89373 0.89464 0.0014038 0.97668 0.52819 0.0018911 0.42657 1.7999 1.7988 16.0084 144.9724 0.00019852 -85.5966 0.54795
3.652 0.98806 5.5019e-005 3.8182 0.011999 4.7867e-005 0.0011571 0.22404 0.00065923 0.22469 0.20708 0 0.032747 0.0389 0 1.135 0.35817 0.10559 0.013755 6.512 0.085847 0.00010661 0.80426 0.0068608 0.0076736 0.001399 0.98678 0.9916 3.0183e-006 1.2073e-005 0.14485 0.89401 0.89477 0.0014038 0.97682 0.52836 0.001891 0.42659 1.8006 1.7995 16.0083 144.9724 0.00019831 -85.5971 0.54895
3.653 0.98806 5.5019e-005 3.8182 0.011999 4.788e-005 0.0011571 0.22405 0.00065923 0.2247 0.20709 0 0.032746 0.0389 0 1.1351 0.35822 0.1056 0.013756 6.5134 0.085857 0.00010662 0.80425 0.0068615 0.0076744 0.0013989 0.98678 0.9916 3.018e-006 1.2072e-005 0.14485 0.89429 0.8949 0.0014037 0.97695 0.52852 0.0018909 0.4266 1.8013 1.8002 16.0083 144.9724 0.00019811 -85.5976 0.54995
3.654 0.98806 5.5019e-005 3.8182 0.011999 4.7894e-005 0.0011571 0.22405 0.00065923 0.22471 0.2071 0 0.032746 0.0389 0 1.1352 0.35827 0.10562 0.013758 6.5148 0.085868 0.00010664 0.80424 0.0068622 0.0076751 0.0013988 0.98678 0.9916 3.0178e-006 1.2071e-005 0.14486 0.89456 0.89503 0.0014037 0.97708 0.52868 0.0018908 0.42661 1.802 1.8009 16.0083 144.9724 0.0001979 -85.5981 0.55095
3.655 0.98806 5.5019e-005 3.8182 0.011999 4.7907e-005 0.0011571 0.22406 0.00065923 0.22472 0.20711 0 0.032745 0.0389 0 1.1353 0.35831 0.10564 0.01376 6.5162 0.085878 0.00010665 0.80423 0.0068629 0.0076759 0.0013987 0.98678 0.9916 3.0175e-006 1.207e-005 0.14486 0.89484 0.89516 0.0014036 0.97721 0.52885 0.0018908 0.42662 1.8027 1.8016 16.0083 144.9724 0.0001977 -85.5986 0.55195
3.656 0.98806 5.5019e-005 3.8182 0.011999 4.792e-005 0.0011571 0.22407 0.00065923 0.22473 0.20712 0 0.032745 0.0389 0 1.1354 0.35836 0.10565 0.013762 6.5176 0.085889 0.00010667 0.80422 0.0068636 0.0076767 0.0013986 0.98679 0.9916 3.0173e-006 1.2069e-005 0.14487 0.89512 0.89529 0.0014035 0.97734 0.52901 0.0018907 0.42664 1.8034 1.8023 16.0083 144.9725 0.0001975 -85.5991 0.55295
3.657 0.98806 5.5018e-005 3.8182 0.011999 4.7933e-005 0.0011571 0.22408 0.00065923 0.22473 0.20712 0 0.032745 0.0389 0 1.1355 0.35841 0.10567 0.013763 6.519 0.0859 0.00010668 0.80421 0.0068644 0.0076774 0.0013985 0.98679 0.9916 3.017e-006 1.2068e-005 0.14487 0.8954 0.89542 0.0014035 0.97747 0.52917 0.0018906 0.42665 1.8041 1.803 16.0082 144.9725 0.00019729 -85.5995 0.55395
3.658 0.98806 5.5018e-005 3.8182 0.011999 4.7946e-005 0.0011571 0.22409 0.00065923 0.22474 0.20713 0 0.032744 0.0389 0 1.1356 0.35845 0.10569 0.013765 6.5205 0.08591 0.00010669 0.8042 0.0068651 0.0076782 0.0013983 0.98679 0.9916 3.0168e-006 1.2067e-005 0.14488 0.89567 0.89555 0.0014034 0.97759 0.52934 0.0018905 0.42666 1.8048 1.8037 16.0082 144.9725 0.00019709 -85.6 0.55495
3.659 0.98806 5.5018e-005 3.8182 0.011999 4.7959e-005 0.0011571 0.2241 0.00065923 0.22475 0.20714 0 0.032744 0.0389 0 1.1357 0.3585 0.1057 0.013767 6.5219 0.085921 0.00010671 0.80419 0.0068658 0.007679 0.0013982 0.98679 0.9916 3.0165e-006 1.2066e-005 0.14489 0.89595 0.89568 0.0014034 0.97772 0.5295 0.0018905 0.42668 1.8055 1.8044 16.0082 144.9725 0.00019689 -85.6005 0.55595
3.66 0.98806 5.5018e-005 3.8182 0.011999 4.7972e-005 0.0011571 0.22411 0.00065923 0.22476 0.20715 0 0.032743 0.0389 0 1.1357 0.35855 0.10572 0.013768 6.5233 0.085931 0.00010672 0.80418 0.0068665 0.0076797 0.0013981 0.98679 0.99161 3.0163e-006 1.2065e-005 0.14489 0.89622 0.89581 0.0014033 0.97785 0.52967 0.0018904 0.42669 1.8062 1.8051 16.0082 144.9725 0.00019669 -85.6009 0.55695
3.661 0.98806 5.5018e-005 3.8182 0.011999 4.7985e-005 0.0011571 0.22412 0.00065923 0.22477 0.20716 0 0.032743 0.0389 0 1.1358 0.35859 0.10573 0.01377 6.5247 0.085942 0.00010674 0.80416 0.0068672 0.0076805 0.001398 0.98679 0.99161 3.016e-006 1.2064e-005 0.1449 0.89649 0.89594 0.0014033 0.97797 0.52983 0.0018903 0.4267 1.8069 1.8058 16.0082 144.9726 0.00019649 -85.6014 0.55795
3.662 0.98806 5.5018e-005 3.8182 0.011999 4.7998e-005 0.0011571 0.22412 0.00065923 0.22478 0.20717 0 0.032742 0.0389 0 1.1359 0.35864 0.10575 0.013772 6.5261 0.085953 0.00010675 0.80415 0.0068679 0.0076813 0.0013979 0.98679 0.99161 3.0158e-006 1.2063e-005 0.1449 0.89676 0.89606 0.0014032 0.9781 0.52999 0.0018902 0.42672 1.8076 1.8065 16.0082 144.9726 0.0001963 -85.6018 0.55895
3.663 0.98806 5.5018e-005 3.8182 0.011999 4.8011e-005 0.0011571 0.22413 0.00065923 0.22479 0.20717 0 0.032742 0.0389 0 1.136 0.35868 0.10577 0.013773 6.5275 0.085963 0.00010677 0.80414 0.0068686 0.007682 0.0013978 0.98679 0.99161 3.0155e-006 1.2062e-005 0.14491 0.89703 0.89619 0.0014032 0.97822 0.53016 0.0018902 0.42673 1.8083 1.8072 16.0081 144.9726 0.0001961 -85.6023 0.55995
3.664 0.98806 5.5018e-005 3.8182 0.011999 4.8024e-005 0.0011571 0.22414 0.00065923 0.2248 0.20718 0 0.032741 0.0389 0 1.1361 0.35873 0.10578 0.013775 6.529 0.085974 0.00010678 0.80413 0.0068694 0.0076828 0.0013977 0.9868 0.99161 3.0153e-006 1.2061e-005 0.14492 0.8973 0.89632 0.0014031 0.97834 0.53032 0.0018901 0.42674 1.809 1.8079 16.0081 144.9726 0.0001959 -85.6028 0.56095
3.665 0.98806 5.5018e-005 3.8182 0.011999 4.8037e-005 0.0011571 0.22415 0.00065923 0.2248 0.20719 0 0.032741 0.0389 0 1.1362 0.35878 0.1058 0.013777 6.5304 0.085984 0.0001068 0.80412 0.0068701 0.0076836 0.0013976 0.9868 0.99161 3.015e-006 1.206e-005 0.14492 0.89757 0.89644 0.0014031 0.97846 0.53048 0.00189 0.42675 1.8097 1.8086 16.0081 144.9726 0.00019571 -85.6032 0.56195
3.666 0.98806 5.5018e-005 3.8182 0.011999 4.805e-005 0.0011571 0.22416 0.00065923 0.22481 0.2072 0 0.03274 0.0389 0 1.1363 0.35882 0.10581 0.013779 6.5318 0.085995 0.00010681 0.80411 0.0068708 0.0076843 0.0013975 0.9868 0.99161 3.0148e-006 1.2059e-005 0.14493 0.89784 0.89657 0.001403 0.97859 0.53065 0.00189 0.42677 1.8104 1.8093 16.0081 144.9727 0.00019551 -85.6037 0.56295
3.667 0.98806 5.5018e-005 3.8182 0.011999 4.8063e-005 0.0011571 0.22417 0.00065923 0.22482 0.20721 0 0.03274 0.0389 0 1.1364 0.35887 0.10583 0.01378 6.5332 0.086005 0.00010683 0.8041 0.0068715 0.0076851 0.0013974 0.9868 0.99161 3.0146e-006 1.2058e-005 0.14493 0.89811 0.89669 0.001403 0.97871 0.53081 0.0018899 0.42678 1.8111 1.81 16.0081 144.9727 0.00019532 -85.6041 0.56395
3.668 0.98806 5.5018e-005 3.8182 0.011999 4.8076e-005 0.0011571 0.22418 0.00065923 0.22483 0.20722 0 0.03274 0.0389 0 1.1365 0.35892 0.10585 0.013782 6.5346 0.086016 0.00010684 0.80409 0.0068722 0.0076858 0.0013973 0.9868 0.99161 3.0143e-006 1.2057e-005 0.14494 0.89838 0.89682 0.0014029 0.97883 0.53097 0.0018898 0.42679 1.8118 1.8107 16.0081 144.9727 0.00019512 -85.6045 0.56495
3.669 0.98806 5.5018e-005 3.8182 0.011999 4.8089e-005 0.0011571 0.22419 0.00065923 0.22484 0.20722 0 0.032739 0.0389 0 1.1366 0.35896 0.10586 0.013784 6.5361 0.086027 0.00010685 0.80408 0.0068729 0.0076866 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.14494 0.89864 0.89694 0.0014028 0.97894 0.53114 0.0018897 0.42681 1.8124 1.8114 16.008 144.9727 0.00019493 -85.605 0.56595
3.67 0.98806 5.5018e-005 3.8182 0.011999 4.8102e-005 0.0011571 0.22419 0.00065923 0.22485 0.20723 0 0.032739 0.0389 0 1.1367 0.35901 0.10588 0.013785 6.5375 0.086037 0.00010687 0.80407 0.0068737 0.0076874 0.0013971 0.9868 0.99161 3.0139e-006 1.2055e-005 0.14495 0.89891 0.89706 0.0014028 0.97906 0.5313 0.0018897 0.42682 1.8131 1.812 16.008 144.9727 0.00019474 -85.6054 0.56695
3.671 0.98806 5.5017e-005 3.8182 0.011999 4.8115e-005 0.0011571 0.2242 0.00065923 0.22486 0.20724 0 0.032738 0.0389 0 1.1368 0.35905 0.10589 0.013787 6.5389 0.086048 0.00010688 0.80406 0.0068744 0.0076881 0.001397 0.98681 0.99161 3.0136e-006 1.2054e-005 0.14496 0.89917 0.89719 0.0014027 0.97918 0.53146 0.0018896 0.42683 1.8138 1.8127 16.008 144.9728 0.00019454 -85.6058 0.56795
3.672 0.98806 5.5017e-005 3.8182 0.011999 4.8128e-005 0.0011571 0.22421 0.00065923 0.22487 0.20725 0 0.032738 0.0389 0 1.1369 0.3591 0.10591 0.013789 6.5403 0.086058 0.0001069 0.80405 0.0068751 0.0076889 0.0013969 0.98681 0.99162 3.0134e-006 1.2054e-005 0.14496 0.89944 0.89731 0.0014027 0.9793 0.53162 0.0018895 0.42685 1.8145 1.8134 16.008 144.9728 0.00019435 -85.6063 0.56895
3.673 0.98806 5.5017e-005 3.8182 0.011999 4.8141e-005 0.0011572 0.22422 0.00065923 0.22487 0.20726 0 0.032737 0.0389 0 1.137 0.35915 0.10593 0.01379 6.5417 0.086069 0.00010691 0.80404 0.0068758 0.0076897 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.14497 0.8997 0.89743 0.0014026 0.97941 0.53179 0.0018895 0.42686 1.8151 1.8141 16.008 144.9728 0.00019416 -85.6067 0.56995
3.674 0.98806 5.5017e-005 3.8182 0.011999 4.8154e-005 0.0011572 0.22423 0.00065923 0.22488 0.20727 0 0.032737 0.0389 0 1.1371 0.35919 0.10594 0.013792 6.5432 0.08608 0.00010693 0.80403 0.0068765 0.0076904 0.0013967 0.98681 0.99162 3.013e-006 1.2052e-005 0.14497 0.89996 0.89755 0.0014026 0.97953 0.53195 0.0018894 0.42687 1.8158 1.8148 16.0079 144.9728 0.00019397 -85.6071 0.57095
3.675 0.98806 5.5017e-005 3.8182 0.011999 4.8167e-005 0.0011572 0.22424 0.00065923 0.22489 0.20727 0 0.032736 0.0389 0 1.1372 0.35924 0.10596 0.013794 6.5446 0.08609 0.00010694 0.80402 0.0068772 0.0076912 0.0013966 0.98681 0.99162 3.0127e-006 1.2051e-005 0.14498 0.90022 0.89767 0.0014025 0.97964 0.53211 0.0018893 0.42688 1.8165 1.8154 16.0079 144.9728 0.00019378 -85.6075 0.57195
3.676 0.98806 5.5017e-005 3.8182 0.011999 4.818e-005 0.0011572 0.22425 0.00065923 0.2249 0.20728 0 0.032736 0.0389 0 1.1373 0.35929 0.10598 0.013796 6.546 0.086101 0.00010696 0.80401 0.0068779 0.007692 0.0013965 0.98681 0.99162 3.0125e-006 1.205e-005 0.14498 0.90048 0.89779 0.0014025 0.97976 0.53228 0.0018893 0.4269 1.8172 1.8161 16.0079 144.9729 0.0001936 -85.608 0.57295
3.677 0.98806 5.5017e-005 3.8182 0.011999 4.8193e-005 0.0011572 0.22425 0.00065923 0.22491 0.20729 0 0.032736 0.0389 0 1.1374 0.35933 0.10599 0.013797 6.5474 0.086111 0.00010697 0.804 0.0068787 0.0076927 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.14499 0.90074 0.89791 0.0014024 0.97987 0.53244 0.0018892 0.42691 1.8178 1.8168 16.0079 144.9729 0.00019341 -85.6084 0.57395
3.678 0.98806 5.5017e-005 3.8182 0.011999 4.8206e-005 0.0011572 0.22426 0.00065923 0.22492 0.2073 0 0.032735 0.0389 0 1.1375 0.35938 0.10601 0.013799 6.5489 0.086122 0.00010699 0.80399 0.0068794 0.0076935 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.145 0.901 0.89803 0.0014023 0.97998 0.5326 0.0018891 0.42692 1.8185 1.8174 16.0079 144.9729 0.00019322 -85.6088 0.57495
3.679 0.98806 5.5017e-005 3.8182 0.011999 4.8219e-005 0.0011572 0.22427 0.00065923 0.22493 0.20731 0 0.032735 0.0389 0 1.1376 0.35943 0.10602 0.013801 6.5503 0.086132 0.000107 0.80397 0.0068801 0.0076943 0.0013962 0.98682 0.99162 3.0119e-006 1.2047e-005 0.145 0.90126 0.89815 0.0014023 0.98009 0.53276 0.0018891 0.42694 1.8192 1.8181 16.0079 144.9729 0.00019304 -85.6092 0.57595
3.68 0.98806 5.5017e-005 3.8182 0.011999 4.8232e-005 0.0011572 0.22428 0.00065923 0.22494 0.20731 0 0.032734 0.0389 0 1.1377 0.35947 0.10604 0.013802 6.5517 0.086143 0.00010701 0.80396 0.0068808 0.007695 0.0013961 0.98682 0.99162 3.0116e-006 1.2046e-005 0.14501 0.90151 0.89827 0.0014023 0.9802 0.53293 0.001889 0.42695 1.8198 1.8188 16.0078 144.9729 0.00019285 -85.6096 0.57695
3.681 0.98806 5.5017e-005 3.8182 0.011999 4.8245e-005 0.0011572 0.22429 0.00065923 0.22494 0.20732 0 0.032734 0.0389 0 1.1378 0.35952 0.10606 0.013804 6.5531 0.086154 0.00010703 0.80395 0.0068815 0.0076958 0.001396 0.98682 0.99162 3.0114e-006 1.2046e-005 0.14501 0.90177 0.89839 0.0014022 0.98031 0.53309 0.0018889 0.42696 1.8205 1.8194 16.0078 144.973 0.00019267 -85.61 0.57795
3.682 0.98806 5.5017e-005 3.8182 0.011999 4.8258e-005 0.0011572 0.2243 0.00065923 0.22495 0.20733 0 0.032733 0.0389 0 1.1379 0.35956 0.10607 0.013806 6.5545 0.086164 0.00010704 0.80394 0.0068822 0.0076966 0.0013959 0.98682 0.99162 3.0112e-006 1.2045e-005 0.14502 0.90203 0.89851 0.0014022 0.98042 0.53325 0.0018889 0.42698 1.8212 1.8201 16.0078 144.973 0.00019248 -85.6104 0.57895
3.683 0.98806 5.5017e-005 3.8182 0.011999 4.8271e-005 0.0011572 0.22431 0.00065923 0.22496 0.20734 0 0.032733 0.0389 0 1.138 0.35961 0.10609 0.013807 6.556 0.086175 0.00010706 0.80393 0.0068829 0.0076973 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.14502 0.90228 0.89863 0.0014021 0.98053 0.53341 0.0018888 0.42699 1.8218 1.8208 16.0078 144.973 0.0001923 -85.6108 0.57995
3.684 0.98806 5.5017e-005 3.8182 0.011999 4.8284e-005 0.0011572 0.22431 0.00065923 0.22497 0.20735 0 0.032733 0.0389 0 1.1381 0.35966 0.1061 0.013809 6.5574 0.086185 0.00010707 0.80392 0.0068837 0.0076981 0.0013957 0.98682 0.99163 3.0108e-006 1.2043e-005 0.14503 0.90253 0.89874 0.0014021 0.98064 0.53358 0.0018887 0.427 1.8225 1.8214 16.0078 144.973 0.00019212 -85.6112 0.58095
3.685 0.98806 5.5017e-005 3.8182 0.011999 4.8297e-005 0.0011572 0.22432 0.00065923 0.22498 0.20736 0 0.032732 0.0389 0 1.1382 0.3597 0.10612 0.013811 6.5588 0.086196 0.00010709 0.80391 0.0068844 0.0076989 0.0013956 0.98682 0.99163 3.0106e-006 1.2042e-005 0.14504 0.90279 0.89886 0.001402 0.98075 0.53374 0.0018887 0.42701 1.8231 1.8221 16.0077 144.973 0.00019193 -85.6116 0.58195
3.686 0.98806 5.5016e-005 3.8182 0.011999 4.831e-005 0.0011572 0.22433 0.00065923 0.22499 0.20736 0 0.032732 0.0389 0 1.1383 0.35975 0.10614 0.013813 6.5603 0.086206 0.0001071 0.8039 0.0068851 0.0076996 0.0013955 0.98682 0.99163 3.0104e-006 1.2041e-005 0.14504 0.90304 0.89898 0.001402 0.98085 0.5339 0.0018886 0.42703 1.8238 1.8228 16.0077 144.9731 0.00019175 -85.612 0.58295
3.687 0.98806 5.5016e-005 3.8182 0.011998 4.8323e-005 0.0011572 0.22434 0.00065923 0.225 0.20737 0 0.032731 0.0389 0 1.1384 0.3598 0.10615 0.013814 6.5617 0.086217 0.00010712 0.80389 0.0068858 0.0077004 0.0013955 0.98683 0.99163 3.0102e-006 1.2041e-005 0.14505 0.90329 0.89909 0.0014019 0.98096 0.53406 0.0018886 0.42704 1.8244 1.8234 16.0077 144.9731 0.00019157 -85.6124 0.58395
3.688 0.98806 5.5016e-005 3.8182 0.011998 4.8336e-005 0.0011572 0.22435 0.00065923 0.225 0.20738 0 0.032731 0.0389 0 1.1385 0.35984 0.10617 0.013816 6.5631 0.086228 0.00010713 0.80388 0.0068865 0.0077011 0.0013954 0.98683 0.99163 3.01e-006 1.204e-005 0.14505 0.90354 0.89921 0.0014019 0.98106 0.53422 0.0018885 0.42705 1.8251 1.8241 16.0077 144.9731 0.00019139 -85.6127 0.58495
3.689 0.98806 5.5016e-005 3.8182 0.011998 4.8349e-005 0.0011572 0.22436 0.00065923 0.22501 0.20739 0 0.03273 0.0389 0 1.1386 0.35989 0.10618 0.013818 6.5645 0.086238 0.00010715 0.80387 0.0068872 0.0077019 0.0013953 0.98683 0.99163 3.0098e-006 1.2039e-005 0.14506 0.90379 0.89932 0.0014019 0.98117 0.53439 0.0018884 0.42707 1.8257 1.8247 16.0077 144.9731 0.00019121 -85.6131 0.58595
3.69 0.98806 5.5016e-005 3.8182 0.011998 4.8362e-005 0.0011572 0.22437 0.00065923 0.22502 0.2074 0 0.03273 0.0389 0 1.1387 0.35994 0.1062 0.013819 6.566 0.086249 0.00010716 0.80386 0.0068879 0.0077027 0.0013952 0.98683 0.99163 3.0096e-006 1.2038e-005 0.14506 0.90404 0.89944 0.0014018 0.98127 0.53455 0.0018884 0.42708 1.8264 1.8254 16.0076 144.9731 0.00019103 -85.6135 0.58695
3.691 0.98806 5.5016e-005 3.8182 0.011998 4.8375e-005 0.0011572 0.22437 0.00065923 0.22503 0.2074 0 0.032729 0.0389 0 1.1388 0.35998 0.10622 0.013821 6.5674 0.086259 0.00010717 0.80385 0.0068887 0.0077034 0.0013951 0.98683 0.99163 3.0094e-006 1.2037e-005 0.14507 0.90429 0.89955 0.0014018 0.98137 0.53471 0.0018883 0.42709 1.827 1.826 16.0076 144.9732 0.00019086 -85.6139 0.58795
3.692 0.98806 5.5016e-005 3.8182 0.011998 4.8388e-005 0.0011572 0.22438 0.00065923 0.22504 0.20741 0 0.032729 0.0389 0 1.1389 0.36003 0.10623 0.013823 6.5688 0.08627 0.00010719 0.80384 0.0068894 0.0077042 0.001395 0.98683 0.99163 3.0092e-006 1.2037e-005 0.14508 0.90454 0.89966 0.0014017 0.98148 0.53487 0.0018883 0.42711 1.8277 1.8267 16.0076 144.9732 0.00019068 -85.6142 0.58895
3.693 0.98806 5.5016e-005 3.8182 0.011998 4.8401e-005 0.0011572 0.22439 0.00065923 0.22505 0.20742 0 0.032729 0.0389 0 1.139 0.36007 0.10625 0.013824 6.5702 0.08628 0.0001072 0.80383 0.0068901 0.007705 0.0013949 0.98683 0.99163 3.009e-006 1.2036e-005 0.14508 0.90478 0.89978 0.0014017 0.98158 0.53503 0.0018882 0.42712 1.8283 1.8273 16.0076 144.9732 0.0001905 -85.6146 0.58995
3.694 0.98806 5.5016e-005 3.8182 0.011998 4.8415e-005 0.0011572 0.2244 0.00065923 0.22506 0.20743 0 0.032728 0.0389 0 1.1391 0.36012 0.10627 0.013826 6.5717 0.086291 0.00010722 0.80382 0.0068908 0.0077057 0.0013948 0.98683 0.99163 3.0088e-006 1.2035e-005 0.14509 0.90503 0.89989 0.0014016 0.98168 0.53519 0.0018881 0.42713 1.829 1.828 16.0076 144.9732 0.00019033 -85.615 0.59095
3.695 0.98806 5.5016e-005 3.8182 0.011998 4.8428e-005 0.0011572 0.22441 0.00065923 0.22506 0.20744 0 0.032728 0.0389 0 1.1392 0.36017 0.10628 0.013828 6.5731 0.086301 0.00010723 0.80381 0.0068915 0.0077065 0.0013948 0.98683 0.99163 3.0086e-006 1.2034e-005 0.14509 0.90527 0.9 0.0014016 0.98178 0.53536 0.0018881 0.42714 1.8296 1.8286 16.0075 144.9732 0.00019015 -85.6154 0.59195
3.696 0.98806 5.5016e-005 3.8182 0.011998 4.8441e-005 0.0011572 0.22442 0.00065923 0.22507 0.20744 0 0.032727 0.0389 0 1.1393 0.36021 0.1063 0.01383 6.5745 0.086312 0.00010725 0.8038 0.0068922 0.0077073 0.0013947 0.98684 0.99163 3.0084e-006 1.2033e-005 0.1451 0.90552 0.90011 0.0014015 0.98188 0.53552 0.001888 0.42716 1.8302 1.8292 16.0075 144.9733 0.00018998 -85.6157 0.59295
3.697 0.98806 5.5016e-005 3.8182 0.011998 4.8454e-005 0.0011572 0.22443 0.00065923 0.22508 0.20745 0 0.032727 0.0389 0 1.1394 0.36026 0.10631 0.013831 6.576 0.086323 0.00010726 0.80378 0.0068929 0.007708 0.0013946 0.98684 0.99163 3.0082e-006 1.2033e-005 0.14511 0.90576 0.90023 0.0014015 0.98198 0.53568 0.001888 0.42717 1.8309 1.8299 16.0075 144.9733 0.0001898 -85.6161 0.59395
3.698 0.98806 5.5016e-005 3.8182 0.011998 4.8467e-005 0.0011572 0.22443 0.00065923 0.22509 0.20746 0 0.032726 0.0389 0 1.1395 0.36031 0.10633 0.013833 6.5774 0.086333 0.00010728 0.80377 0.0068936 0.0077088 0.0013945 0.98684 0.99164 3.008e-006 1.2032e-005 0.14511 0.906 0.90034 0.0014014 0.98208 0.53584 0.0018879 0.42718 1.8315 1.8305 16.0075 144.9733 0.00018963 -85.6164 0.59495
3.699 0.98806 5.5016e-005 3.8182 0.011998 4.848e-005 0.0011572 0.22444 0.00065923 0.2251 0.20747 0 0.032726 0.0389 0 1.1396 0.36035 0.10635 0.013835 6.5788 0.086344 0.00010729 0.80376 0.0068944 0.0077096 0.0013944 0.98684 0.99164 3.0078e-006 1.2031e-005 0.14512 0.90625 0.90045 0.0014014 0.98218 0.536 0.0018878 0.4272 1.8321 1.8311 16.0075 144.9733 0.00018945 -85.6168 0.59595
3.7 0.98806 5.5015e-005 3.8182 0.011998 4.8493e-005 0.0011572 0.22445 0.00065923 0.22511 0.20748 0 0.032726 0.0389 0 1.1397 0.3604 0.10636 0.013836 6.5803 0.086354 0.00010731 0.80375 0.0068951 0.0077103 0.0013943 0.98684 0.99164 3.0076e-006 1.203e-005 0.14512 0.90649 0.90056 0.0014013 0.98227 0.53616 0.0018878 0.42721 1.8328 1.8318 16.0074 144.9733 0.00018928 -85.6172 0.59695
3.701 0.98806 5.5015e-005 3.8182 0.011998 4.8506e-005 0.0011572 0.22446 0.00065923 0.22511 0.20749 0 0.032725 0.0389 0 1.1398 0.36045 0.10638 0.013838 6.5817 0.086365 0.00010732 0.80374 0.0068958 0.0077111 0.0013943 0.98684 0.99164 3.0074e-006 1.203e-005 0.14513 0.90673 0.90067 0.0014013 0.98237 0.53633 0.0018877 0.42722 1.8334 1.8324 16.0074 144.9734 0.00018911 -85.6175 0.59795
3.702 0.98806 5.5015e-005 3.8182 0.011998 4.8519e-005 0.0011572 0.22447 0.00065923 0.22512 0.20749 0 0.032725 0.0389 0 1.1399 0.36049 0.10639 0.01384 6.5831 0.086375 0.00010733 0.80373 0.0068965 0.0077118 0.0013942 0.98684 0.99164 3.0072e-006 1.2029e-005 0.14513 0.90697 0.90078 0.0014012 0.98247 0.53649 0.0018877 0.42724 1.834 1.8331 16.0074 144.9734 0.00018894 -85.6179 0.59895
3.703 0.98806 5.5015e-005 3.8182 0.011998 4.8532e-005 0.0011572 0.22448 0.00065923 0.22513 0.2075 0 0.032724 0.0389 0 1.14 0.36054 0.10641 0.013841 6.5846 0.086386 0.00010735 0.80372 0.0068972 0.0077126 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.14514 0.90721 0.90089 0.0014012 0.98256 0.53665 0.0018876 0.42725 1.8347 1.8337 16.0074 144.9734 0.00018877 -85.6182 0.59995
3.704 0.98806 5.5015e-005 3.8182 0.011998 4.8545e-005 0.0011572 0.22449 0.00065923 0.22514 0.20751 0 0.032724 0.0389 0 1.1401 0.36058 0.10643 0.013843 6.586 0.086396 0.00010736 0.80371 0.0068979 0.0077134 0.001394 0.98684 0.99164 3.0069e-006 1.2027e-005 0.14515 0.90745 0.901 0.0014012 0.98266 0.53681 0.0018876 0.42726 1.8353 1.8343 16.0074 144.9734 0.0001886 -85.6185 0.60095
3.705 0.98806 5.5015e-005 3.8182 0.011998 4.8558e-005 0.0011572 0.22449 0.00065923 0.22515 0.20752 0 0.032723 0.0389 0 1.1402 0.36063 0.10644 0.013845 6.5874 0.086407 0.00010738 0.8037 0.0068986 0.0077141 0.0013939 0.98684 0.99164 3.0067e-006 1.2027e-005 0.14515 0.90768 0.9011 0.0014011 0.98275 0.53697 0.0018875 0.42727 1.8359 1.8349 16.0073 144.9734 0.00018843 -85.6189 0.60195
3.706 0.98806 5.5015e-005 3.8182 0.011998 4.8571e-005 0.0011572 0.2245 0.00065923 0.22516 0.20753 0 0.032723 0.0389 0 1.1403 0.36068 0.10646 0.013847 6.5889 0.086418 0.00010739 0.80369 0.0068994 0.0077149 0.0013939 0.98685 0.99164 3.0065e-006 1.2026e-005 0.14516 0.90792 0.90121 0.0014011 0.98284 0.53713 0.0018875 0.42729 1.8365 1.8356 16.0073 144.9735 0.00018826 -85.6192 0.60295
3.707 0.98806 5.5015e-005 3.8182 0.011998 4.8584e-005 0.0011572 0.22451 0.00065923 0.22517 0.20753 0 0.032722 0.0389 0 1.1404 0.36072 0.10647 0.013848 6.5903 0.086428 0.00010741 0.80368 0.0069001 0.0077157 0.0013938 0.98685 0.99164 3.0063e-006 1.2025e-005 0.14516 0.90816 0.90132 0.001401 0.98294 0.53729 0.0018874 0.4273 1.8372 1.8362 16.0073 144.9735 0.00018809 -85.6196 0.60395
3.708 0.98806 5.5015e-005 3.8182 0.011998 4.8597e-005 0.0011572 0.22452 0.00065923 0.22517 0.20754 0 0.032722 0.0389 0 1.1405 0.36077 0.10649 0.01385 6.5917 0.086439 0.00010742 0.80367 0.0069008 0.0077164 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.14517 0.90839 0.90143 0.001401 0.98303 0.53745 0.0018873 0.42731 1.8378 1.8368 16.0073 144.9735 0.00018793 -85.6199 0.60495
3.709 0.98806 5.5015e-005 3.8182 0.011998 4.861e-005 0.0011572 0.22453 0.00065923 0.22518 0.20755 0 0.032722 0.0389 0 1.1406 0.36082 0.10651 0.013852 6.5932 0.086449 0.00010744 0.80366 0.0069015 0.0077172 0.0013936 0.98685 0.99164 3.006e-006 1.2024e-005 0.14517 0.90863 0.90153 0.001401 0.98312 0.53761 0.0018873 0.42733 1.8384 1.8374 16.0073 144.9735 0.00018776 -85.6202 0.60595
3.71 0.98806 5.5015e-005 3.8182 0.011998 4.8623e-005 0.0011572 0.22454 0.00065923 0.22519 0.20756 0 0.032721 0.0389 0 1.1407 0.36086 0.10652 0.013853 6.5946 0.08646 0.00010745 0.80365 0.0069022 0.007718 0.0013936 0.98685 0.99164 3.0058e-006 1.2023e-005 0.14518 0.90886 0.90164 0.0014009 0.98321 0.53777 0.0018872 0.42734 1.839 1.8381 16.0072 144.9736 0.0001876 -85.6206 0.60695
3.711 0.98806 5.5015e-005 3.8182 0.011998 4.8636e-005 0.0011572 0.22454 0.00065923 0.2252 0.20757 0 0.032721 0.0389 0 1.1408 0.36091 0.10654 0.013855 6.596 0.08647 0.00010746 0.80364 0.0069029 0.0077187 0.0013935 0.98685 0.99164 3.0056e-006 1.2022e-005 0.14519 0.90909 0.90175 0.0014009 0.9833 0.53794 0.0018872 0.42735 1.8396 1.8387 16.0072 144.9736 0.00018743 -85.6209 0.60795
3.712 0.98806 5.5015e-005 3.8182 0.011998 4.8649e-005 0.0011572 0.22455 0.00065923 0.22521 0.20757 0 0.03272 0.0389 0 1.1409 0.36096 0.10656 0.013857 6.5975 0.086481 0.00010748 0.80363 0.0069036 0.0077195 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.14519 0.90933 0.90185 0.0014008 0.98339 0.5381 0.0018871 0.42736 1.8402 1.8393 16.0072 144.9736 0.00018726 -85.6212 0.60895
3.713 0.98806 5.5015e-005 3.8182 0.011998 4.8662e-005 0.0011572 0.22456 0.00065923 0.22522 0.20758 0 0.03272 0.0389 0 1.141 0.361 0.10657 0.013858 6.5989 0.086491 0.00010749 0.80362 0.0069043 0.0077202 0.0013933 0.98685 0.99165 3.0053e-006 1.2021e-005 0.1452 0.90956 0.90196 0.0014008 0.98348 0.53826 0.0018871 0.42738 1.8409 1.8399 16.0072 144.9736 0.0001871 -85.6215 0.60995
3.714 0.98806 5.5014e-005 3.8182 0.011998 4.8675e-005 0.0011572 0.22457 0.00065924 0.22522 0.20759 0 0.032719 0.0389 0 1.1411 0.36105 0.10659 0.01386 6.6003 0.086502 0.00010751 0.80361 0.0069051 0.007721 0.0013932 0.98685 0.99165 3.0051e-006 1.202e-005 0.1452 0.90979 0.90206 0.0014008 0.98357 0.53842 0.001887 0.42739 1.8415 1.8405 16.0072 144.9736 0.00018694 -85.6219 0.61095
3.715 0.98806 5.5014e-005 3.8182 0.011998 4.8688e-005 0.0011572 0.22458 0.00065924 0.22523 0.2076 0 0.032719 0.0389 0 1.1412 0.36109 0.1066 0.013862 6.6018 0.086512 0.00010752 0.8036 0.0069058 0.0077218 0.0013932 0.98685 0.99165 3.0049e-006 1.202e-005 0.14521 0.91002 0.90217 0.0014007 0.98366 0.53858 0.001887 0.4274 1.8421 1.8411 16.0071 144.9737 0.00018677 -85.6222 0.61195
3.716 0.98806 5.5014e-005 3.8182 0.011998 4.8701e-005 0.0011572 0.22459 0.00065924 0.22524 0.2076 0 0.032719 0.0389 0 1.1413 0.36114 0.10662 0.013863 6.6032 0.086523 0.00010754 0.80358 0.0069065 0.0077225 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.14521 0.91025 0.90227 0.0014007 0.98375 0.53874 0.0018869 0.42742 1.8427 1.8417 16.0071 144.9737 0.00018661 -85.6225 0.61295
3.717 0.98806 5.5014e-005 3.8182 0.011998 4.8714e-005 0.0011572 0.22459 0.00065924 0.22525 0.20761 0 0.032718 0.0389 0 1.1414 0.36119 0.10664 0.013865 6.6046 0.086534 0.00010755 0.80357 0.0069072 0.0077233 0.001393 0.98686 0.99165 3.0046e-006 1.2018e-005 0.14522 0.91048 0.90237 0.0014007 0.98383 0.5389 0.0018869 0.42743 1.8433 1.8424 16.0071 144.9737 0.00018645 -85.6228 0.61395
3.718 0.98806 5.5014e-005 3.8182 0.011998 4.8727e-005 0.0011572 0.2246 0.00065924 0.22526 0.20762 0 0.032718 0.0389 0 1.1415 0.36123 0.10665 0.013867 6.6061 0.086544 0.00010757 0.80356 0.0069079 0.0077241 0.001393 0.98686 0.99165 3.0044e-006 1.2018e-005 0.14523 0.91071 0.90248 0.0014006 0.98392 0.53906 0.0018868 0.42744 1.8439 1.843 16.0071 144.9737 0.00018629 -85.6231 0.61495
3.719 0.98806 5.5014e-005 3.8182 0.011998 4.874e-005 0.0011572 0.22461 0.00065924 0.22527 0.20763 0 0.032717 0.0389 0 1.1416 0.36128 0.10667 0.013869 6.6075 0.086555 0.00010758 0.80355 0.0069086 0.0077248 0.0013929 0.98686 0.99165 3.0043e-006 1.2017e-005 0.14523 0.91093 0.90258 0.0014006 0.98401 0.53922 0.0018868 0.42746 1.8445 1.8436 16.0071 144.9737 0.00018613 -85.6234 0.61595
3.72 0.98806 5.5014e-005 3.8182 0.011998 4.8753e-005 0.0011572 0.22462 0.00065924 0.22527 0.20764 0 0.032717 0.0389 0 1.1417 0.36133 0.10668 0.01387 6.609 0.086565 0.0001076 0.80354 0.0069093 0.0077256 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.14524 0.91116 0.90268 0.0014005 0.98409 0.53938 0.0018867 0.42747 1.8451 1.8442 16.007 144.9738 0.00018597 -85.6238 0.61695
3.721 0.98806 5.5014e-005 3.8182 0.011998 4.8766e-005 0.0011572 0.22463 0.00065924 0.22528 0.20764 0 0.032716 0.0389 0 1.1418 0.36137 0.1067 0.013872 6.6104 0.086576 0.00010761 0.80353 0.0069101 0.0077264 0.0013927 0.98686 0.99165 3.0039e-006 1.2016e-005 0.14524 0.91139 0.90278 0.0014005 0.98418 0.53954 0.0018867 0.42748 1.8457 1.8448 16.007 144.9738 0.00018581 -85.6241 0.61795
3.722 0.98806 5.5014e-005 3.8182 0.011998 4.8779e-005 0.0011573 0.22464 0.00065924 0.22529 0.20765 0 0.032716 0.0389 0 1.1419 0.36142 0.10672 0.013874 6.6118 0.086586 0.00010762 0.80352 0.0069108 0.0077271 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.14525 0.91161 0.90289 0.0014005 0.98426 0.5397 0.0018866 0.42749 1.8463 1.8454 16.007 144.9738 0.00018565 -85.6244 0.61895
3.723 0.98806 5.5014e-005 3.8182 0.011998 4.8792e-005 0.0011573 0.22464 0.00065924 0.2253 0.20766 0 0.032716 0.0389 0 1.142 0.36147 0.10673 0.013875 6.6133 0.086597 0.00010764 0.80351 0.0069115 0.0077279 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.14525 0.91184 0.90299 0.0014004 0.98435 0.53986 0.0018866 0.42751 1.8469 1.846 16.007 144.9738 0.00018549 -85.6247 0.61995
3.724 0.98806 5.5014e-005 3.8182 0.011998 4.8805e-005 0.0011573 0.22465 0.00065924 0.22531 0.20767 0 0.032715 0.0389 0 1.1421 0.36151 0.10675 0.013877 6.6147 0.086607 0.00010765 0.8035 0.0069122 0.0077286 0.0013925 0.98686 0.99165 3.0035e-006 1.2014e-005 0.14526 0.91206 0.90309 0.0014004 0.98443 0.54002 0.0018865 0.42752 1.8475 1.8466 16.0069 144.9738 0.00018533 -85.625 0.62095
3.725 0.98806 5.5014e-005 3.8182 0.011998 4.8818e-005 0.0011573 0.22466 0.00065924 0.22532 0.20768 0 0.032715 0.0389 0 1.1422 0.36156 0.10676 0.013879 6.6162 0.086618 0.00010767 0.80349 0.0069129 0.0077294 0.0013925 0.98686 0.99165 3.0033e-006 1.2013e-005 0.14527 0.91228 0.90319 0.0014004 0.98451 0.54018 0.0018865 0.42753 1.8481 1.8472 16.0069 144.9739 0.00018518 -85.6253 0.62195
3.726 0.98806 5.5014e-005 3.8182 0.011998 4.8831e-005 0.0011573 0.22467 0.00065924 0.22532 0.20768 0 0.032714 0.0389 0 1.1423 0.3616 0.10678 0.01388 6.6176 0.086628 0.00010768 0.80348 0.0069136 0.0077302 0.0013924 0.98686 0.99165 3.0031e-006 1.2012e-005 0.14527 0.91251 0.90329 0.0014003 0.98459 0.54034 0.0018864 0.42755 1.8487 1.8478 16.0069 144.9739 0.00018502 -85.6256 0.62295
3.727 0.98806 5.5014e-005 3.8182 0.011998 4.8844e-005 0.0011573 0.22468 0.00065924 0.22533 0.20769 0 0.032714 0.0389 0 1.1424 0.36165 0.1068 0.013882 6.619 0.086639 0.0001077 0.80347 0.0069143 0.0077309 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.14528 0.91273 0.90339 0.0014003 0.98468 0.5405 0.0018864 0.42756 1.8493 1.8484 16.0069 144.9739 0.00018486 -85.6259 0.62395
3.728 0.98806 5.5013e-005 3.8182 0.011998 4.8857e-005 0.0011573 0.22469 0.00065924 0.22534 0.2077 0 0.032714 0.0389 0 1.1425 0.3617 0.10681 0.013884 6.6205 0.086649 0.00010771 0.80346 0.006915 0.0077317 0.0013923 0.98687 0.99165 3.0028e-006 1.2011e-005 0.14528 0.91295 0.90349 0.0014002 0.98476 0.54066 0.0018863 0.42757 1.8499 1.849 16.0069 144.9739 0.00018471 -85.6262 0.62495
3.729 0.98806 5.5013e-005 3.8182 0.011998 4.887e-005 0.0011573 0.22469 0.00065924 0.22535 0.20771 0 0.032713 0.0389 0 1.1426 0.36174 0.10683 0.013885 6.6219 0.08666 0.00010773 0.80345 0.0069158 0.0077325 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.14529 0.91317 0.90359 0.0014002 0.98484 0.54082 0.0018863 0.42758 1.8505 1.8496 16.0068 144.9739 0.00018455 -85.6264 0.62595
3.73 0.98806 5.5013e-005 3.8182 0.011998 4.8883e-005 0.0011573 0.2247 0.00065924 0.22536 0.20772 0 0.032713 0.0389 0 1.1427 0.36179 0.10685 0.013887 6.6234 0.086671 0.00010774 0.80344 0.0069165 0.0077332 0.0013921 0.98687 0.99166 3.0025e-006 1.201e-005 0.14529 0.91339 0.90369 0.0014001 0.98492 0.54098 0.0018863 0.4276 1.8511 1.8502 16.0068 144.974 0.0001844 -85.6267 0.62695
3.731 0.98806 5.5013e-005 3.8182 0.011998 4.8896e-005 0.0011573 0.22471 0.00065924 0.22537 0.20772 0 0.032712 0.0389 0 1.1428 0.36184 0.10686 0.013889 6.6248 0.086681 0.00010776 0.80343 0.0069172 0.007734 0.0013921 0.98687 0.99166 3.0024e-006 1.2009e-005 0.1453 0.91361 0.90379 0.0014001 0.985 0.54114 0.0018862 0.42761 1.8517 1.8508 16.0068 144.974 0.00018425 -85.627 0.62795
3.732 0.98806 5.5013e-005 3.8182 0.011998 4.8909e-005 0.0011573 0.22472 0.00065924 0.22537 0.20773 0 0.032712 0.0389 0 1.1429 0.36188 0.10688 0.013891 6.6263 0.086692 0.00010777 0.80342 0.0069179 0.0077348 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.14531 0.91383 0.90388 0.0014001 0.98508 0.5413 0.0018862 0.42762 1.8523 1.8513 16.0068 144.974 0.00018409 -85.6273 0.62895
3.733 0.98806 5.5013e-005 3.8182 0.011998 4.8922e-005 0.0011573 0.22473 0.00065924 0.22538 0.20774 0 0.032711 0.0389 0 1.143 0.36193 0.10689 0.013892 6.6277 0.086702 0.00010778 0.80341 0.0069186 0.0077355 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.14531 0.91405 0.90398 0.0014 0.98515 0.54146 0.0018861 0.42764 1.8528 1.8519 16.0067 144.974 0.00018394 -85.6276 0.62995
3.734 0.98806 5.5013e-005 3.8182 0.011998 4.8935e-005 0.0011573 0.22474 0.00065924 0.22539 0.20775 0 0.032711 0.0389 0 1.1431 0.36198 0.10691 0.013894 6.6291 0.086713 0.0001078 0.8034 0.0069193 0.0077363 0.0013919 0.98687 0.99166 3.0019e-006 1.2008e-005 0.14532 0.91426 0.90408 0.0014 0.98523 0.54162 0.0018861 0.42765 1.8534 1.8525 16.0067 144.974 0.00018379 -85.6279 0.63095
3.735 0.98806 5.5013e-005 3.8182 0.011998 4.8948e-005 0.0011573 0.22474 0.00065924 0.2254 0.20775 0 0.032711 0.0389 0 1.1432 0.36202 0.10693 0.013896 6.6306 0.086723 0.00010781 0.80338 0.00692 0.007737 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.14532 0.91448 0.90418 0.0014 0.98531 0.54178 0.001886 0.42766 1.854 1.8531 16.0067 144.9741 0.00018364 -85.6282 0.63195
3.736 0.98806 5.5013e-005 3.8182 0.011998 4.8961e-005 0.0011573 0.22475 0.00065924 0.22541 0.20776 0 0.03271 0.0389 0 1.1433 0.36207 0.10694 0.013897 6.632 0.086734 0.00010783 0.80337 0.0069207 0.0077378 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.14533 0.9147 0.90427 0.0013999 0.98539 0.54194 0.001886 0.42767 1.8546 1.8537 16.0067 144.9741 0.00018348 -85.6284 0.63295
3.737 0.98806 5.5013e-005 3.8182 0.011998 4.8975e-005 0.0011573 0.22476 0.00065924 0.22542 0.20777 0 0.03271 0.0389 0 1.1434 0.36212 0.10696 0.013899 6.6335 0.086744 0.00010784 0.80336 0.0069214 0.0077386 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.14533 0.91491 0.90437 0.0013999 0.98546 0.5421 0.0018859 0.42769 1.8552 1.8543 16.0067 144.9741 0.00018333 -85.6287 0.63395
3.738 0.98806 5.5013e-005 3.8182 0.011998 4.8988e-005 0.0011573 0.22477 0.00065924 0.22542 0.20778 0 0.032709 0.0389 0 1.1435 0.36216 0.10697 0.013901 6.6349 0.086755 0.00010786 0.80335 0.0069222 0.0077393 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.14534 0.91512 0.90446 0.0013999 0.98554 0.54226 0.0018859 0.4277 1.8557 1.8548 16.0066 144.9741 0.00018318 -85.629 0.63495
3.739 0.98806 5.5013e-005 3.8182 0.011998 4.9001e-005 0.0011573 0.22478 0.00065924 0.22543 0.20779 0 0.032709 0.0389 0 1.1436 0.36221 0.10699 0.013902 6.6364 0.086765 0.00010787 0.80334 0.0069229 0.0077401 0.0013915 0.98688 0.99166 3.0012e-006 1.2005e-005 0.14535 0.91534 0.90456 0.0013999 0.98562 0.54242 0.0018858 0.42771 1.8563 1.8554 16.0066 144.9741 0.00018303 -85.6293 0.63595
3.74 0.98806 5.5013e-005 3.8182 0.011998 4.9014e-005 0.0011573 0.22479 0.00065924 0.22544 0.20779 0 0.032708 0.0389 0 1.1437 0.36225 0.10701 0.013904 6.6378 0.086776 0.00010789 0.80333 0.0069236 0.0077409 0.0013915 0.98688 0.99166 3.001e-006 1.2004e-005 0.14535 0.91555 0.90466 0.0013998 0.98569 0.54258 0.0018858 0.42773 1.8569 1.856 16.0066 144.9742 0.00018289 -85.6295 0.63695
3.741 0.98806 5.5013e-005 3.8182 0.011998 4.9027e-005 0.0011573 0.22479 0.00065924 0.22545 0.2078 0 0.032708 0.0389 0 1.1438 0.3623 0.10702 0.013906 6.6393 0.086786 0.0001079 0.80332 0.0069243 0.0077416 0.0013914 0.98688 0.99166 3.0009e-006 1.2003e-005 0.14536 0.91576 0.90475 0.0013998 0.98577 0.54273 0.0018858 0.42774 1.8575 1.8566 16.0066 144.9742 0.00018274 -85.6298 0.63795
3.742 0.98806 5.5013e-005 3.8182 0.011998 4.904e-005 0.0011573 0.2248 0.00065924 0.22546 0.20781 0 0.032708 0.0389 0 1.1439 0.36235 0.10704 0.013907 6.6407 0.086797 0.00010791 0.80331 0.006925 0.0077424 0.0013913 0.98688 0.99166 3.0008e-006 1.2003e-005 0.14536 0.91598 0.90485 0.0013998 0.98584 0.54289 0.0018857 0.42775 1.858 1.8572 16.0065 144.9742 0.00018259 -85.6301 0.63895
3.743 0.98806 5.5012e-005 3.8182 0.011998 4.9053e-005 0.0011573 0.22481 0.00065924 0.22546 0.20782 0 0.032707 0.0389 0 1.144 0.36239 0.10705 0.013909 6.6422 0.086807 0.00010793 0.8033 0.0069257 0.0077431 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.14537 0.91619 0.90494 0.0013997 0.98591 0.54305 0.0018857 0.42776 1.8586 1.8577 16.0065 144.9742 0.00018244 -85.6303 0.63995
3.744 0.98806 5.5012e-005 3.8182 0.011998 4.9066e-005 0.0011573 0.22482 0.00065924 0.22547 0.20782 0 0.032707 0.0389 0 1.1441 0.36244 0.10707 0.013911 6.6436 0.086818 0.00010794 0.80329 0.0069264 0.0077439 0.0013912 0.98688 0.99166 3.0005e-006 1.2002e-005 0.14537 0.9164 0.90503 0.0013997 0.98599 0.54321 0.0018856 0.42778 1.8592 1.8583 16.0065 144.9742 0.0001823 -85.6306 0.64095
3.745 0.98806 5.5012e-005 3.8182 0.011998 4.9079e-005 0.0011573 0.22483 0.00065924 0.22548 0.20783 0 0.032706 0.0389 0 1.1442 0.36249 0.10709 0.013913 6.6451 0.086828 0.00010796 0.80328 0.0069271 0.0077447 0.0013912 0.98688 0.99166 3.0003e-006 1.2001e-005 0.14538 0.91661 0.90513 0.0013997 0.98606 0.54337 0.0018856 0.42779 1.8598 1.8589 16.0065 144.9743 0.00018215 -85.6308 0.64195
3.746 0.98806 5.5012e-005 3.8182 0.011998 4.9092e-005 0.0011573 0.22483 0.00065924 0.22549 0.20784 0 0.032706 0.0389 0 1.1443 0.36253 0.1071 0.013914 6.6465 0.086839 0.00010797 0.80327 0.0069279 0.0077454 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.14539 0.91682 0.90522 0.0013996 0.98613 0.54353 0.0018856 0.4278 1.8603 1.8595 16.0065 144.9743 0.000182 -85.6311 0.64295
3.747 0.98806 5.5012e-005 3.8182 0.011998 4.9105e-005 0.0011573 0.22484 0.00065924 0.2255 0.20785 0 0.032706 0.0389 0 1.1444 0.36258 0.10712 0.013916 6.648 0.086849 0.00010799 0.80326 0.0069286 0.0077462 0.001391 0.98688 0.99166 3.0001e-006 1.2e-005 0.14539 0.91702 0.90531 0.0013996 0.9862 0.54369 0.0018855 0.42782 1.8609 1.86 16.0064 144.9743 0.00018186 -85.6314 0.64395
3.748 0.98806 5.5012e-005 3.8182 0.011998 4.9118e-005 0.0011573 0.22485 0.00065924 0.22551 0.20786 0 0.032705 0.0389 0 1.1445 0.36263 0.10713 0.013918 6.6494 0.08686 0.000108 0.80325 0.0069293 0.007747 0.001391 0.98688 0.99166 2.9999e-006 1.2e-005 0.1454 0.91723 0.90541 0.0013996 0.98627 0.54385 0.0018855 0.42783 1.8615 1.8606 16.0064 144.9743 0.00018171 -85.6316 0.64495
3.749 0.98806 5.5012e-005 3.8182 0.011998 4.9131e-005 0.0011573 0.22486 0.00065924 0.22551 0.20786 0 0.032705 0.0389 0 1.1446 0.36267 0.10715 0.013919 6.6509 0.08687 0.00010802 0.80324 0.00693 0.0077477 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.1454 0.91744 0.9055 0.0013995 0.98634 0.54401 0.0018854 0.42784 1.862 1.8612 16.0064 144.9743 0.00018157 -85.6319 0.64595
3.75 0.98806 5.5012e-005 3.8182 0.011998 4.9144e-005 0.0011573 0.22487 0.00065924 0.22552 0.20787 0 0.032704 0.0389 0 1.1447 0.36272 0.10717 0.013921 6.6523 0.086881 0.00010803 0.80323 0.0069307 0.0077485 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.14541 0.91765 0.90559 0.0013995 0.98642 0.54416 0.0018854 0.42785 1.8626 1.8617 16.0064 144.9744 0.00018143 -85.6321 0.64695
3.751 0.98806 5.5012e-005 3.8182 0.011998 4.9157e-005 0.0011573 0.22487 0.00065924 0.22553 0.20788 0 0.032704 0.0389 0 1.1448 0.36276 0.10718 0.013923 6.6538 0.086891 0.00010804 0.80322 0.0069314 0.0077492 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.14541 0.91785 0.90568 0.0013995 0.98649 0.54432 0.0018853 0.42787 1.8632 1.8623 16.0063 144.9744 0.00018128 -85.6324 0.64795
3.752 0.98806 5.5012e-005 3.8182 0.011998 4.917e-005 0.0011573 0.22488 0.00065924 0.22554 0.20789 0 0.032703 0.0389 0 1.1449 0.36281 0.1072 0.013924 6.6552 0.086902 0.00010806 0.80321 0.0069321 0.00775 0.0013907 0.98689 0.99167 2.9994e-006 1.1997e-005 0.14542 0.91806 0.90577 0.0013994 0.98655 0.54448 0.0018853 0.42788 1.8637 1.8628 16.0063 144.9744 0.00018114 -85.6326 0.64895
3.753 0.98806 5.5012e-005 3.8182 0.011998 4.9183e-005 0.0011573 0.22489 0.00065924 0.22555 0.20789 0 0.032703 0.0389 0 1.145 0.36286 0.10722 0.013926 6.6567 0.086913 0.00010807 0.8032 0.0069328 0.0077508 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.14543 0.91826 0.90586 0.0013994 0.98662 0.54464 0.0018853 0.42789 1.8643 1.8634 16.0063 144.9744 0.000181 -85.6329 0.64995
3.754 0.98806 5.5012e-005 3.8182 0.011997 4.9196e-005 0.0011573 0.2249 0.00065924 0.22555 0.2079 0 0.032703 0.0389 0 1.145 0.3629 0.10723 0.013928 6.6581 0.086923 0.00010809 0.80319 0.0069335 0.0077515 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.14543 0.91847 0.90595 0.0013994 0.98669 0.5448 0.0018852 0.42791 1.8648 1.864 16.0063 144.9744 0.00018086 -85.6331 0.65095
3.755 0.98806 5.5012e-005 3.8182 0.011997 4.9209e-005 0.0011573 0.22491 0.00065924 0.22556 0.20791 0 0.032702 0.0389 0 1.1451 0.36295 0.10725 0.013929 6.6596 0.086934 0.0001081 0.80317 0.0069343 0.0077523 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.14544 0.91867 0.90604 0.0013993 0.98676 0.54496 0.0018852 0.42792 1.8654 1.8645 16.0062 144.9745 0.00018072 -85.6334 0.65195
3.756 0.98806 5.5012e-005 3.8182 0.011997 4.9222e-005 0.0011573 0.22492 0.00065924 0.22557 0.20792 0 0.032702 0.0389 0 1.1452 0.363 0.10726 0.013931 6.661 0.086944 0.00010812 0.80316 0.006935 0.0077531 0.0013905 0.98689 0.99167 2.9989e-006 1.1995e-005 0.14544 0.91887 0.90613 0.0013993 0.98683 0.54512 0.0018851 0.42793 1.8659 1.8651 16.0062 144.9745 0.00018058 -85.6336 0.65295
3.757 0.98806 5.5011e-005 3.8182 0.011997 4.9235e-005 0.0011573 0.22492 0.00065924 0.22558 0.20792 0 0.032701 0.0389 0 1.1453 0.36304 0.10728 0.013933 6.6625 0.086955 0.00010813 0.80315 0.0069357 0.0077538 0.0013905 0.98689 0.99167 2.9987e-006 1.1995e-005 0.14545 0.91907 0.90622 0.0013993 0.9869 0.54527 0.0018851 0.42794 1.8665 1.8656 16.0062 144.9745 0.00018044 -85.6339 0.65395
3.758 0.98806 5.5011e-005 3.8182 0.011997 4.9248e-005 0.0011573 0.22493 0.00065924 0.22559 0.20793 0 0.032701 0.0389 0 1.1454 0.36309 0.1073 0.013935 6.6639 0.086965 0.00010815 0.80314 0.0069364 0.0077546 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.14546 0.91927 0.90631 0.0013993 0.98696 0.54543 0.0018851 0.42796 1.867 1.8662 16.0062 144.9745 0.0001803 -85.6341 0.65495
3.759 0.98806 5.5011e-005 3.8182 0.011997 4.9261e-005 0.0011573 0.22494 0.00065924 0.22559 0.20794 0 0.032701 0.0389 0 1.1455 0.36314 0.10731 0.013936 6.6654 0.086976 0.00010816 0.80313 0.0069371 0.0077553 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.14546 0.91948 0.9064 0.0013992 0.98703 0.54559 0.001885 0.42797 1.8676 1.8668 16.0062 144.9745 0.00018016 -85.6343 0.65595
3.76 0.98806 5.5011e-005 3.8182 0.011997 4.9274e-005 0.0011573 0.22495 0.00065924 0.2256 0.20795 0 0.0327 0.0389 0 1.1456 0.36318 0.10733 0.013938 6.6668 0.086986 0.00010818 0.80312 0.0069378 0.0077561 0.0013903 0.98689 0.99167 2.9984e-006 1.1993e-005 0.14547 0.91968 0.90649 0.0013992 0.98709 0.54575 0.001885 0.42798 1.8682 1.8673 16.0061 144.9746 0.00018002 -85.6346 0.65695
3.761 0.98806 5.5011e-005 3.8182 0.011997 4.9287e-005 0.0011573 0.22496 0.00065924 0.22561 0.20796 0 0.0327 0.0389 0 1.1457 0.36323 0.10734 0.01394 6.6683 0.086997 0.00010819 0.80311 0.0069385 0.0077569 0.0013902 0.98689 0.99167 2.9982e-006 1.1993e-005 0.14547 0.91988 0.90658 0.0013992 0.98716 0.54591 0.001885 0.42799 1.8687 1.8679 16.0061 144.9746 0.00017988 -85.6348 0.65795
3.762 0.98806 5.5011e-005 3.8182 0.011997 4.93e-005 0.0011573 0.22496 0.00065924 0.22562 0.20796 0 0.032699 0.0389 0 1.1458 0.36328 0.10736 0.013941 6.6697 0.087007 0.0001082 0.8031 0.0069392 0.0077576 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.14548 0.92007 0.90667 0.0013992 0.98722 0.54606 0.0018849 0.42801 1.8692 1.8684 16.0061 144.9746 0.00017974 -85.635 0.65895
3.763 0.98806 5.5011e-005 3.8182 0.011997 4.9313e-005 0.0011573 0.22497 0.00065924 0.22563 0.20797 0 0.032699 0.0389 0 1.1459 0.36332 0.10738 0.013943 6.6712 0.087018 0.00010822 0.80309 0.0069399 0.0077584 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.14548 0.92027 0.90676 0.0013991 0.98729 0.54622 0.0018849 0.42802 1.8698 1.869 16.0061 144.9746 0.00017961 -85.6353 0.65995
3.764 0.98806 5.5011e-005 3.8182 0.011997 4.9326e-005 0.0011573 0.22498 0.00065924 0.22563 0.20798 0 0.032699 0.0389 0 1.146 0.36337 0.10739 0.013945 6.6726 0.087028 0.00010823 0.80308 0.0069407 0.0077591 0.0013901 0.98689 0.99167 2.9979e-006 1.1991e-005 0.14549 0.92047 0.90684 0.0013991 0.98735 0.54638 0.0018848 0.42803 1.8703 1.8695 16.006 144.9746 0.00017947 -85.6355 0.66095
3.765 0.98806 5.5011e-005 3.8182 0.011997 4.9339e-005 0.0011573 0.22499 0.00065924 0.22564 0.20799 0 0.032698 0.0389 0 1.1461 0.36341 0.10741 0.013946 6.6741 0.087039 0.00010825 0.80307 0.0069414 0.0077599 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.1455 0.92067 0.90693 0.0013991 0.98742 0.54654 0.0018848 0.42805 1.8709 1.8701 16.006 144.9747 0.00017933 -85.6357 0.66195
3.766 0.98806 5.5011e-005 3.8182 0.011997 4.9352e-005 0.0011573 0.225 0.00065924 0.22565 0.20799 0 0.032698 0.0389 0 1.1462 0.36346 0.10742 0.013948 6.6756 0.087049 0.00010826 0.80306 0.0069421 0.0077607 0.00139 0.9869 0.99167 2.9976e-006 1.199e-005 0.1455 0.92086 0.90702 0.0013991 0.98748 0.5467 0.0018848 0.42806 1.8714 1.8706 16.006 144.9747 0.0001792 -85.6359 0.66295
3.767 0.98806 5.5011e-005 3.8182 0.011997 4.9365e-005 0.0011573 0.225 0.00065924 0.22566 0.208 0 0.032697 0.0389 0 1.1463 0.36351 0.10744 0.01395 6.677 0.08706 0.00010828 0.80305 0.0069428 0.0077614 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.14551 0.92106 0.9071 0.001399 0.98754 0.54685 0.0018847 0.42807 1.872 1.8711 16.006 144.9747 0.00017906 -85.6362 0.66395
3.768 0.98806 5.5011e-005 3.8182 0.011997 4.9378e-005 0.0011573 0.22501 0.00065924 0.22567 0.20801 0 0.032697 0.0389 0 1.1464 0.36355 0.10746 0.013951 6.6785 0.08707 0.00010829 0.80304 0.0069435 0.0077622 0.0013899 0.9869 0.99167 2.9974e-006 1.1989e-005 0.14551 0.92125 0.90719 0.001399 0.98761 0.54701 0.0018847 0.42808 1.8725 1.8717 16.0059 144.9747 0.00017893 -85.6364 0.66495
3.769 0.98806 5.5011e-005 3.8182 0.011997 4.9391e-005 0.0011573 0.22502 0.00065924 0.22567 0.20802 0 0.032696 0.0389 0 1.1465 0.3636 0.10747 0.013953 6.6799 0.087081 0.00010831 0.80303 0.0069442 0.007763 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.14552 0.92145 0.90728 0.001399 0.98767 0.54717 0.0018847 0.4281 1.8731 1.8722 16.0059 144.9747 0.00017879 -85.6366 0.66595
3.77 0.98806 5.5011e-005 3.8182 0.011997 4.9404e-005 0.0011574 0.22503 0.00065924 0.22568 0.20802 0 0.032696 0.0389 0 1.1466 0.36365 0.10749 0.013955 6.6814 0.087091 0.00010832 0.80302 0.0069449 0.0077637 0.0013898 0.9869 0.99167 2.9972e-006 1.1989e-005 0.14552 0.92164 0.90736 0.0013989 0.98773 0.54733 0.0018846 0.42811 1.8736 1.8728 16.0059 144.9748 0.00017866 -85.6368 0.66695
3.771 0.98806 5.501e-005 3.8182 0.011997 4.9417e-005 0.0011574 0.22504 0.00065924 0.22569 0.20803 0 0.032696 0.0389 0 1.1467 0.36369 0.10751 0.013956 6.6828 0.087102 0.00010833 0.80301 0.0069456 0.0077645 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.14553 0.92184 0.90745 0.0013989 0.98779 0.54748 0.0018846 0.42812 1.8741 1.8733 16.0059 144.9748 0.00017853 -85.6371 0.66795
3.772 0.98806 5.501e-005 3.8182 0.011997 4.943e-005 0.0011574 0.22504 0.00065924 0.2257 0.20804 0 0.032695 0.0389 0 1.1468 0.36374 0.10752 0.013958 6.6843 0.087112 0.00010835 0.803 0.0069463 0.0077652 0.0013897 0.9869 0.99168 2.9969e-006 1.1988e-005 0.14554 0.92203 0.90753 0.0013989 0.98785 0.54764 0.0018846 0.42814 1.8747 1.8738 16.0058 144.9748 0.00017839 -85.6373 0.66895
3.773 0.98806 5.501e-005 3.8182 0.011997 4.9443e-005 0.0011574 0.22505 0.00065924 0.22571 0.20805 0 0.032695 0.0389 0 1.1469 0.36379 0.10754 0.01396 6.6858 0.087123 0.00010836 0.80299 0.0069471 0.007766 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.14554 0.92222 0.90762 0.0013988 0.98791 0.5478 0.0018845 0.42815 1.8752 1.8744 16.0058 144.9748 0.00017826 -85.6375 0.66995
3.774 0.98806 5.501e-005 3.8182 0.011997 4.9456e-005 0.0011574 0.22506 0.00065924 0.22571 0.20805 0 0.032694 0.0389 0 1.147 0.36383 0.10755 0.013962 6.6872 0.087133 0.00010838 0.80298 0.0069478 0.0077668 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.14555 0.92241 0.9077 0.0013988 0.98797 0.54796 0.0018845 0.42816 1.8757 1.8749 16.0058 144.9748 0.00017813 -85.6377 0.67095
3.775 0.98806 5.501e-005 3.8182 0.011997 4.9469e-005 0.0011574 0.22507 0.00065924 0.22572 0.20806 0 0.032694 0.0389 0 1.1471 0.36388 0.10757 0.013963 6.6887 0.087144 0.00010839 0.80296 0.0069485 0.0077675 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.14555 0.9226 0.90778 0.0013988 0.98803 0.54811 0.0018845 0.42817 1.8763 1.8755 16.0058 144.9749 0.000178 -85.6379 0.67195
3.776 0.98806 5.501e-005 3.8182 0.011997 4.9482e-005 0.0011574 0.22508 0.00065924 0.22573 0.20807 0 0.032694 0.0389 0 1.1472 0.36393 0.10759 0.013965 6.6901 0.087154 0.00010841 0.80295 0.0069492 0.0077683 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.14556 0.92279 0.90787 0.0013988 0.98809 0.54827 0.0018844 0.42819 1.8768 1.876 16.0057 144.9749 0.00017787 -85.6381 0.67295
3.777 0.98806 5.501e-005 3.8182 0.011997 4.9495e-005 0.0011574 0.22508 0.00065924 0.22574 0.20808 0 0.032693 0.0389 0 1.1473 0.36397 0.1076 0.013967 6.6916 0.087165 0.00010842 0.80294 0.0069499 0.007769 0.0013894 0.9869 0.99168 2.9964e-006 1.1985e-005 0.14556 0.92298 0.90795 0.0013987 0.98815 0.54843 0.0018844 0.4282 1.8773 1.8765 16.0057 144.9749 0.00017774 -85.6383 0.67395
3.778 0.98806 5.501e-005 3.8182 0.011997 4.9508e-005 0.0011574 0.22509 0.00065924 0.22575 0.20808 0 0.032693 0.0389 0 1.1474 0.36402 0.10762 0.013968 6.6931 0.087175 0.00010844 0.80293 0.0069506 0.0077698 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.14557 0.92317 0.90804 0.0013987 0.98821 0.54859 0.0018844 0.42821 1.8779 1.877 16.0057 144.9749 0.00017761 -85.6385 0.67495
3.779 0.98806 5.501e-005 3.8182 0.011997 4.9521e-005 0.0011574 0.2251 0.00065924 0.22575 0.20809 0 0.032692 0.0389 0 1.1475 0.36406 0.10763 0.01397 6.6945 0.087186 0.00010845 0.80292 0.0069513 0.0077706 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.14558 0.92336 0.90812 0.0013987 0.98827 0.54874 0.0018843 0.42822 1.8784 1.8776 16.0057 144.975 0.00017748 -85.6388 0.67595
3.78 0.98806 5.501e-005 3.8182 0.011997 4.9534e-005 0.0011574 0.22511 0.00065924 0.22576 0.2081 0 0.032692 0.0389 0 1.1476 0.36411 0.10765 0.013972 6.696 0.087196 0.00010846 0.80291 0.006952 0.0077713 0.0013893 0.9869 0.99168 2.996e-006 1.1984e-005 0.14558 0.92355 0.9082 0.0013987 0.98833 0.5489 0.0018843 0.42824 1.8789 1.8781 16.0056 144.975 0.00017735 -85.639 0.67695
3.781 0.98806 5.501e-005 3.8182 0.011997 4.9547e-005 0.0011574 0.22512 0.00065924 0.22577 0.20811 0 0.032692 0.0389 0 1.1477 0.36416 0.10767 0.013973 6.6975 0.087206 0.00010848 0.8029 0.0069527 0.0077721 0.0013892 0.98691 0.99168 2.9959e-006 1.1984e-005 0.14559 0.92374 0.90828 0.0013986 0.98838 0.54906 0.0018843 0.42825 1.8794 1.8786 16.0056 144.975 0.00017722 -85.6392 0.67795
3.782 0.98806 5.501e-005 3.8182 0.011997 4.956e-005 0.0011574 0.22512 0.00065924 0.22578 0.20811 0 0.032691 0.0389 0 1.1478 0.3642 0.10768 0.013975 6.6989 0.087217 0.00010849 0.80289 0.0069534 0.0077729 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.14559 0.92392 0.90836 0.0013986 0.98844 0.54921 0.0018842 0.42826 1.88 1.8792 16.0056 144.975 0.00017709 -85.6394 0.67895
3.783 0.98806 5.501e-005 3.8182 0.011997 4.9573e-005 0.0011574 0.22513 0.00065924 0.22579 0.20812 0 0.032691 0.0389 0 1.1479 0.36425 0.1077 0.013977 6.7004 0.087227 0.00010851 0.80288 0.0069542 0.0077736 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.1456 0.92411 0.90845 0.0013986 0.9885 0.54937 0.0018842 0.42828 1.8805 1.8797 16.0056 144.975 0.00017696 -85.6396 0.67995
3.784 0.98806 5.501e-005 3.8182 0.011997 4.9587e-005 0.0011574 0.22514 0.00065924 0.22579 0.20813 0 0.03269 0.0389 0 1.148 0.3643 0.10771 0.013978 6.7018 0.087238 0.00010852 0.80287 0.0069549 0.0077744 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.1456 0.9243 0.90853 0.0013986 0.98855 0.54953 0.0018842 0.42829 1.881 1.8802 16.0056 144.9751 0.00017684 -85.6398 0.68095
3.785 0.98806 5.5009e-005 3.8182 0.011997 4.96e-005 0.0011574 0.22515 0.00065924 0.2258 0.20814 0 0.03269 0.0389 0 1.1481 0.36434 0.10773 0.01398 6.7033 0.087248 0.00010854 0.80286 0.0069556 0.0077751 0.001389 0.98691 0.99168 2.9955e-006 1.1982e-005 0.14561 0.92448 0.90861 0.0013986 0.98861 0.54968 0.0018841 0.4283 1.8815 1.8807 16.0055 144.9751 0.00017671 -85.64 0.68195
3.786 0.98806 5.5009e-005 3.8182 0.011997 4.9613e-005 0.0011574 0.22516 0.00065924 0.22581 0.20814 0 0.03269 0.0389 0 1.1482 0.36439 0.10775 0.013982 6.7048 0.087259 0.00010855 0.80285 0.0069563 0.0077759 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.14562 0.92467 0.90869 0.0013985 0.98867 0.54984 0.0018841 0.42831 1.882 1.8813 16.0055 144.9751 0.00017658 -85.6402 0.68295
3.787 0.98806 5.5009e-005 3.8182 0.011997 4.9626e-005 0.0011574 0.22516 0.00065924 0.22582 0.20815 0 0.032689 0.0389 0 1.1483 0.36444 0.10776 0.013983 6.7062 0.087269 0.00010857 0.80284 0.006957 0.0077767 0.001389 0.98691 0.99168 2.9953e-006 1.1981e-005 0.14562 0.92485 0.90877 0.0013985 0.98872 0.55 0.0018841 0.42833 1.8826 1.8818 16.0055 144.9751 0.00017646 -85.6404 0.68395
3.788 0.98806 5.5009e-005 3.8182 0.011997 4.9639e-005 0.0011574 0.22517 0.00065924 0.22583 0.20816 0 0.032689 0.0389 0 1.1484 0.36448 0.10778 0.013985 6.7077 0.08728 0.00010858 0.80283 0.0069577 0.0077774 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.14563 0.92503 0.90885 0.0013985 0.98878 0.55015 0.001884 0.42834 1.8831 1.8823 16.0055 144.9751 0.00017633 -85.6406 0.68495
3.789 0.98806 5.5009e-005 3.8182 0.011997 4.9652e-005 0.0011574 0.22518 0.00065924 0.22583 0.20817 0 0.032688 0.0389 0 1.1485 0.36453 0.10779 0.013987 6.7092 0.08729 0.00010859 0.80282 0.0069584 0.0077782 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.14563 0.92522 0.90893 0.0013985 0.98883 0.55031 0.001884 0.42835 1.8836 1.8828 16.0054 144.9752 0.00017621 -85.6408 0.68595
3.79 0.98806 5.5009e-005 3.8182 0.011997 4.9665e-005 0.0011574 0.22519 0.00065924 0.22584 0.20817 0 0.032688 0.0389 0 1.1486 0.36458 0.10781 0.013989 6.7106 0.087301 0.00010861 0.80281 0.0069591 0.0077789 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.14564 0.9254 0.90901 0.0013984 0.98889 0.55047 0.001884 0.42836 1.8841 1.8833 16.0054 144.9752 0.00017608 -85.6409 0.68695
3.791 0.98806 5.5009e-005 3.8182 0.011997 4.9678e-005 0.0011574 0.22519 0.00065924 0.22585 0.20818 0 0.032688 0.0389 0 1.1487 0.36462 0.10783 0.01399 6.7121 0.087311 0.00010862 0.8028 0.0069598 0.0077797 0.0013888 0.98691 0.99168 2.9949e-006 1.1979e-005 0.14564 0.92558 0.90909 0.0013984 0.98894 0.55062 0.0018839 0.42838 1.8846 1.8838 16.0054 144.9752 0.00017596 -85.6411 0.68795
3.792 0.98806 5.5009e-005 3.8182 0.011997 4.9691e-005 0.0011574 0.2252 0.00065924 0.22586 0.20819 0 0.032687 0.0389 0 1.1488 0.36467 0.10784 0.013992 6.7136 0.087322 0.00010864 0.80279 0.0069605 0.0077805 0.0013887 0.98691 0.99168 2.9948e-006 1.1979e-005 0.14565 0.92576 0.90917 0.0013984 0.98899 0.55078 0.0018839 0.42839 1.8851 1.8844 16.0054 144.9752 0.00017583 -85.6413 0.68895
3.793 0.98806 5.5009e-005 3.8182 0.011997 4.9704e-005 0.0011574 0.22521 0.00065924 0.22587 0.2082 0 0.032687 0.0389 0 1.1489 0.36471 0.10786 0.013994 6.715 0.087332 0.00010865 0.80278 0.0069613 0.0077812 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.14566 0.92594 0.90925 0.0013984 0.98905 0.55094 0.0018839 0.4284 1.8857 1.8849 16.0053 144.9752 0.00017571 -85.6415 0.68995
3.794 0.98806 5.5009e-005 3.8182 0.011997 4.9717e-005 0.0011574 0.22522 0.00065924 0.22587 0.2082 0 0.032686 0.0389 0 1.149 0.36476 0.10788 0.013995 6.7165 0.087343 0.00010867 0.80277 0.006962 0.007782 0.0013886 0.98691 0.99168 2.9946e-006 1.1978e-005 0.14566 0.92612 0.90933 0.0013983 0.9891 0.55109 0.0018839 0.42842 1.8862 1.8854 16.0053 144.9753 0.00017559 -85.6417 0.69095
3.795 0.98806 5.5009e-005 3.8182 0.011997 4.973e-005 0.0011574 0.22523 0.00065924 0.22588 0.20821 0 0.032686 0.0389 0 1.1491 0.36481 0.10789 0.013997 6.718 0.087353 0.00010868 0.80276 0.0069627 0.0077827 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.14567 0.9263 0.9094 0.0013983 0.98915 0.55125 0.0018838 0.42843 1.8867 1.8859 16.0053 144.9753 0.00017546 -85.6419 0.69195
3.796 0.98806 5.5009e-005 3.8182 0.011997 4.9743e-005 0.0011574 0.22523 0.00065924 0.22589 0.20822 0 0.032686 0.0389 0 1.1492 0.36485 0.10791 0.013999 6.7194 0.087364 0.0001087 0.80275 0.0069634 0.0077835 0.0013886 0.98691 0.99168 2.9944e-006 1.1977e-005 0.14567 0.92648 0.90948 0.0013983 0.9892 0.55141 0.0018838 0.42844 1.8872 1.8864 16.0052 144.9753 0.00017534 -85.6421 0.69295
3.797 0.98806 5.5009e-005 3.8182 0.011997 4.9756e-005 0.0011574 0.22524 0.00065924 0.2259 0.20823 0 0.032685 0.0389 0 1.1493 0.3649 0.10792 0.014 6.7209 0.087374 0.00010871 0.80273 0.0069641 0.0077843 0.0013885 0.98691 0.99169 2.9943e-006 1.1977e-005 0.14568 0.92666 0.90956 0.0013982 0.98926 0.55156 0.0018838 0.42845 1.8877 1.8869 16.0052 144.9753 0.00017522 -85.6423 0.69395
3.798 0.98806 5.5009e-005 3.8182 0.011997 4.9769e-005 0.0011574 0.22525 0.00065924 0.2259 0.20823 0 0.032685 0.0389 0 1.1494 0.36495 0.10794 0.014002 6.7224 0.087385 0.00010872 0.80272 0.0069648 0.007785 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.14568 0.92684 0.90964 0.0013982 0.98931 0.55172 0.0018837 0.42847 1.8882 1.8874 16.0052 144.9753 0.0001751 -85.6424 0.69495
3.799 0.98806 5.5009e-005 3.8182 0.011997 4.9782e-005 0.0011574 0.22526 0.00065924 0.22591 0.20824 0 0.032684 0.0389 0 1.1495 0.36499 0.10796 0.014004 6.7238 0.087395 0.00010874 0.80271 0.0069655 0.0077858 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.14569 0.92701 0.90972 0.0013982 0.98936 0.55187 0.0018837 0.42848 1.8887 1.8879 16.0052 144.9754 0.00017498 -85.6426 0.69595
3.8 0.98806 5.5008e-005 3.8182 0.011997 4.9795e-005 0.0011574 0.22527 0.00065924 0.22592 0.20825 0 0.032684 0.0389 0 1.1496 0.36504 0.10797 0.014005 6.7253 0.087406 0.00010875 0.8027 0.0069662 0.0077865 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.1457 0.92719 0.90979 0.0013982 0.98941 0.55203 0.0018837 0.42849 1.8892 1.8884 16.0051 144.9754 0.00017486 -85.6428 0.69695
3.801 0.98806 5.5008e-005 3.8182 0.011997 4.9808e-005 0.0011574 0.22527 0.00065924 0.22593 0.20826 0 0.032684 0.0389 0 1.1497 0.36509 0.10799 0.014007 6.7268 0.087416 0.00010877 0.80269 0.0069669 0.0077873 0.0013883 0.98692 0.99169 2.9939e-006 1.1976e-005 0.1457 0.92737 0.90987 0.0013981 0.98946 0.55219 0.0018836 0.4285 1.8897 1.8889 16.0051 144.9754 0.00017474 -85.643 0.69795
3.802 0.98806 5.5008e-005 3.8182 0.011997 4.9821e-005 0.0011574 0.22528 0.00065924 0.22594 0.20826 0 0.032683 0.0389 0 1.1498 0.36513 0.108 0.014009 6.7282 0.087427 0.00010878 0.80268 0.0069676 0.0077881 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.14571 0.92754 0.90995 0.0013981 0.98951 0.55234 0.0018836 0.42852 1.8902 1.8895 16.0051 144.9754 0.00017462 -85.6432 0.69895
3.803 0.98806 5.5008e-005 3.8182 0.011997 4.9834e-005 0.0011574 0.22529 0.00065924 0.22594 0.20827 0 0.032683 0.0389 0 1.1499 0.36518 0.10802 0.01401 6.7297 0.087437 0.0001088 0.80267 0.0069683 0.0077888 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.14571 0.92772 0.91002 0.0013981 0.98956 0.5525 0.0018836 0.42853 1.8907 1.89 16.0051 144.9754 0.0001745 -85.6433 0.69995
3.804 0.98806 5.5008e-005 3.8182 0.011997 4.9847e-005 0.0011574 0.2253 0.00065924 0.22595 0.20828 0 0.032682 0.0389 0 1.15 0.36523 0.10804 0.014012 6.7312 0.087447 0.00010881 0.80266 0.0069691 0.0077896 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.14572 0.92789 0.9101 0.0013981 0.98961 0.55265 0.0018836 0.42854 1.8912 1.8905 16.005 144.9755 0.00017438 -85.6435 0.70095
3.805 0.98806 5.5008e-005 3.8182 0.011997 4.986e-005 0.0011574 0.2253 0.00065924 0.22596 0.20829 0 0.032682 0.0389 0 1.1501 0.36527 0.10805 0.014014 6.7327 0.087458 0.00010883 0.80265 0.0069698 0.0077903 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.14572 0.92806 0.91017 0.0013981 0.98966 0.55281 0.0018835 0.42855 1.8917 1.891 16.005 144.9755 0.00017426 -85.6437 0.70195
3.806 0.98806 5.5008e-005 3.8182 0.011997 4.9873e-005 0.0011574 0.22531 0.00065924 0.22597 0.20829 0 0.032682 0.0389 0 1.1502 0.36532 0.10807 0.014015 6.7341 0.087468 0.00010884 0.80264 0.0069705 0.0077911 0.0013881 0.98692 0.99169 2.9934e-006 1.1974e-005 0.14573 0.92824 0.91025 0.0013981 0.98971 0.55296 0.0018835 0.42857 1.8922 1.8915 16.005 144.9755 0.00017415 -85.6439 0.70295
3.807 0.98806 5.5008e-005 3.8182 0.011997 4.9886e-005 0.0011574 0.22532 0.00065924 0.22597 0.2083 0 0.032681 0.0389 0 1.1503 0.36536 0.10808 0.014017 6.7356 0.087479 0.00010885 0.80263 0.0069712 0.0077919 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.14574 0.92841 0.91032 0.0013981 0.98976 0.55312 0.0018835 0.42858 1.8927 1.892 16.005 144.9755 0.00017403 -85.644 0.70395
3.808 0.98806 5.5008e-005 3.8182 0.011997 4.9899e-005 0.0011574 0.22533 0.00065924 0.22598 0.20831 0 0.032681 0.0389 0 1.1504 0.36541 0.1081 0.014019 6.7371 0.087489 0.00010887 0.80262 0.0069719 0.0077926 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.14574 0.92858 0.9104 0.001398 0.9898 0.55328 0.0018835 0.42859 1.8932 1.8925 16.0049 144.9755 0.00017391 -85.6442 0.70495
3.809 0.98806 5.5008e-005 3.8182 0.011997 4.9912e-005 0.0011574 0.22534 0.00065924 0.22599 0.20832 0 0.03268 0.0389 0 1.1505 0.36546 0.10812 0.014021 6.7385 0.0875 0.00010888 0.80261 0.0069726 0.0077934 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.14575 0.92875 0.91047 0.001398 0.98985 0.55343 0.0018834 0.4286 1.8937 1.893 16.0049 144.9756 0.00017379 -85.6444 0.70595
3.81 0.98806 5.5008e-005 3.8182 0.011997 4.9925e-005 0.0011574 0.22534 0.00065924 0.226 0.20832 0 0.03268 0.0389 0 1.1506 0.3655 0.10813 0.014022 6.74 0.08751 0.0001089 0.8026 0.0069733 0.0077941 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.14575 0.92893 0.91055 0.001398 0.9899 0.55359 0.0018834 0.42862 1.8942 1.8934 16.0049 144.9756 0.00017368 -85.6445 0.70695
3.811 0.98806 5.5008e-005 3.8182 0.011997 4.9938e-005 0.0011574 0.22535 0.00065924 0.22601 0.20833 0 0.03268 0.0389 0 1.1507 0.36555 0.10815 0.014024 6.7415 0.087521 0.00010891 0.80259 0.006974 0.0077949 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.14576 0.9291 0.91062 0.001398 0.98995 0.55374 0.0018834 0.42863 1.8947 1.8939 16.0049 144.9756 0.00017356 -85.6447 0.70795
3.812 0.98806 5.5008e-005 3.8182 0.011997 4.9951e-005 0.0011574 0.22536 0.00065924 0.22601 0.20834 0 0.032679 0.0389 0 1.1508 0.3656 0.10816 0.014026 6.743 0.087531 0.00010893 0.80258 0.0069747 0.0077957 0.0013879 0.98692 0.99169 2.9929e-006 1.1972e-005 0.14576 0.92927 0.91069 0.001398 0.98999 0.5539 0.0018833 0.42864 1.8952 1.8944 16.0048 144.9756 0.00017345 -85.6449 0.70895
3.813 0.98806 5.5008e-005 3.8182 0.011997 4.9964e-005 0.0011574 0.22537 0.00065924 0.22602 0.20835 0 0.032679 0.0389 0 1.1509 0.36564 0.10818 0.014027 6.7444 0.087542 0.00010894 0.80257 0.0069754 0.0077964 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.14577 0.92944 0.91077 0.001398 0.99004 0.55405 0.0018833 0.42866 1.8957 1.8949 16.0048 144.9756 0.00017333 -85.645 0.70995
3.814 0.98806 5.5007e-005 3.8182 0.011997 4.9977e-005 0.0011574 0.22537 0.00065924 0.22603 0.20835 0 0.032678 0.0389 0 1.151 0.36569 0.1082 0.014029 6.7459 0.087552 0.00010896 0.80256 0.0069761 0.0077972 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.14577 0.9296 0.91084 0.0013979 0.99009 0.55421 0.0018833 0.42867 1.8962 1.8954 16.0048 144.9757 0.00017322 -85.6452 0.71095
3.815 0.98806 5.5007e-005 3.8182 0.011997 4.999e-005 0.0011574 0.22538 0.00065924 0.22604 0.20836 0 0.032678 0.0389 0 1.1511 0.36574 0.10821 0.014031 6.7474 0.087563 0.00010897 0.80255 0.0069769 0.0077979 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.14578 0.92977 0.91091 0.0013979 0.99013 0.55436 0.0018833 0.42868 1.8967 1.8959 16.0048 144.9757 0.0001731 -85.6454 0.71195
3.816 0.98806 5.5007e-005 3.8182 0.011997 5.0003e-005 0.0011574 0.22539 0.00065924 0.22604 0.20837 0 0.032678 0.0389 0 1.1512 0.36578 0.10823 0.014032 6.7489 0.087573 0.00010898 0.80254 0.0069776 0.0077987 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.14579 0.92994 0.91099 0.0013979 0.99018 0.55452 0.0018832 0.42869 1.8971 1.8964 16.0047 144.9757 0.00017299 -85.6455 0.71295
3.817 0.98806 5.5007e-005 3.8182 0.011997 5.0016e-005 0.0011574 0.2254 0.00065924 0.22605 0.20837 0 0.032677 0.0389 0 1.1513 0.36583 0.10825 0.014034 6.7503 0.087583 0.000109 0.80253 0.0069783 0.0077995 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.14579 0.93011 0.91106 0.0013979 0.99022 0.55467 0.0018832 0.42871 1.8976 1.8969 16.0047 144.9757 0.00017288 -85.6457 0.71395
3.818 0.98806 5.5007e-005 3.8182 0.011997 5.0029e-005 0.0011575 0.2254 0.00065924 0.22606 0.20838 0 0.032677 0.0389 0 1.1514 0.36588 0.10826 0.014036 6.7518 0.087594 0.00010901 0.80252 0.006979 0.0078002 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.1458 0.93028 0.91113 0.0013978 0.99027 0.55483 0.0018832 0.42872 1.8981 1.8974 16.0047 144.9757 0.00017276 -85.6458 0.71495
3.819 0.98806 5.5007e-005 3.8182 0.011997 5.0042e-005 0.0011575 0.22541 0.00065924 0.22607 0.20839 0 0.032676 0.0389 0 1.1515 0.36592 0.10828 0.014037 6.7533 0.087604 0.00010903 0.8025 0.0069797 0.007801 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.1458 0.93044 0.9112 0.0013978 0.99031 0.55498 0.0018832 0.42873 1.8986 1.8979 16.0047 144.9758 0.00017265 -85.646 0.71595
3.82 0.98806 5.5007e-005 3.8182 0.011996 5.0055e-005 0.0011575 0.22542 0.00065924 0.22607 0.2084 0 0.032676 0.0389 0 1.1516 0.36597 0.10829 0.014039 6.7548 0.087615 0.00010904 0.80249 0.0069804 0.0078017 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.14581 0.93061 0.91128 0.0013978 0.99036 0.55514 0.0018831 0.42874 1.8991 1.8983 16.0046 144.9758 0.00017254 -85.6462 0.71695
3.821 0.98806 5.5007e-005 3.8182 0.011996 5.0068e-005 0.0011575 0.22543 0.00065924 0.22608 0.2084 0 0.032676 0.0389 0 1.1517 0.36601 0.10831 0.014041 6.7562 0.087625 0.00010906 0.80248 0.0069811 0.0078025 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.14581 0.93077 0.91135 0.0013978 0.9904 0.55529 0.0018831 0.42876 1.8996 1.8988 16.0046 144.9758 0.00017243 -85.6463 0.71795
3.822 0.98806 5.5007e-005 3.8182 0.011996 5.0081e-005 0.0011575 0.22544 0.00065924 0.22609 0.20841 0 0.032675 0.0389 0 1.1518 0.36606 0.10833 0.014042 6.7577 0.087636 0.00010907 0.80247 0.0069818 0.0078033 0.0013875 0.98693 0.99169 2.9921e-006 1.1968e-005 0.14582 0.93094 0.91142 0.0013978 0.99045 0.55545 0.0018831 0.42877 1.9 1.8993 16.0046 144.9758 0.00017232 -85.6465 0.71895
3.823 0.98806 5.5007e-005 3.8182 0.011996 5.0094e-005 0.0011575 0.22544 0.00065924 0.2261 0.20842 0 0.032675 0.0389 0 1.1519 0.36611 0.10834 0.014044 6.7592 0.087646 0.00010909 0.80246 0.0069825 0.007804 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.14583 0.9311 0.91149 0.0013977 0.99049 0.5556 0.0018831 0.42878 1.9005 1.8998 16.0045 144.9758 0.0001722 -85.6466 0.71995
3.824 0.98806 5.5007e-005 3.8182 0.011996 5.0107e-005 0.0011575 0.22545 0.00065924 0.22611 0.20843 0 0.032675 0.0389 0 1.152 0.36615 0.10836 0.014046 6.7607 0.087657 0.0001091 0.80245 0.0069832 0.0078048 0.0013875 0.98693 0.99169 2.9919e-006 1.1967e-005 0.14583 0.93127 0.91156 0.0013977 0.99053 0.55576 0.001883 0.42879 1.901 1.9003 16.0045 144.9759 0.00017209 -85.6468 0.72095
3.825 0.98806 5.5007e-005 3.8182 0.011996 5.012e-005 0.0011575 0.22546 0.00065924 0.22611 0.20843 0 0.032674 0.0389 0 1.1521 0.3662 0.10837 0.014047 6.7621 0.087667 0.00010911 0.80244 0.0069839 0.0078055 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.14584 0.93143 0.91163 0.0013977 0.99058 0.55591 0.001883 0.42881 1.9015 1.9008 16.0045 144.9759 0.00017198 -85.6469 0.72195
3.826 0.98806 5.5007e-005 3.8182 0.011996 5.0133e-005 0.0011575 0.22547 0.00065924 0.22612 0.20844 0 0.032674 0.0389 0 1.1522 0.36625 0.10839 0.014049 6.7636 0.087678 0.00010913 0.80243 0.0069846 0.0078063 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.14584 0.93159 0.9117 0.0013977 0.99062 0.55607 0.001883 0.42882 1.902 1.9012 16.0045 144.9759 0.00017187 -85.6471 0.72295
3.827 0.98806 5.5007e-005 3.8182 0.011996 5.0146e-005 0.0011575 0.22547 0.00065924 0.22613 0.20845 0 0.032673 0.0389 0 1.1523 0.36629 0.10841 0.014051 6.7651 0.087688 0.00010914 0.80242 0.0069853 0.0078071 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.14585 0.93176 0.91177 0.0013977 0.99066 0.55622 0.001883 0.42883 1.9024 1.9017 16.0044 144.9759 0.00017176 -85.6472 0.72395
3.828 0.98807 5.5006e-005 3.8182 0.011996 5.0159e-005 0.0011575 0.22548 0.00065924 0.22614 0.20845 0 0.032673 0.0389 0 1.1524 0.36634 0.10842 0.014052 6.7666 0.087698 0.00010916 0.80241 0.0069861 0.0078078 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.14585 0.93192 0.91184 0.0013976 0.99071 0.55638 0.0018829 0.42884 1.9029 1.9022 16.0044 144.976 0.00017165 -85.6474 0.72495
3.829 0.98807 5.5006e-005 3.8182 0.011996 5.0172e-005 0.0011575 0.22549 0.00065924 0.22614 0.20846 0 0.032673 0.0389 0 1.1525 0.36639 0.10844 0.014054 6.7681 0.087709 0.00010917 0.8024 0.0069868 0.0078086 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.14586 0.93208 0.91191 0.0013976 0.99075 0.55653 0.0018829 0.42886 1.9034 1.9027 16.0044 144.976 0.00017155 -85.6475 0.72595
3.83 0.98807 5.5006e-005 3.8182 0.011996 5.0185e-005 0.0011575 0.2255 0.00065924 0.22615 0.20847 0 0.032672 0.0389 0 1.1526 0.36643 0.10845 0.014056 6.7695 0.087719 0.00010919 0.80239 0.0069875 0.0078093 0.0013873 0.98693 0.9917 2.9914e-006 1.1966e-005 0.14587 0.93224 0.91198 0.0013976 0.99079 0.55668 0.0018829 0.42887 1.9039 1.9031 16.0044 144.976 0.00017144 -85.6477 0.72695
3.831 0.98807 5.5006e-005 3.8182 0.011996 5.0198e-005 0.0011575 0.2255 0.00065924 0.22616 0.20848 0 0.032672 0.0389 0 1.1527 0.36648 0.10847 0.014058 6.771 0.08773 0.0001092 0.80238 0.0069882 0.0078101 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.14587 0.9324 0.91205 0.0013976 0.99083 0.55684 0.0018829 0.42888 1.9043 1.9036 16.0043 144.976 0.00017133 -85.6478 0.72795
3.832 0.98807 5.5006e-005 3.8182 0.011996 5.0211e-005 0.0011575 0.22551 0.00065924 0.22617 0.20848 0 0.032671 0.0389 0 1.1528 0.36653 0.10849 0.014059 6.7725 0.08774 0.00010922 0.80237 0.0069889 0.0078108 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.14588 0.93256 0.91212 0.0013976 0.99087 0.55699 0.0018829 0.42889 1.9048 1.9041 16.0043 144.976 0.00017122 -85.648 0.72895
3.833 0.98807 5.5006e-005 3.8182 0.011996 5.0224e-005 0.0011575 0.22552 0.00065924 0.22617 0.20849 0 0.032671 0.0389 0 1.1529 0.36657 0.1085 0.014061 6.774 0.087751 0.00010923 0.80236 0.0069896 0.0078116 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.14588 0.93272 0.91218 0.0013975 0.99091 0.55715 0.0018828 0.42891 1.9053 1.9046 16.0043 144.9761 0.00017111 -85.6481 0.72995
3.834 0.98807 5.5006e-005 3.8182 0.011996 5.0237e-005 0.0011575 0.22553 0.00065924 0.22618 0.2085 0 0.032671 0.0389 0 1.153 0.36662 0.10852 0.014063 6.7755 0.087761 0.00010924 0.80235 0.0069903 0.0078124 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.14589 0.93288 0.91225 0.0013975 0.99095 0.5573 0.0018828 0.42892 1.9057 1.905 16.0043 144.9761 0.00017101 -85.6482 0.73095
3.835 0.98807 5.5006e-005 3.8182 0.011996 5.025e-005 0.0011575 0.22553 0.00065924 0.22619 0.2085 0 0.03267 0.0389 0 1.1531 0.36667 0.10853 0.014064 6.777 0.087772 0.00010926 0.80234 0.006991 0.0078131 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.14589 0.93304 0.91232 0.0013975 0.99099 0.55746 0.0018828 0.42893 1.9062 1.9055 16.0042 144.9761 0.0001709 -85.6484 0.73195
3.836 0.98807 5.5006e-005 3.8182 0.011996 5.0263e-005 0.0011575 0.22554 0.00065924 0.2262 0.20851 0 0.03267 0.0389 0 1.1532 0.36671 0.10855 0.014066 6.7784 0.087782 0.00010927 0.80233 0.0069917 0.0078139 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.1459 0.93319 0.91239 0.0013975 0.99103 0.55761 0.0018828 0.42894 1.9067 1.906 16.0042 144.9761 0.00017079 -85.6485 0.73295
3.837 0.98807 5.5006e-005 3.8182 0.011996 5.0277e-005 0.0011575 0.22555 0.00065924 0.2262 0.20852 0 0.032669 0.0389 0 1.1533 0.36676 0.10857 0.014068 6.7799 0.087792 0.00010929 0.80232 0.0069924 0.0078146 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.14591 0.93335 0.91246 0.0013975 0.99107 0.55776 0.0018827 0.42896 1.9071 1.9064 16.0042 144.9761 0.00017069 -85.6487 0.73395
3.838 0.98807 5.5006e-005 3.8182 0.011996 5.029e-005 0.0011575 0.22556 0.00065924 0.22621 0.20853 0 0.032669 0.0389 0 1.1534 0.3668 0.10858 0.014069 6.7814 0.087803 0.0001093 0.80231 0.0069931 0.0078154 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.14591 0.93351 0.91252 0.0013975 0.99111 0.55792 0.0018827 0.42897 1.9076 1.9069 16.0041 144.9762 0.00017058 -85.6488 0.73495
3.839 0.98807 5.5006e-005 3.8182 0.011996 5.0303e-005 0.0011575 0.22556 0.00065924 0.22622 0.20853 0 0.032669 0.0389 0 1.1535 0.36685 0.1086 0.014071 6.7829 0.087813 0.00010932 0.8023 0.0069938 0.0078162 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.14592 0.93366 0.91259 0.0013974 0.99115 0.55807 0.0018827 0.42898 1.9081 1.9074 16.0041 144.9762 0.00017048 -85.6489 0.73595
3.84 0.98807 5.5006e-005 3.8182 0.011996 5.0316e-005 0.0011575 0.22557 0.00065924 0.22623 0.20854 0 0.032668 0.0389 0 1.1536 0.3669 0.10862 0.014073 6.7844 0.087824 0.00010933 0.80229 0.0069945 0.0078169 0.0013869 0.98694 0.9917 2.9907e-006 1.1963e-005 0.14592 0.93382 0.91266 0.0013974 0.99119 0.55823 0.0018827 0.42899 1.9085 1.9078 16.0041 144.9762 0.00017037 -85.6491 0.73695
3.841 0.98807 5.5006e-005 3.8182 0.011996 5.0329e-005 0.0011575 0.22558 0.00065924 0.22623 0.20855 0 0.032668 0.0389 0 1.1536 0.36694 0.10863 0.014074 6.7859 0.087834 0.00010934 0.80228 0.0069953 0.0078177 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.14593 0.93398 0.91272 0.0013974 0.99123 0.55838 0.0018827 0.42901 1.909 1.9083 16.0041 144.9762 0.00017027 -85.6492 0.73795
3.842 0.98807 5.5005e-005 3.8182 0.011996 5.0342e-005 0.0011575 0.22559 0.00065924 0.22624 0.20855 0 0.032668 0.0389 0 1.1537 0.36699 0.10865 0.014076 6.7873 0.087845 0.00010936 0.80226 0.006996 0.0078184 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.14593 0.93413 0.91279 0.0013974 0.99127 0.55853 0.0018826 0.42902 1.9095 1.9088 16.004 144.9762 0.00017017 -85.6493 0.73895
3.843 0.98807 5.5005e-005 3.8182 0.011996 5.0355e-005 0.0011575 0.22559 0.00065924 0.22625 0.20856 0 0.032667 0.0389 0 1.1538 0.36704 0.10866 0.014078 6.7888 0.087855 0.00010937 0.80225 0.0069967 0.0078192 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.14594 0.93428 0.91286 0.0013974 0.99131 0.55869 0.0018826 0.42903 1.9099 1.9092 16.004 144.9763 0.00017006 -85.6495 0.73995
3.844 0.98807 5.5005e-005 3.8182 0.011996 5.0368e-005 0.0011575 0.2256 0.00065924 0.22626 0.20857 0 0.032667 0.0389 0 1.1539 0.36708 0.10868 0.014079 6.7903 0.087865 0.00010939 0.80224 0.0069974 0.0078199 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.14595 0.93444 0.91292 0.0013974 0.99135 0.55884 0.0018826 0.42904 1.9104 1.9097 16.004 144.9763 0.00016996 -85.6496 0.74095
3.845 0.98807 5.5005e-005 3.8182 0.011996 5.0381e-005 0.0011575 0.22561 0.00065924 0.22626 0.20858 0 0.032666 0.0389 0 1.154 0.36713 0.1087 0.014081 6.7918 0.087876 0.0001094 0.80223 0.0069981 0.0078207 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.14595 0.93459 0.91299 0.0013973 0.99139 0.55899 0.0018826 0.42906 1.9108 1.9102 16.004 144.9763 0.00016986 -85.6497 0.74195
3.846 0.98807 5.5005e-005 3.8182 0.011996 5.0394e-005 0.0011575 0.22562 0.00065924 0.22627 0.20858 0 0.032666 0.0389 0 1.1541 0.36718 0.10871 0.014083 6.7933 0.087886 0.00010942 0.80222 0.0069988 0.0078215 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.14596 0.93474 0.91305 0.0013973 0.99142 0.55915 0.0018825 0.42907 1.9113 1.9106 16.0039 144.9763 0.00016975 -85.6499 0.74295
3.847 0.98807 5.5005e-005 3.8182 0.011996 5.0407e-005 0.0011575 0.22563 0.00065924 0.22628 0.20859 0 0.032666 0.0389 0 1.1542 0.36722 0.10873 0.014084 6.7948 0.087897 0.00010943 0.80221 0.0069995 0.0078222 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.14596 0.9349 0.91312 0.0013973 0.99146 0.5593 0.0018825 0.42908 1.9118 1.9111 16.0039 144.9763 0.00016965 -85.65 0.74395
3.848 0.98807 5.5005e-005 3.8182 0.011996 5.042e-005 0.0011575 0.22563 0.00065924 0.22629 0.2086 0 0.032665 0.0389 0 1.1543 0.36727 0.10874 0.014086 6.7963 0.087907 0.00010945 0.8022 0.0070002 0.007823 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.14597 0.93505 0.91318 0.0013973 0.9915 0.55945 0.0018825 0.42909 1.9122 1.9115 16.0039 144.9764 0.00016955 -85.6501 0.74495
3.849 0.98807 5.5005e-005 3.8182 0.011996 5.0433e-005 0.0011575 0.22564 0.00065924 0.22629 0.2086 0 0.032665 0.0389 0 1.1544 0.36732 0.10876 0.014088 6.7977 0.087918 0.00010946 0.80219 0.0070009 0.0078237 0.0013867 0.98694 0.9917 2.99e-006 1.196e-005 0.14597 0.9352 0.91325 0.0013973 0.99153 0.55961 0.0018825 0.42911 1.9127 1.912 16.0038 144.9764 0.00016945 -85.6503 0.74595
3.85 0.98807 5.5005e-005 3.8182 0.011996 5.0446e-005 0.0011575 0.22565 0.00065924 0.2263 0.20861 0 0.032664 0.0389 0 1.1545 0.36736 0.10878 0.014089 6.7992 0.087928 0.00010947 0.80218 0.0070016 0.0078245 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.14598 0.93535 0.91331 0.0013973 0.99157 0.55976 0.0018825 0.42912 1.9131 1.9124 16.0038 144.9764 0.00016935 -85.6504 0.74695
3.851 0.98807 5.5005e-005 3.8182 0.011996 5.0459e-005 0.0011575 0.22566 0.00065924 0.22631 0.20862 0 0.032664 0.0389 0 1.1546 0.36741 0.10879 0.014091 6.8007 0.087938 0.00010949 0.80217 0.0070023 0.0078253 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.14599 0.9355 0.91338 0.0013972 0.99161 0.55991 0.0018824 0.42913 1.9136 1.9129 16.0038 144.9764 0.00016925 -85.6505 0.74795
3.852 0.98807 5.5005e-005 3.8182 0.011996 5.0472e-005 0.0011575 0.22566 0.00065924 0.22632 0.20863 0 0.032664 0.0389 0 1.1547 0.36745 0.10881 0.014093 6.8022 0.087949 0.0001095 0.80216 0.007003 0.007826 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.14599 0.93565 0.91344 0.0013972 0.99164 0.56007 0.0018824 0.42914 1.914 1.9134 16.0038 144.9764 0.00016914 -85.6506 0.74895
3.853 0.98807 5.5005e-005 3.8182 0.011996 5.0485e-005 0.0011575 0.22567 0.00065924 0.22632 0.20863 0 0.032663 0.0389 0 1.1548 0.3675 0.10882 0.014094 6.8037 0.087959 0.00010952 0.80215 0.0070037 0.0078268 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.146 0.9358 0.91351 0.0013972 0.99168 0.56022 0.0018824 0.42916 1.9145 1.9138 16.0037 144.9765 0.00016904 -85.6508 0.74995
3.854 0.98807 5.5005e-005 3.8182 0.011996 5.0498e-005 0.0011575 0.22568 0.00065924 0.22633 0.20864 0 0.032663 0.0389 0 1.1549 0.36755 0.10884 0.014096 6.8052 0.08797 0.00010953 0.80214 0.0070044 0.0078275 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.146 0.93595 0.91357 0.0013972 0.99172 0.56037 0.0018824 0.42917 1.9149 1.9143 16.0037 144.9765 0.00016894 -85.6509 0.75095
3.855 0.98807 5.5005e-005 3.8182 0.011996 5.0511e-005 0.0011575 0.22568 0.00065924 0.22634 0.20865 0 0.032663 0.0389 0 1.155 0.36759 0.10886 0.014098 6.8067 0.08798 0.00010955 0.80213 0.0070051 0.0078283 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.14601 0.9361 0.91363 0.0013972 0.99175 0.56053 0.0018824 0.42918 1.9154 1.9147 16.0037 144.9765 0.00016885 -85.651 0.75195
3.856 0.98807 5.5004e-005 3.8182 0.011996 5.0524e-005 0.0011575 0.22569 0.00065924 0.22635 0.20865 0 0.032662 0.0389 0 1.1551 0.36764 0.10887 0.014099 6.8082 0.087991 0.00010956 0.80212 0.0070059 0.007829 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.14601 0.93625 0.9137 0.0013972 0.99179 0.56068 0.0018823 0.42919 1.9158 1.9152 16.0037 144.9765 0.00016875 -85.6511 0.75295
3.857 0.98807 5.5004e-005 3.8182 0.011996 5.0537e-005 0.0011575 0.2257 0.00065924 0.22635 0.20866 0 0.032662 0.0389 0 1.1552 0.36769 0.10889 0.014101 6.8097 0.088001 0.00010958 0.80211 0.0070066 0.0078298 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.14602 0.9364 0.91376 0.0013972 0.99182 0.56083 0.0018823 0.4292 1.9163 1.9156 16.0036 144.9765 0.00016865 -85.6513 0.75395
3.858 0.98807 5.5004e-005 3.8182 0.011996 5.055e-005 0.0011575 0.22571 0.00065924 0.22636 0.20867 0 0.032661 0.0389 0 1.1553 0.36773 0.1089 0.014103 6.8111 0.088011 0.00010959 0.8021 0.0070073 0.0078306 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.14603 0.93654 0.91382 0.0013971 0.99186 0.56099 0.0018823 0.42922 1.9167 1.9161 16.0036 144.9766 0.00016855 -85.6514 0.75495
3.859 0.98807 5.5004e-005 3.8182 0.011996 5.0563e-005 0.0011575 0.22571 0.00065924 0.22637 0.20868 0 0.032661 0.0389 0 1.1554 0.36778 0.10892 0.014104 6.8126 0.088022 0.0001096 0.80209 0.007008 0.0078313 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.14603 0.93669 0.91389 0.0013971 0.99189 0.56114 0.0018823 0.42923 1.9172 1.9165 16.0036 144.9766 0.00016845 -85.6515 0.75595
3.86 0.98807 5.5004e-005 3.8182 0.011996 5.0576e-005 0.0011575 0.22572 0.00065924 0.22638 0.20868 0 0.032661 0.0389 0 1.1555 0.36783 0.10894 0.014106 6.8141 0.088032 0.00010962 0.80208 0.0070087 0.0078321 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.14604 0.93684 0.91395 0.0013971 0.99193 0.56129 0.0018823 0.42924 1.9176 1.917 16.0035 144.9766 0.00016835 -85.6516 0.75695
3.861 0.98807 5.5004e-005 3.8182 0.011996 5.0589e-005 0.0011575 0.22573 0.00065924 0.22638 0.20869 0 0.03266 0.0389 0 1.1556 0.36787 0.10895 0.014108 6.8156 0.088043 0.00010963 0.80207 0.0070094 0.0078328 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.14604 0.93698 0.91401 0.0013971 0.99196 0.56144 0.0018822 0.42925 1.9181 1.9174 16.0035 144.9766 0.00016826 -85.6517 0.75795
3.862 0.98807 5.5004e-005 3.8182 0.011996 5.0602e-005 0.0011575 0.22574 0.00065924 0.22639 0.2087 0 0.03266 0.0389 0 1.1557 0.36792 0.10897 0.01411 6.8171 0.088053 0.00010965 0.80206 0.0070101 0.0078336 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.14605 0.93713 0.91407 0.0013971 0.99199 0.5616 0.0018822 0.42927 1.9185 1.9178 16.0035 144.9766 0.00016816 -85.6519 0.75895
3.863 0.98807 5.5004e-005 3.8182 0.011996 5.0615e-005 0.0011575 0.22574 0.00065925 0.2264 0.2087 0 0.03266 0.0389 0 1.1558 0.36797 0.10898 0.014111 6.8186 0.088063 0.00010966 0.80205 0.0070108 0.0078343 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.14605 0.93727 0.91413 0.0013971 0.99203 0.56175 0.0018822 0.42928 1.919 1.9183 16.0035 144.9767 0.00016806 -85.652 0.75995
3.864 0.98807 5.5004e-005 3.8182 0.011996 5.0628e-005 0.0011576 0.22575 0.00065925 0.22641 0.20871 0 0.032659 0.0389 0 1.1559 0.36801 0.109 0.014113 6.8201 0.088074 0.00010968 0.80204 0.0070115 0.0078351 0.0013862 0.98694 0.9917 2.9891e-006 1.1956e-005 0.14606 0.93742 0.9142 0.0013971 0.99206 0.5619 0.0018822 0.42929 1.9194 1.9187 16.0034 144.9767 0.00016797 -85.6521 0.76095
3.865 0.98807 5.5004e-005 3.8182 0.011996 5.0641e-005 0.0011576 0.22576 0.00065925 0.22641 0.20872 0 0.032659 0.0389 0 1.156 0.36806 0.10902 0.014115 6.8216 0.088084 0.00010969 0.80203 0.0070122 0.0078359 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.14607 0.93756 0.91426 0.001397 0.99209 0.56205 0.0018822 0.4293 1.9198 1.9192 16.0034 144.9767 0.00016787 -85.6522 0.76195
3.866 0.98807 5.5004e-005 3.8182 0.011996 5.0654e-005 0.0011576 0.22577 0.00065925 0.22642 0.20872 0 0.032658 0.0389 0 1.1561 0.36811 0.10903 0.014116 6.8231 0.088095 0.0001097 0.80201 0.0070129 0.0078366 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.14607 0.93771 0.91432 0.001397 0.99213 0.56221 0.0018822 0.42932 1.9203 1.9196 16.0034 144.9767 0.00016777 -85.6523 0.76295
3.867 0.98807 5.5004e-005 3.8182 0.011996 5.0667e-005 0.0011576 0.22577 0.00065925 0.22643 0.20873 0 0.032658 0.0389 0 1.1562 0.36815 0.10905 0.014118 6.8246 0.088105 0.00010972 0.802 0.0070136 0.0078374 0.0013861 0.98695 0.9917 2.9889e-006 1.1956e-005 0.14608 0.93785 0.91438 0.001397 0.99216 0.56236 0.0018821 0.42933 1.9207 1.9201 16.0033 144.9767 0.00016768 -85.6524 0.76395
3.868 0.98807 5.5004e-005 3.8182 0.011996 5.068e-005 0.0011576 0.22578 0.00065925 0.22644 0.20874 0 0.032658 0.0389 0 1.1563 0.3682 0.10907 0.01412 6.8261 0.088116 0.00010973 0.80199 0.0070143 0.0078381 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.14608 0.93799 0.91444 0.001397 0.99219 0.56251 0.0018821 0.42934 1.9212 1.9205 16.0033 144.9768 0.00016758 -85.6525 0.76495
3.869 0.98807 5.5004e-005 3.8182 0.011996 5.0693e-005 0.0011576 0.22579 0.00065925 0.22644 0.20875 0 0.032657 0.0389 0 1.1564 0.36824 0.10908 0.014121 6.8276 0.088126 0.00010975 0.80198 0.007015 0.0078389 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.14609 0.93813 0.9145 0.001397 0.99222 0.56266 0.0018821 0.42935 1.9216 1.9209 16.0033 144.9768 0.00016749 -85.6527 0.76595
3.87 0.98807 5.5003e-005 3.8182 0.011996 5.0706e-005 0.0011576 0.2258 0.00065925 0.22645 0.20875 0 0.032657 0.0389 0 1.1565 0.36829 0.1091 0.014123 6.8291 0.088136 0.00010976 0.80197 0.0070157 0.0078396 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.14609 0.93828 0.91456 0.001397 0.99226 0.56282 0.0018821 0.42937 1.922 1.9214 16.0033 144.9768 0.00016739 -85.6528 0.76695
3.871 0.98807 5.5003e-005 3.8182 0.011996 5.0719e-005 0.0011576 0.2258 0.00065925 0.22646 0.20876 0 0.032657 0.0389 0 1.1566 0.36834 0.10911 0.014125 6.8306 0.088147 0.00010978 0.80196 0.0070164 0.0078404 0.001386 0.98695 0.99171 2.9887e-006 1.1955e-005 0.1461 0.93842 0.91462 0.001397 0.99229 0.56297 0.0018821 0.42938 1.9225 1.9218 16.0032 144.9768 0.0001673 -85.6529 0.76795
3.872 0.98807 5.5003e-005 3.8182 0.011996 5.0732e-005 0.0011576 0.22581 0.00065925 0.22647 0.20877 0 0.032656 0.0389 0 1.1567 0.36838 0.10913 0.014126 6.8321 0.088157 0.00010979 0.80195 0.0070172 0.0078412 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.1461 0.93856 0.91468 0.0013969 0.99232 0.56312 0.001882 0.42939 1.9229 1.9222 16.0032 144.9769 0.00016721 -85.653 0.76895
3.873 0.98807 5.5003e-005 3.8183 0.011996 5.0745e-005 0.0011576 0.22582 0.00065925 0.22647 0.20877 0 0.032656 0.0389 0 1.1568 0.36843 0.10915 0.014128 6.8336 0.088168 0.00010981 0.80194 0.0070179 0.0078419 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.14611 0.9387 0.91474 0.0013969 0.99235 0.56327 0.001882 0.4294 1.9233 1.9227 16.0032 144.9769 0.00016711 -85.6531 0.76995
3.874 0.98807 5.5003e-005 3.8183 0.011996 5.0758e-005 0.0011576 0.22583 0.00065925 0.22648 0.20878 0 0.032655 0.0389 0 1.1569 0.36848 0.10916 0.01413 6.8351 0.088178 0.00010982 0.80193 0.0070186 0.0078427 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.14612 0.93884 0.9148 0.0013969 0.99238 0.56342 0.001882 0.42942 1.9238 1.9231 16.0031 144.9769 0.00016702 -85.6532 0.77095
3.875 0.98807 5.5003e-005 3.8183 0.011996 5.0771e-005 0.0011576 0.22583 0.00065925 0.22649 0.20879 0 0.032655 0.0389 0 1.157 0.36852 0.10918 0.014131 6.8365 0.088188 0.00010983 0.80192 0.0070193 0.0078434 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.14612 0.93898 0.91486 0.0013969 0.99241 0.56358 0.001882 0.42943 1.9242 1.9235 16.0031 144.9769 0.00016693 -85.6533 0.77195
3.876 0.98807 5.5003e-005 3.8183 0.011996 5.0784e-005 0.0011576 0.22584 0.00065925 0.22649 0.20879 0 0.032655 0.0389 0 1.1571 0.36857 0.10919 0.014133 6.838 0.088199 0.00010985 0.80191 0.00702 0.0078442 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.14613 0.93912 0.91492 0.0013969 0.99245 0.56373 0.001882 0.42944 1.9246 1.924 16.0031 144.9769 0.00016683 -85.6534 0.77295
3.877 0.98807 5.5003e-005 3.8183 0.011996 5.0797e-005 0.0011576 0.22585 0.00065925 0.2265 0.2088 0 0.032654 0.0389 0 1.1572 0.36862 0.10921 0.014135 6.8395 0.088209 0.00010986 0.8019 0.0070207 0.0078449 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.14613 0.93926 0.91498 0.0013969 0.99248 0.56388 0.001882 0.42945 1.9251 1.9244 16.0031 144.977 0.00016674 -85.6535 0.77395
3.878 0.98807 5.5003e-005 3.8183 0.011996 5.081e-005 0.0011576 0.22585 0.00065925 0.22651 0.20881 0 0.032654 0.0389 0 1.1573 0.36866 0.10923 0.014136 6.841 0.08822 0.00010988 0.80189 0.0070214 0.0078457 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.14614 0.9394 0.91504 0.0013969 0.99251 0.56403 0.0018819 0.42946 1.9255 1.9248 16.003 144.977 0.00016665 -85.6536 0.77495
3.879 0.98807 5.5003e-005 3.8183 0.011996 5.0823e-005 0.0011576 0.22586 0.00065925 0.22652 0.20882 0 0.032654 0.0389 0 1.1574 0.36871 0.10924 0.014138 6.8425 0.08823 0.00010989 0.80188 0.0070221 0.0078465 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.14614 0.93953 0.91509 0.0013969 0.99254 0.56418 0.0018819 0.42948 1.9259 1.9253 16.003 144.977 0.00016656 -85.6537 0.77595
3.88 0.98807 5.5003e-005 3.8183 0.011996 5.0836e-005 0.0011576 0.22587 0.00065925 0.22652 0.20882 0 0.032653 0.0389 0 1.1575 0.36876 0.10926 0.01414 6.844 0.08824 0.00010991 0.80187 0.0070228 0.0078472 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.14615 0.93967 0.91515 0.0013969 0.99257 0.56434 0.0018819 0.42949 1.9263 1.9257 16.003 144.977 0.00016647 -85.6538 0.77695
3.881 0.98807 5.5003e-005 3.8183 0.011996 5.0849e-005 0.0011576 0.22588 0.00065925 0.22653 0.20883 0 0.032653 0.0389 0 1.1576 0.3688 0.10927 0.014141 6.8455 0.088251 0.00010992 0.80186 0.0070235 0.007848 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.14616 0.93981 0.91521 0.0013968 0.9926 0.56449 0.0018819 0.4295 1.9268 1.9261 16.0029 144.977 0.00016638 -85.6539 0.77795
3.882 0.98807 5.5003e-005 3.8183 0.011996 5.0862e-005 0.0011576 0.22588 0.00065925 0.22654 0.20884 0 0.032652 0.0389 0 1.1577 0.36885 0.10929 0.014143 6.847 0.088261 0.00010994 0.80185 0.0070242 0.0078487 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.14616 0.93994 0.91527 0.0013968 0.99263 0.56464 0.0018819 0.42951 1.9272 1.9266 16.0029 144.9771 0.00016628 -85.654 0.77895
3.883 0.98807 5.5003e-005 3.8183 0.011996 5.0875e-005 0.0011576 0.22589 0.00065925 0.22655 0.20884 0 0.032652 0.0389 0 1.1578 0.3689 0.10931 0.014145 6.8485 0.088272 0.00010995 0.80184 0.0070249 0.0078495 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.14617 0.94008 0.91533 0.0013968 0.99266 0.56479 0.0018819 0.42953 1.9276 1.927 16.0029 144.9771 0.00016619 -85.6541 0.77995
3.884 0.98807 5.5003e-005 3.8183 0.011996 5.0888e-005 0.0011576 0.2259 0.00065925 0.22655 0.20885 0 0.032652 0.0389 0 1.1579 0.36894 0.10932 0.014146 6.85 0.088282 0.00010996 0.80183 0.0070256 0.0078502 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.14617 0.94022 0.91538 0.0013968 0.99269 0.56494 0.0018818 0.42954 1.928 1.9274 16.0029 144.9771 0.0001661 -85.6542 0.78095
3.885 0.98807 5.5002e-005 3.8183 0.011996 5.0901e-005 0.0011576 0.22591 0.00065925 0.22656 0.20886 0 0.032651 0.0389 0 1.158 0.36899 0.10934 0.014148 6.8515 0.088292 0.00010998 0.80182 0.0070263 0.007851 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.14618 0.94035 0.91544 0.0013968 0.99272 0.56509 0.0018818 0.42955 1.9285 1.9278 16.0028 144.9771 0.00016601 -85.6543 0.78195
3.886 0.98807 5.5002e-005 3.8183 0.011995 5.0914e-005 0.0011576 0.22591 0.00065925 0.22657 0.20886 0 0.032651 0.0389 0 1.1581 0.36904 0.10935 0.01415 6.853 0.088303 0.00010999 0.80181 0.007027 0.0078518 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.14618 0.94049 0.9155 0.0013968 0.99274 0.56524 0.0018818 0.42956 1.9289 1.9283 16.0028 144.9771 0.00016592 -85.6544 0.78295
3.887 0.98807 5.5002e-005 3.8183 0.011995 5.0927e-005 0.0011576 0.22592 0.00065925 0.22657 0.20887 0 0.032651 0.0389 0 1.1582 0.36908 0.10937 0.014151 6.8545 0.088313 0.00011001 0.8018 0.0070277 0.0078525 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.14619 0.94062 0.91555 0.0013967 0.99277 0.5654 0.0018818 0.42957 1.9293 1.9287 16.0028 144.9772 0.00016584 -85.6545 0.78395
3.888 0.98807 5.5002e-005 3.8183 0.011995 5.094e-005 0.0011576 0.22593 0.00065925 0.22658 0.20888 0 0.03265 0.0389 0 1.1583 0.36913 0.10939 0.014153 6.856 0.088324 0.00011002 0.80179 0.0070284 0.0078533 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.1462 0.94076 0.91561 0.0013967 0.9928 0.56555 0.0018818 0.42959 1.9297 1.9291 16.0027 144.9772 0.00016575 -85.6546 0.78495
3.889 0.98807 5.5002e-005 3.8183 0.011995 5.0953e-005 0.0011576 0.22593 0.00065925 0.22659 0.20888 0 0.03265 0.0389 0 1.1584 0.36917 0.1094 0.014155 6.8575 0.088334 0.00011004 0.80178 0.0070291 0.007854 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.1462 0.94089 0.91567 0.0013967 0.99283 0.5657 0.0018818 0.4296 1.9302 1.9295 16.0027 144.9772 0.00016566 -85.6547 0.78595
3.89 0.98807 5.5002e-005 3.8183 0.011995 5.0966e-005 0.0011576 0.22594 0.00065925 0.2266 0.20889 0 0.032649 0.0389 0 1.1585 0.36922 0.10942 0.014156 6.8591 0.088344 0.00011005 0.80177 0.0070298 0.0078548 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.14621 0.94102 0.91572 0.0013967 0.99286 0.56585 0.0018818 0.42961 1.9306 1.93 16.0027 144.9772 0.00016557 -85.6548 0.78695
3.891 0.98807 5.5002e-005 3.8183 0.011995 5.0979e-005 0.0011576 0.22595 0.00065925 0.2266 0.2089 0 0.032649 0.0389 0 1.1586 0.36927 0.10943 0.014158 6.8606 0.088355 0.00011006 0.80176 0.0070306 0.0078555 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.14621 0.94116 0.91578 0.0013967 0.99289 0.566 0.0018817 0.42962 1.931 1.9304 16.0027 144.9772 0.00016548 -85.6549 0.78795
3.892 0.98807 5.5002e-005 3.8183 0.011995 5.0992e-005 0.0011576 0.22596 0.00065925 0.22661 0.20891 0 0.032649 0.0389 0 1.1587 0.36931 0.10945 0.01416 6.8621 0.088365 0.00011008 0.80174 0.0070313 0.0078563 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.14622 0.94129 0.91584 0.0013967 0.99291 0.56615 0.0018817 0.42964 1.9314 1.9308 16.0026 144.9773 0.00016539 -85.655 0.78895
3.893 0.98807 5.5002e-005 3.8183 0.011995 5.1005e-005 0.0011576 0.22596 0.00065925 0.22662 0.20891 0 0.032648 0.0389 0 1.1588 0.36936 0.10947 0.014161 6.8636 0.088376 0.00011009 0.80173 0.007032 0.007857 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.14622 0.94142 0.91589 0.0013967 0.99294 0.5663 0.0018817 0.42965 1.9318 1.9312 16.0026 144.9773 0.00016531 -85.6551 0.78995
3.894 0.98807 5.5002e-005 3.8183 0.011995 5.1018e-005 0.0011576 0.22597 0.00065925 0.22663 0.20892 0 0.032648 0.0389 0 1.1589 0.36941 0.10948 0.014163 6.8651 0.088386 0.00011011 0.80172 0.0070327 0.0078578 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.14623 0.94155 0.91595 0.0013967 0.99297 0.56645 0.0018817 0.42966 1.9323 1.9316 16.0026 144.9773 0.00016522 -85.6552 0.79095
3.895 0.98807 5.5002e-005 3.8183 0.011995 5.1031e-005 0.0011576 0.22598 0.00065925 0.22663 0.20893 0 0.032648 0.0389 0 1.159 0.36945 0.1095 0.014165 6.8666 0.088396 0.00011012 0.80171 0.0070334 0.0078586 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.14624 0.94168 0.916 0.0013967 0.993 0.56661 0.0018817 0.42967 1.9327 1.932 16.0025 144.9773 0.00016513 -85.6553 0.79195
3.896 0.98807 5.5002e-005 3.8183 0.011995 5.1044e-005 0.0011576 0.22599 0.00065925 0.22664 0.20893 0 0.032647 0.0389 0 1.1591 0.3695 0.10952 0.014166 6.8681 0.088407 0.00011014 0.8017 0.0070341 0.0078593 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.14624 0.94181 0.91606 0.0013967 0.99302 0.56676 0.0018817 0.42969 1.9331 1.9325 16.0025 144.9773 0.00016505 -85.6554 0.79295
3.897 0.98807 5.5002e-005 3.8183 0.011995 5.1057e-005 0.0011576 0.22599 0.00065925 0.22665 0.20894 0 0.032647 0.0389 0 1.1592 0.36955 0.10953 0.014168 6.8696 0.088417 0.00011015 0.80169 0.0070348 0.0078601 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.14625 0.94194 0.91611 0.0013967 0.99305 0.56691 0.0018816 0.4297 1.9335 1.9329 16.0025 144.9774 0.00016496 -85.6555 0.79395
3.898 0.98807 5.5002e-005 3.8183 0.011995 5.1071e-005 0.0011576 0.226 0.00065925 0.22665 0.20895 0 0.032647 0.0389 0 1.1593 0.36959 0.10955 0.01417 6.8711 0.088427 0.00011016 0.80168 0.0070355 0.0078608 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.14625 0.94207 0.91617 0.0013967 0.99308 0.56706 0.0018816 0.42971 1.9339 1.9333 16.0024 144.9774 0.00016487 -85.6556 0.79495
3.899 0.98807 5.5001e-005 3.8183 0.011995 5.1084e-005 0.0011576 0.22601 0.00065925 0.22666 0.20895 0 0.032646 0.0389 0 1.1594 0.36964 0.10956 0.014171 6.8726 0.088438 0.00011018 0.80167 0.0070362 0.0078616 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.14626 0.9422 0.91622 0.0013966 0.99311 0.56721 0.0018816 0.42972 1.9343 1.9337 16.0024 144.9774 0.00016479 -85.6557 0.79595
3.9 0.98807 5.5001e-005 3.8183 0.011995 5.1097e-005 0.0011576 0.22601 0.00065925 0.22667 0.20896 0 0.032646 0.0389 0 1.1595 0.36969 0.10958 0.014173 6.8741 0.088448 0.00011019 0.80166 0.0070369 0.0078623 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.14626 0.94233 0.91628 0.0013966 0.99313 0.56736 0.0018816 0.42973 1.9347 1.9341 16.0024 144.9774 0.0001647 -85.6558 0.79695
3.901 0.98807 5.5001e-005 3.8183 0.011995 5.111e-005 0.0011576 0.22602 0.00065925 0.22668 0.20897 0 0.032645 0.0389 0 1.1596 0.36973 0.1096 0.014175 6.8756 0.088459 0.00011021 0.80165 0.0070376 0.0078631 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.14627 0.94246 0.91633 0.0013966 0.99316 0.56751 0.0018816 0.42975 1.9351 1.9345 16.0024 144.9774 0.00016462 -85.6558 0.79795
3.902 0.98807 5.5001e-005 3.8183 0.011995 5.1123e-005 0.0011576 0.22603 0.00065925 0.22668 0.20897 0 0.032645 0.0389 0 1.1597 0.36978 0.10961 0.014176 6.8771 0.088469 0.00011022 0.80164 0.0070383 0.0078638 0.0013854 0.98696 0.99171 2.987e-006 1.1948e-005 0.14627 0.94259 0.91639 0.0013966 0.99318 0.56766 0.0018816 0.42976 1.9356 1.9349 16.0023 144.9775 0.00016453 -85.6559 0.79895
3.903 0.98807 5.5001e-005 3.8183 0.011995 5.1136e-005 0.0011576 0.22604 0.00065925 0.22669 0.20898 0 0.032645 0.0389 0 1.1598 0.36983 0.10963 0.014178 6.8786 0.088479 0.00011024 0.80163 0.007039 0.0078646 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.14628 0.94272 0.91644 0.0013966 0.99321 0.56781 0.0018816 0.42977 1.936 1.9354 16.0023 144.9775 0.00016445 -85.656 0.79995
3.904 0.98807 5.5001e-005 3.8183 0.011995 5.1149e-005 0.0011576 0.22604 0.00065925 0.2267 0.20899 0 0.032644 0.0389 0 1.1599 0.36987 0.10964 0.01418 6.8801 0.08849 0.00011025 0.80162 0.0070397 0.0078654 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.14629 0.94285 0.91649 0.0013966 0.99324 0.56796 0.0018815 0.42978 1.9364 1.9358 16.0023 144.9775 0.00016436 -85.6561 0.80095
3.905 0.98807 5.5001e-005 3.8183 0.011995 5.1162e-005 0.0011576 0.22605 0.00065925 0.2267 0.20899 0 0.032644 0.0389 0 1.16 0.36992 0.10966 0.014181 6.8816 0.0885 0.00011027 0.80161 0.0070404 0.0078661 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.14629 0.94297 0.91655 0.0013965 0.99326 0.56811 0.0018815 0.42979 1.9368 1.9362 16.0022 144.9775 0.00016428 -85.6562 0.80195
3.906 0.98807 5.5001e-005 3.8183 0.011995 5.1175e-005 0.0011576 0.22606 0.00065925 0.22671 0.209 0 0.032644 0.0389 0 1.1601 0.36996 0.10968 0.014183 6.8831 0.088511 0.00011028 0.8016 0.0070411 0.0078669 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.1463 0.9431 0.9166 0.0013965 0.99329 0.56826 0.0018815 0.42981 1.9372 1.9366 16.0022 144.9775 0.0001642 -85.6563 0.80295
3.907 0.98807 5.5001e-005 3.8183 0.011995 5.1188e-005 0.0011576 0.22606 0.00065925 0.22672 0.20901 0 0.032643 0.0389 0 1.1602 0.37001 0.10969 0.014185 6.8847 0.088521 0.00011029 0.80159 0.0070418 0.0078676 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.1463 0.94323 0.91665 0.0013965 0.99331 0.56841 0.0018815 0.42982 1.9376 1.937 16.0022 144.9776 0.00016411 -85.6564 0.80395
3.908 0.98807 5.5001e-005 3.8183 0.011995 5.1201e-005 0.0011576 0.22607 0.00065925 0.22673 0.20901 0 0.032643 0.0389 0 1.1603 0.37006 0.10971 0.014186 6.8862 0.088531 0.00011031 0.80158 0.0070425 0.0078684 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.14631 0.94335 0.91671 0.0013965 0.99334 0.56856 0.0018815 0.42983 1.938 1.9374 16.0022 144.9776 0.00016403 -85.6565 0.80495
3.909 0.98807 5.5001e-005 3.8183 0.011995 5.1214e-005 0.0011576 0.22608 0.00065925 0.22673 0.20902 0 0.032643 0.0389 0 1.1604 0.3701 0.10972 0.014188 6.8877 0.088542 0.00011032 0.80157 0.0070432 0.0078691 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.14631 0.94348 0.91676 0.0013965 0.99336 0.56871 0.0018815 0.42984 1.9384 1.9378 16.0021 144.9776 0.00016395 -85.6565 0.80595
3.91 0.98807 5.5001e-005 3.8183 0.011995 5.1227e-005 0.0011577 0.22609 0.00065925 0.22674 0.20903 0 0.032642 0.0389 0 1.1605 0.37015 0.10974 0.01419 6.8892 0.088552 0.00011034 0.80156 0.0070439 0.0078699 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.14632 0.9436 0.91681 0.0013965 0.99339 0.56886 0.0018815 0.42986 1.9388 1.9382 16.0021 144.9776 0.00016387 -85.6566 0.80695
3.911 0.98807 5.5001e-005 3.8183 0.011995 5.124e-005 0.0011577 0.22609 0.00065925 0.22675 0.20903 0 0.032642 0.0389 0 1.1606 0.3702 0.10976 0.014191 6.8907 0.088562 0.00011035 0.80155 0.0070446 0.0078706 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.14633 0.94373 0.91686 0.0013965 0.99341 0.56901 0.0018815 0.42987 1.9392 1.9386 16.0021 144.9776 0.00016378 -85.6567 0.80795
3.912 0.98807 5.5001e-005 3.8183 0.011995 5.1253e-005 0.0011577 0.2261 0.00065925 0.22675 0.20904 0 0.032641 0.0389 0 1.1607 0.37024 0.10977 0.014193 6.8922 0.088573 0.00011037 0.80154 0.0070453 0.0078714 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.14633 0.94385 0.91692 0.0013965 0.99344 0.56916 0.0018814 0.42988 1.9396 1.939 16.002 144.9777 0.0001637 -85.6568 0.80895
3.913 0.98807 5.5e-005 3.8183 0.011995 5.1266e-005 0.0011577 0.22611 0.00065925 0.22676 0.20905 0 0.032641 0.0389 0 1.1608 0.37029 0.10979 0.014195 6.8937 0.088583 0.00011038 0.80153 0.007046 0.0078722 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.14634 0.94398 0.91697 0.0013965 0.99346 0.56931 0.0018814 0.42989 1.94 1.9394 16.002 144.9777 0.00016362 -85.6569 0.80995
3.914 0.98807 5.5e-005 3.8183 0.011995 5.1279e-005 0.0011577 0.22611 0.00065925 0.22677 0.20905 0 0.032641 0.0389 0 1.1609 0.37034 0.1098 0.014196 6.8952 0.088593 0.00011039 0.80152 0.0070467 0.0078729 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.14634 0.9441 0.91702 0.0013965 0.99348 0.56946 0.0018814 0.4299 1.9404 1.9398 16.002 144.9777 0.00016354 -85.6569 0.81095
3.915 0.98807 5.5e-005 3.8183 0.011995 5.1292e-005 0.0011577 0.22612 0.00065925 0.22678 0.20906 0 0.03264 0.0389 0 1.161 0.37038 0.10982 0.014198 6.8967 0.088604 0.00011041 0.80151 0.0070474 0.0078737 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.14635 0.94422 0.91707 0.0013965 0.99351 0.56961 0.0018814 0.42992 1.9408 1.9402 16.0019 144.9777 0.00016346 -85.657 0.81195
3.916 0.98807 5.5e-005 3.8183 0.011995 5.1305e-005 0.0011577 0.22613 0.00065925 0.22678 0.20907 0 0.03264 0.0389 0 1.1611 0.37043 0.10984 0.0142 6.8983 0.088614 0.00011042 0.8015 0.0070482 0.0078744 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.14635 0.94435 0.91712 0.0013964 0.99353 0.56976 0.0018814 0.42993 1.9412 1.9406 16.0019 144.9778 0.00016338 -85.6571 0.81295
3.917 0.98807 5.5e-005 3.8183 0.011995 5.1318e-005 0.0011577 0.22614 0.00065925 0.22679 0.20908 0 0.03264 0.0389 0 1.1612 0.37048 0.10985 0.014202 6.8998 0.088625 0.00011044 0.80149 0.0070489 0.0078752 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.14636 0.94447 0.91717 0.0013964 0.99356 0.56991 0.0018814 0.42994 1.9416 1.941 16.0019 144.9778 0.0001633 -85.6572 0.81395
3.918 0.98807 5.5e-005 3.8183 0.011995 5.1331e-005 0.0011577 0.22614 0.00065925 0.2268 0.20908 0 0.032639 0.0389 0 1.1613 0.37052 0.10987 0.014203 6.9013 0.088635 0.00011045 0.80148 0.0070496 0.0078759 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.14637 0.94459 0.91723 0.0013964 0.99358 0.57006 0.0018814 0.42995 1.942 1.9414 16.0019 144.9778 0.00016322 -85.6573 0.81495
3.919 0.98807 5.5e-005 3.8183 0.011995 5.1344e-005 0.0011577 0.22615 0.00065925 0.2268 0.20909 0 0.032639 0.0389 0 1.1614 0.37057 0.10988 0.014205 6.9028 0.088645 0.00011047 0.80147 0.0070503 0.0078767 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.14637 0.94471 0.91728 0.0013964 0.9936 0.57021 0.0018814 0.42996 1.9424 1.9418 16.0018 144.9778 0.00016314 -85.6573 0.81595
3.92 0.98807 5.5e-005 3.8183 0.011995 5.1357e-005 0.0011577 0.22616 0.00065925 0.22681 0.2091 0 0.032639 0.0389 0 1.1614 0.37062 0.1099 0.014207 6.9043 0.088656 0.00011048 0.80145 0.007051 0.0078774 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.14638 0.94483 0.91733 0.0013964 0.99363 0.57036 0.0018813 0.42998 1.9428 1.9422 16.0018 144.9778 0.00016306 -85.6574 0.81695
3.921 0.98807 5.5e-005 3.8183 0.011995 5.137e-005 0.0011577 0.22616 0.00065925 0.22682 0.2091 0 0.032638 0.0389 0 1.1615 0.37066 0.10992 0.014208 6.9058 0.088666 0.00011049 0.80144 0.0070517 0.0078782 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.14638 0.94495 0.91738 0.0013964 0.99365 0.57051 0.0018813 0.42999 1.9432 1.9426 16.0018 144.9779 0.00016298 -85.6575 0.81795
3.922 0.98807 5.5e-005 3.8183 0.011995 5.1383e-005 0.0011577 0.22617 0.00065925 0.22683 0.20911 0 0.032638 0.0389 0 1.1616 0.37071 0.10993 0.01421 6.9073 0.088676 0.00011051 0.80143 0.0070524 0.0078789 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.14639 0.94507 0.91743 0.0013964 0.99367 0.57066 0.0018813 0.43 1.9436 1.943 16.0017 144.9779 0.0001629 -85.6576 0.81895
3.923 0.98807 5.5e-005 3.8183 0.011995 5.1396e-005 0.0011577 0.22618 0.00065925 0.22683 0.20912 0 0.032637 0.0389 0 1.1617 0.37076 0.10995 0.014212 6.9089 0.088687 0.00011052 0.80142 0.0070531 0.0078797 0.001385 0.98696 0.99171 2.9861e-006 1.1944e-005 0.14639 0.9452 0.91748 0.0013964 0.9937 0.57081 0.0018813 0.43001 1.944 1.9434 16.0017 144.9779 0.00016282 -85.6577 0.81995
3.924 0.98807 5.5e-005 3.8183 0.011995 5.1409e-005 0.0011577 0.22618 0.00065925 0.22684 0.20912 0 0.032637 0.0389 0 1.1618 0.3708 0.10996 0.014213 6.9104 0.088697 0.00011054 0.80141 0.0070538 0.0078805 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.1464 0.94531 0.91753 0.0013964 0.99372 0.57096 0.0018813 0.43003 1.9444 1.9438 16.0017 144.9779 0.00016274 -85.6577 0.82095
3.925 0.98807 5.5e-005 3.8183 0.011995 5.1422e-005 0.0011577 0.22619 0.00065925 0.22685 0.20913 0 0.032637 0.0389 0 1.1619 0.37085 0.10998 0.014215 6.9119 0.088708 0.00011055 0.8014 0.0070545 0.0078812 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.1464 0.94543 0.91758 0.0013964 0.99374 0.57111 0.0018813 0.43004 1.9448 1.9442 16.0016 144.9779 0.00016266 -85.6578 0.82195
3.926 0.98807 5.5e-005 3.8183 0.011995 5.1435e-005 0.0011577 0.2262 0.00065925 0.22685 0.20914 0 0.032636 0.0389 0 1.162 0.37089 0.11 0.014217 6.9134 0.088718 0.00011057 0.80139 0.0070552 0.007882 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.14641 0.94555 0.91763 0.0013964 0.99376 0.57126 0.0018813 0.43005 1.9452 1.9446 16.0016 144.978 0.00016258 -85.6579 0.82295
3.927 0.98807 5.4999e-005 3.8183 0.011995 5.1448e-005 0.0011577 0.22621 0.00065925 0.22686 0.20914 0 0.032636 0.0389 0 1.1621 0.37094 0.11001 0.014218 6.9149 0.088728 0.00011058 0.80138 0.0070559 0.0078827 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.14642 0.94567 0.91768 0.0013964 0.99379 0.57141 0.0018813 0.43006 1.9456 1.945 16.0016 144.978 0.0001625 -85.658 0.82395
3.928 0.98807 5.4999e-005 3.8183 0.011995 5.1461e-005 0.0011577 0.22621 0.00065925 0.22687 0.20915 0 0.032636 0.0389 0 1.1622 0.37099 0.11003 0.01422 6.9164 0.088739 0.0001106 0.80137 0.0070566 0.0078835 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.14642 0.94579 0.91773 0.0013963 0.99381 0.57156 0.0018812 0.43007 1.946 1.9454 16.0016 144.978 0.00016243 -85.658 0.82495
3.929 0.98807 5.4999e-005 3.8183 0.011995 5.1474e-005 0.0011577 0.22622 0.00065925 0.22687 0.20916 0 0.032635 0.0389 0 1.1623 0.37103 0.11005 0.014222 6.918 0.088749 0.00011061 0.80136 0.0070573 0.0078842 0.0013849 0.98696 0.99172 2.9859e-006 1.1943e-005 0.14643 0.94591 0.91778 0.0013963 0.99383 0.57171 0.0018812 0.43009 1.9464 1.9458 16.0015 144.978 0.00016235 -85.6581 0.82595
3.93 0.98807 5.4999e-005 3.8183 0.011995 5.1487e-005 0.0011577 0.22623 0.00065925 0.22688 0.20916 0 0.032635 0.0389 0 1.1624 0.37108 0.11006 0.014223 6.9195 0.088759 0.00011062 0.80135 0.007058 0.007885 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.14643 0.94603 0.91783 0.0013963 0.99385 0.57186 0.0018812 0.4301 1.9467 1.9462 16.0015 144.978 0.00016227 -85.6582 0.82695
3.931 0.98807 5.4999e-005 3.8183 0.011995 5.15e-005 0.0011577 0.22623 0.00065925 0.22689 0.20917 0 0.032635 0.0389 0 1.1625 0.37113 0.11008 0.014225 6.921 0.08877 0.00011064 0.80134 0.0070587 0.0078857 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.14644 0.94614 0.91788 0.0013963 0.99387 0.572 0.0018812 0.43011 1.9471 1.9466 16.0015 144.9781 0.0001622 -85.6582 0.82795
3.932 0.98807 5.4999e-005 3.8183 0.011995 5.1513e-005 0.0011577 0.22624 0.00065925 0.2269 0.20918 0 0.032634 0.0389 0 1.1626 0.37117 0.11009 0.014227 6.9225 0.08878 0.00011065 0.80133 0.0070594 0.0078865 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.14644 0.94626 0.91792 0.0013963 0.99389 0.57215 0.0018812 0.43012 1.9475 1.9469 16.0014 144.9781 0.00016212 -85.6583 0.82895
3.933 0.98807 5.4999e-005 3.8183 0.011995 5.1526e-005 0.0011577 0.22625 0.00065925 0.2269 0.20918 0 0.032634 0.0389 0 1.1627 0.37122 0.11011 0.014228 6.924 0.08879 0.00011067 0.80132 0.0070601 0.0078872 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.14645 0.94638 0.91797 0.0013963 0.99392 0.5723 0.0018812 0.43013 1.9479 1.9473 16.0014 144.9781 0.00016204 -85.6584 0.82995
3.934 0.98807 5.4999e-005 3.8183 0.011995 5.1539e-005 0.0011577 0.22625 0.00065925 0.22691 0.20919 0 0.032634 0.0389 0 1.1628 0.37127 0.11013 0.01423 6.9255 0.088801 0.00011068 0.80131 0.0070608 0.007888 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.14646 0.94649 0.91802 0.0013963 0.99394 0.57245 0.0018812 0.43015 1.9483 1.9477 16.0014 144.9781 0.00016197 -85.6585 0.83095
3.935 0.98807 5.4999e-005 3.8183 0.011995 5.1552e-005 0.0011577 0.22626 0.00065925 0.22692 0.2092 0 0.032633 0.0389 0 1.1629 0.37131 0.11014 0.014232 6.9271 0.088811 0.0001107 0.8013 0.0070615 0.0078888 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.14646 0.94661 0.91807 0.0013963 0.99396 0.5726 0.0018812 0.43016 1.9487 1.9481 16.0013 144.9781 0.00016189 -85.6585 0.83195
3.936 0.98807 5.4999e-005 3.8183 0.011995 5.1565e-005 0.0011577 0.22627 0.00065925 0.22692 0.2092 0 0.032633 0.0389 0 1.163 0.37136 0.11016 0.014233 6.9286 0.088821 0.00011071 0.80129 0.0070622 0.0078895 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.14647 0.94672 0.91812 0.0013963 0.99398 0.57275 0.0018812 0.43017 1.9491 1.9485 16.0013 144.9782 0.00016181 -85.6586 0.83295
3.937 0.98807 5.4999e-005 3.8183 0.011995 5.1578e-005 0.0011577 0.22628 0.00065925 0.22693 0.20921 0 0.032633 0.0389 0 1.1631 0.37141 0.11017 0.014235 6.9301 0.088832 0.00011072 0.80128 0.0070629 0.0078903 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.14647 0.94684 0.91817 0.0013963 0.994 0.5729 0.0018811 0.43018 1.9495 1.9489 16.0013 144.9782 0.00016174 -85.6587 0.83395
3.938 0.98807 5.4999e-005 3.8183 0.011995 5.1591e-005 0.0011577 0.22628 0.00065925 0.22694 0.20922 0 0.032632 0.0389 0 1.1632 0.37145 0.11019 0.014237 6.9316 0.088842 0.00011074 0.80127 0.0070636 0.007891 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.14648 0.94695 0.91821 0.0013962 0.99402 0.57305 0.0018811 0.43019 1.9498 1.9493 16.0013 144.9782 0.00016166 -85.6587 0.83495
3.939 0.98807 5.4999e-005 3.8183 0.011995 5.1604e-005 0.0011577 0.22629 0.00065925 0.22694 0.20922 0 0.032632 0.0389 0 1.1633 0.3715 0.11021 0.014238 6.9331 0.088852 0.00011075 0.80126 0.0070643 0.0078918 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.14648 0.94707 0.91826 0.0013962 0.99404 0.57319 0.0018811 0.43021 1.9502 1.9497 16.0012 144.9782 0.00016159 -85.6588 0.83595
3.94 0.98807 5.4999e-005 3.8183 0.011995 5.1617e-005 0.0011577 0.2263 0.00065925 0.22695 0.20923 0 0.032631 0.0389 0 1.1634 0.37155 0.11022 0.01424 6.9347 0.088863 0.00011077 0.80125 0.007065 0.0078925 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.14649 0.94718 0.91831 0.0013962 0.99406 0.57334 0.0018811 0.43022 1.9506 1.95 16.0012 144.9782 0.00016151 -85.6589 0.83695
3.941 0.98807 5.4998e-005 3.8183 0.011995 5.163e-005 0.0011577 0.2263 0.00065925 0.22696 0.20923 0 0.032631 0.0389 0 1.1635 0.37159 0.11024 0.014242 6.9362 0.088873 0.00011078 0.80124 0.0070657 0.0078933 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.14649 0.9473 0.91836 0.0013962 0.99408 0.57349 0.0018811 0.43023 1.951 1.9504 16.0012 144.9783 0.00016144 -85.6589 0.83795
3.942 0.98807 5.4998e-005 3.8183 0.011995 5.1643e-005 0.0011577 0.22631 0.00065925 0.22697 0.20924 0 0.032631 0.0389 0 1.1636 0.37164 0.11025 0.014243 6.9377 0.088883 0.0001108 0.80123 0.0070664 0.007894 0.0013847 0.98696 0.99172 2.9854e-006 1.1942e-005 0.1465 0.94741 0.9184 0.0013962 0.9941 0.57364 0.0018811 0.43024 1.9514 1.9508 16.0011 144.9783 0.00016137 -85.659 0.83895
3.943 0.98807 5.4998e-005 3.8183 0.011995 5.1656e-005 0.0011577 0.22632 0.00065925 0.22697 0.20925 0 0.03263 0.0389 0 1.1637 0.37169 0.11027 0.014245 6.9392 0.088894 0.00011081 0.80122 0.0070671 0.0078948 0.0013846 0.98696 0.99172 2.9854e-006 1.1941e-005 0.14651 0.94752 0.91845 0.0013962 0.99412 0.57379 0.0018811 0.43025 1.9517 1.9512 16.0011 144.9783 0.00016129 -85.6591 0.83995
3.944 0.98807 5.4998e-005 3.8183 0.011995 5.1669e-005 0.0011577 0.22632 0.00065925 0.22698 0.20925 0 0.03263 0.0389 0 1.1638 0.37173 0.11029 0.014247 6.9408 0.088904 0.00011082 0.80121 0.0070678 0.0078955 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.14651 0.94763 0.9185 0.0013962 0.99414 0.57394 0.0018811 0.43027 1.9521 1.9516 16.0011 144.9783 0.00016122 -85.6591 0.84095
3.945 0.98807 5.4998e-005 3.8183 0.011995 5.1682e-005 0.0011577 0.22633 0.00065925 0.22699 0.20926 0 0.03263 0.0389 0 1.1639 0.37178 0.1103 0.014248 6.9423 0.088915 0.00011084 0.8012 0.0070685 0.0078963 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.14652 0.94775 0.91855 0.0013962 0.99416 0.57409 0.0018811 0.43028 1.9525 1.9519 16.001 144.9783 0.00016114 -85.6592 0.84195
3.946 0.98807 5.4998e-005 3.8183 0.011995 5.1695e-005 0.0011577 0.22634 0.00065925 0.22699 0.20927 0 0.032629 0.0389 0 1.164 0.37183 0.11032 0.01425 6.9438 0.088925 0.00011085 0.80119 0.0070692 0.007897 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.14652 0.94786 0.91859 0.0013962 0.99418 0.57423 0.001881 0.43029 1.9529 1.9523 16.001 144.9784 0.00016107 -85.6593 0.84295
3.947 0.98807 5.4998e-005 3.8183 0.011995 5.1708e-005 0.0011577 0.22635 0.00065925 0.227 0.20927 0 0.032629 0.0389 0 1.1641 0.37187 0.11033 0.014252 6.9453 0.088935 0.00011087 0.80118 0.0070699 0.0078978 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.14653 0.94797 0.91864 0.0013962 0.9942 0.57438 0.001881 0.4303 1.9533 1.9527 16.001 144.9784 0.000161 -85.6593 0.84395
3.948 0.98807 5.4998e-005 3.8183 0.011995 5.1721e-005 0.0011577 0.22635 0.00065925 0.22701 0.20928 0 0.032629 0.0389 0 1.1642 0.37192 0.11035 0.014253 6.9469 0.088946 0.00011088 0.80117 0.0070706 0.0078985 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.14653 0.94808 0.91868 0.0013962 0.99422 0.57453 0.001881 0.43031 1.9536 1.9531 16.0009 144.9784 0.00016093 -85.6594 0.84495
3.949 0.98807 5.4998e-005 3.8183 0.011995 5.1734e-005 0.0011577 0.22636 0.00065925 0.22701 0.20929 0 0.032628 0.0389 0 1.1643 0.37196 0.11037 0.014255 6.9484 0.088956 0.0001109 0.80116 0.0070713 0.0078993 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.14654 0.94819 0.91873 0.0013962 0.99424 0.57468 0.001881 0.43033 1.954 1.9535 16.0009 144.9784 0.00016085 -85.6595 0.84595
3.95 0.98807 5.4998e-005 3.8183 0.011995 5.1747e-005 0.0011577 0.22637 0.00065925 0.22702 0.20929 0 0.032628 0.0389 0 1.1644 0.37201 0.11038 0.014257 6.9499 0.088966 0.00011091 0.80114 0.007072 0.0079001 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.14655 0.9483 0.91878 0.0013962 0.99426 0.57483 0.001881 0.43034 1.9544 1.9538 16.0009 144.9784 0.00016078 -85.6595 0.84695
3.951 0.98807 5.4998e-005 3.8183 0.011994 5.176e-005 0.0011577 0.22637 0.00065925 0.22703 0.2093 0 0.032628 0.0389 0 1.1645 0.37206 0.1104 0.014258 6.9514 0.088977 0.00011092 0.80113 0.0070727 0.0079008 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.14655 0.94841 0.91882 0.0013961 0.99428 0.57497 0.001881 0.43035 1.9548 1.9542 16.0009 144.9785 0.00016071 -85.6596 0.84795
3.952 0.98807 5.4998e-005 3.8183 0.011994 5.1773e-005 0.0011577 0.22638 0.00065925 0.22703 0.20931 0 0.032627 0.0389 0 1.1646 0.3721 0.11041 0.01426 6.953 0.088987 0.00011094 0.80112 0.0070734 0.0079016 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.14656 0.94852 0.91887 0.0013961 0.9943 0.57512 0.001881 0.43036 1.9551 1.9546 16.0008 144.9785 0.00016064 -85.6596 0.84895
3.953 0.98807 5.4998e-005 3.8183 0.011994 5.1786e-005 0.0011577 0.22639 0.00065925 0.22704 0.20931 0 0.032627 0.0389 0 1.1647 0.37215 0.11043 0.014262 6.9545 0.088997 0.00011095 0.80111 0.0070741 0.0079023 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.14656 0.94863 0.91891 0.0013961 0.99431 0.57527 0.001881 0.43037 1.9555 1.955 16.0008 144.9785 0.00016057 -85.6597 0.84995
3.954 0.98807 5.4998e-005 3.8183 0.011994 5.1799e-005 0.0011577 0.22639 0.00065925 0.22705 0.20932 0 0.032627 0.0389 0 1.1648 0.3722 0.11045 0.014263 6.956 0.089008 0.00011097 0.8011 0.0070748 0.0079031 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.14657 0.94874 0.91896 0.0013961 0.99433 0.57542 0.001881 0.43039 1.9559 1.9553 16.0008 144.9785 0.0001605 -85.6598 0.85095
3.955 0.98807 5.4997e-005 3.8183 0.011994 5.1812e-005 0.0011578 0.2264 0.00065925 0.22705 0.20933 0 0.032626 0.0389 0 1.1649 0.37224 0.11046 0.014265 6.9575 0.089018 0.00011098 0.80109 0.0070755 0.0079038 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.14657 0.94885 0.919 0.0013961 0.99435 0.57557 0.001881 0.4304 1.9563 1.9557 16.0007 144.9786 0.00016042 -85.6598 0.85195
3.956 0.98807 5.4997e-005 3.8183 0.011994 5.1825e-005 0.0011578 0.22641 0.00065925 0.22706 0.20933 0 0.032626 0.0389 0 1.165 0.37229 0.11048 0.014266 6.9591 0.089028 0.000111 0.80108 0.0070762 0.0079046 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.14658 0.94896 0.91905 0.0013961 0.99437 0.57571 0.0018809 0.43041 1.9566 1.9561 16.0007 144.9786 0.00016035 -85.6599 0.85295
3.957 0.98807 5.4997e-005 3.8183 0.011994 5.1838e-005 0.0011578 0.22641 0.00065925 0.22707 0.20934 0 0.032625 0.0389 0 1.1651 0.37234 0.11049 0.014268 6.9606 0.089039 0.00011101 0.80107 0.0070769 0.0079053 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.14659 0.94907 0.91909 0.0013961 0.99439 0.57586 0.0018809 0.43042 1.957 1.9565 16.0007 144.9786 0.00016028 -85.6599 0.85395
3.958 0.98807 5.4997e-005 3.8183 0.011994 5.1851e-005 0.0011578 0.22642 0.00065925 0.22708 0.20935 0 0.032625 0.0389 0 1.1652 0.37238 0.11051 0.01427 6.9621 0.089049 0.00011102 0.80106 0.0070776 0.0079061 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.14659 0.94917 0.91914 0.0013961 0.99441 0.57601 0.0018809 0.43043 1.9574 1.9568 16.0006 144.9786 0.00016021 -85.66 0.85495
3.959 0.98807 5.4997e-005 3.8183 0.011994 5.1864e-005 0.0011578 0.22643 0.00065925 0.22708 0.20935 0 0.032625 0.0389 0 1.1653 0.37243 0.11053 0.014271 6.9636 0.089059 0.00011104 0.80105 0.0070783 0.0079068 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.1466 0.94928 0.91918 0.0013961 0.99442 0.57616 0.0018809 0.43045 1.9577 1.9572 16.0006 144.9786 0.00016014 -85.6601 0.85595
3.96 0.98807 5.4997e-005 3.8183 0.011994 5.1877e-005 0.0011578 0.22643 0.00065925 0.22709 0.20936 0 0.032624 0.0389 0 1.1654 0.37248 0.11054 0.014273 6.9652 0.08907 0.00011105 0.80104 0.007079 0.0079076 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.1466 0.94939 0.91923 0.0013961 0.99444 0.5763 0.0018809 0.43046 1.9581 1.9576 16.0006 144.9787 0.00016007 -85.6601 0.85695
3.961 0.98807 5.4997e-005 3.8183 0.011994 5.189e-005 0.0011578 0.22644 0.00065925 0.2271 0.20937 0 0.032624 0.0389 0 1.1655 0.37252 0.11056 0.014275 6.9667 0.08908 0.00011107 0.80103 0.0070797 0.0079083 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.14661 0.9495 0.91927 0.0013961 0.99446 0.57645 0.0018809 0.43047 1.9585 1.9579 16.0005 144.9787 0.00016 -85.6602 0.85795
3.962 0.98807 5.4997e-005 3.8183 0.011994 5.1903e-005 0.0011578 0.22645 0.00065925 0.2271 0.20937 0 0.032624 0.0389 0 1.1656 0.37257 0.11057 0.014276 6.9682 0.08909 0.00011108 0.80102 0.0070804 0.0079091 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.14661 0.9496 0.91932 0.0013961 0.99448 0.5766 0.0018809 0.43048 1.9588 1.9583 16.0005 144.9787 0.00015993 -85.6602 0.85895
3.963 0.98807 5.4997e-005 3.8183 0.011994 5.1916e-005 0.0011578 0.22646 0.00065925 0.22711 0.20938 0 0.032623 0.0389 0 1.1657 0.37262 0.11059 0.014278 6.9698 0.089101 0.0001111 0.80101 0.0070811 0.0079098 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.14662 0.94971 0.91936 0.0013961 0.99449 0.57675 0.0018809 0.43049 1.9592 1.9587 16.0005 144.9787 0.00015986 -85.6603 0.85995
3.964 0.98807 5.4997e-005 3.8183 0.011994 5.1929e-005 0.0011578 0.22646 0.00065925 0.22712 0.20938 0 0.032623 0.0389 0 1.1658 0.37266 0.11061 0.01428 6.9713 0.089111 0.00011111 0.801 0.0070818 0.0079106 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.14662 0.94981 0.9194 0.0013961 0.99451 0.57689 0.0018809 0.4305 1.9596 1.959 16.0004 144.9787 0.0001598 -85.6603 0.86095
3.965 0.98807 5.4997e-005 3.8183 0.011994 5.1942e-005 0.0011578 0.22647 0.00065925 0.22712 0.20939 0 0.032623 0.0389 0 1.1659 0.37271 0.11062 0.014281 6.9728 0.089121 0.00011113 0.80099 0.0070825 0.0079113 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.14663 0.94992 0.91945 0.0013961 0.99453 0.57704 0.0018809 0.43052 1.9599 1.9594 16.0004 144.9788 0.00015973 -85.6604 0.86195
3.966 0.98807 5.4997e-005 3.8183 0.011994 5.1955e-005 0.0011578 0.22648 0.00065925 0.22713 0.2094 0 0.032622 0.0389 0 1.166 0.37276 0.11064 0.014283 6.9744 0.089132 0.00011114 0.80098 0.0070832 0.0079121 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.14664 0.95002 0.91949 0.001396 0.99455 0.57719 0.0018809 0.43053 1.9603 1.9598 16.0004 144.9788 0.00015966 -85.6605 0.86295
3.967 0.98807 5.4997e-005 3.8183 0.011994 5.1968e-005 0.0011578 0.22648 0.00065925 0.22714 0.2094 0 0.032622 0.0389 0 1.1661 0.3728 0.11066 0.014285 6.9759 0.089142 0.00011115 0.80097 0.0070839 0.0079128 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.14664 0.95013 0.91954 0.001396 0.99456 0.57734 0.0018808 0.43054 1.9607 1.9601 16.0004 144.9788 0.00015959 -85.6605 0.86395
3.968 0.98807 5.4997e-005 3.8183 0.011994 5.1981e-005 0.0011578 0.22649 0.00065925 0.22714 0.20941 0 0.032622 0.0389 0 1.1662 0.37285 0.11067 0.014286 6.9774 0.089152 0.00011117 0.80096 0.0070847 0.0079136 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.14665 0.95023 0.91958 0.001396 0.99458 0.57748 0.0018808 0.43055 1.961 1.9605 16.0003 144.9788 0.00015952 -85.6606 0.86495
3.969 0.98807 5.4996e-005 3.8183 0.011994 5.1994e-005 0.0011578 0.2265 0.00065925 0.22715 0.20942 0 0.032621 0.0389 0 1.1663 0.3729 0.11069 0.014288 6.9789 0.089162 0.00011118 0.80095 0.0070854 0.0079144 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.14665 0.95034 0.91962 0.001396 0.9946 0.57763 0.0018808 0.43056 1.9614 1.9609 16.0003 144.9788 0.00015945 -85.6606 0.86595
3.97 0.98807 5.4996e-005 3.8183 0.011994 5.2007e-005 0.0011578 0.2265 0.00065925 0.22716 0.20942 0 0.032621 0.0389 0 1.1664 0.37294 0.1107 0.01429 6.9805 0.089173 0.0001112 0.80094 0.0070861 0.0079151 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14666 0.95044 0.91966 0.001396 0.99461 0.57778 0.0018808 0.43058 1.9618 1.9612 16.0003 144.9789 0.00015939 -85.6607 0.86695
3.971 0.98807 5.4996e-005 3.8183 0.011994 5.202e-005 0.0011578 0.22651 0.00065925 0.22716 0.20943 0 0.032621 0.0389 0 1.1665 0.37299 0.11072 0.014291 6.982 0.089183 0.00011121 0.80093 0.0070868 0.0079159 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14666 0.95054 0.91971 0.001396 0.99463 0.57792 0.0018808 0.43059 1.9621 1.9616 16.0002 144.9789 0.00015932 -85.6607 0.86795
3.972 0.98807 5.4996e-005 3.8183 0.011994 5.2033e-005 0.0011578 0.22652 0.00065925 0.22717 0.20944 0 0.03262 0.0389 0 1.1666 0.37303 0.11074 0.014293 6.9835 0.089193 0.00011123 0.80092 0.0070875 0.0079166 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14667 0.95065 0.91975 0.001396 0.99465 0.57807 0.0018808 0.4306 1.9625 1.962 16.0002 144.9789 0.00015925 -85.6608 0.86895
3.973 0.98807 5.4996e-005 3.8183 0.011994 5.2047e-005 0.0011578 0.22652 0.00065925 0.22718 0.20944 0 0.03262 0.0389 0 1.1667 0.37308 0.11075 0.014295 6.9851 0.089204 0.00011124 0.80091 0.0070882 0.0079174 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.14668 0.95075 0.91979 0.001396 0.99466 0.57822 0.0018808 0.43061 1.9629 1.9623 16.0002 144.9789 0.00015919 -85.6608 0.86995
3.974 0.98807 5.4996e-005 3.8183 0.011994 5.206e-005 0.0011578 0.22653 0.00065925 0.22718 0.20945 0 0.03262 0.0389 0 1.1668 0.37313 0.11077 0.014296 6.9866 0.089214 0.00011125 0.8009 0.0070889 0.0079181 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.14668 0.95085 0.91984 0.001396 0.99468 0.57837 0.0018808 0.43062 1.9632 1.9627 16.0001 144.9789 0.00015912 -85.6609 0.87095
3.975 0.98807 5.4996e-005 3.8183 0.011994 5.2073e-005 0.0011578 0.22654 0.00065925 0.22719 0.20946 0 0.032619 0.0389 0 1.1669 0.37317 0.11078 0.014298 6.9882 0.089224 0.00011127 0.80089 0.0070896 0.0079189 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.14669 0.95095 0.91988 0.001396 0.9947 0.57851 0.0018808 0.43064 1.9636 1.963 16.0001 144.979 0.00015905 -85.6609 0.87195
3.976 0.98807 5.4996e-005 3.8183 0.011994 5.2086e-005 0.0011578 0.22654 0.00065925 0.2272 0.20946 0 0.032619 0.0389 0 1.167 0.37322 0.1108 0.0143 6.9897 0.089235 0.00011128 0.80088 0.0070903 0.0079196 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.14669 0.95106 0.91992 0.001396 0.99471 0.57866 0.0018808 0.43065 1.9639 1.9634 16.0001 144.979 0.00015899 -85.661 0.87295
3.977 0.98807 5.4996e-005 3.8183 0.011994 5.2099e-005 0.0011578 0.22655 0.00065925 0.2272 0.20947 0 0.032619 0.0389 0 1.1671 0.37327 0.11082 0.014301 6.9912 0.089245 0.0001113 0.80087 0.007091 0.0079204 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.1467 0.95116 0.91996 0.001396 0.99473 0.57881 0.0018808 0.43066 1.9643 1.9638 16 144.979 0.00015892 -85.661 0.87395
3.978 0.98807 5.4996e-005 3.8183 0.011994 5.2112e-005 0.0011578 0.22656 0.00065925 0.22721 0.20947 0 0.032618 0.0389 0 1.1672 0.37331 0.11083 0.014303 6.9928 0.089255 0.00011131 0.80086 0.0070917 0.0079211 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.1467 0.95126 0.92 0.001396 0.99474 0.57895 0.0018808 0.43067 1.9646 1.9641 16 144.979 0.00015886 -85.6611 0.87495
3.979 0.98807 5.4996e-005 3.8183 0.011994 5.2125e-005 0.0011578 0.22656 0.00065925 0.22722 0.20948 0 0.032618 0.0389 0 1.1673 0.37336 0.11085 0.014305 6.9943 0.089266 0.00011133 0.80085 0.0070924 0.0079219 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.14671 0.95136 0.92005 0.0013959 0.99476 0.5791 0.0018807 0.43068 1.965 1.9645 16 144.979 0.00015879 -85.6611 0.87595
3.98 0.98807 5.4996e-005 3.8183 0.011994 5.2138e-005 0.0011578 0.22657 0.00065925 0.22722 0.20949 0 0.032618 0.0389 0 1.1674 0.37341 0.11086 0.014306 6.9958 0.089276 0.00011134 0.80084 0.0070931 0.0079226 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.14671 0.95146 0.92009 0.0013959 0.99478 0.57925 0.0018807 0.43069 1.9654 1.9648 15.9999 144.9791 0.00015872 -85.6612 0.87695
3.981 0.98807 5.4996e-005 3.8183 0.011994 5.2151e-005 0.0011578 0.22658 0.00065925 0.22723 0.20949 0 0.032617 0.0389 0 1.1675 0.37345 0.11088 0.014308 6.9974 0.089286 0.00011135 0.80083 0.0070938 0.0079234 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14672 0.95156 0.92013 0.0013959 0.99479 0.57939 0.0018807 0.43071 1.9657 1.9652 15.9999 144.9791 0.00015866 -85.6612 0.87795
3.982 0.98807 5.4996e-005 3.8183 0.011994 5.2164e-005 0.0011578 0.22658 0.00065925 0.22724 0.2095 0 0.032617 0.0389 0 1.1676 0.3735 0.1109 0.01431 6.9989 0.089297 0.00011137 0.80081 0.0070945 0.0079241 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14673 0.95166 0.92017 0.0013959 0.99481 0.57954 0.0018807 0.43072 1.9661 1.9655 15.9999 144.9791 0.00015859 -85.6613 0.87895
3.983 0.98807 5.4995e-005 3.8183 0.011994 5.2177e-005 0.0011578 0.22659 0.00065925 0.22724 0.20951 0 0.032617 0.0389 0 1.1677 0.37355 0.11091 0.014311 7.0004 0.089307 0.00011138 0.8008 0.0070952 0.0079249 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14673 0.95176 0.92021 0.0013959 0.99482 0.57968 0.0018807 0.43073 1.9664 1.9659 15.9999 144.9791 0.00015853 -85.6613 0.87995
3.984 0.98807 5.4995e-005 3.8183 0.011994 5.219e-005 0.0011578 0.2266 0.00065925 0.22725 0.20951 0 0.032616 0.0389 0 1.1678 0.37359 0.11093 0.014313 7.002 0.089317 0.0001114 0.80079 0.0070959 0.0079256 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.14674 0.95186 0.92025 0.0013959 0.99484 0.57983 0.0018807 0.43074 1.9668 1.9663 15.9998 144.9791 0.00015847 -85.6614 0.88095
3.985 0.98807 5.4995e-005 3.8183 0.011994 5.2203e-005 0.0011578 0.2266 0.00065925 0.22726 0.20952 0 0.032616 0.0389 0 1.1679 0.37364 0.11094 0.014315 7.0035 0.089327 0.00011141 0.80078 0.0070965 0.0079264 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.14674 0.95196 0.92029 0.0013959 0.99485 0.57998 0.0018807 0.43075 1.9671 1.9666 15.9998 144.9792 0.0001584 -85.6614 0.88195
3.986 0.98807 5.4995e-005 3.8183 0.011994 5.2216e-005 0.0011578 0.22661 0.00065925 0.22726 0.20953 0 0.032616 0.0389 0 1.168 0.37369 0.11096 0.014316 7.0051 0.089338 0.00011143 0.80077 0.0070972 0.0079271 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.14675 0.95206 0.92033 0.0013959 0.99487 0.58012 0.0018807 0.43077 1.9675 1.967 15.9998 144.9792 0.00015834 -85.6615 0.88295
3.987 0.98807 5.4995e-005 3.8183 0.011994 5.2229e-005 0.0011578 0.22662 0.00065925 0.22727 0.20953 0 0.032615 0.0389 0 1.1681 0.37373 0.11098 0.014318 7.0066 0.089348 0.00011144 0.80076 0.0070979 0.0079279 0.001384 0.98697 0.99172 2.9841e-006 1.1936e-005 0.14675 0.95216 0.92037 0.0013959 0.99488 0.58027 0.0018807 0.43078 1.9678 1.9673 15.9997 144.9792 0.00015827 -85.6615 0.88395
3.988 0.98807 5.4995e-005 3.8183 0.011994 5.2242e-005 0.0011578 0.22662 0.00065925 0.22728 0.20954 0 0.032615 0.0389 0 1.1682 0.37378 0.11099 0.01432 7.0081 0.089358 0.00011145 0.80075 0.0070986 0.0079286 0.001384 0.98697 0.99172 2.9841e-006 1.1936e-005 0.14676 0.95225 0.92041 0.0013959 0.9949 0.58042 0.0018807 0.43079 1.9682 1.9677 15.9997 144.9792 0.00015821 -85.6616 0.88495
3.989 0.98807 5.4995e-005 3.8183 0.011994 5.2255e-005 0.0011578 0.22663 0.00065925 0.22728 0.20954 0 0.032615 0.0389 0 1.1683 0.37383 0.11101 0.014321 7.0097 0.089369 0.00011147 0.80074 0.0070993 0.0079294 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14676 0.95235 0.92045 0.0013959 0.99491 0.58056 0.0018807 0.4308 1.9685 1.968 15.9997 144.9792 0.00015815 -85.6616 0.88595
3.99 0.98807 5.4995e-005 3.8183 0.011994 5.2268e-005 0.0011578 0.22664 0.00065925 0.22729 0.20955 0 0.032614 0.0389 0 1.1684 0.37387 0.11102 0.014323 7.0112 0.089379 0.00011148 0.80073 0.0071 0.0079301 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14677 0.95245 0.9205 0.0013959 0.99493 0.58071 0.0018807 0.43081 1.9689 1.9684 15.9996 144.9793 0.00015808 -85.6617 0.88695
3.991 0.98807 5.4995e-005 3.8183 0.011994 5.2281e-005 0.0011578 0.22664 0.00065925 0.2273 0.20956 0 0.032614 0.0389 0 1.1685 0.37392 0.11104 0.014325 7.0128 0.089389 0.0001115 0.80072 0.0071007 0.0079309 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14678 0.95255 0.92054 0.0013959 0.99494 0.58085 0.0018807 0.43082 1.9692 1.9687 15.9996 144.9793 0.00015802 -85.6617 0.88795
3.992 0.98807 5.4995e-005 3.8183 0.011994 5.2294e-005 0.0011578 0.22665 0.00065925 0.2273 0.20956 0 0.032613 0.0389 0 1.1686 0.37397 0.11106 0.014326 7.0143 0.0894 0.00011151 0.80071 0.0071014 0.0079316 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.14678 0.95264 0.92058 0.0013959 0.99496 0.581 0.0018806 0.43084 1.9696 1.9691 15.9996 144.9793 0.00015796 -85.6618 0.88895
3.993 0.98807 5.4995e-005 3.8183 0.011994 5.2307e-005 0.0011578 0.22666 0.00065925 0.22731 0.20957 0 0.032613 0.0389 0 1.1687 0.37401 0.11107 0.014328 7.0158 0.08941 0.00011153 0.8007 0.0071021 0.0079324 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.14679 0.95274 0.92062 0.0013959 0.99497 0.58115 0.0018806 0.43085 1.9699 1.9694 15.9995 144.9793 0.00015789 -85.6618 0.88995
3.994 0.98807 5.4995e-005 3.8183 0.011994 5.232e-005 0.0011578 0.22666 0.00065925 0.22732 0.20958 0 0.032613 0.0389 0 1.1687 0.37406 0.11109 0.01433 7.0174 0.08942 0.00011154 0.80069 0.0071028 0.0079331 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.14679 0.95284 0.92065 0.0013959 0.99499 0.58129 0.0018806 0.43086 1.9703 1.9698 15.9995 144.9794 0.00015783 -85.6618 0.89095
3.995 0.98807 5.4995e-005 3.8183 0.011994 5.2333e-005 0.0011578 0.22667 0.00065925 0.22732 0.20958 0 0.032612 0.0389 0 1.1688 0.37411 0.1111 0.014331 7.0189 0.08943 0.00011155 0.80068 0.0071035 0.0079339 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.1468 0.95293 0.92069 0.0013959 0.995 0.58144 0.0018806 0.43087 1.9706 1.9701 15.9995 144.9794 0.00015777 -85.6619 0.89195
3.996 0.98807 5.4995e-005 3.8183 0.011994 5.2346e-005 0.0011578 0.22668 0.00065925 0.22733 0.20959 0 0.032612 0.0389 0 1.1689 0.37415 0.11112 0.014333 7.0205 0.089441 0.00011157 0.80067 0.0071042 0.0079346 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.1468 0.95303 0.92073 0.0013958 0.99501 0.58158 0.0018806 0.43088 1.971 1.9705 15.9994 144.9794 0.00015771 -85.6619 0.89295
3.997 0.98807 5.4994e-005 3.8183 0.011994 5.2359e-005 0.0011578 0.22668 0.00065925 0.22734 0.2096 0 0.032612 0.0389 0 1.169 0.3742 0.11114 0.014335 7.022 0.089451 0.00011158 0.80066 0.0071049 0.0079354 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.14681 0.95312 0.92077 0.0013958 0.99503 0.58173 0.0018806 0.43089 1.9713 1.9708 15.9994 144.9794 0.00015765 -85.662 0.89395
3.998 0.98807 5.4994e-005 3.8183 0.011994 5.2372e-005 0.0011578 0.22669 0.00065925 0.22734 0.2096 0 0.032611 0.0389 0 1.1691 0.37424 0.11115 0.014336 7.0235 0.089461 0.0001116 0.80065 0.0071056 0.0079361 0.001384 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14682 0.95322 0.92081 0.0013958 0.99504 0.58187 0.0018806 0.43091 1.9717 1.9712 15.9994 144.9794 0.00015758 -85.662 0.89495
3.999 0.98807 5.4994e-005 3.8183 0.011994 5.2385e-005 0.0011578 0.2267 0.00065925 0.22735 0.20961 0 0.032611 0.0389 0 1.1692 0.37429 0.11117 0.014338 7.0251 0.089472 0.00011161 0.80064 0.0071063 0.0079369 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14682 0.95331 0.92085 0.0013958 0.99506 0.58202 0.0018806 0.43092 1.972 1.9715 15.9993 144.9795 0.00015752 -85.6621 0.89595
4 0.98807 5.4994e-005 3.8183 0.011994 5.2398e-005 0.0011579 0.2267 0.00065925 0.22736 0.20961 0 0.032611 0.0389 0 1.1693 0.37434 0.11118 0.01434 7.0266 0.089482 0.00011163 0.80063 0.007107 0.0079376 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14683 0.95341 0.92089 0.0013958 0.99507 0.58217 0.0018806 0.43093 1.9724 1.9719 15.9993 144.9795 0.00015746 -85.6621 0.89695
4.001 0.98807 5.4994e-005 3.8183 0.011994 5.2411e-005 0.0011579 0.22671 0.00065925 0.22736 0.20962 0 0.03261 0.0389 0 1.1694 0.37438 0.1112 0.014341 7.0282 0.089492 0.00011164 0.80062 0.0071077 0.0079384 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.14683 0.9535 0.92093 0.0013958 0.99508 0.58231 0.0018806 0.43094 1.9727 1.9722 15.9993 144.9795 0.0001574 -85.6622 0.89795
4.002 0.98807 5.4994e-005 3.8183 0.011994 5.2424e-005 0.0011579 0.22672 0.00065925 0.22737 0.20963 0 0.03261 0.0389 0 1.1695 0.37443 0.11122 0.014343 7.0297 0.089503 0.00011165 0.80061 0.0071084 0.0079391 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14684 0.9536 0.92097 0.0013958 0.9951 0.58246 0.0018806 0.43095 1.9731 1.9726 15.9992 144.9795 0.00015734 -85.6622 0.89895
4.003 0.98807 5.4994e-005 3.8183 0.011994 5.2437e-005 0.0011579 0.22672 0.00065925 0.22738 0.20963 0 0.03261 0.0389 0 1.1696 0.37448 0.11123 0.014345 7.0313 0.089513 0.00011167 0.8006 0.0071091 0.0079399 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14684 0.95369 0.92101 0.0013958 0.99511 0.5826 0.0018806 0.43096 1.9734 1.9729 15.9992 144.9795 0.00015728 -85.6622 0.89995
4.004 0.98807 5.4994e-005 3.8183 0.011994 5.245e-005 0.0011579 0.22673 0.00065925 0.22738 0.20964 0 0.032609 0.0389 0 1.1697 0.37452 0.11125 0.014346 7.0328 0.089523 0.00011168 0.80059 0.0071098 0.0079406 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14685 0.95378 0.92104 0.0013958 0.99512 0.58275 0.0018806 0.43098 1.9737 1.9732 15.9992 144.9796 0.00015722 -85.6623 0.90095
4.005 0.98807 5.4994e-005 3.8183 0.011994 5.2463e-005 0.0011579 0.22674 0.00065925 0.22739 0.20965 0 0.032609 0.0389 0 1.1698 0.37457 0.11126 0.014348 7.0344 0.089533 0.0001117 0.80058 0.0071105 0.0079414 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.14685 0.95388 0.92108 0.0013958 0.99514 0.58289 0.0018806 0.43099 1.9741 1.9736 15.9991 144.9796 0.00015716 -85.6623 0.90195
4.006 0.98807 5.4994e-005 3.8183 0.011994 5.2476e-005 0.0011579 0.22674 0.00065925 0.2274 0.20965 0 0.032609 0.0389 0 1.1699 0.37462 0.11128 0.01435 7.0359 0.089544 0.00011171 0.80057 0.0071112 0.0079421 0.0013839 0.98697 0.99172 2.9836e-006 1.1934e-005 0.14686 0.95397 0.92112 0.0013958 0.99515 0.58304 0.0018806 0.431 1.9744 1.9739 15.9991 144.9796 0.0001571 -85.6624 0.90295
4.007 0.98807 5.4994e-005 3.8183 0.011994 5.2489e-005 0.0011579 0.22675 0.00065925 0.2274 0.20966 0 0.032608 0.0389 0 1.17 0.37466 0.1113 0.014351 7.0374 0.089554 0.00011172 0.80056 0.0071119 0.0079429 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.14687 0.95406 0.92116 0.0013958 0.99516 0.58318 0.0018805 0.43101 1.9748 1.9743 15.9991 144.9796 0.00015704 -85.6624 0.90395
4.008 0.98807 5.4994e-005 3.8183 0.011994 5.2502e-005 0.0011579 0.22676 0.00065925 0.22741 0.20966 0 0.032608 0.0389 0 1.1701 0.37471 0.11131 0.014353 7.039 0.089564 0.00011174 0.80055 0.0071126 0.0079436 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.14687 0.95415 0.9212 0.0013958 0.99518 0.58333 0.0018805 0.43102 1.9751 1.9746 15.9991 144.9796 0.00015698 -85.6624 0.90495
4.009 0.98807 5.4994e-005 3.8183 0.011994 5.2515e-005 0.0011579 0.22676 0.00065925 0.22742 0.20967 0 0.032608 0.0389 0 1.1702 0.37476 0.11133 0.014354 7.0405 0.089575 0.00011175 0.80054 0.0071133 0.0079444 0.0013838 0.98698 0.99172 2.9836e-006 1.1934e-005 0.14688 0.95424 0.92123 0.0013958 0.99519 0.58347 0.0018805 0.43103 1.9754 1.9749 15.999 144.9797 0.00015692 -85.6625 0.90595
4.01 0.98807 5.4994e-005 3.8183 0.011994 5.2528e-005 0.0011579 0.22677 0.00065925 0.22742 0.20968 0 0.032607 0.0389 0 1.1703 0.3748 0.11134 0.014356 7.0421 0.089585 0.00011177 0.80053 0.007114 0.0079451 0.0013838 0.98698 0.99172 2.9836e-006 1.1934e-005 0.14688 0.95434 0.92127 0.0013958 0.9952 0.58362 0.0018805 0.43105 1.9758 1.9753 15.999 144.9797 0.00015686 -85.6625 0.90695
4.011 0.98807 5.4994e-005 3.8183 0.011994 5.2541e-005 0.0011579 0.22678 0.00065925 0.22743 0.20968 0 0.032607 0.0389 0 1.1704 0.37485 0.11136 0.014358 7.0436 0.089595 0.00011178 0.80052 0.0071147 0.0079459 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14689 0.95443 0.92131 0.0013958 0.99522 0.58376 0.0018805 0.43106 1.9761 1.9756 15.999 144.9797 0.0001568 -85.6626 0.90795
4.012 0.98807 5.4993e-005 3.8183 0.011994 5.2554e-005 0.0011579 0.22678 0.00065925 0.22744 0.20969 0 0.032607 0.0389 0 1.1705 0.3749 0.11138 0.014359 7.0452 0.089605 0.0001118 0.80051 0.0071154 0.0079466 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14689 0.95452 0.92135 0.0013958 0.99523 0.58391 0.0018805 0.43107 1.9765 1.976 15.9989 144.9797 0.00015674 -85.6626 0.90895
4.013 0.98807 5.4993e-005 3.8183 0.011994 5.2567e-005 0.0011579 0.22679 0.00065925 0.22744 0.2097 0 0.032606 0.0389 0 1.1706 0.37494 0.11139 0.014361 7.0467 0.089616 0.00011181 0.8005 0.0071161 0.0079474 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.1469 0.95461 0.92138 0.0013958 0.99524 0.58405 0.0018805 0.43108 1.9768 1.9763 15.9989 144.9797 0.00015668 -85.6626 0.90995
4.014 0.98807 5.4993e-005 3.8183 0.011994 5.258e-005 0.0011579 0.2268 0.00065925 0.22745 0.2097 0 0.032606 0.0389 0 1.1707 0.37499 0.11141 0.014363 7.0483 0.089626 0.00011182 0.80049 0.0071168 0.0079481 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14691 0.9547 0.92142 0.0013958 0.99525 0.5842 0.0018805 0.43109 1.9771 1.9766 15.9989 144.9798 0.00015663 -85.6627 0.91095
4.015 0.98807 5.4993e-005 3.8183 0.011994 5.2593e-005 0.0011579 0.2268 0.00065925 0.22746 0.20971 0 0.032606 0.0389 0 1.1708 0.37504 0.11142 0.014364 7.0498 0.089636 0.00011184 0.80048 0.0071175 0.0079489 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.14691 0.95479 0.92146 0.0013958 0.99527 0.58434 0.0018805 0.4311 1.9775 1.977 15.9988 144.9798 0.00015657 -85.6627 0.91195
4.016 0.98807 5.4993e-005 3.8183 0.011994 5.2606e-005 0.0011579 0.22681 0.00065925 0.22746 0.20971 0 0.032605 0.0389 0 1.1709 0.37508 0.11144 0.014366 7.0514 0.089647 0.00011185 0.80047 0.0071182 0.0079496 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.14692 0.95488 0.9215 0.0013958 0.99528 0.58449 0.0018805 0.43112 1.9778 1.9773 15.9988 144.9798 0.00015651 -85.6627 0.91295
4.017 0.98807 5.4993e-005 3.8183 0.011993 5.2619e-005 0.0011579 0.22681 0.00065925 0.22747 0.20972 0 0.032605 0.0389 0 1.171 0.37513 0.11146 0.014368 7.0529 0.089657 0.00011187 0.80046 0.0071189 0.0079504 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.14692 0.95497 0.92153 0.0013958 0.99529 0.58463 0.0018805 0.43113 1.9781 1.9777 15.9988 144.9798 0.00015645 -85.6628 0.91395
4.018 0.98807 5.4993e-005 3.8183 0.011993 5.2632e-005 0.0011579 0.22682 0.00065925 0.22748 0.20973 0 0.032605 0.0389 0 1.1711 0.37518 0.11147 0.014369 7.0545 0.089667 0.00011188 0.80044 0.0071196 0.0079511 0.0013838 0.98698 0.99172 2.9834e-006 1.1934e-005 0.14693 0.95506 0.92157 0.0013957 0.9953 0.58478 0.0018805 0.43114 1.9785 1.978 15.9987 144.9798 0.00015639 -85.6628 0.91495
4.019 0.98807 5.4993e-005 3.8183 0.011993 5.2645e-005 0.0011579 0.22683 0.00065925 0.22748 0.20973 0 0.032604 0.0389 0 1.1712 0.37522 0.11149 0.014371 7.056 0.089677 0.0001119 0.80043 0.0071203 0.0079519 0.0013838 0.98698 0.99173 2.9834e-006 1.1933e-005 0.14693 0.95515 0.92161 0.0013957 0.99532 0.58492 0.0018805 0.43115 1.9788 1.9783 15.9987 144.9799 0.00015634 -85.6629 0.91595
4.02 0.98807 5.4993e-005 3.8183 0.011993 5.2658e-005 0.0011579 0.22683 0.00065925 0.22749 0.20974 0 0.032604 0.0389 0 1.1713 0.37527 0.11151 0.014373 7.0576 0.089688 0.00011191 0.80042 0.007121 0.0079526 0.0013837 0.98698 0.99173 2.9834e-006 1.1933e-005 0.14694 0.95524 0.92164 0.0013957 0.99533 0.58507 0.0018805 0.43116 1.9791 1.9787 15.9987 144.9799 0.00015628 -85.6629 0.91695
4.021 0.98807 5.4993e-005 3.8183 0.011993 5.2671e-005 0.0011579 0.22684 0.00065925 0.2275 0.20974 0 0.032604 0.0389 0 1.1714 0.37532 0.11152 0.014374 7.0591 0.089698 0.00011192 0.80041 0.0071217 0.0079534 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14694 0.95532 0.92168 0.0013957 0.99534 0.58521 0.0018805 0.43117 1.9795 1.979 15.9986 144.9799 0.00015622 -85.6629 0.91795
4.022 0.98807 5.4993e-005 3.8183 0.011993 5.2684e-005 0.0011579 0.22685 0.00065925 0.2275 0.20975 0 0.032603 0.0389 0 1.1715 0.37536 0.11154 0.014376 7.0607 0.089708 0.00011194 0.8004 0.0071224 0.0079541 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14695 0.95541 0.92171 0.0013957 0.99535 0.58535 0.0018805 0.43119 1.9798 1.9793 15.9986 144.9799 0.00015617 -85.663 0.91895
4.023 0.98807 5.4993e-005 3.8183 0.011993 5.2697e-005 0.0011579 0.22685 0.00065925 0.22751 0.20976 0 0.032603 0.0389 0 1.1716 0.37541 0.11155 0.014378 7.0622 0.089718 0.00011195 0.80039 0.0071231 0.0079549 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14696 0.9555 0.92175 0.0013957 0.99536 0.5855 0.0018804 0.4312 1.9801 1.9797 15.9986 144.9799 0.00015611 -85.663 0.91995
4.024 0.98807 5.4993e-005 3.8183 0.011993 5.271e-005 0.0011579 0.22686 0.00065925 0.22751 0.20976 0 0.032603 0.0389 0 1.1717 0.37545 0.11157 0.014379 7.0638 0.089729 0.00011197 0.80038 0.0071238 0.0079556 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14696 0.95559 0.92179 0.0013957 0.99537 0.58564 0.0018804 0.43121 1.9805 1.98 15.9985 144.98 0.00015605 -85.663 0.92095
4.025 0.98807 5.4993e-005 3.8183 0.011993 5.2723e-005 0.0011579 0.22687 0.00065925 0.22752 0.20977 0 0.032602 0.0389 0 1.1718 0.3755 0.11159 0.014381 7.0653 0.089739 0.00011198 0.80037 0.0071245 0.0079564 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14697 0.95568 0.92182 0.0013957 0.99539 0.58579 0.0018804 0.43122 1.9808 1.9803 15.9985 144.98 0.000156 -85.6631 0.92195
4.026 0.98807 5.4992e-005 3.8183 0.011993 5.2736e-005 0.0011579 0.22687 0.00065925 0.22753 0.20978 0 0.032602 0.0389 0 1.1719 0.37555 0.1116 0.014383 7.0669 0.089749 0.000112 0.80036 0.0071252 0.0079571 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.14697 0.95576 0.92186 0.0013957 0.9954 0.58593 0.0018804 0.43123 1.9811 1.9807 15.9985 144.98 0.00015594 -85.6631 0.92295
4.027 0.98807 5.4992e-005 3.8183 0.011993 5.2749e-005 0.0011579 0.22688 0.00065925 0.22753 0.20978 0 0.032602 0.0389 0 1.172 0.37559 0.11162 0.014384 7.0685 0.08976 0.00011201 0.80035 0.0071259 0.0079579 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14698 0.95585 0.92189 0.0013957 0.99541 0.58608 0.0018804 0.43124 1.9815 1.981 15.9984 144.98 0.00015588 -85.6631 0.92395
4.028 0.98807 5.4992e-005 3.8183 0.011993 5.2762e-005 0.0011579 0.22689 0.00065925 0.22754 0.20979 0 0.032602 0.0389 0 1.1721 0.37564 0.11163 0.014386 7.07 0.08977 0.00011202 0.80034 0.0071266 0.0079586 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14698 0.95594 0.92193 0.0013957 0.99542 0.58622 0.0018804 0.43126 1.9818 1.9813 15.9984 144.9801 0.00015583 -85.6632 0.92495
4.029 0.98807 5.4992e-005 3.8183 0.011993 5.2775e-005 0.0011579 0.22689 0.00065925 0.22755 0.20979 0 0.032601 0.0389 0 1.1722 0.37569 0.11165 0.014388 7.0716 0.08978 0.00011204 0.80033 0.0071273 0.0079594 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14699 0.95602 0.92196 0.0013957 0.99543 0.58636 0.0018804 0.43127 1.9821 1.9816 15.9984 144.9801 0.00015577 -85.6632 0.92595
4.03 0.98807 5.4992e-005 3.8183 0.011993 5.2788e-005 0.0011579 0.2269 0.00065925 0.22755 0.2098 0 0.032601 0.0389 0 1.1723 0.37573 0.11167 0.014389 7.0731 0.08979 0.00011205 0.80032 0.007128 0.0079601 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.14699 0.95611 0.922 0.0013957 0.99544 0.58651 0.0018804 0.43128 1.9825 1.982 15.9983 144.9801 0.00015572 -85.6632 0.92695
4.031 0.98807 5.4992e-005 3.8183 0.011993 5.2801e-005 0.0011579 0.22691 0.00065925 0.22756 0.20981 0 0.032601 0.0389 0 1.1724 0.37578 0.11168 0.014391 7.0747 0.089801 0.00011207 0.80031 0.0071287 0.0079609 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.147 0.95619 0.92204 0.0013957 0.99546 0.58665 0.0018804 0.43129 1.9828 1.9823 15.9983 144.9801 0.00015566 -85.6633 0.92795
4.032 0.98807 5.4992e-005 3.8183 0.011993 5.2814e-005 0.0011579 0.22691 0.00065925 0.22757 0.20981 0 0.0326 0.0389 0 1.1725 0.37583 0.1117 0.014393 7.0762 0.089811 0.00011208 0.8003 0.0071294 0.0079616 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14701 0.95628 0.92207 0.0013957 0.99547 0.5868 0.0018804 0.4313 1.9831 1.9826 15.9983 144.9801 0.00015561 -85.6633 0.92895
4.033 0.98807 5.4992e-005 3.8183 0.011993 5.2827e-005 0.0011579 0.22692 0.00065925 0.22757 0.20982 0 0.0326 0.0389 0 1.1726 0.37587 0.11171 0.014394 7.0778 0.089821 0.0001121 0.80029 0.0071301 0.0079624 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14701 0.95636 0.92211 0.0013957 0.99548 0.58694 0.0018804 0.43131 1.9834 1.983 15.9982 144.9802 0.00015555 -85.6633 0.92995
4.034 0.98807 5.4992e-005 3.8183 0.011993 5.284e-005 0.0011579 0.22692 0.00065925 0.22758 0.20982 0 0.0326 0.0389 0 1.1727 0.37592 0.11173 0.014396 7.0793 0.089831 0.00011211 0.80028 0.0071308 0.0079631 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14702 0.95645 0.92214 0.0013957 0.99549 0.58708 0.0018804 0.43132 1.9838 1.9833 15.9982 144.9802 0.0001555 -85.6634 0.93095
4.035 0.98807 5.4992e-005 3.8183 0.011993 5.2853e-005 0.0011579 0.22693 0.00065925 0.22759 0.20983 0 0.032599 0.0389 0 1.1728 0.37597 0.11175 0.014398 7.0809 0.089842 0.00011212 0.80027 0.0071315 0.0079639 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14702 0.95653 0.92217 0.0013957 0.9955 0.58723 0.0018804 0.43134 1.9841 1.9836 15.9982 144.9802 0.00015544 -85.6634 0.93195
4.036 0.98807 5.4992e-005 3.8183 0.011993 5.2866e-005 0.0011579 0.22694 0.00065926 0.22759 0.20984 0 0.032599 0.0389 0 1.1729 0.37601 0.11176 0.014399 7.0825 0.089852 0.00011214 0.80026 0.0071321 0.0079646 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14703 0.95662 0.92221 0.0013957 0.99551 0.58737 0.0018804 0.43135 1.9844 1.9839 15.9981 144.9802 0.00015539 -85.6634 0.93295
4.037 0.98807 5.4992e-005 3.8183 0.011993 5.2879e-005 0.0011579 0.22694 0.00065926 0.2276 0.20984 0 0.032599 0.0389 0 1.173 0.37606 0.11178 0.014401 7.084 0.089862 0.00011215 0.80025 0.0071328 0.0079654 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.14703 0.9567 0.92224 0.0013957 0.99552 0.58751 0.0018804 0.43136 1.9847 1.9843 15.9981 144.9802 0.00015533 -85.6635 0.93395
4.038 0.98807 5.4992e-005 3.8183 0.011993 5.2892e-005 0.0011579 0.22695 0.00065926 0.22761 0.20985 0 0.032598 0.0389 0 1.1731 0.37611 0.11179 0.014402 7.0856 0.089872 0.00011217 0.80024 0.0071335 0.0079661 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14704 0.95679 0.92228 0.0013957 0.99553 0.58766 0.0018804 0.43137 1.9851 1.9846 15.9981 144.9803 0.00015528 -85.6635 0.93495
4.039 0.98807 5.4992e-005 3.8183 0.011993 5.2905e-005 0.0011579 0.22696 0.00065926 0.22761 0.20985 0 0.032598 0.0389 0 1.1732 0.37615 0.11181 0.014404 7.0871 0.089883 0.00011218 0.80023 0.0071342 0.0079669 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14704 0.95687 0.92231 0.0013957 0.99554 0.5878 0.0018804 0.43138 1.9854 1.9849 15.998 144.9803 0.00015523 -85.6635 0.93595
4.04 0.98807 5.4991e-005 3.8183 0.011993 5.2918e-005 0.0011579 0.22696 0.00065926 0.22762 0.20986 0 0.032598 0.0389 0 1.1733 0.3762 0.11183 0.014406 7.0887 0.089893 0.0001122 0.80022 0.0071349 0.0079676 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14705 0.95695 0.92235 0.0013957 0.99555 0.58794 0.0018804 0.43139 1.9857 1.9852 15.998 144.9803 0.00015517 -85.6636 0.93695
4.041 0.98807 5.4991e-005 3.8183 0.011993 5.2931e-005 0.0011579 0.22697 0.00065926 0.22762 0.20987 0 0.032597 0.0389 0 1.1734 0.37625 0.11184 0.014407 7.0902 0.089903 0.00011221 0.80021 0.0071356 0.0079684 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14706 0.95704 0.92238 0.0013957 0.99556 0.58809 0.0018804 0.43141 1.986 1.9856 15.998 144.9803 0.00015512 -85.6636 0.93795
4.042 0.98807 5.4991e-005 3.8183 0.011993 5.2944e-005 0.0011579 0.22698 0.00065926 0.22763 0.20987 0 0.032597 0.0389 0 1.1735 0.37629 0.11186 0.014409 7.0918 0.089913 0.00011222 0.8002 0.0071363 0.0079691 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14706 0.95712 0.92241 0.0013957 0.99557 0.58823 0.0018803 0.43142 1.9864 1.9859 15.9979 144.9803 0.00015507 -85.6636 0.93895
4.043 0.98807 5.4991e-005 3.8183 0.011993 5.2957e-005 0.0011579 0.22698 0.00065926 0.22764 0.20988 0 0.032597 0.0389 0 1.1736 0.37634 0.11187 0.014411 7.0934 0.089924 0.00011224 0.80019 0.007137 0.0079698 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.14707 0.9572 0.92245 0.0013957 0.99558 0.58837 0.0018803 0.43143 1.9867 1.9862 15.9979 144.9804 0.00015501 -85.6637 0.93995
4.044 0.98807 5.4991e-005 3.8183 0.011993 5.297e-005 0.001158 0.22699 0.00065926 0.22764 0.20989 0 0.032596 0.0389 0 1.1737 0.37639 0.11189 0.014412 7.0949 0.089934 0.00011225 0.80018 0.0071377 0.0079706 0.0013836 0.98698 0.99173 2.9829e-006 1.1932e-005 0.14707 0.95728 0.92248 0.0013957 0.99559 0.58852 0.0018803 0.43144 1.987 1.9865 15.9979 144.9804 0.00015496 -85.6637 0.94095
4.045 0.98807 5.4991e-005 3.8183 0.011993 5.2983e-005 0.001158 0.227 0.00065926 0.22765 0.20989 0 0.032596 0.0389 0 1.1738 0.37643 0.11191 0.014414 7.0965 0.089944 0.00011227 0.80017 0.0071384 0.0079713 0.0013836 0.98698 0.99173 2.9829e-006 1.1932e-005 0.14708 0.95737 0.92252 0.0013956 0.99561 0.58866 0.0018803 0.43145 1.9873 1.9869 15.9978 144.9804 0.00015491 -85.6637 0.94195
4.046 0.98807 5.4991e-005 3.8183 0.011993 5.2996e-005 0.001158 0.227 0.00065926 0.22766 0.2099 0 0.032596 0.0389 0 1.1739 0.37648 0.11192 0.014416 7.098 0.089954 0.00011228 0.80016 0.0071391 0.0079721 0.0013836 0.98698 0.99173 2.9829e-006 1.1932e-005 0.14708 0.95745 0.92255 0.0013956 0.99562 0.5888 0.0018803 0.43146 1.9876 1.9872 15.9978 144.9804 0.00015486 -85.6637 0.94295
4.047 0.98807 5.4991e-005 3.8183 0.011993 5.3009e-005 0.001158 0.22701 0.00065926 0.22766 0.2099 0 0.032595 0.0389 0 1.174 0.37653 0.11194 0.014417 7.0996 0.089965 0.00011229 0.80015 0.0071398 0.0079728 0.0013835 0.98698 0.99173 2.9829e-006 1.1932e-005 0.14709 0.95753 0.92258 0.0013956 0.99563 0.58895 0.0018803 0.43147 1.988 1.9875 15.9978 144.9804 0.0001548 -85.6638 0.94395
4.048 0.98807 5.4991e-005 3.8183 0.011993 5.3022e-005 0.001158 0.22701 0.00065926 0.22767 0.20991 0 0.032595 0.0389 0 1.1741 0.37657 0.11195 0.014419 7.1012 0.089975 0.00011231 0.80014 0.0071405 0.0079736 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.1471 0.95761 0.92262 0.0013956 0.99564 0.58909 0.0018803 0.43149 1.9883 1.9878 15.9977 144.9805 0.00015475 -85.6638 0.94495
4.049 0.98807 5.4991e-005 3.8183 0.011993 5.3035e-005 0.001158 0.22702 0.00065926 0.22768 0.20992 0 0.032595 0.0389 0 1.1742 0.37662 0.11197 0.014421 7.1027 0.089985 0.00011232 0.80013 0.0071412 0.0079743 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.1471 0.95769 0.92265 0.0013956 0.99565 0.58923 0.0018803 0.4315 1.9886 1.9881 15.9977 144.9805 0.0001547 -85.6638 0.94595
4.05 0.98807 5.4991e-005 3.8183 0.011993 5.3048e-005 0.001158 0.22703 0.00065926 0.22768 0.20992 0 0.032594 0.0389 0 1.1743 0.37667 0.11199 0.014422 7.1043 0.089995 0.00011234 0.80012 0.0071419 0.0079751 0.0013835 0.98698 0.99173 2.9829e-006 1.1931e-005 0.14711 0.95777 0.92268 0.0013956 0.99566 0.58938 0.0018803 0.43151 1.9889 1.9885 15.9977 144.9805 0.00015465 -85.6639 0.94695
4.051 0.98807 5.4991e-005 3.8183 0.011993 5.3061e-005 0.001158 0.22703 0.00065926 0.22769 0.20993 0 0.032594 0.0389 0 1.1744 0.37671 0.112 0.014424 7.1059 0.090006 0.00011235 0.80011 0.0071426 0.0079758 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14711 0.95785 0.92271 0.0013956 0.99567 0.58952 0.0018803 0.43152 1.9892 1.9888 15.9976 144.9805 0.00015459 -85.6639 0.94795
4.052 0.98807 5.4991e-005 3.8183 0.011993 5.3074e-005 0.001158 0.22704 0.00065926 0.22769 0.20993 0 0.032594 0.0389 0 1.1745 0.37676 0.11202 0.014426 7.1074 0.090016 0.00011237 0.8001 0.0071433 0.0079766 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14712 0.95793 0.92275 0.0013956 0.99568 0.58966 0.0018803 0.43153 1.9895 1.9891 15.9976 144.9805 0.00015454 -85.6639 0.94895
4.053 0.98807 5.4991e-005 3.8183 0.011993 5.3087e-005 0.001158 0.22705 0.00065926 0.2277 0.20994 0 0.032593 0.0389 0 1.1746 0.3768 0.11203 0.014427 7.109 0.090026 0.00011238 0.80009 0.007144 0.0079773 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14712 0.95801 0.92278 0.0013956 0.99568 0.58981 0.0018803 0.43154 1.9899 1.9894 15.9976 144.9806 0.00015449 -85.6639 0.94995
4.054 0.98807 5.499e-005 3.8183 0.011993 5.31e-005 0.001158 0.22705 0.00065926 0.22771 0.20995 0 0.032593 0.0389 0 1.1747 0.37685 0.11205 0.014429 7.1105 0.090036 0.00011239 0.80008 0.0071447 0.0079781 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14713 0.95809 0.92281 0.0013956 0.99569 0.58995 0.0018803 0.43155 1.9902 1.9897 15.9975 144.9806 0.00015444 -85.664 0.95095
4.055 0.98807 5.499e-005 3.8183 0.011993 5.3113e-005 0.001158 0.22706 0.00065926 0.22771 0.20995 0 0.032593 0.0389 0 1.1748 0.3769 0.11207 0.014431 7.1121 0.090047 0.00011241 0.80007 0.0071454 0.0079788 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14713 0.95817 0.92284 0.0013956 0.9957 0.59009 0.0018803 0.43157 1.9905 1.99 15.9975 144.9806 0.00015439 -85.664 0.95195
4.056 0.98807 5.499e-005 3.8183 0.011993 5.3126e-005 0.001158 0.22706 0.00065926 0.22772 0.20996 0 0.032592 0.0389 0 1.1749 0.37694 0.11208 0.014432 7.1137 0.090057 0.00011242 0.80006 0.0071461 0.0079796 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14714 0.95825 0.92288 0.0013956 0.99571 0.59023 0.0018803 0.43158 1.9908 1.9904 15.9975 144.9806 0.00015434 -85.664 0.95295
4.057 0.98807 5.499e-005 3.8183 0.011993 5.3139e-005 0.001158 0.22707 0.00065926 0.22773 0.20996 0 0.032592 0.0389 0 1.175 0.37699 0.1121 0.014434 7.1152 0.090067 0.00011244 0.80005 0.0071468 0.0079803 0.0013835 0.98698 0.99173 2.9828e-006 1.1931e-005 0.14715 0.95833 0.92291 0.0013956 0.99572 0.59038 0.0018803 0.43159 1.9911 1.9907 15.9974 144.9806 0.00015429 -85.6641 0.95395
4.058 0.98807 5.499e-005 3.8183 0.011993 5.3152e-005 0.001158 0.22708 0.00065926 0.22773 0.20997 0 0.032592 0.0389 0 1.1751 0.37704 0.11211 0.014435 7.1168 0.090077 0.00011245 0.80004 0.0071475 0.0079811 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14715 0.95841 0.92294 0.0013956 0.99573 0.59052 0.0018803 0.4316 1.9914 1.991 15.9974 144.9807 0.00015424 -85.6641 0.95495
4.059 0.98807 5.499e-005 3.8183 0.011993 5.3165e-005 0.001158 0.22708 0.00065926 0.22774 0.20998 0 0.032591 0.0389 0 1.1752 0.37708 0.11213 0.014437 7.1184 0.090088 0.00011247 0.80002 0.0071482 0.0079818 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14716 0.95849 0.92297 0.0013956 0.99574 0.59066 0.0018803 0.43161 1.9918 1.9913 15.9974 144.9807 0.00015419 -85.6641 0.95595
4.06 0.98807 5.499e-005 3.8183 0.011993 5.3178e-005 0.001158 0.22709 0.00065926 0.22774 0.20998 0 0.032591 0.0389 0 1.1753 0.37713 0.11215 0.014439 7.1199 0.090098 0.00011248 0.80001 0.0071488 0.0079826 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14716 0.95857 0.92301 0.0013956 0.99575 0.5908 0.0018803 0.43162 1.9921 1.9916 15.9973 144.9807 0.00015414 -85.6641 0.95695
4.061 0.98807 5.499e-005 3.8183 0.011993 5.3191e-005 0.001158 0.2271 0.00065926 0.22775 0.20999 0 0.032591 0.0389 0 1.1754 0.37718 0.11216 0.01444 7.1215 0.090108 0.00011249 0.8 0.0071495 0.0079833 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14717 0.95865 0.92304 0.0013956 0.99576 0.59095 0.0018803 0.43163 1.9924 1.9919 15.9973 144.9807 0.00015409 -85.6642 0.95795
4.062 0.98807 5.499e-005 3.8183 0.011993 5.3204e-005 0.001158 0.2271 0.00065926 0.22776 0.20999 0 0.032591 0.0389 0 1.1754 0.37722 0.11218 0.014442 7.1231 0.090118 0.00011251 0.79999 0.0071502 0.007984 0.0013835 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14717 0.95872 0.92307 0.0013956 0.99577 0.59109 0.0018803 0.43165 1.9927 1.9922 15.9973 144.9807 0.00015404 -85.6642 0.95895
4.063 0.98807 5.499e-005 3.8183 0.011993 5.3217e-005 0.001158 0.22711 0.00065926 0.22776 0.21 0 0.03259 0.0389 0 1.1755 0.37727 0.11219 0.014444 7.1246 0.090129 0.00011252 0.79998 0.0071509 0.0079848 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14718 0.9588 0.9231 0.0013956 0.99578 0.59123 0.0018803 0.43166 1.993 1.9926 15.9972 144.9808 0.00015399 -85.6642 0.95995
4.064 0.98807 5.499e-005 3.8183 0.011993 5.323e-005 0.001158 0.22712 0.00065926 0.22777 0.21 0 0.03259 0.0389 0 1.1756 0.37732 0.11221 0.014445 7.1262 0.090139 0.00011254 0.79997 0.0071516 0.0079855 0.0013834 0.98698 0.99173 2.9827e-006 1.1931e-005 0.14718 0.95888 0.92313 0.0013956 0.99579 0.59137 0.0018803 0.43167 1.9933 1.9929 15.9972 144.9808 0.00015394 -85.6642 0.96095
4.065 0.98807 5.499e-005 3.8183 0.011993 5.3243e-005 0.001158 0.22712 0.00065926 0.22778 0.21001 0 0.03259 0.0389 0 1.1757 0.37736 0.11223 0.014447 7.1278 0.090149 0.00011255 0.79996 0.0071523 0.0079863 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14719 0.95895 0.92316 0.0013956 0.9958 0.59152 0.0018802 0.43168 1.9936 1.9932 15.9972 144.9808 0.00015389 -85.6643 0.96195
4.066 0.98807 5.499e-005 3.8183 0.011993 5.3256e-005 0.001158 0.22713 0.00065926 0.22778 0.21002 0 0.032589 0.0389 0 1.1758 0.37741 0.11224 0.014449 7.1293 0.090159 0.00011256 0.79995 0.007153 0.007987 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.1472 0.95903 0.9232 0.0013956 0.99581 0.59166 0.0018802 0.43169 1.9939 1.9935 15.9971 144.9808 0.00015384 -85.6643 0.96295
4.067 0.98807 5.499e-005 3.8183 0.011993 5.3269e-005 0.001158 0.22713 0.00065926 0.22779 0.21002 0 0.032589 0.0389 0 1.1759 0.37746 0.11226 0.01445 7.1309 0.090169 0.00011258 0.79994 0.0071537 0.0079878 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.1472 0.95911 0.92323 0.0013956 0.99581 0.5918 0.0018802 0.4317 1.9943 1.9938 15.9971 144.9809 0.00015379 -85.6643 0.96395
4.068 0.98807 5.4989e-005 3.8183 0.011993 5.3282e-005 0.001158 0.22714 0.00065926 0.22779 0.21003 0 0.032589 0.0389 0 1.176 0.3775 0.11227 0.014452 7.1325 0.09018 0.00011259 0.79993 0.0071544 0.0079885 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14721 0.95918 0.92326 0.0013956 0.99582 0.59194 0.0018802 0.43171 1.9946 1.9941 15.9971 144.9809 0.00015374 -85.6643 0.96495
4.069 0.98807 5.4989e-005 3.8183 0.011993 5.3295e-005 0.001158 0.22715 0.00065926 0.2278 0.21003 0 0.032588 0.0389 0 1.1761 0.37755 0.11229 0.014454 7.134 0.09019 0.00011261 0.79992 0.0071551 0.0079893 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14721 0.95926 0.92329 0.0013956 0.99583 0.59208 0.0018802 0.43172 1.9949 1.9944 15.997 144.9809 0.00015369 -85.6644 0.96595
4.07 0.98807 5.4989e-005 3.8183 0.011993 5.3308e-005 0.001158 0.22715 0.00065926 0.22781 0.21004 0 0.032588 0.0389 0 1.1762 0.3776 0.11231 0.014455 7.1356 0.0902 0.00011262 0.79991 0.0071558 0.00799 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14722 0.95934 0.92332 0.0013956 0.99584 0.59223 0.0018802 0.43174 1.9952 1.9947 15.997 144.9809 0.00015364 -85.6644 0.96695
4.071 0.98807 5.4989e-005 3.8183 0.011993 5.3321e-005 0.001158 0.22716 0.00065926 0.22781 0.21005 0 0.032588 0.0389 0 1.1763 0.37764 0.11232 0.014457 7.1372 0.09021 0.00011264 0.7999 0.0071565 0.0079908 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14722 0.95941 0.92335 0.0013956 0.99585 0.59237 0.0018802 0.43175 1.9955 1.995 15.997 144.9809 0.00015359 -85.6644 0.96795
4.072 0.98807 5.4989e-005 3.8183 0.011993 5.3334e-005 0.001158 0.22716 0.00065926 0.22782 0.21005 0 0.032587 0.0389 0 1.1764 0.37769 0.11234 0.014459 7.1388 0.090221 0.00011265 0.79989 0.0071572 0.0079915 0.0013834 0.98698 0.99173 2.9826e-006 1.193e-005 0.14723 0.95949 0.92338 0.0013955 0.99586 0.59251 0.0018802 0.43176 1.9958 1.9953 15.9969 144.981 0.00015355 -85.6644 0.96895
4.073 0.98807 5.4989e-005 3.8183 0.011993 5.3347e-005 0.001158 0.22717 0.00065926 0.22783 0.21006 0 0.032587 0.0389 0 1.1765 0.37774 0.11235 0.01446 7.1403 0.090231 0.00011266 0.79988 0.0071579 0.0079923 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14723 0.95956 0.92341 0.0013955 0.99587 0.59265 0.0018802 0.43177 1.9961 1.9957 15.9969 144.981 0.0001535 -85.6644 0.96995
4.074 0.98807 5.4989e-005 3.8183 0.011993 5.336e-005 0.001158 0.22718 0.00065926 0.22783 0.21006 0 0.032587 0.0389 0 1.1766 0.37778 0.11237 0.014462 7.1419 0.090241 0.00011268 0.79987 0.0071586 0.007993 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14724 0.95964 0.92344 0.0013955 0.99588 0.59279 0.0018802 0.43178 1.9964 1.996 15.9969 144.981 0.00015345 -85.6645 0.97095
4.075 0.98807 5.4989e-005 3.8183 0.011993 5.3373e-005 0.001158 0.22718 0.00065926 0.22784 0.21007 0 0.032586 0.0389 0 1.1767 0.37783 0.11239 0.014464 7.1435 0.090251 0.00011269 0.79986 0.0071593 0.0079937 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14725 0.95971 0.92347 0.0013955 0.99588 0.59294 0.0018802 0.43179 1.9967 1.9963 15.9968 144.981 0.0001534 -85.6645 0.97195
4.076 0.98807 5.4989e-005 3.8183 0.011993 5.3386e-005 0.001158 0.22719 0.00065926 0.22784 0.21008 0 0.032586 0.0389 0 1.1768 0.37788 0.1124 0.014465 7.145 0.090262 0.00011271 0.79985 0.00716 0.0079945 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14725 0.95979 0.9235 0.0013955 0.99589 0.59308 0.0018802 0.4318 1.997 1.9966 15.9968 144.981 0.00015335 -85.6645 0.97295
4.077 0.98807 5.4989e-005 3.8183 0.011993 5.3399e-005 0.001158 0.2272 0.00065926 0.22785 0.21008 0 0.032586 0.0389 0 1.1769 0.37792 0.11242 0.014467 7.1466 0.090272 0.00011272 0.79984 0.0071607 0.0079952 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14726 0.95986 0.92353 0.0013955 0.9959 0.59322 0.0018802 0.43182 1.9973 1.9969 15.9968 144.9811 0.00015331 -85.6645 0.97395
4.078 0.98807 5.4989e-005 3.8183 0.011993 5.3412e-005 0.001158 0.2272 0.00065926 0.22786 0.21009 0 0.032585 0.0389 0 1.177 0.37797 0.11243 0.014468 7.1482 0.090282 0.00011274 0.79983 0.0071613 0.007996 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14726 0.95994 0.92356 0.0013955 0.99591 0.59336 0.0018802 0.43183 1.9976 1.9972 15.9967 144.9811 0.00015326 -85.6646 0.97495
4.079 0.98807 5.4989e-005 3.8183 0.011993 5.3425e-005 0.001158 0.22721 0.00065926 0.22786 0.21009 0 0.032585 0.0389 0 1.1771 0.37802 0.11245 0.01447 7.1498 0.090292 0.00011275 0.79982 0.007162 0.0079967 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14727 0.96001 0.92359 0.0013955 0.99592 0.5935 0.0018802 0.43184 1.9979 1.9975 15.9967 144.9811 0.00015321 -85.6646 0.97595
4.08 0.98807 5.4989e-005 3.8183 0.011993 5.3438e-005 0.001158 0.22721 0.00065926 0.22787 0.2101 0 0.032585 0.0389 0 1.1772 0.37806 0.11247 0.014472 7.1513 0.090302 0.00011276 0.79981 0.0071627 0.0079975 0.0013834 0.98698 0.99173 2.9825e-006 1.193e-005 0.14727 0.96008 0.92362 0.0013955 0.99593 0.59364 0.0018802 0.43185 1.9982 1.9978 15.9967 144.9811 0.00015317 -85.6646 0.97695
4.081 0.98807 5.4989e-005 3.8183 0.011993 5.3451e-005 0.001158 0.22722 0.00065926 0.22788 0.21011 0 0.032585 0.0389 0 1.1773 0.37811 0.11248 0.014473 7.1529 0.090313 0.00011278 0.7998 0.0071634 0.0079982 0.0013833 0.98698 0.99173 2.9825e-006 1.193e-005 0.14728 0.96016 0.92365 0.0013955 0.99593 0.59379 0.0018802 0.43186 1.9985 1.9981 15.9966 144.9811 0.00015312 -85.6646 0.97795
4.082 0.98807 5.4988e-005 3.8183 0.011992 5.3465e-005 0.001158 0.22723 0.00065926 0.22788 0.21011 0 0.032584 0.0389 0 1.1774 0.37816 0.1125 0.014475 7.1545 0.090323 0.00011279 0.79979 0.0071641 0.007999 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.14728 0.96023 0.92368 0.0013955 0.99594 0.59393 0.0018802 0.43187 1.9988 1.9984 15.9966 144.9812 0.00015307 -85.6646 0.97895
4.083 0.98807 5.4988e-005 3.8183 0.011992 5.3478e-005 0.001158 0.22723 0.00065926 0.22789 0.21012 0 0.032584 0.0389 0 1.1775 0.3782 0.11251 0.014477 7.1561 0.090333 0.00011281 0.79978 0.0071648 0.0079997 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.14729 0.9603 0.92371 0.0013955 0.99595 0.59407 0.0018802 0.43188 1.9992 1.9987 15.9966 144.9812 0.00015303 -85.6647 0.97995
4.084 0.98807 5.4988e-005 3.8183 0.011992 5.3491e-005 0.001158 0.22724 0.00065926 0.22789 0.21012 0 0.032584 0.0389 0 1.1776 0.37825 0.11253 0.014478 7.1576 0.090343 0.00011282 0.79977 0.0071655 0.0080005 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.1473 0.96037 0.92374 0.0013955 0.99596 0.59421 0.0018802 0.43189 1.9995 1.999 15.9965 144.9812 0.00015298 -85.6647 0.98095
4.085 0.98807 5.4988e-005 3.8183 0.011992 5.3504e-005 0.001158 0.22725 0.00065926 0.2279 0.21013 0 0.032583 0.0389 0 1.1777 0.3783 0.11255 0.01448 7.1592 0.090353 0.00011283 0.79976 0.0071662 0.0080012 0.0013833 0.98698 0.99173 2.9824e-006 1.193e-005 0.1473 0.96045 0.92377 0.0013955 0.99597 0.59435 0.0018802 0.43191 1.9998 1.9993 15.9965 144.9812 0.00015293 -85.6647 0.98195
4.086 0.98807 5.4988e-005 3.8183 0.011992 5.3517e-005 0.001158 0.22725 0.00065926 0.22791 0.21013 0 0.032583 0.0389 0 1.1778 0.37834 0.11256 0.014482 7.1608 0.090364 0.00011285 0.79975 0.0071669 0.0080019 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14731 0.96052 0.9238 0.0013955 0.99597 0.59449 0.0018802 0.43192 2.0001 1.9996 15.9965 144.9812 0.00015289 -85.6647 0.98295
4.087 0.98807 5.4988e-005 3.8183 0.011992 5.353e-005 0.001158 0.22726 0.00065926 0.22791 0.21014 0 0.032583 0.0389 0 1.1779 0.37839 0.11258 0.014483 7.1624 0.090374 0.00011286 0.79974 0.0071676 0.0080027 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14731 0.96059 0.92383 0.0013955 0.99598 0.59463 0.0018802 0.43193 2.0004 1.9999 15.9964 144.9813 0.00015284 -85.6647 0.98395
4.088 0.98807 5.4988e-005 3.8183 0.011992 5.3543e-005 0.0011581 0.22726 0.00065926 0.22792 0.21015 0 0.032582 0.0389 0 1.178 0.37843 0.11259 0.014485 7.1639 0.090384 0.00011288 0.79973 0.0071683 0.0080034 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14732 0.96066 0.92386 0.0013955 0.99599 0.59477 0.0018802 0.43194 2.0007 2.0002 15.9964 144.9813 0.00015279 -85.6648 0.98495
4.089 0.98807 5.4988e-005 3.8183 0.011992 5.3556e-005 0.0011581 0.22727 0.00065926 0.22792 0.21015 0 0.032582 0.0389 0 1.1781 0.37848 0.11261 0.014487 7.1655 0.090394 0.00011289 0.79972 0.007169 0.0080042 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14732 0.96073 0.92389 0.0013955 0.996 0.59492 0.0018802 0.43195 2.001 2.0005 15.9964 144.9813 0.00015275 -85.6648 0.98595
4.09 0.98807 5.4988e-005 3.8183 0.011992 5.3569e-005 0.0011581 0.22728 0.00065926 0.22793 0.21016 0 0.032582 0.0389 0 1.1782 0.37853 0.11263 0.014488 7.1671 0.090405 0.00011291 0.79971 0.0071697 0.0080049 0.0013833 0.98698 0.99173 2.9824e-006 1.1929e-005 0.14733 0.96081 0.92392 0.0013955 0.996 0.59506 0.0018802 0.43196 2.0013 2.0008 15.9963 144.9813 0.0001527 -85.6648 0.98695
4.091 0.98807 5.4988e-005 3.8183 0.011992 5.3582e-005 0.0011581 0.22728 0.00065926 0.22794 0.21016 0 0.032581 0.0389 0 1.1783 0.37857 0.11264 0.01449 7.1687 0.090415 0.00011292 0.7997 0.0071704 0.0080057 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14733 0.96088 0.92395 0.0013955 0.99601 0.5952 0.0018802 0.43197 2.0016 2.0011 15.9963 144.9813 0.00015266 -85.6648 0.98795
4.092 0.98807 5.4988e-005 3.8183 0.011992 5.3595e-005 0.0011581 0.22729 0.00065926 0.22794 0.21017 0 0.032581 0.0389 0 1.1784 0.37862 0.11266 0.014492 7.1702 0.090425 0.00011293 0.79969 0.0071711 0.0080064 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14734 0.96095 0.92397 0.0013955 0.99602 0.59534 0.0018802 0.43198 2.0019 2.0014 15.9963 144.9814 0.00015261 -85.6648 0.98895
4.093 0.98807 5.4988e-005 3.8183 0.011992 5.3608e-005 0.0011581 0.22729 0.00065926 0.22795 0.21018 0 0.032581 0.0389 0 1.1785 0.37867 0.11267 0.014493 7.1718 0.090435 0.00011295 0.79968 0.0071718 0.0080072 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14735 0.96102 0.924 0.0013955 0.99603 0.59548 0.0018801 0.432 2.0022 2.0017 15.9962 144.9814 0.00015257 -85.6649 0.98995
4.094 0.98807 5.4988e-005 3.8183 0.011992 5.3621e-005 0.0011581 0.2273 0.00065926 0.22796 0.21018 0 0.03258 0.0389 0 1.1786 0.37871 0.11269 0.014495 7.1734 0.090445 0.00011296 0.79967 0.0071724 0.0080079 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14735 0.96109 0.92403 0.0013955 0.99603 0.59562 0.0018801 0.43201 2.0025 2.002 15.9962 144.9814 0.00015252 -85.6649 0.99095
4.095 0.98807 5.4988e-005 3.8183 0.011992 5.3634e-005 0.0011581 0.22731 0.00065926 0.22796 0.21019 0 0.03258 0.0389 0 1.1787 0.37876 0.11271 0.014496 7.175 0.090456 0.00011298 0.79966 0.0071731 0.0080087 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14736 0.96116 0.92406 0.0013955 0.99604 0.59576 0.0018801 0.43202 2.0028 2.0023 15.9962 144.9814 0.00015248 -85.6649 0.99195
4.096 0.98807 5.4987e-005 3.8183 0.011992 5.3647e-005 0.0011581 0.22731 0.00065926 0.22797 0.21019 0 0.03258 0.0389 0 1.1788 0.37881 0.11272 0.014498 7.1766 0.090466 0.00011299 0.79965 0.0071738 0.0080094 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14736 0.96123 0.92409 0.0013955 0.99605 0.5959 0.0018801 0.43203 2.0031 2.0026 15.9961 144.9814 0.00015243 -85.6649 0.99295
4.097 0.98807 5.4987e-005 3.8183 0.011992 5.366e-005 0.0011581 0.22732 0.00065926 0.22797 0.2102 0 0.03258 0.0389 0 1.1789 0.37885 0.11274 0.0145 7.1781 0.090476 0.000113 0.79964 0.0071745 0.0080101 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14737 0.9613 0.92412 0.0013955 0.99606 0.59604 0.0018801 0.43204 2.0033 2.0029 15.9961 144.9815 0.00015239 -85.6649 0.99395
4.098 0.98807 5.4987e-005 3.8183 0.011992 5.3673e-005 0.0011581 0.22732 0.00065926 0.22798 0.2102 0 0.032579 0.0389 0 1.179 0.3789 0.11275 0.014501 7.1797 0.090486 0.00011302 0.79963 0.0071752 0.0080109 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14737 0.96137 0.92415 0.0013955 0.99606 0.59618 0.0018801 0.43205 2.0036 2.0032 15.9961 144.9815 0.00015234 -85.665 0.99495
4.099 0.98807 5.4987e-005 3.8183 0.011992 5.3686e-005 0.0011581 0.22733 0.00065926 0.22799 0.21021 0 0.032579 0.0389 0 1.1791 0.37895 0.11277 0.014503 7.1813 0.090496 0.00011303 0.79962 0.0071759 0.0080116 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14738 0.96144 0.92417 0.0013955 0.99607 0.59632 0.0018801 0.43206 2.0039 2.0035 15.996 144.9815 0.0001523 -85.665 0.99595
4.1 0.98807 5.4987e-005 3.8183 0.011992 5.3699e-005 0.0011581 0.22734 0.00065926 0.22799 0.21022 0 0.032579 0.0389 0 1.1792 0.37899 0.11279 0.014505 7.1829 0.090507 0.00011305 0.79961 0.0071766 0.0080124 0.0013833 0.98698 0.99173 2.9823e-006 1.1929e-005 0.14738 0.96151 0.9242 0.0013955 0.99608 0.59646 0.0018801 0.43207 2.0042 2.0038 15.996 144.9815 0.00015226 -85.6636 0.99695
4.101 0.98807 5.4987e-005 3.8183 0.011992 5.3712e-005 0.0011581 0.22734 0.00065926 0.228 0.21022 0 0.032578 0.0389 0 1.1793 0.37904 0.1128 0.014506 7.1845 0.090517 0.00011306 0.7996 0.0071773 0.0080131 0.0064733 0.98323 0.991 1.4518e-005 5.3336e-005 0.14739 0.96152 0.92423 0.0027732 0.99607 0.59659 0.0023954 0.43203 2.0045 2.0041 15.9959 144.9815 0.00015222 -76.1605 0.99795
4.102 0.98807 5.4987e-005 3.8183 0.011992 5.3725e-005 0.0011581 0.22735 0.00065926 0.228 0.21023 0 0.032578 0.0389 0 1.1794 0.37909 0.11282 0.014508 7.186 0.090527 0.00011308 0.79959 0.007178 0.0080139 0.026222 0.97171 0.98767 6.5982e-005 0.00022951 0.1474 0.96132 0.92426 0.0053008 0.99602 0.59669 0.0033361 0.43191 2.0048 2.0044 15.9959 144.9815 0.00015221 -67.1465 0.99895
4.103 0.98807 5.4987e-005 3.8183 0.011992 5.3738e-005 0.0011581 0.22736 0.00065926 0.22801 0.21023 0 0.032578 0.0389 0 1.1795 0.37913 0.11283 0.01451 7.1876 0.090537 0.00011309 0.79958 0.0071787 0.0080146 0.094879 0.94722 0.97733 0.00028442 0.00091318 0.1474 0.96057 0.92428 0.0092477 0.99575 0.59678 0.0044249 0.43175 2.0051 2.0047 15.9958 144.9815 0.00015222 -58.0148 0.99995
4.104 0.98807 5.4987e-005 3.8183 0.011992 5.3751e-005 0.0011581 0.22736 0.00065926 0.22802 0.21024 0 0.032577 0.0389 0 1.1796 0.37918 0.11285 0.014511 7.1892 0.090547 0.0001131 0.79957 0.0071794 0.0080154 0.48812 0.85628 0.93873 0.0021798 0.0054769 0.14741 0.95856 0.92431 0.015753 0.99165 0.5968 0.0056239 0.43156 2.0054 2.005 15.9966 144.9815 0.00015225 -37.2126 0.15598
4.105 0.98807 5.4987e-005 3.8183 0.011992 5.3764e-005 0.0011581 0.22737 0.00065926 0.22802 0.21024 0 0.032577 0.0389 0 1.1797 0.37923 0.11287 0.014513 7.1908 0.090558 0.00011312 0.79956 0.0071801 0.0080161 0.99961 0.0021706 0.71211 0.93945 0.99615 0.14741 0.9251 0.92132 0.33367 0.96423 0.58369 0.044223 0.43135 1.9592 0.94838 16.0004 144.9811 0.00023814 24.4562 0.0019435
4.106 0.98807 5.4987e-005 3.8183 0.011992 5.3777e-005 0.0011581 0.22737 0.00065926 0.22803 0.21025 0 0.032577 0.0389 0 1.1798 0.37927 0.11288 0.014515 7.1924 0.090568 0.00011313 0.79955 0.0071808 0.0080168 0.9994 1.3709e-006 0.52823 0.99735 0.99942 0.14742 0.88507 0.90333 0.61155 0.93707 0.56739 0.097105 0.43115 1.769 0.58942 16.0001 144.9798 0.00034855 19.8557 0.0029435
4.107 0.98807 5.4987e-005 3.8183 0.011992 5.379e-005 0.0011581 0.22738 0.00065926 0.22803 0.21026 0 0.032576 0.0389 0 1.1799 0.37932 0.1129 0.014516 7.1939 0.090578 0.00011315 0.79954 0.0071814 0.0080176 0.99894 4.4697e-010 0.3922 0.99502 0.99857 0.14742 0.84749 0.88009 0.73123 0.91068 0.55178 0.13695 0.43094 1.5885 0.56592 15.9997 144.9781 0.00041854 14.4402 0.0039435
4.108 0.98807 5.4987e-005 3.8183 0.011992 5.3803e-005 0.0011581 0.22739 0.00065926 0.22804 0.21026 0 0.032576 0.0389 0 1.18 0.37937 0.11291 0.014518 7.1955 0.090588 0.00011316 0.79953 0.0071821 0.0080183 0.99841 -8.1231e-011 0.29157 0.99056 0.99725 0.14743 0.81287 0.85427 0.78311 0.88503 0.53706 0.16786 0.43074 1.4381 0.60475 15.9994 144.9763 0.0004709 10.7634 0.0049435
4.109 0.98807 5.4987e-005 3.8183 0.011992 5.3816e-005 0.0011581 0.22739 0.00065926 0.22805 0.21027 0 0.032576 0.0389 0 1.1801 0.37941 0.11293 0.014519 7.1971 0.090598 0.00011318 0.79951 0.0071828 0.0080191 0.99792 3.9373e-011 0.21701 0.9852 0.99571 0.14743 0.78106 0.82713 0.80492 0.86011 0.52324 0.19348 0.43053 1.3185 0.66343 15.999 144.9746 0.00051114 8.3281 0.0059435
4.11 0.98807 5.4986e-005 3.8183 0.011992 5.3829e-005 0.0011581 0.2274 0.00065926 0.22805 0.21027 0 0.032576 0.0389 0 1.1802 0.37946 0.11295 0.014521 7.1987 0.090609 0.00011319 0.7995 0.0071835 0.0080198 0.99747 -8.9597e-011 0.16169 0.97935 0.99404 0.14744 0.75168 0.79954 0.81175 0.8359 0.51027 0.21561 0.43033 1.2266 0.7267 15.9987 144.9729 0.00054197 6.5151 0.0069435
4.111 0.98807 5.4986e-005 3.8183 0.011992 5.3842e-005 0.0011581 0.2274 0.00065926 0.22806 0.21028 0 0.032575 0.0389 0 1.1803 0.37951 0.11296 0.014523 7.2003 0.090619 0.0001132 0.79949 0.0071842 0.0080206 0.99701 4.7174e-011 0.12059 0.973 0.99221 0.14745 0.72444 0.77211 0.81026 0.81237 0.49808 0.23511 0.43012 1.1583 0.78673 15.9984 144.9713 0.00056548 5.0017 0.0079435
4.112 0.98807 5.4986e-005 3.8183 0.011992 5.3855e-005 0.0011581 0.22741 0.00065926 0.22806 0.21028 0 0.032575 0.0389 0 1.1804 0.37955 0.11298 0.014524 7.2019 0.090629 0.00011322 0.79948 0.0071849 0.0080213 0.99653 -4.2599e-010 0.090032 0.96599 0.99015 0.14745 0.69915 0.7453 0.80375 0.78951 0.48665 0.25247 0.42992 1.1091 0.83928 15.9981 144.9698 0.00058342 3.6333 0.0089435
4.113 0.98807 5.4986e-005 3.8183 0.011992 5.3868e-005 0.0011581 0.22742 0.00065926 0.22807 0.21029 0 0.032575 0.0389 0 1.1805 0.3796 0.11299 0.014526 7.2035 0.090639 0.00011323 0.79947 0.0071856 0.008022 0.99599 -3.1908e-010 0.067288 0.95807 0.98776 0.14746 0.67566 0.71941 0.79393 0.7673 0.47597 0.26795 0.42971 1.0747 0.88262 15.9978 144.9683 0.00059727 2.3288 0.0099435
4.114 0.98807 5.4986e-005 3.8183 0.011992 5.3881e-005 0.0011581 0.22742 0.00065926 0.22808 0.2103 0 0.032574 0.0389 0 1.1806 0.37965 0.11301 0.014528 7.205 0.090649 0.00011325 0.79946 0.0071863 0.0080228 0.99538 1.1945e-010 0.050349 0.94892 0.98491 0.14746 0.65388 0.69466 0.7817 0.74572 0.46603 0.28176 0.42951 1.0514 0.91677 15.9976 144.9669 0.00060818 1.0392 0.010943
4.115 0.98807 5.4986e-005 3.8183 0.011992 5.3894e-005 0.0011581 0.22743 0.00065926 0.22808 0.2103 0 0.032574 0.0389 0 1.1807 0.37969 0.11303 0.014529 7.2066 0.090659 0.00011326 0.79945 0.007187 0.0080235 0.99466 -4.3003e-011 0.037724 0.93819 0.98144 0.14747 0.63373 0.67123 0.76756 0.72475 0.45684 0.29402 0.4293 1.0363 0.94278 15.9973 144.9656 0.00061696 -0.27123 0.011943
4.116 0.98807 5.4986e-005 3.8183 0.011992 5.3907e-005 0.0011581 0.22743 0.00065926 0.22809 0.21031 0 0.032574 0.0389 0 1.1808 0.37974 0.11304 0.014531 7.2082 0.09067 0.00011327 0.79944 0.0071877 0.0080243 0.9938 -1.3439e-011 0.028309 0.92539 0.97715 0.14747 0.61517 0.64924 0.75169 0.70438 0.44841 0.30483 0.4291 1.0269 0.96216 15.997 144.9644 0.00062421 -1.6354 0.012943
4.117 0.98807 5.4986e-005 3.8183 0.011992 5.392e-005 0.0011581 0.22744 0.00065926 0.22809 0.21031 0 0.032573 0.0389 0 1.1809 0.37979 0.11306 0.014533 7.2098 0.09068 0.00011329 0.79943 0.0071884 0.008025 0.99271 2.5154e-011 0.021283 0.90987 0.97173 0.14748 0.59816 0.62881 0.73412 0.68459 0.44076 0.31424 0.42889 1.0215 0.97647 15.9968 144.9633 0.00063029 -3.089 0.013943
4.118 0.98807 5.4986e-005 3.8183 0.011992 5.3933e-005 0.0011581 0.22745 0.00065926 0.2281 0.21032 0 0.032573 0.0389 0 1.181 0.37983 0.11307 0.014534 7.2114 0.09069 0.0001133 0.79942 0.0071891 0.0080258 0.99131 -1.921e-011 0.016037 0.89076 0.96471 0.14748 0.5827 0.61008 0.71472 0.66538 0.43394 0.32229 0.42869 1.0187 0.98704 15.9965 144.9623 0.00063545 -4.6763 0.014943
4.119 0.98807 5.4986e-005 3.8183 0.011992 5.3946e-005 0.0011581 0.22745 0.00065926 0.22811 0.21032 0 0.032573 0.0389 0 1.1811 0.37988 0.11309 0.014536 7.213 0.0907 0.00011332 0.79941 0.0071897 0.0080265 0.98942 2.5255e-011 0.012119 0.8668 0.95539 0.14749 0.56881 0.59316 0.69324 0.64672 0.42796 0.329 0.42849 1.0178 0.99496 15.9963 144.9613 0.00063982 -6.4573 0.015943
4.12 0.98807 5.4986e-005 3.8183 0.011992 5.3959e-005 0.0011581 0.22746 0.00065926 0.22811 0.21033 0 0.032573 0.0389 0 1.1812 0.37993 0.11311 0.014538 7.2146 0.09071 0.00011333 0.7994 0.0071904 0.0080272 0.9867 -2.8129e-011 0.009194 0.83613 0.94265 0.1475 0.55652 0.57823 0.66931 0.62862 0.42288 0.33436 0.42828 1.0181 1.0011 15.996 144.9604 0.00064344 -8.5158 0.016943
4.121 0.98807 5.4986e-005 3.8183 0.011992 5.3972e-005 0.0011581 0.22746 0.00065926 0.22812 0.21034 0 0.032572 0.0389 0 1.1813 0.37997 0.11312 0.014539 7.2162 0.090721 0.00011335 0.79939 0.0071911 0.008028 0.98252 4.1447e-011 0.0070128 0.796 0.92465 0.1475 0.54591 0.56546 0.64247 0.61108 0.41873 0.33833 0.42808 1.0192 1.0059 15.9958 144.9596 0.00064632 -10.9713 0.017943
4.122 0.98807 5.4986e-005 3.8183 0.011992 5.3985e-005 0.0011581 0.22747 0.00065926 0.22812 0.21034 0 0.032572 0.0389 0 1.1814 0.38002 0.11314 0.014541 7.2177 0.090731 0.00011336 0.79938 0.0071918 0.0080287 0.97554 -5.7307e-011 0.0053922 0.74232 0.89833 0.14751 0.53705 0.55505 0.61222 0.5941 0.41553 0.34088 0.42788 1.0208 1.01 15.9956 144.9588 0.00064838 -13.9875 0.018943
4.123 0.98807 5.4986e-005 3.8183 0.011992 5.3998e-005 0.0011581 0.22748 0.00065926 0.22813 0.21035 0 0.032572 0.0389 0 1.1815 0.38007 0.11315 0.014542 7.2193 0.090741 0.00011337 0.79937 0.0071925 0.0080295 0.96275 1.4989e-011 0.0041984 0.66925 0.85863 0.14751 0.52999 0.54716 0.57821 0.57776 0.41324 0.34202 0.42767 1.0227 1.0135 15.9954 144.9582 0.00064953 -17.7636 0.019943
4.124 0.98807 5.4985e-005 3.8183 0.011992 5.4011e-005 0.0011581 0.22748 0.00065926 0.22814 0.21035 0 0.032571 0.0389 0 1.1816 0.38011 0.11317 0.014544 7.2209 0.090751 0.00011339 0.79936 0.0071932 0.0080302 0.93722 8.5838e-012 0.0033353 0.56959 0.79753 0.14752 0.52467 0.54181 0.54044 0.5622 0.41177 0.34182 0.42747 1.0249 1.0167 15.9952 144.9577 0.00064967 -22.4576 0.020943
4.125 0.98807 5.4985e-005 3.8183 0.011992 5.4024e-005 0.0011581 0.22749 0.00065926 0.22814 0.21036 0 0.032571 0.0389 0 1.1816 0.38016 0.11319 0.014546 7.2225 0.090761 0.0001134 0.79935 0.0071939 0.008031 0.88481 -7.3995e-011 0.0027332 0.4388 0.7045 0.14752 0.52085 0.53869 0.49904 0.54786 0.41093 0.34043 0.42727 1.0272 1.0196 15.9951 144.9572 0.00064883 -27.9753 0.021943
4.126 0.98807 5.4985e-005 3.8183 0.011992 5.4037e-005 0.0011581 0.22749 0.00065926 0.22815 0.21036 0 0.032571 0.0389 0 1.1817 0.3802 0.1132 0.014547 7.2241 0.090771 0.00011342 0.79934 0.0071946 0.0080317 0.78775 -3.9266e-011 0.0023329 0.28676 0.57247 0.14753 0.51812 0.53708 0.45311 0.53573 0.4105 0.33798 0.42707 1.0295 1.0224 15.995 144.9568 0.00064731 -33.742 0.022943
4.127 0.98807 5.4985e-005 3.8183 0.011992 5.405e-005 0.0011581 0.2275 0.00065926 0.22815 0.21037 0 0.03257 0.0389 0 1.1818 0.38025 0.11322 0.014549 7.2257 0.090782 0.00011343 0.79933 0.0071953 0.0080324 0.64848 -1.3987e-011 0.0020743 0.1477 0.41181 0.14753 0.5161 0.53623 0.40029 0.52736 0.41031 0.33436 0.42687 1.032 1.0251 15.9949 144.9565 0.00064547 -38.9831 0.023943
4.128 0.98807 5.4985e-005 3.8183 0.011992 5.4063e-005 0.0011581 0.22751 0.00065926 0.22816 0.21038 0 0.03257 0.0389 0 1.1819 0.3803 0.11323 0.014551 7.2273 0.090792 0.00011344 0.79932 0.007196 0.0080332 0.49992 0.00035428 0.0020277 0.057038 0.25433 0.14754 0.51459 0.53596 0.33929 0.52351 0.41028 0.32922 0.42667 1.0344 1.0277 15.9948 144.9563 0.00064353 -43.3659 0.024943
4.129 0.98807 5.4985e-005 3.8183 0.011992 5.4076e-005 0.0011581 0.22751 0.00065926 0.22817 0.21038 0 0.03257 0.0389 0 1.182 0.38034 0.11325 0.014552 7.2289 0.090802 0.00011346 0.79931 0.0071967 0.0080339 0.37384 0.0010792 0.002276 0.016764 0.13276 0.14755 0.51348 0.53657 0.27247 0.523 0.41032 0.32221 0.42647 1.0369 1.0302 15.9947 144.9561 0.00064155 -46.9372 0.025943
4.13 0.98807 5.4985e-005 3.8183 0.011992 5.4089e-005 0.0011581 0.22752 0.00065926 0.22817 0.21039 0 0.03257 0.0389 0 1.1821 0.38039 0.11327 0.014554 7.2305 0.090812 0.00011347 0.7993 0.0071974 0.0080347 0.28094 0.0022415 0.0028333 0.0044853 0.058953 0.14755 0.5127 0.53814 0.20577 0.52408 0.41041 0.31313 0.42628 1.0393 1.0328 15.9947 144.956 0.00063953 -49.8191 0.026943
4.131 0.98807 5.4985e-005 3.8183 0.011992 5.4102e-005 0.0011582 0.22752 0.00065926 0.22818 0.21039 0 0.032569 0.0389 0 1.1822 0.38044 0.11328 0.014556 7.2321 0.090822 0.00011349 0.79929 0.007198 0.0080354 0.21663 0.003941 0.0037132 0.0016402 0.023258 0.14756 0.51221 0.54038 0.1462 0.52569 0.41052 0.30197 0.42609 1.0418 1.0353 15.9946 144.9559 0.00063749 -52.1428 0.027943
4.132 0.98807 5.4985e-005 3.8183 0.011992 5.4115e-005 0.0011582 0.22753 0.00065926 0.22818 0.2104 0 0.032569 0.0389 0 1.1823 0.38048 0.1133 0.014557 7.2336 0.090832 0.0001135 0.79928 0.0071987 0.0080362 0.17228 0.0062471 0.0049165 0.00094335 0.009081 0.14756 0.51196 0.54294 0.098647 0.52741 0.41065 0.28891 0.4259 1.0443 1.0378 15.9946 144.9558 0.00063543 -54.0423 0.028943
4.133 0.98807 5.4985e-005 3.8183 0.011992 5.4128e-005 0.0011582 0.22753 0.00065926 0.22819 0.2104 0 0.032569 0.0389 0 1.1824 0.38053 0.11331 0.014559 7.2352 0.090843 0.00011351 0.79927 0.0071994 0.0080369 0.14069 0.0092097 0.0064392 0.0006689 0.00416 0.14757 0.51191 0.54561 0.064439 0.52909 0.41079 0.27422 0.42572 1.0467 1.0403 15.9946 144.9558 0.00063335 -55.6409 0.029943
4.134 0.98807 5.4985e-005 3.8183 0.011992 5.4141e-005 0.0011582 0.22754 0.00065926 0.2282 0.21041 0 0.032568 0.0389 0 1.1825 0.38058 0.11333 0.014561 7.2368 0.090853 0.00011353 0.79926 0.0072001 0.0080376 0.11711 0.012877 0.0082797 0.00050934 0.0024677 0.14757 0.51202 0.5483 0.041969 0.5307 0.41092 0.25819 0.42554 1.0492 1.0428 15.9946 144.9558 0.00063127 -57.0386 0.030943
4.135 0.98807 5.4985e-005 3.8183 0.011992 5.4154e-005 0.0011582 0.22755 0.00065926 0.2282 0.21041 0 0.032568 0.0389 0 1.1826 0.38062 0.11335 0.014562 7.2384 0.090863 0.00011354 0.79925 0.0072008 0.0080384 0.098695 0.017308 0.010444 0.000401 0.0017659 0.14758 0.51227 0.55098 0.028266 0.53224 0.41107 0.24112 0.42536 1.0517 1.0453 15.9946 144.9557 0.00062918 -58.3079 0.031943
4.136 0.98807 5.4985e-005 3.8183 0.011992 5.4167e-005 0.0011582 0.22755 0.00065926 0.22821 0.21042 0 0.032568 0.0389 0 1.1827 0.38067 0.11336 0.014564 7.24 0.090873 0.00011356 0.79924 0.0072015 0.0080391 0.083789 0.022585 0.012945 0.00032177 0.0013734 0.14758 0.51264 0.55363 0.020332 0.53369 0.41121 0.22326 0.42519 1.0542 1.0478 15.9946 144.9557 0.00062708 -59.4956 0.032943
4.137 0.98807 5.4985e-005 3.8183 0.011992 5.418e-005 0.0011582 0.22756 0.00065926 0.22821 0.21043 0 0.032567 0.0389 0 1.1828 0.38072 0.11338 0.014565 7.2416 0.090883 0.00011357 0.79923 0.0072022 0.0080399 0.071445 0.028809 0.015804 0.00026128 0.0011021 0.14759 0.51313 0.55626 0.015815 0.53507 0.41135 0.20486 0.42502 1.0566 1.0502 15.9946 144.9557 0.00062498 -60.6297 0.033943
4.138 0.98807 5.4984e-005 3.8183 0.011992 5.4193e-005 0.0011582 0.22756 0.00065926 0.22822 0.21043 0 0.032567 0.0389 0 1.1829 0.38076 0.11339 0.014567 7.2432 0.090893 0.00011359 0.79922 0.0072029 0.0080406 0.06109 0.036102 0.019049 0.0002145 0.00089663 0.1476 0.51371 0.55887 0.013152 0.5364 0.4115 0.18616 0.42485 1.0591 1.0527 15.9946 144.9557 0.00062288 -61.7252 0.034943
4.139 0.98807 5.4984e-005 3.8183 0.011992 5.4206e-005 0.0011582 0.22757 0.00065926 0.22822 0.21044 0 0.032567 0.0389 0 1.183 0.38081 0.11341 0.014569 7.2448 0.090904 0.0001136 0.79921 0.0072036 0.0080414 0.052347 0.044599 0.022709 0.00017682 0.00073556 0.1476 0.51439 0.56145 0.011433 0.53766 0.41164 0.16742 0.42468 1.0615 1.0552 15.9947 144.9556 0.00062077 -62.79 0.035943
4.14 0.98807 5.4984e-005 3.8183 0.011992 5.4219e-005 0.0011582 0.22758 0.00065926 0.22823 0.21044 0 0.032567 0.0389 0 1.1831 0.38086 0.11343 0.01457 7.2464 0.090914 0.00011361 0.7992 0.0072043 0.0080421 0.044942 0.05445 0.026819 0.00014673 0.00060728 0.14761 0.51515 0.564 0.010188 0.53889 0.41179 0.1489 0.42452 1.064 1.0577 15.9947 144.9556 0.00061866 -63.8279 0.036943
4.141 0.98807 5.4984e-005 3.8183 0.011992 5.4232e-005 0.0011582 0.22758 0.00065926 0.22824 0.21045 0 0.032566 0.0389 0 1.1832 0.3809 0.11344 0.014572 7.248 0.090924 0.00011363 0.79919 0.0072049 0.0080428 0.038659 0.065811 0.031418 0.00012221 0.00050416 0.14761 0.51599 0.56653 0.009195 0.54007 0.41194 0.13087 0.42437 1.0665 1.0602 15.9947 144.9556 0.00061655 -64.8408 0.037943
4.142 0.98807 5.4984e-005 3.8183 0.011992 5.4245e-005 0.0011582 0.22759 0.00065926 0.22824 0.21045 0 0.032566 0.0389 0 1.1833 0.38095 0.11346 0.014574 7.2496 0.090934 0.00011364 0.79918 0.0072056 0.0080436 0.033323 0.078846 0.036544 0.00010234 0.00042072 0.14762 0.51689 0.56903 0.0083547 0.54123 0.41208 0.11358 0.42421 1.0689 1.0626 15.9947 144.9555 0.00061444 -65.8296 0.038943
4.143 0.98807 5.4984e-005 3.8183 0.011992 5.4258e-005 0.0011582 0.22759 0.00065926 0.22825 0.21046 0 0.032566 0.0389 0 1.1834 0.381 0.11347 0.014575 7.2512 0.090944 0.00011366 0.79917 0.0072063 0.0080443 0.028787 0.093716 0.042244 8.6035e-005 0.00035282 0.14762 0.51785 0.57151 0.0076243 0.54236 0.41223 0.097284 0.42407 1.0714 1.0651 15.9948 144.9555 0.00061232 -66.7945 0.039943
4.144 0.98807 5.4984e-005 3.8183 0.011992 5.4271e-005 0.0011582 0.2276 0.00065926 0.22825 0.21046 0 0.032565 0.0389 0 1.1835 0.38104 0.11349 0.014577 7.2528 0.090954 0.00011367 0.79916 0.007207 0.0080451 0.024929 0.11058 0.048566 7.2699e-005 0.0002973 0.14763 0.51887 0.57396 0.0069809 0.54348 0.41238 0.082191 0.42392 1.0738 1.0676 15.9948 144.9555 0.00061021 -67.7357 0.040943
4.145 0.98807 5.4984e-005 3.8183 0.011992 5.4284e-005 0.0011582 0.22761 0.00065926 0.22826 0.21047 0 0.032565 0.0389 0 1.1836 0.38109 0.11351 0.014579 7.2544 0.090965 0.00011368 0.79915 0.0072077 0.0080458 0.021645 0.12958 0.055563 6.1644e-005 0.00025171 0.14763 0.51993 0.57639 0.0064108 0.54459 0.41253 0.068471 0.42378 1.0763 1.07 15.9949 144.9555 0.0006081 -68.6529 0.041943
4.146 0.98807 5.4984e-005 3.8183 0.011992 5.4297e-005 0.0011582 0.22761 0.00065926 0.22827 0.21048 0 0.032565 0.0389 0 1.1837 0.38114 0.11352 0.01458 7.256 0.090975 0.0001137 0.79914 0.0072084 0.0080465 0.018848 0.15084 0.063296 5.2561e-005 0.00021414 0.14764 0.52103 0.57879 0.0059041 0.5457 0.41268 0.056244 0.42365 1.0787 1.0725 15.9949 144.9554 0.00060598 -69.5454 0.042943
4.147 0.98807 5.4984e-005 3.8183 0.011992 5.431e-005 0.0011582 0.22762 0.00065926 0.22827 0.21048 0 0.032564 0.0389 0 1.1838 0.38118 0.11354 0.014582 7.2576 0.090985 0.00011371 0.79913 0.0072091 0.0080473 0.016463 0.17446 0.071829 4.5032e-005 0.00018306 0.14764 0.52217 0.58117 0.0054525 0.5468 0.41283 0.045573 0.42352 1.0811 1.075 15.995 144.9554 0.00060387 -70.4125 0.043943
4.148 0.98807 5.4984e-005 3.8183 0.011991 5.4323e-005 0.0011582 0.22762 0.00065926 0.22828 0.21049 0 0.032564 0.0389 0 1.1839 0.38123 0.11355 0.014583 7.2592 0.090995 0.00011373 0.79912 0.0072098 0.008048 0.014428 0.2005 0.081231 3.873e-005 0.00015728 0.14765 0.52333 0.58352 0.0050494 0.54792 0.41298 0.03646 0.4234 1.0836 1.0774 15.9951 144.9554 0.00060176 -71.2532 0.044943
4.149 0.98807 5.4984e-005 3.8183 0.011991 5.4336e-005 0.0011582 0.22763 0.00065926 0.22828 0.21049 0 0.032564 0.0389 0 1.184 0.38128 0.11357 0.014585 7.2608 0.091005 0.00011374 0.79911 0.0072105 0.0080488 0.012692 0.22897 0.091578 3.3508e-005 0.00013583 0.14766 0.52453 0.58585 0.0046893 0.54905 0.41313 0.02885 0.42328 1.086 1.0799 15.9951 144.9553 0.00059965 -72.0664 0.045943
4.15 0.98807 5.4984e-005 3.8183 0.011991 5.4349e-005 0.0011582 0.22763 0.00065926 0.22829 0.2105 0 0.032564 0.0389 0 1.1841 0.38132 0.11359 0.014587 7.2624 0.091015 0.00011376 0.7991 0.0072112 0.0080495 0.011209 0.25981 0.10294 2.9134e-005 0.00011793 0.14766 0.52575 0.58815 0.0043673 0.5502 0.41328 0.022642 0.42317 1.0884 1.0823 15.9952 144.9553 0.00059754 -72.8507 0.046943
4.151 0.98807 5.4984e-005 3.8183 0.011991 5.4362e-005 0.0011582 0.22764 0.00065926 0.2283 0.2105 0 0.032563 0.0389 0 1.1842 0.38137 0.1136 0.014588 7.264 0.091026 0.00011377 0.79909 0.0072118 0.0080503 0.0099411 0.2929 0.1154 2.5445e-005 0.00010296 0.14767 0.52699 0.59044 0.0040793 0.55137 0.41344 0.017695 0.42306 1.0909 1.0848 15.9953 144.9553 0.00059543 -73.605 0.047943
4.152 0.98807 5.4983e-005 3.8183 0.011991 5.4375e-005 0.0011582 0.22765 0.00065926 0.2283 0.21051 0 0.032563 0.0389 0 1.1843 0.38142 0.11362 0.01459 7.2656 0.091036 0.00011378 0.79908 0.0072125 0.008051 0.0088576 0.32805 0.129 2.2375e-005 9.0414e-005 0.14767 0.52825 0.5927 0.0038217 0.55257 0.41359 0.013842 0.42296 1.0933 1.0872 15.9953 144.9553 0.00059333 -74.3279 0.048943
4.153 0.98807 5.4983e-005 3.8183 0.011991 5.4388e-005 0.0011582 0.22765 0.00065926 0.22831 0.21051 0 0.032563 0.0389 0 1.1844 0.38146 0.11363 0.014592 7.2672 0.091046 0.0001138 0.79907 0.0072132 0.0080517 0.0079291 0.365 0.14381 1.9791e-005 7.9861e-005 0.14768 0.52952 0.59493 0.0035914 0.5538 0.41375 0.010908 0.42287 1.0957 1.0897 15.9954 144.9552 0.00059123 -75.0183 0.049943
4.154 0.98807 5.4983e-005 3.8183 0.011991 5.4401e-005 0.0011582 0.22766 0.00065926 0.22831 0.21052 0 0.032562 0.0389 0 1.1845 0.38151 0.11365 0.014593 7.2688 0.091056 0.00011381 0.79906 0.0072139 0.0080525 0.0071345 0.4034 0.15985 1.7601e-005 7.0976e-005 0.14768 0.5308 0.59715 0.0033855 0.55506 0.41391 0.0087194 0.42278 1.0982 1.0921 15.9955 144.9552 0.00058913 -75.6752 0.050943
4.155 0.98807 5.4983e-005 3.8183 0.011991 5.4414e-005 0.0011582 0.22766 0.00065926 0.22832 0.21053 0 0.032562 0.0389 0 1.1846 0.38156 0.11367 0.014595 7.2704 0.091066 0.00011383 0.79905 0.0072146 0.0080532 0.0064528 0.44286 0.17713 1.5755e-005 6.3474e-005 0.14769 0.5321 0.59934 0.0032016 0.55636 0.41407 0.0071165 0.4227 1.1006 1.0945 15.9956 144.9552 0.00058704 -76.2977 0.051943
4.156 0.98807 5.4983e-005 3.8183 0.011991 5.4427e-005 0.0011582 0.22767 0.00065926 0.22832 0.21053 0 0.032562 0.0389 0 1.1847 0.3816 0.11368 0.014597 7.272 0.091076 0.00011384 0.79904 0.0072153 0.008054 0.0058677 0.48291 0.1956 1.4187e-005 5.7121e-005 0.14769 0.5334 0.60151 0.0030374 0.55769 0.41423 0.0059583 0.42262 1.103 1.097 15.9957 144.9551 0.00058495 -76.8855 0.052943
4.157 0.98807 5.4983e-005 3.8183 0.011991 5.444e-005 0.0011582 0.22768 0.00065926 0.22833 0.21054 0 0.032562 0.0389 0 1.1848 0.38165 0.1137 0.014598 7.2736 0.091086 0.00011385 0.79903 0.007216 0.0080547 0.0053648 0.52309 0.21521 1.2856e-005 5.1731e-005 0.1477 0.53471 0.60366 0.0028908 0.55907 0.41439 0.0051282 0.42254 1.1054 1.0994 15.9957 144.9551 0.00058287 -77.4384 0.053943
4.158 0.98807 5.4983e-005 3.8183 0.011991 5.4453e-005 0.0011582 0.22768 0.00065926 0.22834 0.21054 0 0.032561 0.0389 0 1.1849 0.3817 0.11371 0.0146 7.2752 0.091097 0.00011387 0.79902 0.0072167 0.0080554 0.0049316 0.56289 0.23587 1.1726e-005 4.7146e-005 0.14771 0.53602 0.60578 0.00276 0.56049 0.41456 0.0045335 0.42248 1.1078 1.1018 15.9958 144.9551 0.00058079 -77.9564 0.054943
4.159 0.98807 5.4983e-005 3.8183 0.011991 5.4466e-005 0.0011582 0.22769 0.00065926 0.22834 0.21055 0 0.032561 0.0389 0 1.185 0.38174 0.11373 0.014601 7.2768 0.091107 0.00011388 0.79901 0.0072174 0.0080562 0.0045581 0.60185 0.25747 1.0758e-005 4.3233e-005 0.14771 0.53734 0.60789 0.0026434 0.56195 0.41472 0.0041041 0.42241 1.1102 1.1043 15.9959 144.9551 0.00057872 -78.44 0.055943
4.16 0.98807 5.4983e-005 3.8183 0.011991 5.4479e-005 0.0011582 0.22769 0.00065926 0.22835 0.21055 0 0.032561 0.0389 0 1.1851 0.38179 0.11375 0.014603 7.2784 0.091117 0.0001139 0.799 0.007218 0.0080569 0.0042358 0.6395 0.27985 9.9286e-006 3.9886e-005 0.14772 0.53867 0.60997 0.0025394 0.56346 0.41489 0.0037885 0.42235 1.1126 1.1067 15.996 144.9551 0.00057666 -78.8899 0.056943
4.161 0.98807 5.4983e-005 3.8183 0.011991 5.4492e-005 0.0011582 0.2277 0.00065926 0.22835 0.21056 0 0.03256 0.0389 0 1.1852 0.38184 0.11376 0.014605 7.28 0.091127 0.00011391 0.79899 0.0072187 0.0080577 0.0039565 0.67546 0.30288 9.2217e-006 3.7016e-005 0.14772 0.53999 0.61204 0.0024467 0.565 0.41506 0.003551 0.4223 1.115 1.1091 15.9961 144.955 0.00057461 -79.3071 0.057943
4.162 0.98807 5.4983e-005 3.8183 0.011991 5.4505e-005 0.0011582 0.2277 0.00065926 0.22836 0.21056 0 0.03256 0.0389 0 1.1853 0.38188 0.11378 0.014606 7.2816 0.091137 0.00011392 0.79898 0.0072194 0.0080584 0.0037145 0.7094 0.32639 8.6081e-006 3.4547e-005 0.14773 0.54132 0.61408 0.0023641 0.56659 0.41523 0.0033669 0.42225 1.1174 1.1115 15.9962 144.955 0.00057256 -79.6929 0.058943
4.163 0.98807 5.4983e-005 3.8183 0.011991 5.4518e-005 0.0011582 0.22771 0.00065926 0.22836 0.21057 0 0.03256 0.0389 0 1.1854 0.38193 0.11379 0.014608 7.2832 0.091147 0.00011394 0.79897 0.0072201 0.0080591 0.0035042 0.74107 0.35021 8.0792e-006 3.2417e-005 0.14773 0.54265 0.61611 0.0022904 0.56822 0.41541 0.0032197 0.4222 1.1198 1.1139 15.9963 144.955 0.00057052 -80.0485 0.059943
4.164 0.98807 5.4983e-005 3.8183 0.011991 5.4531e-005 0.0011582 0.22772 0.00065926 0.22837 0.21058 0 0.032559 0.0389 0 1.1855 0.38198 0.11381 0.01461 7.2848 0.091157 0.00011395 0.79896 0.0072208 0.0080599 0.0033211 0.7703 0.37421 7.6233e-006 3.0575e-005 0.14774 0.54398 0.61811 0.0022248 0.56988 0.41558 0.0030987 0.42216 1.1222 1.1163 15.9964 144.955 0.00056848 -80.3756 0.060943
4.165 0.98807 5.4983e-005 3.8183 0.011991 5.4544e-005 0.0011582 0.22772 0.00065926 0.22838 0.21058 0 0.032559 0.0389 0 1.1856 0.38202 0.11383 0.014611 7.2864 0.091168 0.00011397 0.79895 0.0072215 0.0080606 0.0031613 0.79701 0.39822 7.2269e-006 2.8977e-005 0.14774 0.54531 0.6201 0.0021662 0.57158 0.41575 0.002997 0.42211 1.1246 1.1188 15.9965 144.955 0.00056646 -80.6757 0.061943
4.166 0.98807 5.4982e-005 3.8183 0.011991 5.4557e-005 0.0011582 0.22773 0.00065926 0.22838 0.21059 0 0.032559 0.0389 0 1.1857 0.38207 0.11384 0.014613 7.288 0.091178 0.00011398 0.79894 0.0072222 0.0080614 0.0030217 0.82116 0.42212 6.8819e-006 2.7588e-005 0.14775 0.54663 0.62207 0.002114 0.57332 0.41593 0.0029101 0.42208 1.127 1.1212 15.9966 144.955 0.00056444 -80.9506 0.062943
4.167 0.98807 5.4982e-005 3.8183 0.011991 5.457e-005 0.0011582 0.22773 0.00065926 0.22839 0.21059 0 0.032559 0.0389 0 1.1858 0.38212 0.11386 0.014615 7.2896 0.091188 0.000114 0.79893 0.0072229 0.0080621 0.0028993 0.8428 0.44578 6.5809e-006 2.6377e-005 0.14776 0.54796 0.62402 0.0020673 0.57508 0.41611 0.0028346 0.42204 1.1294 1.1236 15.9967 144.955 0.00056243 -81.2018 0.063943
4.168 0.98807 5.4982e-005 3.8183 0.011991 5.4583e-005 0.0011582 0.22774 0.00065926 0.22839 0.2106 0 0.032558 0.0389 0 1.1859 0.38216 0.11387 0.014616 7.2912 0.091198 0.00011401 0.79892 0.0072236 0.0080628 0.0027918 0.86202 0.4691 6.3187e-006 2.5318e-005 0.14776 0.54929 0.62594 0.0020257 0.57688 0.41629 0.0027687 0.42201 1.1317 1.126 15.9968 144.955 0.00056044 -81.4311 0.064943
4.169 0.98807 5.4982e-005 3.8183 0.011991 5.4596e-005 0.0011582 0.22774 0.00065926 0.2284 0.2106 0 0.032558 0.0389 0 1.186 0.38221 0.11389 0.014618 7.2928 0.091208 0.00011402 0.79891 0.0072242 0.0080636 0.0026972 0.87896 0.49199 6.0883e-006 2.439e-005 0.14777 0.55061 0.62786 0.0019885 0.5787 0.41647 0.0027106 0.42198 1.1341 1.1283 15.9969 144.955 0.00055845 -81.6402 0.065943
4.17 0.98807 5.4982e-005 3.8183 0.011991 5.4609e-005 0.0011582 0.22775 0.00065926 0.2284 0.21061 0 0.032558 0.0389 0 1.1861 0.38225 0.11391 0.014619 7.2944 0.091218 0.00011404 0.7989 0.0072249 0.0080643 0.0026139 0.89377 0.51437 5.8853e-006 2.3574e-005 0.14777 0.55193 0.62975 0.0019552 0.58055 0.41665 0.0026594 0.42195 1.1365 1.1307 15.997 144.955 0.00055647 -81.8306 0.066943
4.171 0.98807 5.4982e-005 3.8183 0.011991 5.4622e-005 0.0011582 0.22776 0.00065926 0.22841 0.21061 0 0.032557 0.0389 0 1.1862 0.3823 0.11392 0.014621 7.296 0.091228 0.00011405 0.79889 0.0072256 0.0080651 0.0025402 0.90664 0.53617 5.7065e-006 2.2856e-005 0.14778 0.55325 0.63162 0.0019254 0.58242 0.41683 0.002614 0.42193 1.1389 1.1331 15.9971 144.9549 0.0005545 -82.0039 0.067943
4.172 0.98807 5.4982e-005 3.8183 0.011991 5.4635e-005 0.0011582 0.22776 0.00065926 0.22842 0.21062 0 0.032557 0.0389 0 1.1863 0.38235 0.11394 0.014623 7.2976 0.091239 0.00011407 0.79888 0.0072263 0.0080658 0.0024748 0.91776 0.55735 5.5493e-006 2.2221e-005 0.14778 0.55457 0.63348 0.0018987 0.58431 0.41701 0.0025736 0.4219 1.1412 1.1355 15.9972 144.9549 0.00055254 -82.1615 0.068943
4.173 0.98807 5.4982e-005 3.8183 0.011991 5.4648e-005 0.0011583 0.22777 0.00065926 0.22842 0.21062 0 0.032557 0.0389 0 1.1864 0.38239 0.11395 0.014624 7.2993 0.091249 0.00011408 0.79887 0.007227 0.0080665 0.0024169 0.9273 0.57787 5.4098e-006 2.166e-005 0.14779 0.55588 0.63532 0.0018747 0.58622 0.41719 0.0025376 0.42188 1.1436 1.1379 15.9973 144.9549 0.00055059 -82.3049 0.069943
4.174 0.98807 5.4982e-005 3.8183 0.011991 5.4661e-005 0.0011583 0.22777 0.00065926 0.22843 0.21063 0 0.032557 0.0389 0 1.1865 0.38244 0.11397 0.014626 7.3009 0.091259 0.00011409 0.79886 0.0072277 0.0080673 0.0023654 0.93546 0.5977 5.2856e-006 2.1162e-005 0.14779 0.55719 0.63715 0.0018532 0.58814 0.41737 0.0025055 0.42186 1.1459 1.1403 15.9974 144.9549 0.00054865 -82.4352 0.070943
4.175 0.98807 5.4982e-005 3.8183 0.011991 5.4674e-005 0.0011583 0.22778 0.00065926 0.22843 0.21063 0 0.032556 0.0389 0 1.1866 0.38249 0.11399 0.014628 7.3025 0.091269 0.00011411 0.79885 0.0072284 0.008068 0.0023195 0.94239 0.61682 5.1752e-006 2.0719e-005 0.1478 0.5585 0.63895 0.0018338 0.59008 0.41756 0.0024767 0.42184 1.1483 1.1426 15.9975 144.9549 0.00054672 -82.5538 0.071943
4.176 0.98807 5.4982e-005 3.8183 0.011991 5.4687e-005 0.0011583 0.22778 0.00065926 0.22844 0.21064 0 0.032556 0.0389 0 1.1867 0.38253 0.114 0.014629 7.3041 0.091279 0.00011412 0.79884 0.0072291 0.0080688 0.0022784 0.94828 0.63522 5.0772e-006 2.0324e-005 0.1478 0.55981 0.64074 0.0018164 0.59203 0.41774 0.002451 0.42182 1.1506 1.145 15.9976 144.9549 0.00054479 -82.6618 0.072943
4.177 0.98807 5.4982e-005 3.8183 0.011991 5.47e-005 0.0011583 0.22779 0.00065926 0.22844 0.21065 0 0.032556 0.0389 0 1.1868 0.38258 0.11402 0.014631 7.3057 0.091289 0.00011414 0.79882 0.0072297 0.0080695 0.0022416 0.95325 0.6529 4.9897e-006 1.9971e-005 0.14781 0.56111 0.64252 0.0018007 0.59399 0.41793 0.0024278 0.4218 1.153 1.1474 15.9977 144.9549 0.00054288 -82.76 0.073943
4.178 0.98807 5.4982e-005 3.8183 0.011991 5.4713e-005 0.0011583 0.2278 0.00065926 0.22845 0.21065 0 0.032555 0.0389 0 1.1869 0.38263 0.11403 0.014633 7.3073 0.091299 0.00011415 0.79881 0.0072304 0.0080702 0.0022086 0.95744 0.66985 4.9109e-006 1.9654e-005 0.14782 0.56241 0.64427 0.0017865 0.59595 0.41811 0.002407 0.42179 1.1553 1.1497 15.9978 144.9549 0.00054098 -82.8496 0.074943
4.179 0.98807 5.4982e-005 3.8183 0.011991 5.4726e-005 0.0011583 0.2278 0.00065926 0.22846 0.21066 0 0.032555 0.0389 0 1.187 0.38267 0.11405 0.014634 7.3089 0.091309 0.00011416 0.7988 0.0072311 0.008071 0.002179 0.96096 0.68609 4.8398e-006 1.937e-005 0.14782 0.56371 0.64601 0.0017736 0.59792 0.4183 0.0023883 0.42177 1.1577 1.1521 15.9979 144.9549 0.00053909 -82.9313 0.075943
4.18 0.98807 5.4981e-005 3.8183 0.011991 5.4739e-005 0.0011583 0.22781 0.00065926 0.22846 0.21066 0 0.032555 0.0389 0 1.1871 0.38272 0.11407 0.014636 7.3105 0.09132 0.00011418 0.79879 0.0072318 0.0080717 0.0021523 0.96392 0.70162 4.7758e-006 1.9114e-005 0.14783 0.565 0.64774 0.001762 0.5999 0.41848 0.0023714 0.42176 1.16 1.1545 15.998 144.9549 0.00053721 -83.0059 0.076943
4.181 0.98807 5.4981e-005 3.8183 0.011991 5.4752e-005 0.0011583 0.22781 0.00065926 0.22847 0.21067 0 0.032555 0.0389 0 1.1872 0.38277 0.11408 0.014637 7.3121 0.09133 0.00011419 0.79878 0.0072325 0.0080725 0.0021281 0.9664 0.71646 4.7184e-006 1.8883e-005 0.14783 0.56629 0.64945 0.0017514 0.60188 0.41867 0.002356 0.42175 1.1624 1.1568 15.9981 144.9549 0.00053534 -83.0742 0.077943
4.182 0.98807 5.4981e-005 3.8183 0.011991 5.4765e-005 0.0011583 0.22782 0.00065926 0.22847 0.21067 0 0.032554 0.0389 0 1.1873 0.38281 0.1141 0.014639 7.3137 0.09134 0.00011421 0.79877 0.0072332 0.0080732 0.002106 0.96849 0.73062 4.6667e-006 1.8673e-005 0.14784 0.56757 0.65114 0.0017417 0.60387 0.41886 0.0023421 0.42173 1.1647 1.1592 15.9982 144.9549 0.00053348 -83.1368 0.078943
4.183 0.98807 5.4981e-005 3.8183 0.011991 5.4778e-005 0.0011583 0.22782 0.00065926 0.22848 0.21068 0 0.032554 0.0389 0 1.1874 0.38286 0.11411 0.014641 7.3154 0.09135 0.00011422 0.79876 0.0072339 0.0080739 0.002086 0.97023 0.74413 4.6194e-006 1.8483e-005 0.14784 0.56886 0.65282 0.0017329 0.60585 0.41904 0.0023295 0.42172 1.167 1.1615 15.9983 144.9549 0.00053164 -83.1943 0.079943
4.184 0.98807 5.4981e-005 3.8183 0.011991 5.4791e-005 0.0011583 0.22783 0.00065926 0.22848 0.21068 0 0.032554 0.0389 0 1.1874 0.38291 0.11413 0.014642 7.317 0.09136 0.00011424 0.79875 0.0072346 0.0080747 0.0020679 0.9717 0.75699 4.576e-006 1.831e-005 0.14785 0.57013 0.65449 0.0017248 0.60784 0.41923 0.0023179 0.42171 1.1693 1.1639 15.9984 144.9549 0.0005298 -83.2471 0.080943
4.185 0.98807 5.4981e-005 3.8183 0.011991 5.4804e-005 0.0011583 0.22784 0.00065926 0.22849 0.21069 0 0.032553 0.0389 0 1.1875 0.38295 0.11415 0.014644 7.3186 0.09137 0.00011425 0.79874 0.0072352 0.0080754 0.0020514 0.97293 0.76924 4.5362e-006 1.8152e-005 0.14785 0.57141 0.65613 0.0017174 0.60982 0.41942 0.0023074 0.4217 1.1717 1.1662 15.9985 144.9549 0.00052797 -83.2959 0.081943
4.186 0.98807 5.4981e-005 3.8183 0.011991 5.4817e-005 0.0011583 0.22784 0.00065926 0.2285 0.21069 0 0.032553 0.0389 0 1.1876 0.383 0.11416 0.014646 7.3202 0.09138 0.00011426 0.79873 0.0072359 0.0080762 0.0020359 0.97397 0.78089 4.5003e-006 1.8007e-005 0.14786 0.57268 0.65777 0.0017106 0.61181 0.41961 0.0022977 0.42169 1.174 1.1685 15.9986 144.955 0.00052615 -83.3409 0.082943
4.187 0.98807 5.4981e-005 3.8183 0.011991 5.483e-005 0.0011583 0.22785 0.00065926 0.2285 0.2107 0 0.032553 0.0389 0 1.1877 0.38305 0.11418 0.014647 7.3218 0.09139 0.00011428 0.79872 0.0072366 0.0080769 0.0020218 0.97485 0.79197 4.4674e-006 1.7873e-005 0.14787 0.57395 0.65939 0.0017043 0.61379 0.41979 0.0022889 0.42168 1.1763 1.1709 15.9987 144.955 0.00052434 -83.3827 0.083943
4.188 0.98807 5.4981e-005 3.8183 0.011991 5.4843e-005 0.0011583 0.22785 0.00065926 0.22851 0.2107 0 0.032553 0.0389 0 1.1878 0.38309 0.11419 0.014649 7.3234 0.091401 0.00011429 0.79871 0.0072373 0.0080776 0.0020091 0.97559 0.8025 4.4364e-006 1.775e-005 0.14787 0.57521 0.66099 0.0016985 0.61577 0.41998 0.0022807 0.42167 1.1786 1.1732 15.9988 144.955 0.00052254 -83.4214 0.084943
4.189 0.98807 5.4981e-005 3.8183 0.011991 5.4856e-005 0.0011583 0.22786 0.00065926 0.22851 0.21071 0 0.032552 0.0389 0 1.1879 0.38314 0.11421 0.01465 7.325 0.091411 0.00011431 0.7987 0.007238 0.0080784 0.0019973 0.97622 0.8125 4.4078e-006 1.7637e-005 0.14788 0.57647 0.66258 0.0016931 0.61775 0.42017 0.0022731 0.42166 1.1809 1.1755 15.9989 144.955 0.00052075 -83.4575 0.085943
4.19 0.98807 5.4981e-005 3.8183 0.011991 5.4869e-005 0.0011583 0.22786 0.00065926 0.22852 0.21072 0 0.032552 0.0389 0 1.188 0.38319 0.11423 0.014652 7.3266 0.091421 0.00011432 0.79869 0.0072387 0.0080791 0.001986 0.97675 0.82199 4.3818e-006 1.7531e-005 0.14788 0.57773 0.66416 0.0016881 0.61972 0.42036 0.0022661 0.42165 1.1832 1.1778 15.999 144.955 0.00051897 -83.4913 0.086943
4.191 0.98807 5.4981e-005 3.8183 0.011991 5.4882e-005 0.0011583 0.22787 0.00065926 0.22852 0.21072 0 0.032552 0.0389 0 1.1881 0.38323 0.11424 0.014654 7.3283 0.091431 0.00011433 0.79868 0.0072394 0.0080798 0.0019755 0.97721 0.831 4.3575e-006 1.7433e-005 0.14789 0.57899 0.66572 0.0016834 0.62169 0.42055 0.0022596 0.42164 1.1855 1.1801 15.9991 144.955 0.0005172 -83.5229 0.087943
4.192 0.98807 5.4981e-005 3.8183 0.011991 5.4895e-005 0.0011583 0.22787 0.00065926 0.22853 0.21073 0 0.032551 0.0389 0 1.1882 0.38328 0.11426 0.014655 7.3299 0.091441 0.00011435 0.79867 0.00724 0.0080806 0.0019657 0.97761 0.83955 4.3346e-006 1.7341e-005 0.14789 0.58023 0.66727 0.001679 0.62366 0.42073 0.0022535 0.42163 1.1878 1.1825 15.9992 144.955 0.00051544 -83.5526 0.088943
4.193 0.98807 5.4981e-005 3.8183 0.011991 5.4908e-005 0.0011583 0.22788 0.00065926 0.22854 0.21073 0 0.032551 0.0389 0 1.1883 0.38333 0.11427 0.014657 7.3315 0.091451 0.00011436 0.79866 0.0072407 0.0080813 0.0019566 0.97795 0.84765 4.3131e-006 1.7255e-005 0.1479 0.58148 0.66881 0.0016749 0.62562 0.42092 0.0022478 0.42163 1.1901 1.1848 15.9993 144.955 0.00051369 -83.5805 0.089943
4.194 0.98807 5.498e-005 3.8183 0.011991 5.4921e-005 0.0011583 0.22789 0.00065926 0.22854 0.21074 0 0.032551 0.0389 0 1.1884 0.38337 0.11429 0.014659 7.3331 0.091461 0.00011438 0.79865 0.0072414 0.0080821 0.0019483 0.97825 0.85533 4.2927e-006 1.7174e-005 0.1479 0.58272 0.67033 0.001671 0.62757 0.42111 0.0022424 0.42162 1.1924 1.1871 15.9994 144.955 0.00051195 -83.607 0.090943
4.195 0.98807 5.498e-005 3.8183 0.011991 5.4934e-005 0.0011583 0.22789 0.00065926 0.22855 0.21074 0 0.032551 0.0389 0 1.1885 0.38342 0.11431 0.01466 7.3347 0.091471 0.00011439 0.79864 0.0072421 0.0080828 0.0019403 0.97851 0.86261 4.2736e-006 1.7098e-005 0.14791 0.58396 0.67184 0.0016673 0.62953 0.4213 0.0022373 0.42161 1.1947 1.1894 15.9995 144.955 0.00051022 -83.632 0.091943
4.196 0.98807 5.498e-005 3.8183 0.011991 5.4947e-005 0.0011583 0.2279 0.00065926 0.22855 0.21075 0 0.03255 0.0389 0 1.1886 0.38347 0.11432 0.014662 7.3363 0.091481 0.0001144 0.79863 0.0072428 0.0080835 0.0019325 0.97874 0.8695 4.2558e-006 1.7026e-005 0.14791 0.5852 0.67334 0.0016638 0.63147 0.42149 0.0022326 0.42161 1.1969 1.1917 15.9996 144.955 0.0005085 -83.6559 0.092943
4.197 0.98807 5.498e-005 3.8183 0.011991 5.496e-005 0.0011583 0.2279 0.00065926 0.22856 0.21075 0 0.03255 0.0389 0 1.1887 0.38351 0.11434 0.014664 7.3379 0.091492 0.00011442 0.79862 0.0072435 0.0080843 0.0019251 0.97894 0.87604 4.2388e-006 1.6957e-005 0.14792 0.58643 0.67482 0.0016605 0.63341 0.42168 0.002228 0.4216 1.1992 1.194 15.9997 144.955 0.00050679 -83.6786 0.093943
4.198 0.98807 5.498e-005 3.8183 0.011991 5.4973e-005 0.0011583 0.22791 0.00065926 0.22856 0.21076 0 0.03255 0.0389 0 1.1888 0.38356 0.11435 0.014665 7.3396 0.091502 0.00011443 0.79861 0.0072442 0.008085 0.001918 0.97912 0.88222 4.2226e-006 1.6892e-005 0.14793 0.58766 0.67629 0.0016573 0.63534 0.42187 0.0022237 0.42159 1.2015 1.1963 15.9997 144.955 0.00050509 -83.7003 0.094943
4.199 0.98807 5.498e-005 3.8183 0.011991 5.4986e-005 0.0011583 0.22791 0.00065926 0.22857 0.21076 0 0.032549 0.0389 0 1.1889 0.38361 0.11437 0.014667 7.3412 0.091512 0.00011445 0.7986 0.0072449 0.0080858 0.0019114 0.97929 0.88808 4.207e-006 1.683e-005 0.14793 0.58888 0.67775 0.0016543 0.63727 0.42206 0.0022196 0.42159 1.2038 1.1986 15.9998 144.955 0.0005034 -83.7211 0.095943
4.2 0.98807 5.498e-005 3.8183 0.011991 5.4999e-005 0.0011583 0.22792 0.00065926 0.22857 0.21077 0 0.032549 0.0389 0 1.189 0.38365 0.11439 0.014668 7.3428 0.091522 0.00011446 0.79859 0.0072455 0.0080865 0.0019052 0.97944 0.89362 4.192e-006 1.677e-005 0.14794 0.5901 0.6792 0.0016514 0.63919 0.42225 0.0022157 0.42158 1.206 1.2008 15.9999 144.955 0.00050171 -83.7411 0.096943
4.201 0.98807 5.498e-005 3.8183 0.011991 5.5012e-005 0.0011583 0.22793 0.00065926 0.22858 0.21077 0 0.032549 0.0389 0 1.1891 0.3837 0.1144 0.01467 7.3444 0.091532 0.00011447 0.79858 0.0072462 0.0080872 0.0018992 0.97957 0.89887 4.1776e-006 1.6713e-005 0.14794 0.59132 0.68063 0.0016486 0.6411 0.42243 0.002212 0.42158 1.2083 1.2031 16 144.955 0.00050004 -83.7603 0.097943
4.202 0.98807 5.498e-005 3.8183 0.011991 5.5025e-005 0.0011583 0.22793 0.00065926 0.22859 0.21078 0 0.032549 0.0389 0 1.1892 0.38375 0.11442 0.014672 7.346 0.091542 0.00011449 0.79857 0.0072469 0.008088 0.0018934 0.9797 0.90384 4.1639e-006 1.6658e-005 0.14795 0.59253 0.68206 0.0016459 0.64301 0.42262 0.0022084 0.42157 1.2106 1.2054 16.0001 144.955 0.00049838 -83.7789 0.098943
4.203 0.98807 5.498e-005 3.8183 0.011991 5.5038e-005 0.0011583 0.22794 0.00065926 0.22859 0.21078 0 0.032548 0.0389 0 1.1893 0.38379 0.11443 0.014673 7.3477 0.091552 0.0001145 0.79856 0.0072476 0.0080887 0.0018878 0.97981 0.90854 4.1508e-006 1.6605e-005 0.14795 0.59374 0.68347 0.0016433 0.64491 0.42281 0.0022049 0.42157 1.2128 1.2077 16.0002 144.955 0.00049672 -83.7969 0.099943
4.204 0.98807 5.498e-005 3.8183 0.011991 5.5051e-005 0.0011583 0.22794 0.00065926 0.2286 0.21079 0 0.032548 0.0389 0 1.1894 0.38384 0.11445 0.014675 7.3493 0.091562 0.00011452 0.79855 0.0072483 0.0080894 0.0018824 0.97992 0.91298 4.138e-006 1.6554e-005 0.14796 0.59495 0.68486 0.0016408 0.64681 0.423 0.0022015 0.42156 1.2151 1.2099 16.0003 144.9551 0.00049507 -83.8144 0.10094
4.205 0.98807 5.498e-005 3.8183 0.011991 5.5064e-005 0.0011583 0.22795 0.00065926 0.2286 0.2108 0 0.032548 0.0389 0 1.1895 0.38389 0.11447 0.014677 7.3509 0.091572 0.00011453 0.79854 0.007249 0.0080902 0.001877 0.98002 0.91718 4.1254e-006 1.6504e-005 0.14796 0.59615 0.68625 0.0016384 0.64869 0.42319 0.0021983 0.42156 1.2173 1.2122 16.0004 144.9551 0.00049344 -83.8313 0.10194
4.206 0.98807 5.498e-005 3.8183 0.011991 5.5077e-005 0.0011583 0.22795 0.00065926 0.22861 0.2108 0 0.032547 0.0389 0 1.1896 0.38393 0.11448 0.014678 7.3525 0.091582 0.00011455 0.79853 0.0072497 0.0080909 0.0018718 0.98012 0.92116 4.1133e-006 1.6456e-005 0.14797 0.59735 0.68763 0.001636 0.65057 0.42338 0.0021951 0.42155 1.2195 1.2145 16.0005 144.9551 0.00049181 -83.8478 0.10294
4.207 0.98807 5.498e-005 3.8183 0.011991 5.509e-005 0.0011583 0.22796 0.00065926 0.22861 0.21081 0 0.032547 0.0389 0 1.1897 0.38398 0.1145 0.01468 7.3541 0.091593 0.00011456 0.79852 0.0072503 0.0080917 0.0018667 0.98021 0.92492 4.1016e-006 1.6409e-005 0.14798 0.59854 0.68899 0.0016337 0.65245 0.42357 0.002192 0.42155 1.2218 1.2167 16.0006 144.9551 0.00049019 -83.8639 0.10394
4.208 0.98807 5.4979e-005 3.8183 0.011991 5.5103e-005 0.0011583 0.22796 0.00065926 0.22862 0.21081 0 0.032547 0.0389 0 1.1898 0.38403 0.11451 0.014681 7.3558 0.091603 0.00011457 0.79851 0.007251 0.0080924 0.0018618 0.98029 0.92848 4.0903e-006 1.6364e-005 0.14798 0.59973 0.69034 0.0016315 0.65431 0.42376 0.002189 0.42154 1.224 1.219 16.0006 144.9551 0.00048858 -83.8796 0.10494
4.209 0.98807 5.4979e-005 3.8183 0.011991 5.5116e-005 0.0011583 0.22797 0.00065926 0.22862 0.21082 0 0.032547 0.0389 0 1.1899 0.38407 0.11453 0.014683 7.3574 0.091613 0.00011459 0.7985 0.0072517 0.0080931 0.0018572 0.98037 0.93184 4.0794e-006 1.6319e-005 0.14799 0.60092 0.69168 0.0016293 0.65617 0.42395 0.0021861 0.42154 1.2263 1.2212 16.0007 144.9551 0.00048698 -83.8949 0.10594
4.21 0.98807 5.4979e-005 3.8183 0.011991 5.5129e-005 0.0011583 0.22798 0.00065926 0.22863 0.21082 0 0.032546 0.0389 0 1.19 0.38412 0.11455 0.014685 7.359 0.091623 0.0001146 0.79849 0.0072524 0.0080939 0.0018525 0.98045 0.93502 4.0686e-006 1.6276e-005 0.14799 0.60211 0.69301 0.0016271 0.65802 0.42414 0.0021833 0.42154 1.2285 1.2235 16.0008 144.9551 0.00048539 -83.91 0.10694
4.211 0.98807 5.4979e-005 3.8183 0.011991 5.5142e-005 0.0011583 0.22798 0.00065926 0.22864 0.21083 0 0.032546 0.0389 0 1.1901 0.38417 0.11456 0.014686 7.3606 0.091633 0.00011462 0.79848 0.0072531 0.0080946 0.001848 0.98053 0.93802 4.058e-006 1.6233e-005 0.148 0.60329 0.69433 0.001625 0.65987 0.42433 0.0021805 0.42153 1.2307 1.2257 16.0009 144.9551 0.0004838 -83.9247 0.10794
4.212 0.98807 5.4979e-005 3.8183 0.011991 5.5155e-005 0.0011583 0.22799 0.00065926 0.22864 0.21083 0 0.032546 0.0389 0 1.1902 0.38421 0.11458 0.014688 7.3622 0.091643 0.00011463 0.79847 0.0072538 0.0080953 0.0018436 0.9806 0.94086 4.0476e-006 1.6191e-005 0.148 0.60446 0.69564 0.001623 0.6617 0.42452 0.0021778 0.42153 1.2329 1.2279 16.001 144.9551 0.00048223 -83.9392 0.10894
4.213 0.98807 5.4979e-005 3.8183 0.01199 5.5168e-005 0.0011583 0.22799 0.00065926 0.22865 0.21084 0 0.032545 0.0389 0 1.1903 0.38426 0.11459 0.01469 7.3639 0.091653 0.00011464 0.79846 0.0072545 0.0080961 0.0018393 0.98067 0.94355 4.0373e-006 1.6151e-005 0.14801 0.60564 0.69694 0.001621 0.66353 0.42471 0.0021751 0.42152 1.2351 1.2302 16.0011 144.9551 0.00048066 -83.9534 0.10994
4.214 0.98807 5.4979e-005 3.8183 0.01199 5.5181e-005 0.0011583 0.228 0.00065926 0.22865 0.21084 0 0.032545 0.0389 0 1.1904 0.38431 0.11461 0.014691 7.3655 0.091663 0.00011466 0.79845 0.0072551 0.0080968 0.001835 0.98074 0.94608 4.0273e-006 1.6111e-005 0.14801 0.60681 0.69823 0.001619 0.66535 0.4249 0.0021725 0.42152 1.2374 1.2324 16.0011 144.9551 0.00047911 -83.9674 0.11094
4.215 0.98807 5.4979e-005 3.8183 0.01199 5.5194e-005 0.0011584 0.228 0.00065926 0.22866 0.21085 0 0.032545 0.0389 0 1.1905 0.38435 0.11462 0.014693 7.3671 0.091673 0.00011467 0.79844 0.0072558 0.0080976 0.0018308 0.98081 0.94848 4.0175e-006 1.6071e-005 0.14802 0.60797 0.6995 0.001617 0.66717 0.42509 0.0021699 0.42152 1.2396 1.2346 16.0012 144.9551 0.00047756 -83.9812 0.11194
4.216 0.98807 5.4979e-005 3.8183 0.01199 5.5207e-005 0.0011584 0.22801 0.00065926 0.22866 0.21085 0 0.032545 0.0389 0 1.1906 0.3844 0.11464 0.014695 7.3687 0.091683 0.00011469 0.79843 0.0072565 0.0080983 0.0018267 0.98087 0.95075 4.0079e-006 1.6033e-005 0.14802 0.60914 0.70077 0.0016151 0.66897 0.42528 0.0021674 0.42152 1.2418 1.2368 16.0013 144.9551 0.00047602 -83.9947 0.11294
4.217 0.98807 5.4979e-005 3.8183 0.01199 5.522e-005 0.0011584 0.22801 0.00065926 0.22867 0.21086 0 0.032544 0.0389 0 1.1907 0.38445 0.11466 0.014696 7.3704 0.091694 0.0001147 0.79842 0.0072572 0.008099 0.0018226 0.98093 0.95289 3.9985e-006 1.5995e-005 0.14803 0.6103 0.70203 0.0016132 0.67077 0.42547 0.0021649 0.42151 1.244 1.2391 16.0014 144.9551 0.00047448 -84.0081 0.11394
4.218 0.98807 5.4979e-005 3.8183 0.01199 5.5233e-005 0.0011584 0.22802 0.00065926 0.22867 0.21086 0 0.032544 0.0389 0 1.1908 0.38449 0.11467 0.014698 7.372 0.091704 0.00011471 0.79841 0.0072579 0.0080998 0.0018186 0.98099 0.95491 3.9891e-006 1.5958e-005 0.14804 0.61145 0.70327 0.0016114 0.67257 0.42566 0.0021625 0.42151 1.2462 1.2413 16.0015 144.9552 0.00047296 -84.0213 0.11494
4.219 0.98807 5.4979e-005 3.8183 0.01199 5.5246e-005 0.0011584 0.22803 0.00065926 0.22868 0.21087 0 0.032544 0.0389 0 1.1909 0.38454 0.11469 0.014699 7.3736 0.091714 0.00011473 0.7984 0.0072586 0.0081005 0.0018147 0.98105 0.95682 3.98e-006 1.5921e-005 0.14804 0.6126 0.70451 0.0016095 0.67435 0.42585 0.0021601 0.42151 1.2484 1.2435 16.0016 144.9552 0.00047144 -84.0343 0.11594
4.22 0.98807 5.4979e-005 3.8183 0.01199 5.5259e-005 0.0011584 0.22803 0.00065926 0.22869 0.21087 0 0.032544 0.0389 0 1.191 0.38459 0.1147 0.014701 7.3752 0.091724 0.00011474 0.79839 0.0072592 0.0081012 0.0018109 0.98111 0.95863 3.9709e-006 1.5885e-005 0.14805 0.61375 0.70574 0.0016077 0.67613 0.42604 0.0021577 0.42151 1.2505 1.2457 16.0016 144.9552 0.00046994 -84.0471 0.11694
4.221 0.98807 5.4979e-005 3.8183 0.01199 5.5272e-005 0.0011584 0.22804 0.00065926 0.22869 0.21088 0 0.032543 0.0389 0 1.1911 0.38463 0.11472 0.014703 7.3768 0.091734 0.00011476 0.79838 0.0072599 0.008102 0.0018071 0.98117 0.96034 3.962e-006 1.5849e-005 0.14805 0.6149 0.70695 0.0016059 0.6779 0.42623 0.0021554 0.4215 1.2527 1.2479 16.0017 144.9552 0.00046844 -84.0598 0.11794
4.222 0.98807 5.4978e-005 3.8183 0.01199 5.5285e-005 0.0011584 0.22804 0.00065926 0.2287 0.21088 0 0.032543 0.0389 0 1.1912 0.38468 0.11474 0.014704 7.3785 0.091744 0.00011477 0.79837 0.0072606 0.0081027 0.0018033 0.98122 0.96195 3.9532e-006 1.5814e-005 0.14806 0.61604 0.70816 0.0016042 0.67966 0.42641 0.002153 0.4215 1.2549 1.2501 16.0018 144.9552 0.00046695 -84.0723 0.11894
4.223 0.98807 5.4978e-005 3.8183 0.01199 5.5298e-005 0.0011584 0.22805 0.00065926 0.2287 0.21089 0 0.032543 0.0389 0 1.1913 0.38473 0.11475 0.014706 7.3801 0.091754 0.00011478 0.79836 0.0072613 0.0081034 0.0017996 0.98128 0.96347 3.9446e-006 1.5779e-005 0.14806 0.61718 0.70936 0.0016024 0.68141 0.4266 0.0021508 0.4215 1.2571 1.2523 16.0019 144.9552 0.00046546 -84.0847 0.11994
4.224 0.98807 5.4978e-005 3.8183 0.01199 5.5311e-005 0.0011584 0.22805 0.00065926 0.22871 0.21089 0 0.032542 0.0389 0 1.1914 0.38477 0.11477 0.014708 7.3817 0.091764 0.0001148 0.79835 0.007262 0.0081042 0.0017959 0.98133 0.96491 3.9361e-006 1.5745e-005 0.14807 0.61831 0.71055 0.0016007 0.68316 0.42679 0.0021485 0.4215 1.2593 1.2545 16.002 144.9552 0.00046399 -84.097 0.12094
4.225 0.98807 5.4978e-005 3.8183 0.01199 5.5324e-005 0.0011584 0.22806 0.00065926 0.22871 0.2109 0 0.032542 0.0389 0 1.1915 0.38482 0.11478 0.014709 7.3834 0.091774 0.00011481 0.79834 0.0072627 0.0081049 0.0017923 0.98139 0.96627 3.9276e-006 1.5711e-005 0.14807 0.61944 0.71173 0.001599 0.6849 0.42698 0.0021463 0.4215 1.2614 1.2567 16.002 144.9552 0.00046252 -84.1091 0.12194
4.226 0.98807 5.4978e-005 3.8183 0.01199 5.5337e-005 0.0011584 0.22806 0.00065926 0.22872 0.21091 0 0.032542 0.0389 0 1.1916 0.38486 0.1148 0.014711 7.385 0.091784 0.00011483 0.79833 0.0072634 0.0081057 0.0017888 0.98144 0.96755 3.9193e-006 1.5678e-005 0.14808 0.62057 0.7129 0.0015973 0.68663 0.42717 0.0021441 0.4215 1.2636 1.2588 16.0021 144.9552 0.00046106 -84.1211 0.12294
4.227 0.98807 5.4978e-005 3.8183 0.01199 5.535e-005 0.0011584 0.22807 0.00065926 0.22872 0.21091 0 0.032542 0.0389 0 1.1917 0.38491 0.11482 0.014712 7.3866 0.091794 0.00011484 0.79832 0.007264 0.0081064 0.0017852 0.98149 0.96876 3.9111e-006 1.5645e-005 0.14808 0.6217 0.71406 0.0015957 0.68836 0.42736 0.0021419 0.42149 1.2657 1.261 16.0022 144.9552 0.00045961 -84.133 0.12394
4.228 0.98807 5.4978e-005 3.8183 0.01199 5.5363e-005 0.0011584 0.22807 0.00065926 0.22873 0.21092 0 0.032541 0.0389 0 1.1918 0.38496 0.11483 0.014714 7.3882 0.091804 0.00011485 0.79831 0.0072647 0.0081071 0.0017818 0.98154 0.96991 3.9029e-006 1.5613e-005 0.14809 0.62282 0.71521 0.001594 0.69007 0.42755 0.0021398 0.42149 1.2679 1.2632 16.0023 144.9552 0.00045817 -84.1447 0.12494
4.229 0.98807 5.4978e-005 3.8183 0.01199 5.5376e-005 0.0011584 0.22808 0.00065926 0.22873 0.21092 0 0.032541 0.0389 0 1.1919 0.385 0.11485 0.014716 7.3899 0.091815 0.00011487 0.7983 0.0072654 0.0081079 0.0017783 0.98159 0.97099 3.8949e-006 1.5581e-005 0.1481 0.62393 0.71636 0.0015924 0.69178 0.42774 0.0021376 0.42149 1.2701 1.2653 16.0023 144.9553 0.00045673 -84.1564 0.12594
4.23 0.98807 5.4978e-005 3.8183 0.01199 5.5389e-005 0.0011584 0.22809 0.00065926 0.22874 0.21093 0 0.032541 0.0389 0 1.192 0.38505 0.11486 0.014717 7.3915 0.091825 0.00011488 0.79829 0.0072661 0.0081086 0.0017749 0.98164 0.97201 3.8869e-006 1.5549e-005 0.1481 0.62505 0.71749 0.0015908 0.69349 0.42793 0.0021355 0.42149 1.2722 1.2675 16.0024 144.9553 0.00045531 -84.1679 0.12694
4.231 0.98807 5.4978e-005 3.8183 0.01199 5.5402e-005 0.0011584 0.22809 0.00065926 0.22875 0.21093 0 0.03254 0.0389 0 1.1921 0.3851 0.11488 0.014719 7.3931 0.091835 0.0001149 0.79828 0.0072668 0.0081093 0.0017715 0.98169 0.97298 3.8791e-006 1.5517e-005 0.14811 0.62616 0.71862 0.0015892 0.69518 0.42812 0.0021335 0.42149 1.2743 1.2697 16.0025 144.9553 0.00045389 -84.1793 0.12794
4.232 0.98807 5.4978e-005 3.8183 0.01199 5.5415e-005 0.0011584 0.2281 0.00065926 0.22875 0.21094 0 0.03254 0.0389 0 1.1922 0.38514 0.1149 0.014721 7.3948 0.091845 0.00011491 0.79827 0.0072675 0.0081101 0.0017682 0.98174 0.97389 3.8713e-006 1.5486e-005 0.14811 0.62727 0.71973 0.0015876 0.69687 0.42831 0.0021314 0.42149 1.2765 1.2718 16.0026 144.9553 0.00045247 -84.1906 0.12894
4.233 0.98807 5.4978e-005 3.8183 0.01199 5.5428e-005 0.0011584 0.2281 0.00065926 0.22876 0.21094 0 0.03254 0.0389 0 1.1923 0.38519 0.11491 0.014722 7.3964 0.091855 0.00011492 0.79826 0.0072681 0.0081108 0.0017649 0.98179 0.97475 3.8637e-006 1.5456e-005 0.14812 0.62837 0.72084 0.0015861 0.69855 0.4285 0.0021294 0.42149 1.2786 1.274 16.0026 144.9553 0.00045107 -84.2018 0.12994
4.234 0.98807 5.4978e-005 3.8183 0.01199 5.5441e-005 0.0011584 0.22811 0.00065926 0.22876 0.21095 0 0.03254 0.0389 0 1.1924 0.38524 0.11493 0.014724 7.398 0.091865 0.00011494 0.79825 0.0072688 0.0081115 0.0017617 0.98183 0.97556 3.8561e-006 1.5425e-005 0.14812 0.62947 0.72194 0.0015845 0.70022 0.42869 0.0021273 0.42149 1.2808 1.2761 16.0027 144.9553 0.00044967 -84.213 0.13094
4.235 0.98807 5.4978e-005 3.8183 0.01199 5.5454e-005 0.0011584 0.22811 0.00065926 0.22877 0.21095 0 0.032539 0.0389 0 1.1925 0.38528 0.11494 0.014725 7.3996 0.091875 0.00011495 0.79824 0.0072695 0.0081123 0.0017584 0.98188 0.97633 3.8486e-006 1.5395e-005 0.14813 0.63057 0.72304 0.001583 0.70188 0.42888 0.0021254 0.42149 1.2829 1.2783 16.0028 144.9553 0.00044828 -84.224 0.13194
4.236 0.98807 5.4977e-005 3.8183 0.01199 5.5467e-005 0.0011584 0.22812 0.00065926 0.22877 0.21096 0 0.032539 0.0389 0 1.1926 0.38533 0.11496 0.014727 7.4013 0.091885 0.00011497 0.79823 0.0072702 0.008113 0.0017553 0.98193 0.97706 3.8411e-006 1.5365e-005 0.14813 0.63166 0.72412 0.0015815 0.70354 0.42907 0.0021234 0.42149 1.285 1.2804 16.0029 144.9553 0.0004469 -84.2349 0.13294
4.237 0.98807 5.4977e-005 3.8183 0.01199 5.548e-005 0.0011584 0.22812 0.00065926 0.22878 0.21096 0 0.032539 0.0389 0 1.1927 0.38538 0.11498 0.014729 7.4029 0.091895 0.00011498 0.79822 0.0072709 0.0081137 0.0017521 0.98197 0.97775 3.8338e-006 1.5336e-005 0.14814 0.63275 0.7252 0.00158 0.70519 0.42926 0.0021214 0.42149 1.2871 1.2825 16.0029 144.9553 0.00044552 -84.2457 0.13394
4.238 0.98807 5.4977e-005 3.8183 0.01199 5.5493e-005 0.0011584 0.22813 0.00065926 0.22878 0.21097 0 0.032539 0.0389 0 1.1928 0.38542 0.11499 0.01473 7.4045 0.091905 0.000115 0.79821 0.0072716 0.0081145 0.001749 0.98202 0.97839 3.8265e-006 1.5307e-005 0.14814 0.63384 0.72626 0.0015785 0.70683 0.42945 0.0021195 0.42149 1.2892 1.2847 16.003 144.9553 0.00044415 -84.2564 0.13494
4.239 0.98807 5.4977e-005 3.8183 0.01199 5.5506e-005 0.0011584 0.22813 0.00065927 0.22879 0.21097 0 0.032538 0.0389 0 1.1928 0.38547 0.11501 0.014732 7.4062 0.091915 0.00011501 0.7982 0.0072722 0.0081152 0.0017459 0.98206 0.97901 3.8193e-006 1.5278e-005 0.14815 0.63493 0.72732 0.0015771 0.70847 0.42964 0.0021176 0.42149 1.2914 1.2868 16.0031 144.9553 0.00044279 -84.2671 0.13594
4.24 0.98807 5.4977e-005 3.8183 0.01199 5.5519e-005 0.0011584 0.22814 0.00065927 0.22879 0.21098 0 0.032538 0.0389 0 1.1929 0.38552 0.11502 0.014734 7.4078 0.091925 0.00011502 0.79819 0.0072729 0.008116 0.0017428 0.9821 0.97959 3.8122e-006 1.525e-005 0.14816 0.63601 0.72837 0.0015756 0.71009 0.42983 0.0021157 0.42149 1.2935 1.2889 16.0031 144.9554 0.00044144 -84.2776 0.13694
4.241 0.98807 5.4977e-005 3.8183 0.01199 5.5532e-005 0.0011584 0.22814 0.00065927 0.2288 0.21098 0 0.032538 0.0389 0 1.193 0.38556 0.11504 0.014735 7.4094 0.091935 0.00011504 0.79818 0.0072736 0.0081167 0.0017398 0.98215 0.98013 3.8051e-006 1.5221e-005 0.14816 0.63708 0.72942 0.0015742 0.71171 0.43002 0.0021138 0.42149 1.2956 1.291 16.0032 144.9554 0.0004401 -84.2881 0.13794
4.242 0.98807 5.4977e-005 3.8183 0.01199 5.5545e-005 0.0011584 0.22815 0.00065927 0.2288 0.21099 0 0.032537 0.0389 0 1.1931 0.38561 0.11506 0.014737 7.4111 0.091945 0.00011505 0.79817 0.0072743 0.0081174 0.0017368 0.98219 0.98065 3.7982e-006 1.5193e-005 0.14817 0.63816 0.73046 0.0015727 0.71332 0.43021 0.0021119 0.42149 1.2977 1.2932 16.0033 144.9554 0.00043876 -84.2985 0.13894
4.243 0.98807 5.4977e-005 3.8183 0.01199 5.5558e-005 0.0011584 0.22816 0.00065927 0.22881 0.21099 0 0.032537 0.0389 0 1.1932 0.38566 0.11507 0.014738 7.4127 0.091956 0.00011507 0.79816 0.007275 0.0081182 0.0017338 0.98223 0.98114 3.7912e-006 1.5166e-005 0.14817 0.63923 0.73148 0.0015713 0.71493 0.4304 0.00211 0.42149 1.2998 1.2953 16.0034 144.9554 0.00043742 -84.3087 0.13994
4.244 0.98807 5.4977e-005 3.8183 0.01199 5.5571e-005 0.0011584 0.22816 0.00065927 0.22882 0.211 0 0.032537 0.0389 0 1.1933 0.3857 0.11509 0.01474 7.4143 0.091966 0.00011508 0.79815 0.0072757 0.0081189 0.0017309 0.98227 0.9816 3.7844e-006 1.5138e-005 0.14818 0.6403 0.73251 0.0015699 0.71653 0.43059 0.0021082 0.42149 1.3018 1.2974 16.0034 144.9554 0.0004361 -84.3189 0.14094
4.245 0.98807 5.4977e-005 3.8183 0.01199 5.5584e-005 0.0011584 0.22817 0.00065927 0.22882 0.211 0 0.032537 0.0389 0 1.1934 0.38575 0.1151 0.014742 7.416 0.091976 0.00011509 0.79814 0.0072763 0.0081196 0.001728 0.98232 0.98203 3.7776e-006 1.5111e-005 0.14818 0.64136 0.73352 0.0015685 0.71812 0.43078 0.0021064 0.42149 1.3039 1.2995 16.0035 144.9554 0.00043478 -84.3291 0.14194
4.246 0.98807 5.4977e-005 3.8183 0.01199 5.5597e-005 0.0011584 0.22817 0.00065927 0.22883 0.21101 0 0.032536 0.0389 0 1.1935 0.3858 0.11512 0.014743 7.4176 0.091986 0.00011511 0.79813 0.007277 0.0081204 0.0017251 0.98236 0.98245 3.7709e-006 1.5085e-005 0.14819 0.64242 0.73453 0.0015672 0.7197 0.43097 0.0021046 0.42149 1.306 1.3016 16.0036 144.9554 0.00043347 -84.3391 0.14294
4.247 0.98807 5.4977e-005 3.8183 0.01199 5.561e-005 0.0011584 0.22818 0.00065927 0.22883 0.21101 0 0.032536 0.0389 0 1.1936 0.38584 0.11514 0.014745 7.4192 0.091996 0.00011512 0.79812 0.0072777 0.0081211 0.0017223 0.9824 0.98284 3.7643e-006 1.5058e-005 0.14819 0.64348 0.73553 0.0015658 0.72128 0.43116 0.0021028 0.4215 1.3081 1.3037 16.0036 144.9554 0.00043217 -84.349 0.14394
4.248 0.98807 5.4977e-005 3.8183 0.01199 5.5623e-005 0.0011584 0.22818 0.00065927 0.22884 0.21102 0 0.032536 0.0389 0 1.1937 0.38589 0.11515 0.014747 7.4209 0.092006 0.00011514 0.79811 0.0072784 0.0081218 0.0017195 0.98244 0.9832 3.7577e-006 1.5032e-005 0.1482 0.64453 0.73652 0.0015644 0.72284 0.43135 0.0021011 0.4215 1.3102 1.3058 16.0037 144.9554 0.00043087 -84.3589 0.14494
4.249 0.98807 5.4977e-005 3.8183 0.01199 5.5636e-005 0.0011584 0.22819 0.00065927 0.22884 0.21102 0 0.032536 0.0389 0 1.1938 0.38594 0.11517 0.014748 7.4225 0.092016 0.00011515 0.7981 0.0072791 0.0081226 0.0017167 0.98248 0.98355 3.7512e-006 1.5006e-005 0.14821 0.64558 0.7375 0.0015631 0.7244 0.43154 0.0020993 0.4215 1.3122 1.3078 16.0038 144.9554 0.00042958 -84.3687 0.14594
4.25 0.98807 5.4976e-005 3.8183 0.01199 5.5649e-005 0.0011584 0.22819 0.00065927 0.22885 0.21103 0 0.032535 0.0389 0 1.1939 0.38598 0.11518 0.01475 7.4241 0.092026 0.00011516 0.79809 0.0072798 0.0081233 0.0017139 0.98252 0.98388 3.7448e-006 1.498e-005 0.14821 0.64663 0.73848 0.0015618 0.72596 0.43173 0.0020976 0.4215 1.3143 1.3099 16.0038 144.9555 0.0004283 -84.3784 0.14694
4.251 0.98807 5.4976e-005 3.8183 0.01199 5.5662e-005 0.0011584 0.2282 0.00065927 0.22885 0.21103 0 0.032535 0.0389 0 1.194 0.38603 0.1152 0.014751 7.4258 0.092036 0.00011518 0.79808 0.0072804 0.008124 0.0017111 0.98255 0.98419 3.7384e-006 1.4954e-005 0.14822 0.64768 0.73945 0.0015605 0.7275 0.43192 0.0020958 0.4215 1.3164 1.312 16.0039 144.9555 0.00042702 -84.388 0.14794
4.252 0.98807 5.4976e-005 3.8183 0.01199 5.5675e-005 0.0011584 0.2282 0.00065927 0.22886 0.21104 0 0.032535 0.0389 0 1.1941 0.38608 0.11522 0.014753 7.4274 0.092046 0.00011519 0.79807 0.0072811 0.0081248 0.0017084 0.98259 0.98449 3.7321e-006 1.4929e-005 0.14822 0.64872 0.74042 0.0015592 0.72904 0.43211 0.0020941 0.4215 1.3184 1.3141 16.004 144.9555 0.00042575 -84.3976 0.14894
4.253 0.98807 5.4976e-005 3.8183 0.01199 5.5688e-005 0.0011584 0.22821 0.00065927 0.22886 0.21104 0 0.032534 0.0389 0 1.1942 0.38612 0.11523 0.014755 7.429 0.092056 0.00011521 0.79806 0.0072818 0.0081255 0.0017057 0.98263 0.98477 3.7259e-006 1.4904e-005 0.14823 0.64976 0.74137 0.0015579 0.73057 0.4323 0.0020925 0.42151 1.3205 1.3161 16.004 144.9555 0.00042449 -84.407 0.14994
4.254 0.98807 5.4976e-005 3.8183 0.01199 5.5701e-005 0.0011584 0.22821 0.00065927 0.22887 0.21105 0 0.032534 0.0389 0 1.1943 0.38617 0.11525 0.014756 7.4307 0.092066 0.00011522 0.79805 0.0072825 0.0081262 0.0017031 0.98267 0.98503 3.7197e-006 1.4879e-005 0.14823 0.65079 0.74232 0.0015566 0.7321 0.43249 0.0020908 0.42151 1.3225 1.3182 16.0041 144.9555 0.00042323 -84.4164 0.15094
4.255 0.98807 5.4976e-005 3.8183 0.01199 5.5714e-005 0.0011584 0.22822 0.00065927 0.22887 0.21105 0 0.032534 0.0389 0 1.1944 0.38622 0.11526 0.014758 7.4323 0.092076 0.00011523 0.79804 0.0072832 0.008127 0.0017004 0.98271 0.98528 3.7135e-006 1.4855e-005 0.14824 0.65183 0.74327 0.0015553 0.73361 0.43268 0.0020891 0.42151 1.3246 1.3203 16.0042 144.9555 0.00042198 -84.4258 0.15194
4.256 0.98807 5.4976e-005 3.8183 0.01199 5.5727e-005 0.0011584 0.22823 0.00065927 0.22888 0.21106 0 0.032534 0.0389 0 1.1945 0.38626 0.11528 0.01476 7.434 0.092086 0.00011525 0.79803 0.0072839 0.0081277 0.0016978 0.98274 0.98551 3.7075e-006 1.4831e-005 0.14824 0.65285 0.7442 0.0015541 0.73512 0.43287 0.0020875 0.42151 1.3266 1.3223 16.0042 144.9555 0.00042074 -84.435 0.15294
4.257 0.98807 5.4976e-005 3.8183 0.01199 5.574e-005 0.0011585 0.22823 0.00065927 0.22889 0.21106 0 0.032533 0.0389 0 1.1946 0.38631 0.1153 0.014761 7.4356 0.092096 0.00011526 0.79802 0.0072845 0.0081284 0.0016952 0.98278 0.98574 3.7015e-006 1.4807e-005 0.14825 0.65388 0.74513 0.0015528 0.73663 0.43306 0.0020858 0.42151 1.3286 1.3244 16.0043 144.9555 0.0004195 -84.4442 0.15394
4.258 0.98807 5.4976e-005 3.8183 0.01199 5.5753e-005 0.0011585 0.22824 0.00065927 0.22889 0.21107 0 0.032533 0.0389 0 1.1947 0.38636 0.11531 0.014763 7.4372 0.092106 0.00011528 0.79801 0.0072852 0.0081292 0.0016927 0.98281 0.98595 3.6955e-006 1.4783e-005 0.14825 0.6549 0.74606 0.0015516 0.73812 0.43325 0.0020842 0.42152 1.3307 1.3264 16.0043 144.9555 0.00041827 -84.4533 0.15494
4.259 0.98807 5.4976e-005 3.8183 0.01199 5.5766e-005 0.0011585 0.22824 0.00065927 0.2289 0.21107 0 0.032533 0.0389 0 1.1948 0.3864 0.11533 0.014764 7.4389 0.092116 0.00011529 0.798 0.0072859 0.0081299 0.0016901 0.98285 0.98615 3.6896e-006 1.4759e-005 0.14826 0.65592 0.74697 0.0015503 0.73961 0.43344 0.0020826 0.42152 1.3327 1.3285 16.0044 144.9556 0.00041704 -84.4623 0.15594
4.26 0.98807 5.4976e-005 3.8183 0.01199 5.5779e-005 0.0011585 0.22825 0.00065927 0.2289 0.21108 0 0.032533 0.0389 0 1.1949 0.38645 0.11534 0.014766 7.4405 0.092127 0.0001153 0.79799 0.0072866 0.0081306 0.0016876 0.98289 0.98634 3.6838e-006 1.4736e-005 0.14827 0.65694 0.74789 0.0015491 0.74109 0.43363 0.002081 0.42152 1.3347 1.3305 16.0045 144.9556 0.00041583 -84.4713 0.15694
4.261 0.98807 5.4976e-005 3.8183 0.01199 5.5792e-005 0.0011585 0.22825 0.00065927 0.22891 0.21108 0 0.032532 0.0389 0 1.195 0.3865 0.11536 0.014768 7.4422 0.092137 0.00011532 0.79798 0.0072873 0.0081314 0.0016851 0.98292 0.98652 3.678e-006 1.4713e-005 0.14827 0.65795 0.74879 0.0015479 0.74256 0.43382 0.0020795 0.42152 1.3367 1.3325 16.0045 144.9556 0.00041462 -84.4801 0.15794
4.262 0.98807 5.4976e-005 3.8183 0.01199 5.5805e-005 0.0011585 0.22826 0.00065927 0.22891 0.21109 0 0.032532 0.0389 0 1.1951 0.38654 0.11537 0.014769 7.4438 0.092147 0.00011533 0.79797 0.0072879 0.0081321 0.0016827 0.98296 0.98669 3.6722e-006 1.469e-005 0.14828 0.65896 0.74969 0.0015467 0.74403 0.43401 0.0020779 0.42153 1.3387 1.3346 16.0046 144.9556 0.00041341 -84.489 0.15894
4.263 0.98807 5.4975e-005 3.8183 0.01199 5.5818e-005 0.0011585 0.22826 0.00065927 0.22892 0.21109 0 0.032532 0.0389 0 1.1952 0.38659 0.11539 0.014771 7.4454 0.092157 0.00011535 0.79796 0.0072886 0.0081328 0.0016802 0.98299 0.98685 3.6666e-006 1.4667e-005 0.14828 0.65997 0.75058 0.0015455 0.74549 0.4342 0.0020764 0.42153 1.3408 1.3366 16.0046 144.9556 0.00041221 -84.4977 0.15994
4.264 0.98807 5.4975e-005 3.8183 0.01199 5.5831e-005 0.0011585 0.22827 0.00065927 0.22892 0.2111 0 0.032532 0.0389 0 1.1953 0.38664 0.11541 0.014773 7.4471 0.092167 0.00011536 0.79795 0.0072893 0.0081336 0.0016778 0.98302 0.98701 3.6609e-006 1.4644e-005 0.14829 0.66097 0.75147 0.0015444 0.74694 0.43439 0.0020748 0.42153 1.3428 1.3386 16.0047 144.9556 0.00041102 -84.5064 0.16094
4.265 0.98807 5.4975e-005 3.8183 0.01199 5.5844e-005 0.0011585 0.22827 0.00065927 0.22893 0.2111 0 0.032531 0.0389 0 1.1954 0.38668 0.11542 0.014774 7.4487 0.092177 0.00011537 0.79794 0.00729 0.0081343 0.0016754 0.98306 0.98715 3.6554e-006 1.4622e-005 0.14829 0.66197 0.75235 0.0015432 0.74839 0.43458 0.0020733 0.42154 1.3448 1.3406 16.0048 144.9556 0.00040983 -84.515 0.16194
4.266 0.98807 5.4975e-005 3.8183 0.01199 5.5857e-005 0.0011585 0.22828 0.00065927 0.22893 0.21111 0 0.032531 0.0389 0 1.1955 0.38673 0.11544 0.014776 7.4504 0.092187 0.00011539 0.79793 0.0072907 0.008135 0.001673 0.98309 0.98729 3.6498e-006 1.46e-005 0.1483 0.66297 0.75322 0.0015421 0.74982 0.43477 0.0020718 0.42154 1.3468 1.3426 16.0048 144.9556 0.00040865 -84.5235 0.16294
4.267 0.98807 5.4975e-005 3.8183 0.01199 5.587e-005 0.0011585 0.22828 0.00065927 0.22894 0.21111 0 0.032531 0.0389 0 1.1956 0.38678 0.11545 0.014777 7.452 0.092197 0.0001154 0.79792 0.0072914 0.0081358 0.0016707 0.98312 0.98742 3.6444e-006 1.4578e-005 0.1483 0.66397 0.75409 0.0015409 0.75126 0.43496 0.0020703 0.42154 1.3488 1.3446 16.0049 144.9557 0.00040748 -84.532 0.16394
4.268 0.98807 5.4975e-005 3.8183 0.01199 5.5883e-005 0.0011585 0.22829 0.00065927 0.22894 0.21112 0 0.03253 0.0389 0 1.1957 0.38682 0.11547 0.014779 7.4536 0.092207 0.00011542 0.79791 0.007292 0.0081365 0.0016683 0.98316 0.98755 3.639e-006 1.4556e-005 0.14831 0.66496 0.75495 0.0015398 0.75268 0.43515 0.0020688 0.42155 1.3507 1.3466 16.0049 144.9557 0.00040631 -84.5404 0.16494
4.269 0.98807 5.4975e-005 3.8183 0.01199 5.5896e-005 0.0011585 0.22829 0.00065927 0.22895 0.21112 0 0.03253 0.0389 0 1.1958 0.38687 0.11549 0.014781 7.4553 0.092217 0.00011543 0.7979 0.0072927 0.0081372 0.001666 0.98319 0.98766 3.6336e-006 1.4535e-005 0.14831 0.66595 0.75581 0.0015387 0.7541 0.43534 0.0020674 0.42155 1.3527 1.3486 16.005 144.9557 0.00040515 -84.5487 0.16594
4.27 0.98807 5.4975e-005 3.8183 0.01199 5.5909e-005 0.0011585 0.2283 0.00065927 0.22895 0.21113 0 0.03253 0.0389 0 1.1959 0.38692 0.1155 0.014782 7.4569 0.092227 0.00011544 0.79789 0.0072934 0.008138 0.0016637 0.98322 0.98778 3.6283e-006 1.4514e-005 0.14832 0.66693 0.75666 0.0015375 0.75551 0.43552 0.0020659 0.42155 1.3547 1.3506 16.0051 144.9557 0.00040399 -84.557 0.16694
4.271 0.98807 5.4975e-005 3.8183 0.01199 5.5922e-005 0.0011585 0.2283 0.00065927 0.22896 0.21113 0 0.03253 0.0389 0 1.196 0.38696 0.11552 0.014784 7.4586 0.092237 0.00011546 0.79788 0.0072941 0.0081387 0.0016614 0.98325 0.98788 3.623e-006 1.4493e-005 0.14833 0.66792 0.7575 0.0015364 0.75691 0.43571 0.0020645 0.42156 1.3567 1.3526 16.0051 144.9557 0.00040284 -84.5652 0.16794
4.272 0.98807 5.4975e-005 3.8183 0.01199 5.5935e-005 0.0011585 0.22831 0.00065927 0.22896 0.21114 0 0.032529 0.0389 0 1.1961 0.38701 0.11553 0.014785 7.4602 0.092247 0.00011547 0.79787 0.0072948 0.0081394 0.0016592 0.98328 0.98798 3.6178e-006 1.4472e-005 0.14833 0.6689 0.75834 0.0015354 0.75831 0.4359 0.002063 0.42156 1.3587 1.3546 16.0052 144.9557 0.0004017 -84.5734 0.16894
4.273 0.98807 5.4975e-005 3.8183 0.01199 5.5948e-005 0.0011585 0.22832 0.00065927 0.22897 0.21114 0 0.032529 0.0389 0 1.1962 0.38706 0.11555 0.014787 7.4619 0.092257 0.00011549 0.79786 0.0072954 0.0081402 0.001657 0.98331 0.98808 3.6126e-006 1.4451e-005 0.14834 0.66987 0.75917 0.0015343 0.75969 0.43609 0.0020616 0.42156 1.3606 1.3566 16.0052 144.9557 0.00040056 -84.5814 0.16994
4.274 0.98807 5.4975e-005 3.8183 0.01199 5.5961e-005 0.0011585 0.22832 0.00065927 0.22898 0.21115 0 0.032529 0.0389 0 1.1963 0.3871 0.11557 0.014789 7.4635 0.092267 0.0001155 0.79785 0.0072961 0.0081409 0.0016548 0.98335 0.98817 3.6075e-006 1.4431e-005 0.14834 0.67085 0.76 0.0015332 0.76108 0.43628 0.0020602 0.42157 1.3626 1.3586 16.0053 144.9557 0.00039943 -84.5895 0.17094
4.275 0.98807 5.4975e-005 3.8183 0.01199 5.5974e-005 0.0011585 0.22833 0.00065927 0.22898 0.21115 0 0.032529 0.0389 0 1.1964 0.38715 0.11558 0.01479 7.4652 0.092277 0.00011551 0.79784 0.0072968 0.0081416 0.0016526 0.98338 0.98826 3.6024e-006 1.441e-005 0.14835 0.67182 0.76082 0.0015321 0.76245 0.43647 0.0020588 0.42157 1.3645 1.3605 16.0053 144.9557 0.0003983 -84.5974 0.17194
4.276 0.98807 5.4975e-005 3.8183 0.01199 5.5987e-005 0.0011585 0.22833 0.00065927 0.22899 0.21116 0 0.032528 0.0389 0 1.1965 0.3872 0.1156 0.014792 7.4668 0.092287 0.00011553 0.79783 0.0072975 0.0081424 0.0016504 0.98341 0.98834 3.5974e-006 1.439e-005 0.14835 0.67278 0.76164 0.0015311 0.76382 0.43666 0.0020574 0.42158 1.3665 1.3625 16.0054 144.9558 0.00039718 -84.6053 0.17294
4.277 0.98807 5.4974e-005 3.8183 0.011989 5.6e-005 0.0011585 0.22834 0.00065927 0.22899 0.21116 0 0.032528 0.0389 0 1.1966 0.38724 0.11561 0.014794 7.4684 0.092297 0.00011554 0.79782 0.0072982 0.0081431 0.0016483 0.98344 0.98842 3.5924e-006 1.437e-005 0.14836 0.67375 0.76245 0.00153 0.76518 0.43685 0.0020561 0.42158 1.3684 1.3645 16.0055 144.9558 0.00039606 -84.6131 0.17394
4.278 0.98807 5.4974e-005 3.8183 0.011989 5.6013e-005 0.0011585 0.22834 0.00065927 0.229 0.21117 0 0.032528 0.0389 0 1.1967 0.38729 0.11563 0.014795 7.4701 0.092307 0.00011556 0.79781 0.0072989 0.0081438 0.0016461 0.98347 0.9885 3.5875e-006 1.435e-005 0.14836 0.67471 0.76326 0.001529 0.76654 0.43704 0.0020547 0.42158 1.3704 1.3664 16.0055 144.9558 0.00039495 -84.6209 0.17494
4.279 0.98807 5.4974e-005 3.8183 0.011989 5.6026e-005 0.0011585 0.22835 0.00065927 0.229 0.21117 0 0.032528 0.0389 0 1.1968 0.38734 0.11565 0.014797 7.4717 0.092317 0.00011557 0.7978 0.0072995 0.0081446 0.001644 0.98349 0.98857 3.5826e-006 1.4331e-005 0.14837 0.67567 0.76406 0.0015279 0.76788 0.43723 0.0020533 0.42159 1.3723 1.3684 16.0056 144.9558 0.00039385 -84.6286 0.17594
4.28 0.98807 5.4974e-005 3.8183 0.011989 5.6039e-005 0.0011585 0.22835 0.00065927 0.22901 0.21118 0 0.032527 0.0389 0 1.1969 0.38738 0.11566 0.014798 7.4734 0.092327 0.00011558 0.79779 0.0073002 0.0081453 0.0016419 0.98352 0.98864 3.5778e-006 1.4312e-005 0.14837 0.67663 0.76486 0.0015269 0.76922 0.43742 0.002052 0.42159 1.3743 1.3703 16.0056 144.9558 0.00039275 -84.6363 0.17694
4.281 0.98807 5.4974e-005 3.8183 0.011989 5.6052e-005 0.0011585 0.22836 0.00065927 0.22901 0.21118 0 0.032527 0.0389 0 1.197 0.38743 0.11568 0.0148 7.475 0.092337 0.0001156 0.79778 0.0073009 0.008146 0.0016398 0.98355 0.98871 3.573e-006 1.4292e-005 0.14838 0.67758 0.76565 0.0015259 0.77056 0.43761 0.0020507 0.4216 1.3762 1.3723 16.0057 144.9558 0.00039166 -84.6438 0.17794
4.282 0.98807 5.4974e-005 3.8183 0.011989 5.6065e-005 0.0011585 0.22836 0.00065927 0.22902 0.21119 0 0.032527 0.0389 0 1.1971 0.38748 0.11569 0.014802 7.4767 0.092347 0.00011561 0.79777 0.0073016 0.0081468 0.0016378 0.98358 0.98877 3.5682e-006 1.4273e-005 0.14838 0.67853 0.76643 0.0015249 0.77189 0.4378 0.0020494 0.4216 1.3781 1.3742 16.0057 144.9558 0.00039057 -84.6514 0.17894
4.283 0.98807 5.4974e-005 3.8183 0.011989 5.6078e-005 0.0011585 0.22837 0.00065927 0.22902 0.21119 0 0.032526 0.0389 0 1.1972 0.38752 0.11571 0.014803 7.4783 0.092357 0.00011563 0.79776 0.0073023 0.0081475 0.0016358 0.98361 0.98883 3.5635e-006 1.4254e-005 0.14839 0.67948 0.76721 0.0015239 0.77321 0.43799 0.0020481 0.42161 1.3801 1.3762 16.0058 144.9558 0.00038949 -84.6588 0.17994
4.284 0.98807 5.4974e-005 3.8183 0.011989 5.6091e-005 0.0011585 0.22837 0.00065927 0.22903 0.2112 0 0.032526 0.0389 0 1.1973 0.38757 0.11573 0.014805 7.48 0.092367 0.00011564 0.79775 0.0073029 0.0081482 0.0016338 0.98364 0.98889 3.5588e-006 1.4236e-005 0.1484 0.68042 0.76799 0.0015229 0.77452 0.43818 0.0020468 0.42161 1.382 1.3781 16.0058 144.9559 0.00038842 -84.6663 0.18094
4.285 0.98807 5.4974e-005 3.8183 0.011989 5.6104e-005 0.0011585 0.22838 0.00065927 0.22903 0.2112 0 0.032526 0.0389 0 1.1974 0.38762 0.11574 0.014807 7.4816 0.092377 0.00011565 0.79774 0.0073036 0.008149 0.0016318 0.98366 0.98894 3.5542e-006 1.4217e-005 0.1484 0.68136 0.76876 0.0015219 0.77583 0.43837 0.0020455 0.42162 1.3839 1.38 16.0059 144.9559 0.00038735 -84.6736 0.18194
4.286 0.98807 5.4974e-005 3.8183 0.011989 5.6117e-005 0.0011585 0.22838 0.00065927 0.22904 0.21121 0 0.032526 0.0389 0 1.1975 0.38766 0.11576 0.014808 7.4833 0.092387 0.00011567 0.79773 0.0073043 0.0081497 0.0016298 0.98369 0.98899 3.5496e-006 1.4199e-005 0.14841 0.6823 0.76952 0.001521 0.77713 0.43856 0.0020442 0.42162 1.3858 1.3819 16.0059 144.9559 0.00038628 -84.6809 0.18294
4.287 0.98807 5.4974e-005 3.8183 0.011989 5.613e-005 0.0011585 0.22839 0.00065927 0.22904 0.21121 0 0.032525 0.0389 0 1.1976 0.38771 0.11577 0.01481 7.4849 0.092398 0.00011568 0.79772 0.007305 0.0081504 0.0016278 0.98372 0.98904 3.5451e-006 1.4181e-005 0.14841 0.68324 0.77028 0.00152 0.77842 0.43875 0.002043 0.42163 1.3877 1.3839 16.006 144.9559 0.00038522 -84.6881 0.18394
4.288 0.98807 5.4974e-005 3.8183 0.011989 5.6143e-005 0.0011585 0.22839 0.00065927 0.22905 0.21122 0 0.032525 0.0389 0 1.1977 0.38776 0.11579 0.014811 7.4866 0.092408 0.0001157 0.79771 0.0073057 0.0081512 0.0016259 0.98375 0.98909 3.5405e-006 1.4163e-005 0.14842 0.68417 0.77104 0.0015191 0.77971 0.43894 0.0020417 0.42163 1.3896 1.3858 16.006 144.9559 0.00038417 -84.6953 0.18494
4.289 0.98807 5.4974e-005 3.8183 0.011989 5.6156e-005 0.0011585 0.2284 0.00065927 0.22905 0.21122 0 0.032525 0.0389 0 1.1978 0.3878 0.11581 0.014813 7.4882 0.092418 0.00011571 0.7977 0.0073063 0.0081519 0.001624 0.98377 0.98914 3.5361e-006 1.4145e-005 0.14842 0.6851 0.77179 0.0015181 0.78099 0.43913 0.0020405 0.42164 1.3915 1.3877 16.0061 144.9559 0.00038312 -84.7025 0.18594
4.29 0.98807 5.4974e-005 3.8183 0.011989 5.6169e-005 0.0011585 0.2284 0.00065927 0.22906 0.21123 0 0.032525 0.0389 0 1.1979 0.38785 0.11582 0.014815 7.4899 0.092428 0.00011572 0.79769 0.007307 0.0081526 0.001622 0.9838 0.98918 3.5317e-006 1.4127e-005 0.14843 0.68603 0.77253 0.0015172 0.78226 0.43931 0.0020393 0.42164 1.3934 1.3896 16.0061 144.9559 0.00038207 -84.7095 0.18694
4.291 0.98807 5.4973e-005 3.8183 0.011989 5.6182e-005 0.0011585 0.22841 0.00065927 0.22906 0.21123 0 0.032524 0.0389 0 1.198 0.3879 0.11584 0.014816 7.4915 0.092438 0.00011574 0.79768 0.0073077 0.0081534 0.0016201 0.98383 0.98923 3.5273e-006 1.411e-005 0.14843 0.68695 0.77328 0.0015162 0.78353 0.4395 0.002038 0.42165 1.3953 1.3915 16.0062 144.956 0.00038104 -84.7165 0.18794
4.292 0.98807 5.4973e-005 3.8183 0.011989 5.6195e-005 0.0011585 0.22841 0.00065927 0.22907 0.21124 0 0.032524 0.0389 0 1.198 0.38794 0.11585 0.014818 7.4932 0.092448 0.00011575 0.79767 0.0073084 0.0081541 0.0016182 0.98385 0.98927 3.5229e-006 1.4092e-005 0.14844 0.68787 0.77401 0.0015153 0.78479 0.43969 0.0020368 0.42165 1.3972 1.3934 16.0062 144.956 0.00038 -84.7235 0.18894
4.293 0.98807 5.4973e-005 3.8183 0.011989 5.6208e-005 0.0011585 0.22842 0.00065927 0.22907 0.21124 0 0.032524 0.0389 0 1.1981 0.38799 0.11587 0.014819 7.4948 0.092458 0.00011577 0.79766 0.0073091 0.0081548 0.0016164 0.98388 0.98931 3.5186e-006 1.4075e-005 0.14844 0.68879 0.77474 0.0015144 0.78605 0.43988 0.0020356 0.42166 1.3991 1.3953 16.0063 144.956 0.00037898 -84.7304 0.18994
4.294 0.98807 5.4973e-005 3.8183 0.011989 5.6221e-005 0.0011585 0.22842 0.00065927 0.22908 0.21125 0 0.032524 0.0389 0 1.1982 0.38804 0.11588 0.014821 7.4965 0.092468 0.00011578 0.79765 0.0073097 0.0081555 0.0016145 0.9839 0.98935 3.5144e-006 1.4058e-005 0.14845 0.6897 0.77547 0.0015135 0.78729 0.44007 0.0020344 0.42166 1.4009 1.3972 16.0063 144.956 0.00037795 -84.7373 0.19094
4.295 0.98807 5.4973e-005 3.8183 0.011989 5.6234e-005 0.0011585 0.22843 0.00065927 0.22908 0.21125 0 0.032523 0.0389 0 1.1983 0.38808 0.1159 0.014823 7.4981 0.092478 0.00011579 0.79764 0.0073104 0.0081563 0.0016128 0.98393 0.98938 3.5101e-006 1.4041e-005 0.14846 0.69062 0.77619 0.0015126 0.78854 0.44026 0.0020333 0.42167 1.4028 1.3991 16.0064 144.956 0.00037694 -84.7441 0.19194
4.296 0.98807 5.4973e-005 3.8183 0.011989 5.6247e-005 0.0011585 0.22843 0.00065927 0.22909 0.21126 0 0.032523 0.0389 0 1.1984 0.38813 0.11592 0.014824 7.4998 0.092488 0.00011581 0.79763 0.0073111 0.008157 0.001611 0.98395 0.98942 3.5059e-006 1.4024e-005 0.14846 0.69153 0.77691 0.0015117 0.78977 0.44045 0.0020321 0.42167 1.4047 1.401 16.0064 144.956 0.00037592 -84.7508 0.19294
4.297 0.98807 5.4973e-005 3.8183 0.011989 5.626e-005 0.0011585 0.22844 0.00065927 0.22909 0.21126 0 0.032523 0.0389 0 1.1985 0.38818 0.11593 0.014826 7.5014 0.092498 0.00011582 0.79762 0.0073118 0.0081577 0.0016092 0.98398 0.98945 3.5018e-006 1.4008e-005 0.14847 0.69243 0.77762 0.0015108 0.791 0.44064 0.0020309 0.42168 1.4065 1.4028 16.0065 144.956 0.00037492 -84.7575 0.19394
4.298 0.98807 5.4973e-005 3.8183 0.011989 5.6273e-005 0.0011586 0.22845 0.00065927 0.2291 0.21127 0 0.032523 0.0389 0 1.1986 0.38822 0.11595 0.014828 7.5031 0.092508 0.00011584 0.79761 0.0073125 0.0081585 0.0016074 0.984 0.98949 3.4977e-006 1.3991e-005 0.14847 0.69334 0.77833 0.0015099 0.79222 0.44083 0.0020298 0.42169 1.4084 1.4047 16.0065 144.956 0.00037391 -84.7642 0.19494
4.299 0.98807 5.4973e-005 3.8183 0.011989 5.6286e-005 0.0011586 0.22845 0.00065927 0.2291 0.21127 0 0.032522 0.0389 0 1.1987 0.38827 0.11596 0.014829 7.5047 0.092518 0.00011585 0.7976 0.0073131 0.0081592 0.0016056 0.98403 0.98952 3.4936e-006 1.3975e-005 0.14848 0.69424 0.77904 0.0015091 0.79344 0.44102 0.0020286 0.42169 1.4103 1.4066 16.0066 144.9561 0.00037292 -84.7708 0.19594
4.3 0.98807 5.4973e-005 3.8183 0.011989 5.6299e-005 0.0011586 0.22846 0.00065927 0.22911 0.21128 0 0.032522 0.0389 0 1.1988 0.38831 0.11598 0.014831 7.5064 0.092528 0.00011586 0.79759 0.0073138 0.0081599 0.0016038 0.98405 0.98955 3.4895e-006 1.3959e-005 0.14848 0.69514 0.77974 0.0015082 0.79465 0.44121 0.0020275 0.4217 1.4121 1.4084 16.0066 144.9561 0.00037192 -84.7773 0.19694
4.301 0.98807 5.4973e-005 3.8183 0.011989 5.6312e-005 0.0011586 0.22846 0.00065927 0.22912 0.21128 0 0.032522 0.0389 0 1.1989 0.38836 0.116 0.014832 7.508 0.092538 0.00011588 0.79758 0.0073145 0.0081607 0.0016021 0.98407 0.98958 3.4855e-006 1.3943e-005 0.14849 0.69604 0.78043 0.0015073 0.79585 0.4414 0.0020264 0.4217 1.4139 1.4103 16.0067 144.9561 0.00037094 -84.7838 0.19794
4.302 0.98807 5.4973e-005 3.8183 0.011989 5.6325e-005 0.0011586 0.22847 0.00065927 0.22912 0.21129 0 0.032522 0.0389 0 1.199 0.38841 0.11601 0.014834 7.5097 0.092548 0.00011589 0.79757 0.0073152 0.0081614 0.0016004 0.9841 0.98961 3.4816e-006 1.3927e-005 0.14849 0.69693 0.78113 0.0015065 0.79705 0.44159 0.0020253 0.42171 1.4158 1.4121 16.0067 144.9561 0.00036995 -84.7903 0.19894
4.303 0.98807 5.4973e-005 3.8183 0.011989 5.6338e-005 0.0011586 0.22847 0.00065927 0.22913 0.21129 0 0.032521 0.0389 0 1.1991 0.38845 0.11603 0.014836 7.5114 0.092558 0.00011591 0.79756 0.0073158 0.0081621 0.0015987 0.98412 0.98963 3.4776e-006 1.3911e-005 0.1485 0.69782 0.78181 0.0015056 0.79824 0.44177 0.0020242 0.42172 1.4176 1.414 16.0068 144.9561 0.00036898 -84.7967 0.19994
4.304 0.98807 5.4973e-005 3.8183 0.011989 5.6351e-005 0.0011586 0.22848 0.00065927 0.22913 0.2113 0 0.032521 0.0389 0 1.1992 0.3885 0.11604 0.014837 7.513 0.092568 0.00011592 0.79755 0.0073165 0.0081629 0.001597 0.98414 0.98966 3.4737e-006 1.3895e-005 0.1485 0.69871 0.7825 0.0015048 0.79942 0.44196 0.0020231 0.42172 1.4195 1.4158 16.0068 144.9561 0.000368 -84.803 0.20094
4.305 0.98807 5.4972e-005 3.8183 0.011989 5.6364e-005 0.0011586 0.22848 0.00065927 0.22914 0.2113 0 0.032521 0.0389 0 1.1993 0.38855 0.11606 0.014839 7.5147 0.092578 0.00011593 0.79754 0.0073172 0.0081636 0.0015953 0.98417 0.98969 3.4698e-006 1.388e-005 0.14851 0.69959 0.78318 0.001504 0.8006 0.44215 0.002022 0.42173 1.4213 1.4177 16.0068 144.9561 0.00036704 -84.8093 0.20194
4.306 0.98807 5.4972e-005 3.8183 0.011989 5.6377e-005 0.0011586 0.22849 0.00065927 0.22914 0.21131 0 0.032521 0.0389 0 1.1994 0.38859 0.11608 0.01484 7.5163 0.092588 0.00011595 0.79753 0.0073179 0.0081643 0.0015937 0.98419 0.98971 3.466e-006 1.3864e-005 0.14852 0.70047 0.78385 0.0015032 0.80177 0.44234 0.0020209 0.42173 1.4231 1.4195 16.0069 144.9562 0.00036607 -84.8156 0.20294
4.307 0.98807 5.4972e-005 3.8183 0.011989 5.639e-005 0.0011586 0.22849 0.00065927 0.22915 0.21131 0 0.03252 0.0389 0 1.1995 0.38864 0.11609 0.014842 7.518 0.092598 0.00011596 0.79752 0.0073186 0.0081651 0.001592 0.98421 0.98974 3.4622e-006 1.3849e-005 0.14852 0.70135 0.78452 0.0015023 0.80293 0.44253 0.0020199 0.42174 1.4249 1.4214 16.0069 144.9562 0.00036512 -84.8218 0.20394
4.308 0.98807 5.4972e-005 3.8183 0.011989 5.6403e-005 0.0011586 0.2285 0.00065927 0.22915 0.21132 0 0.03252 0.0389 0 1.1996 0.38869 0.11611 0.014844 7.5196 0.092608 0.00011598 0.79751 0.0073192 0.0081658 0.0015904 0.98423 0.98976 3.4584e-006 1.3834e-005 0.14853 0.70223 0.78519 0.0015015 0.80409 0.44272 0.0020188 0.42175 1.4268 1.4232 16.007 144.9562 0.00036416 -84.8279 0.20494
4.309 0.98807 5.4972e-005 3.8183 0.011989 5.6416e-005 0.0011586 0.2285 0.00065927 0.22916 0.21132 0 0.03252 0.0389 0 1.1997 0.38873 0.11612 0.014845 7.5213 0.092618 0.00011599 0.7975 0.0073199 0.0081665 0.0015888 0.98426 0.98978 3.4547e-006 1.3819e-005 0.14853 0.70311 0.78585 0.0015007 0.80524 0.44291 0.0020178 0.42175 1.4286 1.425 16.007 144.9562 0.00036321 -84.834 0.20594
4.31 0.98807 5.4972e-005 3.8183 0.011989 5.6429e-005 0.0011586 0.22851 0.00065927 0.22916 0.21133 0 0.032519 0.0389 0 1.1998 0.38878 0.11614 0.014847 7.523 0.092628 0.000116 0.79749 0.0073206 0.0081672 0.0015872 0.98428 0.98981 3.451e-006 1.3804e-005 0.14854 0.70398 0.78651 0.0014999 0.80639 0.4431 0.0020167 0.42176 1.4304 1.4268 16.0071 144.9562 0.00036227 -84.8401 0.20694
4.311 0.98807 5.4972e-005 3.8183 0.011989 5.6442e-005 0.0011586 0.22851 0.00065927 0.22917 0.21133 0 0.032519 0.0389 0 1.1999 0.38883 0.11616 0.014849 7.5246 0.092638 0.00011602 0.79748 0.0073213 0.008168 0.0015856 0.9843 0.98983 3.4473e-006 1.379e-005 0.14854 0.70485 0.78716 0.0014991 0.80753 0.44329 0.0020157 0.42177 1.4322 1.4286 16.0071 144.9562 0.00036133 -84.8461 0.20794
4.312 0.98807 5.4972e-005 3.8183 0.011989 5.6455e-005 0.0011586 0.22852 0.00065927 0.22917 0.21134 0 0.032519 0.0389 0 1.2 0.38887 0.11617 0.01485 7.5263 0.092648 0.00011603 0.79747 0.007322 0.0081687 0.001584 0.98432 0.98985 3.4437e-006 1.3775e-005 0.14855 0.70571 0.78782 0.0014984 0.80867 0.44347 0.0020147 0.42177 1.434 1.4305 16.0072 144.9562 0.0003604 -84.8521 0.20894
4.313 0.98807 5.4972e-005 3.8183 0.011989 5.6468e-005 0.0011586 0.22852 0.00065927 0.22918 0.21134 0 0.032519 0.0389 0 1.2001 0.38892 0.11619 0.014852 7.5279 0.092658 0.00011605 0.79746 0.0073226 0.0081694 0.0015824 0.98434 0.98987 3.4401e-006 1.3761e-005 0.14855 0.70658 0.78846 0.0014976 0.80979 0.44366 0.0020137 0.42178 1.4358 1.4323 16.0072 144.9563 0.00035947 -84.858 0.20994
4.314 0.98807 5.4972e-005 3.8183 0.011989 5.6481e-005 0.0011586 0.22853 0.00065927 0.22918 0.21135 0 0.032518 0.0389 0 1.2002 0.38897 0.1162 0.014853 7.5296 0.092668 0.00011606 0.79745 0.0073233 0.0081702 0.0015809 0.98436 0.98989 3.4365e-006 1.3746e-005 0.14856 0.70744 0.78911 0.0014968 0.81092 0.44385 0.0020126 0.42179 1.4376 1.4341 16.0072 144.9563 0.00035854 -84.8639 0.21094
4.315 0.98807 5.4972e-005 3.8183 0.011989 5.6494e-005 0.0011586 0.22853 0.00065927 0.22919 0.21135 0 0.032518 0.0389 0 1.2003 0.38901 0.11622 0.014855 7.5312 0.092678 0.00011607 0.79744 0.007324 0.0081709 0.0015794 0.98438 0.98991 3.433e-006 1.3732e-005 0.14856 0.70829 0.78974 0.0014961 0.81203 0.44404 0.0020116 0.42179 1.4393 1.4359 16.0073 144.9563 0.00035762 -84.8697 0.21194
4.316 0.98807 5.4972e-005 3.8183 0.011989 5.6507e-005 0.0011586 0.22854 0.00065927 0.22919 0.21135 0 0.032518 0.0389 0 1.2004 0.38906 0.11624 0.014857 7.5329 0.092688 0.00011609 0.79743 0.0073247 0.0081716 0.0015779 0.98441 0.98993 3.4294e-006 1.3718e-005 0.14857 0.70915 0.79038 0.0014953 0.81314 0.44423 0.0020107 0.4218 1.4411 1.4377 16.0073 144.9563 0.00035671 -84.8755 0.21294
4.317 0.98807 5.4972e-005 3.8183 0.011989 5.652e-005 0.0011586 0.22854 0.00065927 0.2292 0.21136 0 0.032518 0.0389 0 1.2005 0.38911 0.11625 0.014858 7.5346 0.092698 0.0001161 0.79742 0.0073253 0.0081724 0.0015764 0.98443 0.98995 3.426e-006 1.3704e-005 0.14857 0.71 0.79101 0.0014945 0.81425 0.44442 0.0020097 0.42181 1.4429 1.4394 16.0074 144.9563 0.00035579 -84.8812 0.21394
4.318 0.98807 5.4972e-005 3.8183 0.011989 5.6533e-005 0.0011586 0.22855 0.00065927 0.2292 0.21136 0 0.032517 0.0389 0 1.2006 0.38915 0.11627 0.01486 7.5362 0.092708 0.00011612 0.79741 0.007326 0.0081731 0.0015749 0.98445 0.98997 3.4225e-006 1.369e-005 0.14858 0.71085 0.79164 0.0014938 0.81535 0.44461 0.0020087 0.42182 1.4447 1.4412 16.0074 144.9563 0.00035489 -84.8869 0.21494
4.319 0.98807 5.4971e-005 3.8183 0.011989 5.6546e-005 0.0011586 0.22855 0.00065927 0.22921 0.21137 0 0.032517 0.0389 0 1.2007 0.3892 0.11628 0.014861 7.5379 0.092718 0.00011613 0.7974 0.0073267 0.0081738 0.0015734 0.98447 0.98999 3.4191e-006 1.3677e-005 0.14859 0.7117 0.79226 0.0014931 0.81644 0.4448 0.0020077 0.42182 1.4464 1.443 16.0074 144.9563 0.00035398 -84.8926 0.21594
4.32 0.98807 5.4971e-005 3.8183 0.011989 5.6559e-005 0.0011586 0.22856 0.00065927 0.22921 0.21137 0 0.032517 0.0389 0 1.2008 0.38925 0.1163 0.014863 7.5395 0.092728 0.00011614 0.79739 0.0073274 0.0081745 0.0015719 0.98449 0.99 3.4157e-006 1.3663e-005 0.14859 0.71255 0.79288 0.0014923 0.81752 0.44498 0.0020068 0.42183 1.4482 1.4448 16.0075 144.9564 0.00035309 -84.8982 0.21694
4.321 0.98807 5.4971e-005 3.8183 0.011989 5.6572e-005 0.0011586 0.22856 0.00065927 0.22922 0.21138 0 0.032517 0.0389 0 1.2009 0.38929 0.11631 0.014865 7.5412 0.092738 0.00011616 0.79738 0.0073281 0.0081753 0.0015704 0.98451 0.99002 3.4123e-006 1.365e-005 0.1486 0.71339 0.7935 0.0014916 0.8186 0.44517 0.0020058 0.42184 1.45 1.4466 16.0075 144.9564 0.00035219 -84.9038 0.21794
4.322 0.98807 5.4971e-005 3.8183 0.011989 5.6585e-005 0.0011586 0.22857 0.00065927 0.22922 0.21138 0 0.032516 0.0389 0 1.201 0.38934 0.11633 0.014866 7.5429 0.092748 0.00011617 0.79737 0.0073287 0.008176 0.0015689 0.98453 0.99004 3.409e-006 1.3636e-005 0.1486 0.71423 0.79411 0.0014909 0.81968 0.44536 0.0020049 0.42185 1.4517 1.4483 16.0076 144.9564 0.0003513 -84.9093 0.21894
4.323 0.98807 5.4971e-005 3.8183 0.011989 5.6598e-005 0.0011586 0.22857 0.00065927 0.22923 0.21139 0 0.032516 0.0389 0 1.2011 0.38939 0.11635 0.014868 7.5445 0.092758 0.00011619 0.79736 0.0073294 0.0081767 0.0015675 0.98455 0.99006 3.4057e-006 1.3623e-005 0.14861 0.71507 0.79472 0.0014902 0.82075 0.44555 0.0020039 0.42185 1.4535 1.4501 16.0076 144.9564 0.00035042 -84.9148 0.21994
4.324 0.98807 5.4971e-005 3.8183 0.011989 5.6611e-005 0.0011586 0.22858 0.00065927 0.22923 0.21139 0 0.032516 0.0389 0 1.2012 0.38943 0.11636 0.01487 7.5462 0.092768 0.0001162 0.79735 0.0073301 0.0081775 0.0015661 0.98456 0.99007 3.4024e-006 1.361e-005 0.14861 0.7159 0.79533 0.0014895 0.82181 0.44574 0.002003 0.42186 1.4552 1.4518 16.0076 144.9564 0.00034954 -84.9202 0.22094
4.325 0.98807 5.4971e-005 3.8183 0.011989 5.6624e-005 0.0011586 0.22858 0.00065927 0.22924 0.2114 0 0.032516 0.0389 0 1.2013 0.38948 0.11638 0.014871 7.5479 0.092778 0.00011621 0.79734 0.0073308 0.0081782 0.0015647 0.98458 0.99009 3.3991e-006 1.3597e-005 0.14862 0.71673 0.79593 0.0014887 0.82287 0.44593 0.0020021 0.42187 1.457 1.4536 16.0077 144.9564 0.00034866 -84.9256 0.22194
4.326 0.98807 5.4971e-005 3.8183 0.011989 5.6637e-005 0.0011586 0.22859 0.00065927 0.22924 0.2114 0 0.032515 0.0389 0 1.2014 0.38953 0.11639 0.014873 7.5495 0.092788 0.00011623 0.79733 0.0073314 0.0081789 0.0015634 0.9846 0.9901 3.3959e-006 1.3584e-005 0.14862 0.71756 0.79653 0.0014881 0.82392 0.44612 0.0020012 0.42188 1.4587 1.4554 16.0077 144.9564 0.00034779 -84.931 0.22294
4.327 0.98807 5.4971e-005 3.8183 0.011989 5.665e-005 0.0011586 0.22859 0.00065927 0.22925 0.21141 0 0.032515 0.0389 0 1.2015 0.38957 0.11641 0.014874 7.5512 0.092798 0.00011624 0.79732 0.0073321 0.0081796 0.001562 0.98462 0.99012 3.3927e-006 1.3571e-005 0.14863 0.71839 0.79713 0.0014874 0.82496 0.4463 0.0020003 0.42188 1.4604 1.4571 16.0077 144.9565 0.00034692 -84.9363 0.22394
4.328 0.98807 5.4971e-005 3.8183 0.011989 5.6663e-005 0.0011586 0.2286 0.00065927 0.22925 0.21141 0 0.032515 0.0389 0 1.2016 0.38962 0.11643 0.014876 7.5529 0.092808 0.00011626 0.79731 0.0073328 0.0081804 0.0015606 0.98464 0.99013 3.3896e-006 1.3559e-005 0.14863 0.71921 0.79772 0.0014867 0.826 0.44649 0.0019994 0.42189 1.4622 1.4588 16.0078 144.9565 0.00034606 -84.9416 0.22494
4.329 0.98807 5.4971e-005 3.8183 0.011989 5.6676e-005 0.0011586 0.2286 0.00065927 0.22926 0.21142 0 0.032515 0.0389 0 1.2017 0.38967 0.11644 0.014878 7.5545 0.092818 0.00011627 0.7973 0.0073335 0.0081811 0.0015592 0.98466 0.99015 3.3864e-006 1.3546e-005 0.14864 0.72004 0.79831 0.001486 0.82704 0.44668 0.0019985 0.4219 1.4639 1.4606 16.0078 144.9565 0.0003452 -84.9468 0.22594
4.33 0.98807 5.4971e-005 3.8183 0.011989 5.6689e-005 0.0011586 0.22861 0.00065927 0.22926 0.21142 0 0.032514 0.0389 0 1.2018 0.38971 0.11646 0.014879 7.5562 0.092828 0.00011628 0.79729 0.0073342 0.0081818 0.0015579 0.98468 0.99016 3.3833e-006 1.3533e-005 0.14865 0.72086 0.7989 0.0014853 0.82807 0.44687 0.0019976 0.42191 1.4656 1.4623 16.0079 144.9565 0.00034434 -84.952 0.22694
4.331 0.98807 5.4971e-005 3.8183 0.011989 5.6702e-005 0.0011586 0.22861 0.00065927 0.22927 0.21143 0 0.032514 0.0389 0 1.2019 0.38976 0.11647 0.014881 7.5578 0.092838 0.0001163 0.79728 0.0073348 0.0081826 0.0015565 0.98469 0.99018 3.3802e-006 1.3521e-005 0.14865 0.72167 0.79948 0.0014846 0.82909 0.44706 0.0019967 0.42191 1.4673 1.464 16.0079 144.9565 0.00034349 -84.9572 0.22794
4.332 0.98807 5.4971e-005 3.8183 0.011989 5.6715e-005 0.0011586 0.22862 0.00065927 0.22927 0.21143 0 0.032514 0.0389 0 1.202 0.38981 0.11649 0.014882 7.5595 0.092848 0.00011631 0.79727 0.0073355 0.0081833 0.0015552 0.98471 0.99019 3.3771e-006 1.3509e-005 0.14866 0.72249 0.80006 0.001484 0.83011 0.44725 0.0019959 0.42192 1.469 1.4658 16.0079 144.9565 0.00034265 -84.9623 0.22894
4.333 0.98807 5.497e-005 3.8183 0.011989 5.6728e-005 0.0011586 0.22862 0.00065927 0.22928 0.21144 0 0.032514 0.0389 0 1.2021 0.38985 0.11651 0.014884 7.5612 0.092858 0.00011633 0.79726 0.0073362 0.008184 0.0015539 0.98473 0.99021 3.3741e-006 1.3497e-005 0.14866 0.7233 0.80063 0.0014833 0.83112 0.44743 0.001995 0.42193 1.4708 1.4675 16.008 144.9565 0.0003418 -84.9674 0.22994
4.334 0.98807 5.497e-005 3.8183 0.011989 5.6741e-005 0.0011586 0.22863 0.00065927 0.22928 0.21144 0 0.032513 0.0389 0 1.2022 0.3899 0.11652 0.014886 7.5628 0.092868 0.00011634 0.79725 0.0073369 0.0081847 0.0015526 0.98475 0.99022 3.3711e-006 1.3485e-005 0.14867 0.72411 0.8012 0.0014827 0.83212 0.44762 0.0019941 0.42194 1.4725 1.4692 16.008 144.9566 0.00034097 -84.9725 0.23094
4.335 0.98807 5.497e-005 3.8183 0.011989 5.6754e-005 0.0011586 0.22863 0.00065927 0.22929 0.21145 0 0.032513 0.0389 0 1.2023 0.38995 0.11654 0.014887 7.5645 0.092878 0.00011635 0.79724 0.0073375 0.0081855 0.0015513 0.98477 0.99023 3.3681e-006 1.3473e-005 0.14867 0.72491 0.80177 0.001482 0.83312 0.44781 0.0019933 0.42195 1.4742 1.4709 16.008 144.9566 0.00034013 -84.9775 0.23194
4.336 0.98807 5.497e-005 3.8183 0.011989 5.6767e-005 0.0011586 0.22864 0.00065927 0.22929 0.21145 0 0.032513 0.0389 0 1.2024 0.38999 0.11655 0.014889 7.5662 0.092887 0.00011637 0.79723 0.0073382 0.0081862 0.00155 0.98478 0.99025 3.3651e-006 1.3461e-005 0.14868 0.72572 0.80234 0.0014814 0.83412 0.448 0.0019924 0.42195 1.4759 1.4726 16.0081 144.9566 0.0003393 -84.9824 0.23294
4.337 0.98807 5.497e-005 3.8183 0.011989 5.678e-005 0.0011586 0.22864 0.00065927 0.2293 0.21146 0 0.032513 0.0389 0 1.2025 0.39004 0.11657 0.014891 7.5678 0.092897 0.00011638 0.79722 0.0073389 0.0081869 0.0015487 0.9848 0.99026 3.3622e-006 1.3449e-005 0.14868 0.72652 0.8029 0.0014807 0.83511 0.44819 0.0019916 0.42196 1.4775 1.4743 16.0081 144.9566 0.00033847 -84.9874 0.23394
4.338 0.98807 5.497e-005 3.8183 0.011989 5.6793e-005 0.0011587 0.22865 0.00065927 0.2293 0.21146 0 0.032512 0.0389 0 1.2026 0.39009 0.11659 0.014892 7.5695 0.092907 0.00011639 0.79721 0.0073396 0.0081877 0.0015474 0.98482 0.99027 3.3593e-006 1.3437e-005 0.14869 0.72732 0.80346 0.0014801 0.83609 0.44837 0.0019908 0.42197 1.4792 1.476 16.0081 144.9566 0.00033765 -84.9923 0.23494
4.339 0.98807 5.497e-005 3.8183 0.011989 5.6806e-005 0.0011587 0.22865 0.00065927 0.22931 0.21146 0 0.032512 0.0389 0 1.2027 0.39013 0.1166 0.014894 7.5712 0.092917 0.00011641 0.7972 0.0073402 0.0081884 0.0015462 0.98483 0.99029 3.3564e-006 1.3426e-005 0.14869 0.72812 0.80402 0.0014795 0.83707 0.44856 0.00199 0.42198 1.4809 1.4777 16.0082 144.9566 0.00033683 -84.9971 0.23594
4.34 0.98807 5.497e-005 3.8183 0.011989 5.6819e-005 0.0011587 0.22866 0.00065927 0.22931 0.21147 0 0.032512 0.0389 0 1.2028 0.39018 0.11662 0.014895 7.5729 0.092927 0.00011642 0.79719 0.0073409 0.0081891 0.0015449 0.98485 0.9903 3.3535e-006 1.3414e-005 0.1487 0.72891 0.80457 0.0014788 0.83804 0.44875 0.0019891 0.42199 1.4826 1.4794 16.0082 144.9567 0.00033602 -85.002 0.23694
4.341 0.98807 5.497e-005 3.8183 0.011989 5.6832e-005 0.0011587 0.22866 0.00065927 0.22932 0.21147 0 0.032512 0.0389 0 1.2028 0.39023 0.11663 0.014897 7.5745 0.092937 0.00011644 0.79718 0.0073416 0.0081898 0.0015437 0.98487 0.99031 3.3507e-006 1.3403e-005 0.1487 0.7297 0.80512 0.0014782 0.83901 0.44894 0.0019883 0.422 1.4843 1.4811 16.0082 144.9567 0.00033521 -85.0067 0.23794
4.342 0.98807 5.497e-005 3.8183 0.011988 5.6845e-005 0.0011587 0.22867 0.00065927 0.22932 0.21148 0 0.032511 0.0389 0 1.2029 0.39027 0.11665 0.014899 7.5762 0.092947 0.00011645 0.79717 0.0073423 0.0081906 0.0015425 0.98488 0.99032 3.3479e-006 1.3392e-005 0.14871 0.73049 0.80567 0.0014776 0.83997 0.44913 0.0019875 0.42201 1.4859 1.4828 16.0083 144.9567 0.0003344 -85.0115 0.23894
4.343 0.98807 5.497e-005 3.8183 0.011988 5.6858e-005 0.0011587 0.22867 0.00065927 0.22933 0.21148 0 0.032511 0.0389 0 1.203 0.39032 0.11667 0.0149 7.5779 0.092957 0.00011646 0.79716 0.007343 0.0081913 0.0015413 0.9849 0.99033 3.3451e-006 1.3381e-005 0.14872 0.73128 0.80621 0.001477 0.84093 0.44931 0.0019867 0.42201 1.4876 1.4845 16.0083 144.9567 0.0003336 -85.0162 0.23994
4.344 0.98807 5.497e-005 3.8183 0.011988 5.6871e-005 0.0011587 0.22868 0.00065927 0.22933 0.21149 0 0.032511 0.0389 0 1.2031 0.39037 0.11668 0.014902 7.5795 0.092967 0.00011648 0.79715 0.0073436 0.008192 0.0015401 0.98492 0.99035 3.3423e-006 1.337e-005 0.14872 0.73206 0.80676 0.0014764 0.84188 0.4495 0.0019859 0.42202 1.4893 1.4861 16.0083 144.9567 0.0003328 -85.0209 0.24094
4.345 0.98807 5.497e-005 3.8183 0.011988 5.6884e-005 0.0011587 0.22868 0.00065927 0.22934 0.21149 0 0.032511 0.0389 0 1.2032 0.39041 0.1167 0.014903 7.5812 0.092977 0.00011649 0.79714 0.0073443 0.0081928 0.0015389 0.98493 0.99036 3.3396e-006 1.3359e-005 0.14873 0.73285 0.80729 0.0014758 0.84283 0.44969 0.0019852 0.42203 1.4909 1.4878 16.0084 144.9567 0.000332 -85.0255 0.24194
4.346 0.98807 5.497e-005 3.8183 0.011988 5.6897e-005 0.0011587 0.22869 0.00065927 0.22934 0.2115 0 0.03251 0.0389 0 1.2033 0.39046 0.11671 0.014905 7.5829 0.092987 0.00011651 0.79713 0.007345 0.0081935 0.0015377 0.98495 0.99037 3.3368e-006 1.3348e-005 0.14873 0.73363 0.80783 0.0014752 0.84377 0.44988 0.0019844 0.42204 1.4926 1.4895 16.0084 144.9567 0.00033121 -85.0301 0.24294
4.347 0.98807 5.4969e-005 3.8183 0.011988 5.691e-005 0.0011587 0.22869 0.00065927 0.22935 0.2115 0 0.03251 0.0389 0 1.2034 0.39051 0.11673 0.014907 7.5845 0.092997 0.00011652 0.79712 0.0073457 0.0081942 0.0015365 0.98496 0.99038 3.3341e-006 1.3337e-005 0.14874 0.7344 0.80836 0.0014746 0.8447 0.45006 0.0019836 0.42205 1.4942 1.4911 16.0084 144.9568 0.00033043 -85.0347 0.24394
4.348 0.98807 5.4969e-005 3.8183 0.011988 5.6923e-005 0.0011587 0.2287 0.00065927 0.22935 0.21151 0 0.03251 0.0389 0 1.2035 0.39055 0.11674 0.014908 7.5862 0.093007 0.00011653 0.79711 0.0073463 0.0081949 0.0015354 0.98498 0.99039 3.3315e-006 1.3326e-005 0.14874 0.73518 0.80889 0.001474 0.84563 0.45025 0.0019828 0.42206 1.4959 1.4928 16.0085 144.9568 0.00032964 -85.0393 0.24494
4.349 0.98807 5.4969e-005 3.8183 0.011988 5.6936e-005 0.0011587 0.2287 0.00065927 0.22936 0.21151 0 0.03251 0.0389 0 1.2036 0.3906 0.11676 0.01491 7.5879 0.093017 0.00011655 0.7971 0.007347 0.0081957 0.0015342 0.985 0.9904 3.3288e-006 1.3315e-005 0.14875 0.73595 0.80942 0.0014734 0.84656 0.45044 0.0019821 0.42207 1.4975 1.4944 16.0085 144.9568 0.00032886 -85.0438 0.24594
4.35 0.98807 5.4969e-005 3.8183 0.011988 5.6949e-005 0.0011587 0.22871 0.00065927 0.22936 0.21152 0 0.032509 0.0389 0 1.2037 0.39065 0.11678 0.014911 7.5896 0.093027 0.00011656 0.79709 0.0073477 0.0081964 0.0015331 0.98501 0.99042 3.3262e-006 1.3305e-005 0.14875 0.73672 0.80994 0.0014729 0.84748 0.45063 0.0019813 0.42207 1.4992 1.4961 16.0085 144.9568 0.00032809 -85.0482 0.24694
4.351 0.98807 5.4969e-005 3.8183 0.011988 5.6962e-005 0.0011587 0.22871 0.00065927 0.22937 0.21152 0 0.032509 0.0389 0 1.2038 0.39069 0.11679 0.014913 7.5912 0.093037 0.00011658 0.79708 0.0073484 0.0081971 0.001532 0.98503 0.99043 3.3236e-006 1.3294e-005 0.14876 0.73749 0.81046 0.0014723 0.84839 0.45082 0.0019806 0.42208 1.5008 1.4977 16.0086 144.9568 0.00032731 -85.0527 0.24794
4.352 0.98807 5.4969e-005 3.8183 0.011988 5.6975e-005 0.0011587 0.22872 0.00065927 0.22937 0.21153 0 0.032509 0.0389 0 1.2039 0.39074 0.11681 0.014915 7.5929 0.093047 0.00011659 0.79707 0.007349 0.0081978 0.0015308 0.98504 0.99044 3.321e-006 1.3284e-005 0.14876 0.73826 0.81098 0.0014717 0.8493 0.451 0.0019798 0.42209 1.5024 1.4994 16.0086 144.9568 0.00032655 -85.0571 0.24894
4.353 0.98807 5.4969e-005 3.8183 0.011988 5.6988e-005 0.0011587 0.22872 0.00065927 0.22938 0.21153 0 0.032509 0.0389 0 1.204 0.39079 0.11682 0.014916 7.5946 0.093057 0.0001166 0.79706 0.0073497 0.0081986 0.0015297 0.98506 0.99045 3.3184e-006 1.3274e-005 0.14877 0.73902 0.81149 0.0014712 0.85021 0.45119 0.0019791 0.4221 1.504 1.501 16.0086 144.9569 0.00032578 -85.0615 0.24994
4.354 0.98807 5.4969e-005 3.8183 0.011988 5.7001e-005 0.0011587 0.22873 0.00065927 0.22938 0.21153 0 0.032508 0.0389 0 1.2041 0.39083 0.11684 0.014918 7.5963 0.093067 0.00011662 0.79705 0.0073504 0.0081993 0.0015286 0.98507 0.99046 3.3159e-006 1.3264e-005 0.14878 0.73978 0.81201 0.0014706 0.85111 0.45138 0.0019784 0.42211 1.5057 1.5026 16.0087 144.9569 0.00032502 -85.0658 0.25094
4.355 0.98807 5.4969e-005 3.8183 0.011988 5.7014e-005 0.0011587 0.22873 0.00065927 0.22939 0.21154 0 0.032508 0.0389 0 1.2042 0.39088 0.11686 0.014919 7.5979 0.093077 0.00011663 0.79704 0.0073511 0.0082 0.0015275 0.98509 0.99047 3.3133e-006 1.3254e-005 0.14878 0.74054 0.81252 0.00147 0.852 0.45157 0.0019776 0.42212 1.5073 1.5043 16.0087 144.9569 0.00032426 -85.0701 0.25194
4.356 0.98807 5.4969e-005 3.8183 0.011988 5.7027e-005 0.0011587 0.22874 0.00065927 0.22939 0.21154 0 0.032508 0.0389 0 1.2043 0.39093 0.11687 0.014921 7.5996 0.093087 0.00011665 0.79703 0.0073517 0.0082008 0.0015264 0.9851 0.99048 3.3108e-006 1.3244e-005 0.14879 0.74129 0.81302 0.0014695 0.85289 0.45175 0.0019769 0.42213 1.5089 1.5059 16.0087 144.9569 0.00032351 -85.0744 0.25294
4.357 0.98807 5.4969e-005 3.8183 0.011988 5.704e-005 0.0011587 0.22874 0.00065927 0.2294 0.21155 0 0.032508 0.0389 0 1.2044 0.39097 0.11689 0.014923 7.6013 0.093097 0.00011666 0.79702 0.0073524 0.0082015 0.0015253 0.98512 0.99049 3.3084e-006 1.3234e-005 0.14879 0.74205 0.81353 0.001469 0.85377 0.45194 0.0019762 0.42214 1.5105 1.5075 16.0087 144.9569 0.00032276 -85.0786 0.25394
4.358 0.98807 5.4969e-005 3.8183 0.011988 5.7053e-005 0.0011587 0.22875 0.00065927 0.2294 0.21155 0 0.032507 0.0389 0 1.2045 0.39102 0.1169 0.014924 7.6029 0.093107 0.00011667 0.79701 0.0073531 0.0082022 0.0015243 0.98513 0.9905 3.3059e-006 1.3224e-005 0.1488 0.7428 0.81403 0.0014684 0.85465 0.45213 0.0019755 0.42215 1.5121 1.5091 16.0088 144.9569 0.00032201 -85.0828 0.25494
4.359 0.98807 5.4969e-005 3.8183 0.011988 5.7066e-005 0.0011587 0.22875 0.00065927 0.22941 0.21156 0 0.032507 0.0389 0 1.2046 0.39107 0.11692 0.014926 7.6046 0.093117 0.00011669 0.797 0.0073538 0.0082029 0.0015232 0.98514 0.99051 3.3034e-006 1.3214e-005 0.1488 0.74355 0.81453 0.0014679 0.85553 0.45231 0.0019748 0.42216 1.5137 1.5107 16.0088 144.957 0.00032127 -85.087 0.25594
4.36 0.98807 5.4969e-005 3.8183 0.011988 5.7079e-005 0.0011587 0.22876 0.00065927 0.22941 0.21156 0 0.032507 0.0389 0 1.2047 0.39111 0.11694 0.014928 7.6063 0.093127 0.0001167 0.79699 0.0073544 0.0082037 0.0015222 0.98516 0.99052 3.301e-006 1.3204e-005 0.14881 0.7443 0.81502 0.0014673 0.8564 0.4525 0.0019741 0.42217 1.5153 1.5123 16.0088 144.957 0.00032053 -85.0911 0.25694
4.361 0.98807 5.4968e-005 3.8183 0.011988 5.7092e-005 0.0011587 0.22876 0.00065927 0.22942 0.21157 0 0.032507 0.0389 0 1.2048 0.39116 0.11695 0.014929 7.608 0.093137 0.00011672 0.79698 0.0073551 0.0082044 0.0015211 0.98517 0.99053 3.2986e-006 1.3195e-005 0.14881 0.74504 0.81551 0.0014668 0.85726 0.45269 0.0019734 0.42218 1.5169 1.5139 16.0089 144.957 0.00031979 -85.0953 0.25794
4.362 0.98807 5.4968e-005 3.8183 0.011988 5.7105e-005 0.0011587 0.22877 0.00065927 0.22942 0.21157 0 0.032506 0.0389 0 1.2049 0.39121 0.11697 0.014931 7.6097 0.093147 0.00011673 0.79697 0.0073558 0.0082051 0.0015201 0.98519 0.99054 3.2962e-006 1.3185e-005 0.14882 0.74578 0.81601 0.0014663 0.85812 0.45288 0.0019727 0.42218 1.5185 1.5155 16.0089 144.957 0.00031906 -85.0994 0.25894
4.363 0.98807 5.4968e-005 3.8183 0.011988 5.7118e-005 0.0011587 0.22877 0.00065927 0.22943 0.21158 0 0.032506 0.0389 0 1.205 0.39125 0.11698 0.014932 7.6113 0.093157 0.00011674 0.79696 0.0073565 0.0082058 0.0015191 0.9852 0.99055 3.2939e-006 1.3176e-005 0.14882 0.74652 0.81649 0.0014658 0.85897 0.45306 0.001972 0.42219 1.5201 1.5171 16.0089 144.957 0.00031833 -85.1034 0.25994
4.364 0.98807 5.4968e-005 3.8183 0.011988 5.7131e-005 0.0011587 0.22878 0.00065927 0.22943 0.21158 0 0.032506 0.0389 0 1.2051 0.3913 0.117 0.014934 7.613 0.093166 0.00011676 0.79695 0.0073571 0.0082066 0.001518 0.98521 0.99056 3.2915e-006 1.3166e-005 0.14883 0.74726 0.81698 0.0014653 0.85982 0.45325 0.0019714 0.4222 1.5216 1.5187 16.0089 144.957 0.0003176 -85.1074 0.26094
4.365 0.98807 5.4968e-005 3.8183 0.011988 5.7144e-005 0.0011587 0.22878 0.00065927 0.22943 0.21159 0 0.032506 0.0389 0 1.2052 0.39135 0.11702 0.014936 7.6147 0.093176 0.00011677 0.79694 0.0073578 0.0082073 0.001517 0.98523 0.99057 3.2892e-006 1.3157e-005 0.14883 0.748 0.81746 0.0014647 0.86067 0.45344 0.0019707 0.42221 1.5232 1.5203 16.009 144.9571 0.00031688 -85.1114 0.26194
4.366 0.98807 5.4968e-005 3.8183 0.011988 5.7157e-005 0.0011587 0.22878 0.00065927 0.22944 0.21159 0 0.032505 0.0389 0 1.2053 0.39139 0.11703 0.014937 7.6164 0.093186 0.00011679 0.79693 0.0073585 0.008208 0.001516 0.98524 0.99058 3.2869e-006 1.3148e-005 0.14884 0.74873 0.81794 0.0014642 0.86151 0.45362 0.00197 0.42222 1.5248 1.5219 16.009 144.9571 0.00031616 -85.1154 0.26294
4.367 0.98807 5.4968e-005 3.8183 0.011988 5.717e-005 0.0011587 0.22879 0.00065927 0.22944 0.21159 0 0.032505 0.0389 0 1.2054 0.39144 0.11705 0.014939 7.618 0.093196 0.0001168 0.79692 0.0073592 0.0082087 0.001515 0.98525 0.99058 3.2846e-006 1.3139e-005 0.14885 0.74946 0.81842 0.0014637 0.86234 0.45381 0.0019694 0.42223 1.5264 1.5235 16.009 144.9571 0.00031545 -85.1193 0.26394
4.368 0.98807 5.4968e-005 3.8183 0.011988 5.7183e-005 0.0011587 0.22879 0.00065927 0.22945 0.2116 0 0.032505 0.0389 0 1.2055 0.39149 0.11706 0.01494 7.6197 0.093206 0.00011681 0.79691 0.0073598 0.0082095 0.001514 0.98527 0.99059 3.2823e-006 1.3129e-005 0.14885 0.75019 0.81889 0.0014632 0.86317 0.454 0.0019687 0.42224 1.5279 1.525 16.009 144.9571 0.00031473 -85.1232 0.26494
4.369 0.98807 5.4968e-005 3.8183 0.011988 5.7196e-005 0.0011587 0.2288 0.00065927 0.22945 0.2116 0 0.032505 0.0389 0 1.2056 0.39153 0.11708 0.014942 7.6214 0.093216 0.00011683 0.7969 0.0073605 0.0082102 0.0015131 0.98528 0.9906 3.2801e-006 1.312e-005 0.14886 0.75091 0.81937 0.0014627 0.86399 0.45419 0.0019681 0.42225 1.5295 1.5266 16.0091 144.9571 0.00031403 -85.1271 0.26594
4.37 0.98807 5.4968e-005 3.8183 0.011988 5.7209e-005 0.0011587 0.2288 0.00065927 0.22946 0.21161 0 0.032504 0.0389 0 1.2057 0.39158 0.11709 0.014944 7.6231 0.093226 0.00011684 0.79689 0.0073612 0.0082109 0.0015121 0.98529 0.99061 3.2778e-006 1.3112e-005 0.14886 0.75164 0.81984 0.0014622 0.86482 0.45437 0.0019674 0.42226 1.531 1.5282 16.0091 144.9571 0.00031332 -85.131 0.26694
4.371 0.98807 5.4968e-005 3.8183 0.011988 5.7222e-005 0.0011587 0.22881 0.00065927 0.22946 0.21161 0 0.032504 0.0389 0 1.2058 0.39163 0.11711 0.014945 7.6248 0.093236 0.00011685 0.79688 0.0073619 0.0082117 0.0015111 0.98531 0.99062 3.2756e-006 1.3103e-005 0.14887 0.75236 0.82031 0.0014617 0.86563 0.45456 0.0019668 0.42227 1.5326 1.5297 16.0091 144.9571 0.00031262 -85.1348 0.26794
4.372 0.98807 5.4968e-005 3.8183 0.011988 5.7235e-005 0.0011587 0.22881 0.00065927 0.22947 0.21162 0 0.032504 0.0389 0 1.2059 0.39167 0.11713 0.014947 7.6264 0.093246 0.00011687 0.79687 0.0073625 0.0082124 0.0015102 0.98532 0.99063 3.2734e-006 1.3094e-005 0.14887 0.75308 0.82077 0.0014613 0.86644 0.45475 0.0019662 0.42228 1.5341 1.5313 16.0091 144.9572 0.00031192 -85.1386 0.26894
4.373 0.98807 5.4968e-005 3.8183 0.011988 5.7248e-005 0.0011587 0.22882 0.00065927 0.22947 0.21162 0 0.032504 0.0389 0 1.206 0.39172 0.11714 0.014948 7.6281 0.093256 0.00011688 0.79686 0.0073632 0.0082131 0.0015092 0.98533 0.99064 3.2712e-006 1.3085e-005 0.14888 0.7538 0.82123 0.0014608 0.86725 0.45493 0.0019655 0.42229 1.5357 1.5328 16.0092 144.9572 0.00031122 -85.1423 0.26994
4.374 0.98807 5.4968e-005 3.8183 0.011988 5.7261e-005 0.0011587 0.22882 0.00065927 0.22948 0.21163 0 0.032503 0.0389 0 1.2061 0.39177 0.11716 0.01495 7.6298 0.093266 0.0001169 0.79685 0.0073639 0.0082138 0.0015083 0.98534 0.99065 3.2691e-006 1.3076e-005 0.14888 0.75451 0.82169 0.0014603 0.86805 0.45512 0.0019649 0.4223 1.5372 1.5344 16.0092 144.9572 0.00031053 -85.1461 0.27094
4.375 0.98807 5.4967e-005 3.8183 0.011988 5.7273e-005 0.0011587 0.22883 0.00065927 0.22948 0.21163 0 0.032503 0.0389 0 1.2062 0.39181 0.11717 0.014952 7.6315 0.093276 0.00011691 0.79684 0.0073646 0.0082146 0.0015074 0.98536 0.99066 3.2669e-006 1.3068e-005 0.14889 0.75522 0.82215 0.0014598 0.86885 0.45531 0.0019643 0.42231 1.5388 1.5359 16.0092 144.9572 0.00030984 -85.1498 0.27194
4.376 0.98807 5.4967e-005 3.8183 0.011988 5.7286e-005 0.0011587 0.22883 0.00065927 0.22949 0.21164 0 0.032503 0.0389 0 1.2063 0.39186 0.11719 0.014953 7.6332 0.093286 0.00011692 0.79683 0.0073652 0.0082153 0.0015064 0.98537 0.99066 3.2648e-006 1.3059e-005 0.14889 0.75594 0.82261 0.0014594 0.86964 0.45549 0.0019637 0.42232 1.5403 1.5375 16.0092 144.9572 0.00030916 -85.1535 0.27294
4.377 0.98807 5.4967e-005 3.8183 0.011988 5.7299e-005 0.0011587 0.22884 0.00065927 0.22949 0.21164 0 0.032503 0.0389 0 1.2064 0.39191 0.11721 0.014955 7.6348 0.093296 0.00011694 0.79682 0.0073659 0.008216 0.0015055 0.98538 0.99067 3.2627e-006 1.3051e-005 0.1489 0.75664 0.82306 0.0014589 0.87043 0.45568 0.0019631 0.42233 1.5418 1.539 16.0093 144.9572 0.00030847 -85.1571 0.27394
4.378 0.98807 5.4967e-005 3.8183 0.011988 5.7312e-005 0.0011588 0.22884 0.00065927 0.2295 0.21165 0 0.032502 0.0389 0 1.2065 0.39195 0.11722 0.014956 7.6365 0.093306 0.00011695 0.79681 0.0073666 0.0082167 0.0015046 0.98539 0.99068 3.2606e-006 1.3043e-005 0.1489 0.75735 0.82351 0.0014584 0.87121 0.45587 0.0019625 0.42234 1.5433 1.5406 16.0093 144.9573 0.0003078 -85.1608 0.27494
4.379 0.98807 5.4967e-005 3.8183 0.011988 5.7325e-005 0.0011588 0.22885 0.00065927 0.2295 0.21165 0 0.032502 0.0389 0 1.2066 0.392 0.11724 0.014958 7.6382 0.093316 0.00011697 0.7968 0.0073672 0.0082175 0.0015037 0.9854 0.99069 3.2585e-006 1.3034e-005 0.14891 0.75805 0.82396 0.001458 0.87199 0.45605 0.0019619 0.42235 1.5449 1.5421 16.0093 144.9573 0.00030712 -85.1644 0.27594
4.38 0.98807 5.4967e-005 3.8183 0.011988 5.7338e-005 0.0011588 0.22885 0.00065927 0.22951 0.21165 0 0.032502 0.0389 0 1.2067 0.39205 0.11725 0.01496 7.6399 0.093326 0.00011698 0.79679 0.0073679 0.0082182 0.0015028 0.98542 0.9907 3.2565e-006 1.3026e-005 0.14892 0.75876 0.82441 0.0014575 0.87276 0.45624 0.0019613 0.42236 1.5464 1.5436 16.0093 144.9573 0.00030645 -85.1679 0.27694
4.381 0.98807 5.4967e-005 3.8183 0.011988 5.7351e-005 0.0011588 0.22886 0.00065927 0.22951 0.21166 0 0.032502 0.0389 0 1.2068 0.39209 0.11727 0.014961 7.6416 0.093335 0.00011699 0.79678 0.0073686 0.0082189 0.0015019 0.98543 0.9907 3.2544e-006 1.3018e-005 0.14892 0.75946 0.82485 0.0014571 0.87353 0.45642 0.0019607 0.42237 1.5479 1.5451 16.0094 144.9573 0.00030578 -85.1715 0.27794
4.382 0.98807 5.4967e-005 3.8183 0.011988 5.7364e-005 0.0011588 0.22886 0.00065927 0.22952 0.21166 0 0.032502 0.0389 0 1.2069 0.39214 0.11729 0.014963 7.6433 0.093345 0.00011701 0.79677 0.0073693 0.0082196 0.001501 0.98544 0.99071 3.2524e-006 1.301e-005 0.14893 0.76015 0.82529 0.0014566 0.8743 0.45661 0.0019601 0.42238 1.5494 1.5466 16.0094 144.9573 0.00030511 -85.175 0.27894
4.383 0.98807 5.4967e-005 3.8183 0.011988 5.7377e-005 0.0011588 0.22887 0.00065927 0.22952 0.21167 0 0.032501 0.0389 0 1.207 0.39219 0.1173 0.014964 7.6449 0.093355 0.00011702 0.79676 0.0073699 0.0082204 0.0015002 0.98545 0.99072 3.2504e-006 1.3002e-005 0.14893 0.76085 0.82573 0.0014562 0.87506 0.4568 0.0019595 0.42239 1.5509 1.5482 16.0094 144.9573 0.00030445 -85.1785 0.27994
4.384 0.98807 5.4967e-005 3.8183 0.011988 5.739e-005 0.0011588 0.22887 0.00065927 0.22953 0.21167 0 0.032501 0.0389 0 1.2071 0.39223 0.11732 0.014966 7.6466 0.093365 0.00011704 0.79675 0.0073706 0.0082211 0.0014993 0.98546 0.99073 3.2484e-006 1.2994e-005 0.14894 0.76154 0.82617 0.0014557 0.87581 0.45698 0.0019589 0.4224 1.5524 1.5497 16.0094 144.9574 0.00030379 -85.182 0.28094
4.385 0.98807 5.4967e-005 3.8183 0.011988 5.7403e-005 0.0011588 0.22888 0.00065927 0.22953 0.21168 0 0.032501 0.0389 0 1.2072 0.39228 0.11733 0.014968 7.6483 0.093375 0.00011705 0.79674 0.0073713 0.0082218 0.0014984 0.98547 0.99074 3.2464e-006 1.2986e-005 0.14894 0.76223 0.82661 0.0014553 0.87657 0.45717 0.0019583 0.42241 1.5539 1.5512 16.0095 144.9574 0.00030313 -85.1854 0.28194
4.386 0.98807 5.4967e-005 3.8183 0.011988 5.7416e-005 0.0011588 0.22888 0.00065927 0.22954 0.21168 0 0.032501 0.0389 0 1.2073 0.39233 0.11735 0.014969 7.65 0.093385 0.00011706 0.79673 0.007372 0.0082225 0.0014976 0.98549 0.99074 3.2445e-006 1.2978e-005 0.14895 0.76292 0.82704 0.0014549 0.87731 0.45736 0.0019578 0.42242 1.5554 1.5527 16.0095 144.9574 0.00030247 -85.1888 0.28294
4.387 0.98807 5.4967e-005 3.8183 0.011988 5.7429e-005 0.0011588 0.22889 0.00065927 0.22954 0.21169 0 0.0325 0.0389 0 1.2074 0.39237 0.11736 0.014971 7.6517 0.093395 0.00011708 0.79672 0.0073726 0.0082233 0.0014967 0.9855 0.99075 3.2425e-006 1.297e-005 0.14895 0.76361 0.82747 0.0014544 0.87806 0.45754 0.0019572 0.42243 1.5569 1.5542 16.0095 144.9574 0.00030182 -85.1922 0.28394
4.388 0.98807 5.4966e-005 3.8183 0.011988 5.7442e-005 0.0011588 0.22889 0.00065927 0.22955 0.21169 0 0.0325 0.0389 0 1.2074 0.39242 0.11738 0.014973 7.6534 0.093405 0.00011709 0.79671 0.0073733 0.008224 0.0014959 0.98551 0.99076 3.2406e-006 1.2962e-005 0.14896 0.76429 0.8279 0.001454 0.8788 0.45773 0.0019566 0.42244 1.5584 1.5557 16.0095 144.9574 0.00030117 -85.1956 0.28494
4.389 0.98807 5.4966e-005 3.8183 0.011988 5.7455e-005 0.0011588 0.2289 0.00065927 0.22955 0.2117 0 0.0325 0.0389 0 1.2075 0.39247 0.1174 0.014974 7.6551 0.093415 0.0001171 0.7967 0.007374 0.0082247 0.0014951 0.98552 0.99077 3.2387e-006 1.2955e-005 0.14896 0.76498 0.82832 0.0014536 0.87953 0.45791 0.0019561 0.42245 1.5598 1.5572 16.0095 144.9574 0.00030053 -85.1989 0.28594
4.39 0.98807 5.4966e-005 3.8183 0.011988 5.7468e-005 0.0011588 0.2289 0.00065927 0.22955 0.2117 0 0.0325 0.0389 0 1.2076 0.39251 0.11741 0.014976 7.6567 0.093425 0.00011712 0.79669 0.0073747 0.0082254 0.0014942 0.98553 0.99077 3.2367e-006 1.2947e-005 0.14897 0.76566 0.82875 0.0014531 0.88026 0.4581 0.0019555 0.42246 1.5613 1.5586 16.0096 144.9575 0.00029989 -85.2022 0.28694
4.391 0.98807 5.4966e-005 3.8183 0.011988 5.7481e-005 0.0011588 0.2289 0.00065927 0.22956 0.2117 0 0.032499 0.0389 0 1.2077 0.39256 0.11743 0.014977 7.6584 0.093435 0.00011713 0.79668 0.0073753 0.0082262 0.0014934 0.98554 0.99078 3.2349e-006 1.294e-005 0.14897 0.76634 0.82917 0.0014527 0.88099 0.45829 0.001955 0.42247 1.5628 1.5601 16.0096 144.9575 0.00029925 -85.2055 0.28794
4.392 0.98807 5.4966e-005 3.8183 0.011988 5.7494e-005 0.0011588 0.22891 0.00065927 0.22956 0.21171 0 0.032499 0.0389 0 1.2078 0.39261 0.11744 0.014979 7.6601 0.093445 0.00011715 0.79667 0.007376 0.0082269 0.0014926 0.98555 0.99079 3.233e-006 1.2932e-005 0.14898 0.76701 0.82959 0.0014523 0.88171 0.45847 0.0019544 0.42249 1.5642 1.5616 16.0096 144.9575 0.00029861 -85.2088 0.28894
4.393 0.98807 5.4966e-005 3.8183 0.011988 5.7507e-005 0.0011588 0.22891 0.00065927 0.22957 0.21171 0 0.032499 0.0389 0 1.2079 0.39265 0.11746 0.014981 7.6618 0.093455 0.00011716 0.79666 0.0073767 0.0082276 0.0014918 0.98556 0.9908 3.2311e-006 1.2925e-005 0.14898 0.76769 0.83001 0.0014519 0.88243 0.45866 0.0019539 0.4225 1.5657 1.5631 16.0096 144.9575 0.00029798 -85.2121 0.28994
4.394 0.98807 5.4966e-005 3.8183 0.011988 5.752e-005 0.0011588 0.22892 0.00065927 0.22957 0.21172 0 0.032499 0.0389 0 1.208 0.3927 0.11748 0.014982 7.6635 0.093465 0.00011717 0.79665 0.0073773 0.0082283 0.001491 0.98557 0.9908 3.2293e-006 1.2917e-005 0.14899 0.76836 0.83042 0.0014515 0.88314 0.45884 0.0019534 0.42251 1.5672 1.5645 16.0096 144.9575 0.00029735 -85.2153 0.29094
4.395 0.98807 5.4966e-005 3.8183 0.011988 5.7533e-005 0.0011588 0.22892 0.00065927 0.22958 0.21172 0 0.032498 0.0389 0 1.2081 0.39275 0.11749 0.014984 7.6652 0.093474 0.00011719 0.79664 0.007378 0.008229 0.0014902 0.98558 0.99081 3.2275e-006 1.291e-005 0.149 0.76903 0.83084 0.0014511 0.88385 0.45903 0.0019528 0.42252 1.5686 1.566 16.0097 144.9576 0.00029672 -85.2185 0.29194
4.396 0.98807 5.4966e-005 3.8183 0.011988 5.7546e-005 0.0011588 0.22893 0.00065927 0.22958 0.21173 0 0.032498 0.0389 0 1.2082 0.39279 0.11751 0.014985 7.6669 0.093484 0.0001172 0.79663 0.0073787 0.0082298 0.0014894 0.98559 0.99082 3.2257e-006 1.2903e-005 0.149 0.7697 0.83125 0.0014507 0.88455 0.45922 0.0019523 0.42253 1.5701 1.5675 16.0097 144.9576 0.00029609 -85.2217 0.29294
4.397 0.98807 5.4966e-005 3.8183 0.011988 5.7559e-005 0.0011588 0.22893 0.00065927 0.22959 0.21173 0 0.032498 0.0389 0 1.2083 0.39284 0.11752 0.014987 7.6686 0.093494 0.00011722 0.79662 0.0073794 0.0082305 0.0014886 0.98561 0.99082 3.2239e-006 1.2896e-005 0.14901 0.77036 0.83166 0.0014503 0.88525 0.4594 0.0019518 0.42254 1.5715 1.5689 16.0097 144.9576 0.00029547 -85.2248 0.29394
4.398 0.98807 5.4966e-005 3.8183 0.011988 5.7572e-005 0.0011588 0.22894 0.00065927 0.22959 0.21174 0 0.032498 0.0389 0 1.2084 0.39289 0.11754 0.014989 7.6703 0.093504 0.00011723 0.79661 0.00738 0.0082312 0.0014879 0.98562 0.99083 3.2221e-006 1.2888e-005 0.14901 0.77103 0.83207 0.0014499 0.88595 0.45959 0.0019513 0.42255 1.573 1.5704 16.0097 144.9576 0.00029485 -85.2279 0.29494
4.399 0.98807 5.4966e-005 3.8183 0.011988 5.7585e-005 0.0011588 0.22894 0.00065927 0.2296 0.21174 0 0.032497 0.0389 0 1.2085 0.39293 0.11756 0.01499 7.6719 0.093514 0.00011724 0.7966 0.0073807 0.0082319 0.0014871 0.98563 0.99084 3.2203e-006 1.2881e-005 0.14902 0.77169 0.83247 0.0014495 0.88664 0.45977 0.0019508 0.42256 1.5744 1.5718 16.0097 144.9576 0.00029424 -85.231 0.29594
4.4 0.98807 5.4966e-005 3.8183 0.011988 5.7598e-005 0.0011588 0.22895 0.00065927 0.2296 0.21174 0 0.032497 0.0389 0 1.2086 0.39298 0.11757 0.014992 7.6736 0.093524 0.00011726 0.79659 0.0073814 0.0082327 0.0014863 0.98564 0.99084 3.2185e-006 1.2874e-005 0.14902 0.77235 0.83288 0.0014491 0.88733 0.45996 0.0019502 0.42257 1.5758 1.5733 16.0098 144.9576 0.00029362 -85.2341 0.29694
4.401 0.98807 5.4966e-005 3.8183 0.011988 5.7611e-005 0.0011588 0.22895 0.00065927 0.22961 0.21175 0 0.032497 0.0389 0 1.2087 0.39303 0.11759 0.014993 7.6753 0.093534 0.00011727 0.79658 0.007382 0.0082334 0.0014855 0.98565 0.99085 3.2168e-006 1.2867e-005 0.14903 0.77301 0.83328 0.0014487 0.88801 0.46014 0.0019497 0.42258 1.5773 1.5747 16.0098 144.9577 0.00029301 -85.2372 0.29794
4.402 0.98807 5.4965e-005 3.8183 0.011988 5.7624e-005 0.0011588 0.22896 0.00065927 0.22961 0.21175 0 0.032497 0.0389 0 1.2088 0.39307 0.1176 0.014995 7.677 0.093544 0.00011729 0.79657 0.0073827 0.0082341 0.0014848 0.98566 0.99086 3.2151e-006 1.286e-005 0.14903 0.77366 0.83368 0.0014483 0.8887 0.46033 0.0019492 0.42259 1.5787 1.5762 16.0098 144.9577 0.00029241 -85.2402 0.29894
4.403 0.98807 5.4965e-005 3.8183 0.011988 5.7637e-005 0.0011588 0.22896 0.00065927 0.22962 0.21176 0 0.032496 0.0389 0 1.2089 0.39312 0.11762 0.014997 7.6787 0.093554 0.0001173 0.79656 0.0073834 0.0082348 0.0014841 0.98567 0.99086 3.2134e-006 1.2854e-005 0.14904 0.77432 0.83408 0.0014479 0.88937 0.46051 0.0019487 0.4226 1.5801 1.5776 16.0098 144.9577 0.0002918 -85.2432 0.29994
4.404 0.98807 5.4965e-005 3.8183 0.011988 5.765e-005 0.0011588 0.22897 0.00065927 0.22962 0.21176 0 0.032496 0.0389 0 1.209 0.39317 0.11764 0.014998 7.6804 0.093564 0.00011731 0.79655 0.0073841 0.0082356 0.0014833 0.98568 0.99087 3.2117e-006 1.2847e-005 0.14904 0.77497 0.83447 0.0014476 0.89004 0.4607 0.0019482 0.42261 1.5816 1.579 16.0098 144.9577 0.0002912 -85.2462 0.30094
4.405 0.98807 5.4965e-005 3.8183 0.011988 5.7663e-005 0.0011588 0.22897 0.00065927 0.22963 0.21177 0 0.032496 0.0389 0 1.2091 0.39321 0.11765 0.015 7.6821 0.093574 0.00011733 0.79654 0.0073847 0.0082363 0.0014826 0.98569 0.99088 3.21e-006 1.284e-005 0.14905 0.77562 0.83486 0.0014472 0.89071 0.46089 0.0019477 0.42262 1.583 1.5804 16.0098 144.9577 0.0002906 -85.2492 0.30194
4.406 0.98807 5.4965e-005 3.8183 0.011988 5.7676e-005 0.0011588 0.22898 0.00065927 0.22963 0.21177 0 0.032496 0.0389 0 1.2092 0.39326 0.11767 0.015001 7.6838 0.093583 0.00011734 0.79653 0.0073854 0.008237 0.0014819 0.9857 0.99088 3.2083e-006 1.2833e-005 0.14905 0.77626 0.83526 0.0014468 0.89138 0.46107 0.0019473 0.42264 1.5844 1.5819 16.0099 144.9577 0.00029 -85.2522 0.30294
4.407 0.98807 5.4965e-005 3.8183 0.011987 5.7689e-005 0.0011588 0.22898 0.00065927 0.22964 0.21178 0 0.032496 0.0389 0 1.2093 0.3933 0.11768 0.015003 7.6855 0.093593 0.00011735 0.79652 0.0073861 0.0082377 0.0014812 0.9857 0.99089 3.2066e-006 1.2827e-005 0.14906 0.77691 0.83565 0.0014464 0.89204 0.46126 0.0019468 0.42265 1.5858 1.5833 16.0099 144.9578 0.00028941 -85.2551 0.30394
4.408 0.98807 5.4965e-005 3.8183 0.011987 5.7702e-005 0.0011588 0.22899 0.00065927 0.22964 0.21178 0 0.032495 0.0389 0 1.2094 0.39335 0.1177 0.015005 7.6872 0.093603 0.00011737 0.79651 0.0073868 0.0082385 0.0014804 0.98571 0.9909 3.205e-006 1.282e-005 0.14907 0.77755 0.83603 0.0014461 0.89269 0.46144 0.0019463 0.42266 1.5872 1.5847 16.0099 144.9578 0.00028882 -85.258 0.30494
4.409 0.98807 5.4965e-005 3.8183 0.011987 5.7715e-005 0.0011588 0.22899 0.00065927 0.22964 0.21178 0 0.032495 0.0389 0 1.2095 0.3934 0.11771 0.015006 7.6889 0.093613 0.00011738 0.7965 0.0073874 0.0082392 0.0014797 0.98572 0.9909 3.2033e-006 1.2813e-005 0.14907 0.77819 0.83642 0.0014457 0.89335 0.46163 0.0019458 0.42267 1.5886 1.5861 16.0099 144.9578 0.00028823 -85.2609 0.30594
4.41 0.98807 5.4965e-005 3.8183 0.011987 5.7728e-005 0.0011588 0.22899 0.00065927 0.22965 0.21179 0 0.032495 0.0389 0 1.2096 0.39344 0.11773 0.015008 7.6906 0.093623 0.0001174 0.79649 0.0073881 0.0082399 0.001479 0.98573 0.99091 3.2017e-006 1.2807e-005 0.14908 0.77883 0.8368 0.0014453 0.89399 0.46181 0.0019453 0.42268 1.59 1.5875 16.0099 144.9578 0.00028764 -85.2637 0.30694
4.411 0.98807 5.4965e-005 3.8183 0.011987 5.7741e-005 0.0011588 0.229 0.00065927 0.22965 0.21179 0 0.032495 0.0389 0 1.2097 0.39349 0.11775 0.015009 7.6923 0.093633 0.00011741 0.79648 0.0073888 0.0082406 0.0014783 0.98574 0.99092 3.2001e-006 1.28e-005 0.14908 0.77947 0.83719 0.001445 0.89464 0.462 0.0019449 0.42269 1.5914 1.5889 16.0099 144.9578 0.00028706 -85.2666 0.30794
4.412 0.98807 5.4965e-005 3.8183 0.011987 5.7754e-005 0.0011588 0.229 0.00065927 0.22966 0.2118 0 0.032494 0.0389 0 1.2098 0.39354 0.11776 0.015011 7.6939 0.093643 0.00011742 0.79647 0.0073894 0.0082413 0.0014776 0.98575 0.99092 3.1985e-006 1.2794e-005 0.14909 0.78011 0.83757 0.0014446 0.89528 0.46218 0.0019444 0.4227 1.5928 1.5903 16.01 144.9578 0.00028648 -85.2694 0.30894
4.413 0.98807 5.4965e-005 3.8183 0.011987 5.7767e-005 0.0011588 0.22901 0.00065927 0.22966 0.2118 0 0.032494 0.0389 0 1.2099 0.39358 0.11778 0.015013 7.6956 0.093653 0.00011744 0.79646 0.0073901 0.0082421 0.0014769 0.98576 0.99093 3.1969e-006 1.2788e-005 0.14909 0.78074 0.83795 0.0014443 0.89592 0.46237 0.0019439 0.42271 1.5942 1.5917 16.01 144.9579 0.0002859 -85.2722 0.30994
4.414 0.98807 5.4965e-005 3.8183 0.011987 5.778e-005 0.0011588 0.22901 0.00065927 0.22967 0.21181 0 0.032494 0.0389 0 1.21 0.39363 0.11779 0.015014 7.6973 0.093663 0.00011745 0.79645 0.0073908 0.0082428 0.0014762 0.98577 0.99093 3.1953e-006 1.2781e-005 0.1491 0.78137 0.83832 0.0014439 0.89655 0.46255 0.0019435 0.42272 1.5956 1.5931 16.01 144.9579 0.00028533 -85.275 0.31094
4.415 0.98807 5.4965e-005 3.8183 0.011987 5.7793e-005 0.0011588 0.22902 0.00065927 0.22967 0.21181 0 0.032494 0.0389 0 1.2101 0.39368 0.11781 0.015016 7.699 0.093673 0.00011747 0.79644 0.0073914 0.0082435 0.0014755 0.98578 0.99094 3.1938e-006 1.2775e-005 0.1491 0.782 0.8387 0.0014436 0.89718 0.46274 0.001943 0.42274 1.5969 1.5945 16.01 144.9579 0.00028476 -85.2778 0.31194
4.416 0.98807 5.4964e-005 3.8183 0.011987 5.7806e-005 0.0011588 0.22902 0.00065927 0.22968 0.21182 0 0.032493 0.0389 0 1.2102 0.39372 0.11783 0.015017 7.7007 0.093683 0.00011748 0.79643 0.0073921 0.0082442 0.0014749 0.98579 0.99095 3.1922e-006 1.2769e-005 0.14911 0.78263 0.83907 0.0014432 0.89781 0.46292 0.0019426 0.42275 1.5983 1.5959 16.01 144.9579 0.00028419 -85.2805 0.31294
4.417 0.98807 5.4964e-005 3.8183 0.011987 5.7819e-005 0.0011588 0.22903 0.00065927 0.22968 0.21182 0 0.032493 0.0389 0 1.2103 0.39377 0.11784 0.015019 7.7024 0.093692 0.00011749 0.79643 0.0073928 0.008245 0.0014742 0.9858 0.99095 3.1907e-006 1.2763e-005 0.14911 0.78326 0.83944 0.0014429 0.89843 0.46311 0.0019421 0.42276 1.5997 1.5973 16.01 144.9579 0.00028362 -85.2832 0.31394
4.418 0.98807 5.4964e-005 3.8183 0.011987 5.7832e-005 0.0011589 0.22903 0.00065927 0.22969 0.21182 0 0.032493 0.0389 0 1.2104 0.39382 0.11786 0.015021 7.7041 0.093702 0.00011751 0.79642 0.0073935 0.0082457 0.0014735 0.98581 0.99096 3.1892e-006 1.2757e-005 0.14912 0.78388 0.83981 0.0014425 0.89905 0.46329 0.0019417 0.42277 1.6011 1.5986 16.01 144.9579 0.00028305 -85.2859 0.31494
4.419 0.98807 5.4964e-005 3.8183 0.011987 5.7845e-005 0.0011589 0.22904 0.00065927 0.22969 0.21183 0 0.032493 0.0389 0 1.2105 0.39386 0.11787 0.015022 7.7058 0.093712 0.00011752 0.79641 0.0073941 0.0082464 0.0014729 0.98581 0.99096 3.1877e-006 1.2751e-005 0.14912 0.7845 0.84018 0.0014422 0.89966 0.46348 0.0019412 0.42278 1.6024 1.6 16.0101 144.958 0.00028249 -85.2886 0.31594
4.42 0.98807 5.4964e-005 3.8183 0.011987 5.7858e-005 0.0011589 0.22904 0.00065927 0.2297 0.21183 0 0.032492 0.0389 0 1.2106 0.39391 0.11789 0.015024 7.7075 0.093722 0.00011754 0.7964 0.0073948 0.0082471 0.0014722 0.98582 0.99097 3.1862e-006 1.2745e-005 0.14913 0.78512 0.84055 0.0014419 0.90027 0.46366 0.0019408 0.42279 1.6038 1.6014 16.0101 144.958 0.00028193 -85.2913 0.31694
4.421 0.98807 5.4964e-005 3.8183 0.011987 5.7871e-005 0.0011589 0.22905 0.00065927 0.2297 0.21184 0 0.032492 0.0389 0 1.2107 0.39396 0.11791 0.015025 7.7092 0.093732 0.00011755 0.79639 0.0073955 0.0082478 0.0014716 0.98583 0.99097 3.1847e-006 1.2739e-005 0.14914 0.78574 0.84091 0.0014415 0.90088 0.46385 0.0019404 0.4228 1.6052 1.6028 16.0101 144.958 0.00028137 -85.2939 0.31794
4.422 0.98807 5.4964e-005 3.8183 0.011987 5.7884e-005 0.0011589 0.22905 0.00065927 0.22971 0.21184 0 0.032492 0.0389 0 1.2108 0.394 0.11792 0.015027 7.7109 0.093742 0.00011756 0.79638 0.0073961 0.0082486 0.0014709 0.98584 0.99098 3.1832e-006 1.2733e-005 0.14914 0.78636 0.84127 0.0014412 0.90148 0.46403 0.0019399 0.42281 1.6065 1.6041 16.0101 144.958 0.00028082 -85.2965 0.31894
4.423 0.98807 5.4964e-005 3.8183 0.011987 5.7897e-005 0.0011589 0.22905 0.00065927 0.22971 0.21185 0 0.032492 0.0389 0 1.2109 0.39405 0.11794 0.015029 7.7126 0.093752 0.00011758 0.79637 0.0073968 0.0082493 0.0014703 0.98585 0.99099 3.1817e-006 1.2727e-005 0.14915 0.78697 0.84163 0.0014409 0.90208 0.46421 0.0019395 0.42283 1.6079 1.6055 16.0101 144.958 0.00028027 -85.2991 0.31994
4.424 0.98807 5.4964e-005 3.8183 0.011987 5.791e-005 0.0011589 0.22906 0.00065927 0.22971 0.21185 0 0.032492 0.0389 0 1.211 0.3941 0.11795 0.01503 7.7143 0.093762 0.00011759 0.79636 0.0073975 0.00825 0.0014697 0.98586 0.99099 3.1803e-006 1.2721e-005 0.14915 0.78758 0.84199 0.0014406 0.90268 0.4644 0.0019391 0.42284 1.6092 1.6068 16.0101 144.9581 0.00027972 -85.3017 0.32094
4.425 0.98807 5.4964e-005 3.8183 0.011987 5.7923e-005 0.0011589 0.22906 0.00065927 0.22972 0.21186 0 0.032491 0.0389 0 1.2111 0.39414 0.11797 0.015032 7.716 0.093772 0.0001176 0.79635 0.0073982 0.0082507 0.001469 0.98586 0.991 3.1788e-006 1.2715e-005 0.14916 0.78819 0.84235 0.0014402 0.90327 0.46458 0.0019386 0.42285 1.6105 1.6082 16.0101 144.9581 0.00027917 -85.3043 0.32194
4.426 0.98807 5.4964e-005 3.8183 0.011987 5.7936e-005 0.0011589 0.22907 0.00065927 0.22972 0.21186 0 0.032491 0.0389 0 1.2112 0.39419 0.11798 0.015033 7.7177 0.093781 0.00011762 0.79634 0.0073988 0.0082515 0.0014684 0.98587 0.991 3.1774e-006 1.271e-005 0.14916 0.7888 0.84271 0.0014399 0.90386 0.46477 0.0019382 0.42286 1.6119 1.6095 16.0102 144.9581 0.00027863 -85.3068 0.32294
4.427 0.98807 5.4964e-005 3.8183 0.011987 5.7949e-005 0.0011589 0.22907 0.00065927 0.22973 0.21186 0 0.032491 0.0389 0 1.2113 0.39424 0.118 0.015035 7.7194 0.093791 0.00011763 0.79633 0.0073995 0.0082522 0.0014678 0.98588 0.99101 3.176e-006 1.2704e-005 0.14917 0.78941 0.84306 0.0014396 0.90445 0.46495 0.0019378 0.42287 1.6132 1.6109 16.0102 144.9581 0.00027808 -85.3094 0.32394
4.428 0.98807 5.4964e-005 3.8183 0.011987 5.7962e-005 0.0011589 0.22908 0.00065927 0.22973 0.21187 0 0.032491 0.0389 0 1.2114 0.39428 0.11802 0.015037 7.7211 0.093801 0.00011765 0.79632 0.0074002 0.0082529 0.0014672 0.98589 0.99101 3.1746e-006 1.2698e-005 0.14917 0.79001 0.84341 0.0014393 0.90503 0.46514 0.0019374 0.42288 1.6146 1.6122 16.0102 144.9581 0.00027754 -85.3119 0.32494
4.429 0.98807 5.4964e-005 3.8183 0.011987 5.7975e-005 0.0011589 0.22908 0.00065927 0.22974 0.21187 0 0.03249 0.0389 0 1.2115 0.39433 0.11803 0.015038 7.7228 0.093811 0.00011766 0.79631 0.0074008 0.0082536 0.0014666 0.9859 0.99102 3.1732e-006 1.2693e-005 0.14918 0.79062 0.84376 0.001439 0.90561 0.46532 0.001937 0.42289 1.6159 1.6136 16.0102 144.9581 0.00027701 -85.3144 0.32594
4.43 0.98807 5.4963e-005 3.8183 0.011987 5.7988e-005 0.0011589 0.22909 0.00065927 0.22974 0.21188 0 0.03249 0.0389 0 1.2116 0.39438 0.11805 0.01504 7.7245 0.093821 0.00011767 0.7963 0.0074015 0.0082543 0.001466 0.98591 0.99102 3.1718e-006 1.2687e-005 0.14918 0.79122 0.84411 0.0014386 0.90619 0.4655 0.0019366 0.42291 1.6172 1.6149 16.0102 144.9582 0.00027647 -85.3169 0.32694
4.431 0.98807 5.4963e-005 3.8183 0.011987 5.8001e-005 0.0011589 0.22909 0.00065927 0.22975 0.21188 0 0.03249 0.0389 0 1.2117 0.39442 0.11806 0.015041 7.7262 0.093831 0.00011769 0.79629 0.0074022 0.0082551 0.0014654 0.98591 0.99103 3.1704e-006 1.2682e-005 0.14919 0.79182 0.84446 0.0014383 0.90676 0.46569 0.0019362 0.42292 1.6185 1.6162 16.0102 144.9582 0.00027594 -85.3193 0.32794
4.432 0.98807 5.4963e-005 3.8183 0.011987 5.8014e-005 0.0011589 0.2291 0.00065927 0.22975 0.21189 0 0.03249 0.0389 0 1.2118 0.39447 0.11808 0.015043 7.7279 0.093841 0.0001177 0.79628 0.0074028 0.0082558 0.0014648 0.98592 0.99103 3.169e-006 1.2676e-005 0.14919 0.79242 0.84481 0.001438 0.90733 0.46587 0.0019358 0.42293 1.6199 1.6175 16.0102 144.9582 0.00027541 -85.3218 0.32894
4.433 0.98807 5.4963e-005 3.8183 0.011987 5.8027e-005 0.0011589 0.2291 0.00065927 0.22976 0.21189 0 0.032489 0.0389 0 1.2118 0.39452 0.1181 0.015045 7.7296 0.093851 0.00011772 0.79627 0.0074035 0.0082565 0.0014642 0.98593 0.99104 3.1677e-006 1.2671e-005 0.1492 0.79301 0.84515 0.0014377 0.90789 0.46606 0.0019354 0.42294 1.6212 1.6189 16.0102 144.9582 0.00027488 -85.3242 0.32994
4.434 0.98807 5.4963e-005 3.8183 0.011987 5.804e-005 0.0011589 0.22911 0.00065927 0.22976 0.21189 0 0.032489 0.0389 0 1.2119 0.39456 0.11811 0.015046 7.7313 0.093861 0.00011773 0.79626 0.0074042 0.0082572 0.0014636 0.98594 0.99104 3.1663e-006 1.2665e-005 0.1492 0.7936 0.84549 0.0014374 0.90845 0.46624 0.001935 0.42295 1.6225 1.6202 16.0103 144.9582 0.00027435 -85.3266 0.33094
4.435 0.98807 5.4963e-005 3.8183 0.011987 5.8053e-005 0.0011589 0.22911 0.00065927 0.22976 0.2119 0 0.032489 0.0389 0 1.212 0.39461 0.11813 0.015048 7.733 0.09387 0.00011774 0.79625 0.0074049 0.0082579 0.001463 0.98594 0.99105 3.165e-006 1.266e-005 0.14921 0.7942 0.84583 0.0014371 0.90901 0.46642 0.0019346 0.42296 1.6238 1.6215 16.0103 144.9583 0.00027383 -85.329 0.33194
4.436 0.98807 5.4963e-005 3.8183 0.011987 5.8066e-005 0.0011589 0.22911 0.00065927 0.22977 0.2119 0 0.032489 0.0389 0 1.2121 0.39466 0.11814 0.015049 7.7347 0.09388 0.00011776 0.79624 0.0074055 0.0082587 0.0014624 0.98595 0.99106 3.1637e-006 1.2655e-005 0.14922 0.79479 0.84617 0.0014368 0.90957 0.46661 0.0019342 0.42298 1.6251 1.6228 16.0103 144.9583 0.00027331 -85.3313 0.33294
4.437 0.98807 5.4963e-005 3.8183 0.011987 5.8079e-005 0.0011589 0.22912 0.00065927 0.22977 0.21191 0 0.032489 0.0389 0 1.2122 0.3947 0.11816 0.015051 7.7364 0.09389 0.00011777 0.79623 0.0074062 0.0082594 0.0014619 0.98596 0.99106 3.1623e-006 1.2649e-005 0.14922 0.79538 0.84651 0.0014365 0.91012 0.46679 0.0019338 0.42299 1.6264 1.6241 16.0103 144.9583 0.00027279 -85.3337 0.33394
4.438 0.98807 5.4963e-005 3.8183 0.011987 5.8092e-005 0.0011589 0.22912 0.00065927 0.22978 0.21191 0 0.032488 0.0389 0 1.2123 0.39475 0.11817 0.015053 7.7381 0.0939 0.00011778 0.79622 0.0074069 0.0082601 0.0014613 0.98597 0.99107 3.161e-006 1.2644e-005 0.14923 0.79596 0.84685 0.0014362 0.91066 0.46698 0.0019334 0.423 1.6277 1.6254 16.0103 144.9583 0.00027228 -85.336 0.33494
4.439 0.98807 5.4963e-005 3.8183 0.011987 5.8105e-005 0.0011589 0.22913 0.00065927 0.22978 0.21192 0 0.032488 0.0389 0 1.2124 0.3948 0.11819 0.015054 7.7398 0.09391 0.0001178 0.79621 0.0074075 0.0082608 0.0014607 0.98597 0.99107 3.1597e-006 1.2639e-005 0.14923 0.79655 0.84718 0.0014359 0.91121 0.46716 0.001933 0.42301 1.629 1.6267 16.0103 144.9583 0.00027176 -85.3383 0.33594
4.44 0.98807 5.4963e-005 3.8183 0.011987 5.8118e-005 0.0011589 0.22913 0.00065927 0.22979 0.21192 0 0.032488 0.0389 0 1.2125 0.39484 0.11821 0.015056 7.7415 0.09392 0.00011781 0.7962 0.0074082 0.0082615 0.0014602 0.98598 0.99107 3.1584e-006 1.2634e-005 0.14924 0.79713 0.84751 0.0014357 0.91175 0.46734 0.0019327 0.42302 1.6303 1.628 16.0103 144.9583 0.00027125 -85.3406 0.33694
4.441 0.98807 5.4963e-005 3.8183 0.011987 5.8131e-005 0.0011589 0.22914 0.00065927 0.22979 0.21193 0 0.032488 0.0389 0 1.2126 0.39489 0.11822 0.015057 7.7433 0.09393 0.00011783 0.79619 0.0074089 0.0082623 0.0014596 0.98599 0.99108 3.1572e-006 1.2629e-005 0.14924 0.79771 0.84785 0.0014354 0.91229 0.46753 0.0019323 0.42303 1.6316 1.6293 16.0103 144.9584 0.00027074 -85.3429 0.33794
4.442 0.98807 5.4963e-005 3.8183 0.011987 5.8144e-005 0.0011589 0.22914 0.00065927 0.2298 0.21193 0 0.032487 0.0389 0 1.2127 0.39494 0.11824 0.015059 7.745 0.09394 0.00011784 0.79618 0.0074095 0.008263 0.001459 0.986 0.99108 3.1559e-006 1.2624e-005 0.14925 0.79829 0.84818 0.0014351 0.91282 0.46771 0.0019319 0.42305 1.6328 1.6306 16.0103 144.9584 0.00027023 -85.3452 0.33894
4.443 0.98807 5.4963e-005 3.8183 0.011987 5.8157e-005 0.0011589 0.22915 0.00065927 0.2298 0.21193 0 0.032487 0.0389 0 1.2128 0.39498 0.11825 0.015061 7.7467 0.093949 0.00011785 0.79617 0.0074102 0.0082637 0.0014585 0.986 0.99109 3.1546e-006 1.2619e-005 0.14925 0.79887 0.8485 0.0014348 0.91336 0.46789 0.0019315 0.42306 1.6341 1.6319 16.0104 144.9584 0.00026973 -85.3475 0.33994
4.444 0.98807 5.4962e-005 3.8183 0.011987 5.817e-005 0.0011589 0.22915 0.00065927 0.22981 0.21194 0 0.032487 0.0389 0 1.2129 0.39503 0.11827 0.015062 7.7484 0.093959 0.00011787 0.79616 0.0074109 0.0082644 0.001458 0.98601 0.99109 3.1534e-006 1.2614e-005 0.14926 0.79944 0.84883 0.0014345 0.91388 0.46808 0.0019312 0.42307 1.6354 1.6332 16.0104 144.9584 0.00026923 -85.3497 0.34094
4.445 0.98807 5.4962e-005 3.8183 0.011987 5.8183e-005 0.0011589 0.22916 0.00065927 0.22981 0.21194 0 0.032487 0.0389 0 1.213 0.39508 0.11829 0.015064 7.7501 0.093969 0.00011788 0.79615 0.0074115 0.0082651 0.0014574 0.98602 0.9911 3.1522e-006 1.2609e-005 0.14926 0.80002 0.84916 0.0014342 0.91441 0.46826 0.0019308 0.42308 1.6367 1.6345 16.0104 144.9584 0.00026873 -85.3519 0.34194
4.446 0.98807 5.4962e-005 3.8183 0.011987 5.8196e-005 0.0011589 0.22916 0.00065927 0.22981 0.21195 0 0.032486 0.0389 0 1.2131 0.39512 0.1183 0.015065 7.7518 0.093979 0.0001179 0.79614 0.0074122 0.0082659 0.0014569 0.98602 0.9911 3.1509e-006 1.2604e-005 0.14927 0.80059 0.84948 0.001434 0.91493 0.46845 0.0019305 0.42309 1.6379 1.6357 16.0104 144.9584 0.00026823 -85.3541 0.34294
4.447 0.98807 5.4962e-005 3.8183 0.011987 5.8209e-005 0.0011589 0.22916 0.00065927 0.22982 0.21195 0 0.032486 0.0389 0 1.2132 0.39517 0.11832 0.015067 7.7535 0.093989 0.00011791 0.79613 0.0074129 0.0082666 0.0014564 0.98603 0.99111 3.1497e-006 1.2599e-005 0.14927 0.80116 0.8498 0.0014337 0.91545 0.46863 0.0019301 0.42311 1.6392 1.637 16.0104 144.9585 0.00026773 -85.3563 0.34394
4.448 0.98807 5.4962e-005 3.8183 0.011987 5.8222e-005 0.0011589 0.22917 0.00065927 0.22982 0.21196 0 0.032486 0.0389 0 1.2133 0.39522 0.11833 0.015068 7.7552 0.093999 0.00011792 0.79612 0.0074135 0.0082673 0.0014558 0.98604 0.99111 3.1485e-006 1.2594e-005 0.14928 0.80173 0.85012 0.0014334 0.91597 0.46881 0.0019297 0.42312 1.6405 1.6383 16.0104 144.9585 0.00026724 -85.3585 0.34494
4.449 0.98807 5.4962e-005 3.8183 0.011987 5.8235e-005 0.0011589 0.22917 0.00065927 0.22983 0.21196 0 0.032486 0.0389 0 1.2134 0.39526 0.11835 0.01507 7.7569 0.094009 0.00011794 0.79611 0.0074142 0.008268 0.0014553 0.98605 0.99112 3.1473e-006 1.2589e-005 0.14928 0.80229 0.85044 0.0014331 0.91648 0.469 0.0019294 0.42313 1.6417 1.6396 16.0104 144.9585 0.00026675 -85.3606 0.34594
4.45 0.98807 5.4962e-005 3.8183 0.011987 5.8248e-005 0.0011589 0.22918 0.00065927 0.22983 0.21196 0 0.032486 0.0389 0 1.2135 0.39531 0.11837 0.015072 7.7586 0.094019 0.00011795 0.7961 0.0074149 0.0082687 0.0014548 0.98605 0.99112 3.1461e-006 1.2584e-005 0.14929 0.80286 0.85076 0.0014329 0.91699 0.46918 0.001929 0.42314 1.643 1.6408 16.0104 144.9585 0.00026626 -85.3628 0.34694
4.451 0.98807 5.4962e-005 3.8183 0.011987 5.8261e-005 0.0011589 0.22918 0.00065927 0.22984 0.21197 0 0.032485 0.0389 0 1.2136 0.39536 0.11838 0.015073 7.7603 0.094028 0.00011796 0.79609 0.0074156 0.0082695 0.0014543 0.98606 0.99113 3.1449e-006 1.258e-005 0.1493 0.80342 0.85108 0.0014326 0.9175 0.46936 0.0019287 0.42315 1.6442 1.6421 16.0104 144.9585 0.00026577 -85.3649 0.34794
4.452 0.98807 5.4962e-005 3.8183 0.011987 5.8274e-005 0.0011589 0.22919 0.00065927 0.22984 0.21197 0 0.032485 0.0389 0 1.2137 0.3954 0.1184 0.015075 7.762 0.094038 0.00011798 0.79608 0.0074162 0.0082702 0.0014537 0.98607 0.99113 3.1437e-006 1.2575e-005 0.1493 0.80398 0.85139 0.0014323 0.918 0.46954 0.0019283 0.42317 1.6455 1.6433 16.0104 144.9586 0.00026529 -85.367 0.34894
4.453 0.98807 5.4962e-005 3.8183 0.011987 5.8287e-005 0.0011589 0.22919 0.00065927 0.22985 0.21198 0 0.032485 0.0389 0 1.2138 0.39545 0.11841 0.015076 7.7637 0.094048 0.00011799 0.79607 0.0074169 0.0082709 0.0014532 0.98607 0.99114 3.1426e-006 1.257e-005 0.14931 0.80454 0.85171 0.0014321 0.9185 0.46973 0.001928 0.42318 1.6467 1.6446 16.0104 144.9586 0.0002648 -85.3691 0.34994
4.454 0.98807 5.4962e-005 3.8183 0.011987 5.83e-005 0.0011589 0.2292 0.00065927 0.22985 0.21198 0 0.032485 0.0389 0 1.2139 0.3955 0.11843 0.015078 7.7655 0.094058 0.00011801 0.79606 0.0074176 0.0082716 0.0014527 0.98608 0.99114 3.1414e-006 1.2566e-005 0.14931 0.8051 0.85202 0.0014318 0.919 0.46991 0.0019277 0.42319 1.648 1.6458 16.0104 144.9586 0.00026432 -85.3712 0.35094
4.455 0.98807 5.4962e-005 3.8183 0.011987 5.8313e-005 0.0011589 0.2292 0.00065927 0.22986 0.21199 0 0.032484 0.0389 0 1.214 0.39554 0.11844 0.01508 7.7672 0.094068 0.00011802 0.79605 0.0074182 0.0082723 0.0014523 0.98609 0.99114 3.1403e-006 1.2561e-005 0.14932 0.80566 0.85233 0.0014316 0.91949 0.47009 0.0019273 0.4232 1.6492 1.6471 16.0105 144.9586 0.00026384 -85.3733 0.35194
4.456 0.98807 5.4962e-005 3.8183 0.011987 5.8326e-005 0.0011589 0.22921 0.00065927 0.22986 0.21199 0 0.032484 0.0389 0 1.2141 0.39559 0.11846 0.015081 7.7689 0.094078 0.00011803 0.79604 0.0074189 0.0082731 0.0014518 0.98609 0.99115 3.1391e-006 1.2557e-005 0.14932 0.80621 0.85264 0.0014313 0.91998 0.47028 0.001927 0.42321 1.6504 1.6483 16.0105 144.9586 0.00026337 -85.3753 0.35294
4.457 0.98807 5.4962e-005 3.8183 0.011987 5.8339e-005 0.001159 0.22921 0.00065927 0.22986 0.21199 0 0.032484 0.0389 0 1.2142 0.39564 0.11848 0.015083 7.7706 0.094088 0.00011805 0.79603 0.0074196 0.0082738 0.0014513 0.9861 0.99115 3.138e-006 1.2552e-005 0.14933 0.80676 0.85295 0.0014311 0.92047 0.47046 0.0019266 0.42323 1.6517 1.6496 16.0105 144.9586 0.00026289 -85.3773 0.35394
4.458 0.98807 5.4961e-005 3.8183 0.011987 5.8352e-005 0.001159 0.22921 0.00065927 0.22987 0.212 0 0.032484 0.0389 0 1.2143 0.39568 0.11849 0.015084 7.7723 0.094097 0.00011806 0.79602 0.0074202 0.0082745 0.0014508 0.98611 0.99116 3.1369e-006 1.2548e-005 0.14933 0.80731 0.85325 0.0014308 0.92096 0.47064 0.0019263 0.42324 1.6529 1.6508 16.0105 144.9587 0.00026242 -85.3794 0.35494
4.459 0.98807 5.4961e-005 3.8183 0.011987 5.8365e-005 0.001159 0.22922 0.00065927 0.22987 0.212 0 0.032484 0.0389 0 1.2144 0.39573 0.11851 0.015086 7.774 0.094107 0.00011808 0.79601 0.0074209 0.0082752 0.0014503 0.98611 0.99116 3.1358e-006 1.2543e-005 0.14934 0.80786 0.85356 0.0014305 0.92144 0.47083 0.001926 0.42325 1.6541 1.652 16.0105 144.9587 0.00026195 -85.3814 0.35594
4.46 0.98807 5.4961e-005 3.8183 0.011987 5.8378e-005 0.001159 0.22922 0.00065927 0.22988 0.21201 0 0.032483 0.0389 0 1.2145 0.39578 0.11852 0.015088 7.7757 0.094117 0.00011809 0.796 0.0074216 0.0082759 0.0014498 0.98612 0.99117 3.1347e-006 1.2539e-005 0.14934 0.80841 0.85386 0.0014303 0.92192 0.47101 0.0019257 0.42326 1.6554 1.6533 16.0105 144.9587 0.00026148 -85.3834 0.35694
4.461 0.98807 5.4961e-005 3.8183 0.011987 5.8391e-005 0.001159 0.22923 0.00065927 0.22988 0.21201 0 0.032483 0.0389 0 1.2146 0.39582 0.11854 0.015089 7.7774 0.094127 0.0001181 0.79599 0.0074222 0.0082767 0.0014493 0.98612 0.99117 3.1336e-006 1.2534e-005 0.14935 0.80896 0.85416 0.00143 0.92239 0.47119 0.0019253 0.42327 1.6566 1.6545 16.0105 144.9587 0.00026102 -85.3853 0.35794
4.462 0.98807 5.4961e-005 3.8183 0.011987 5.8404e-005 0.001159 0.22923 0.00065927 0.22989 0.21202 0 0.032483 0.0389 0 1.2147 0.39587 0.11856 0.015091 7.7791 0.094137 0.00011812 0.79598 0.0074229 0.0082774 0.0014488 0.98613 0.99117 3.1325e-006 1.253e-005 0.14935 0.8095 0.85447 0.0014298 0.92287 0.47137 0.001925 0.42329 1.6578 1.6557 16.0105 144.9587 0.00026055 -85.3873 0.35894
4.463 0.98807 5.4961e-005 3.8183 0.011987 5.8417e-005 0.001159 0.22924 0.00065927 0.22989 0.21202 0 0.032483 0.0389 0 1.2148 0.39592 0.11857 0.015092 7.7809 0.094147 0.00011813 0.79597 0.0074236 0.0082781 0.0014484 0.98614 0.99118 3.1314e-006 1.2526e-005 0.14936 0.81004 0.85477 0.0014296 0.92334 0.47156 0.0019247 0.4233 1.659 1.6569 16.0105 144.9588 0.00026009 -85.3893 0.35994
4.464 0.98807 5.4961e-005 3.8183 0.011987 5.843e-005 0.001159 0.22924 0.00065927 0.2299 0.21202 0 0.032482 0.0389 0 1.2149 0.39596 0.11859 0.015094 7.7826 0.094157 0.00011814 0.79596 0.0074242 0.0082788 0.0014479 0.98614 0.99118 3.1303e-006 1.2521e-005 0.14936 0.81059 0.85506 0.0014293 0.9238 0.47174 0.0019244 0.42331 1.6602 1.6581 16.0105 144.9588 0.00025963 -85.3912 0.36094
4.465 0.98807 5.4961e-005 3.8183 0.011987 5.8443e-005 0.001159 0.22925 0.00065927 0.2299 0.21203 0 0.032482 0.0389 0 1.215 0.39601 0.1186 0.015096 7.7843 0.094166 0.00011816 0.79595 0.0074249 0.0082795 0.0014474 0.98615 0.99119 3.1293e-006 1.2517e-005 0.14937 0.81112 0.85536 0.0014291 0.92427 0.47192 0.0019241 0.42332 1.6614 1.6594 16.0105 144.9588 0.00025917 -85.3931 0.36194
4.466 0.98807 5.4961e-005 3.8183 0.011987 5.8456e-005 0.001159 0.22925 0.00065927 0.2299 0.21203 0 0.032482 0.0389 0 1.2151 0.39606 0.11862 0.015097 7.786 0.094176 0.00011817 0.79594 0.0074256 0.0082803 0.001447 0.98615 0.99119 3.1282e-006 1.2513e-005 0.14938 0.81166 0.85566 0.0014288 0.92473 0.4721 0.0019238 0.42334 1.6626 1.6606 16.0105 144.9588 0.00025872 -85.395 0.36294
4.467 0.98807 5.4961e-005 3.8183 0.011987 5.8469e-005 0.001159 0.22925 0.00065927 0.22991 0.21204 0 0.032482 0.0389 0 1.2152 0.3961 0.11864 0.015099 7.7877 0.094186 0.00011819 0.79593 0.0074262 0.008281 0.0014465 0.98616 0.99119 3.1271e-006 1.2509e-005 0.14938 0.8122 0.85595 0.0014286 0.92519 0.47229 0.0019234 0.42335 1.6638 1.6618 16.0105 144.9588 0.00025826 -85.3969 0.36394
4.468 0.98807 5.4961e-005 3.8183 0.011987 5.8482e-005 0.001159 0.22926 0.00065927 0.22991 0.21204 0 0.032482 0.0389 0 1.2153 0.39615 0.11865 0.0151 7.7894 0.094196 0.0001182 0.79592 0.0074269 0.0082817 0.0014461 0.98617 0.9912 3.1261e-006 1.2504e-005 0.14939 0.81273 0.85624 0.0014284 0.92565 0.47247 0.0019231 0.42336 1.665 1.663 16.0105 144.9589 0.00025781 -85.3988 0.36494
4.469 0.98807 5.4961e-005 3.8183 0.011987 5.8495e-005 0.001159 0.22926 0.00065927 0.22992 0.21204 0 0.032481 0.0389 0 1.2154 0.3962 0.11867 0.015102 7.7911 0.094206 0.00011821 0.79591 0.0074276 0.0082824 0.0014456 0.98617 0.9912 3.1251e-006 1.25e-005 0.14939 0.81326 0.85654 0.0014281 0.9261 0.47265 0.0019228 0.42337 1.6662 1.6642 16.0105 144.9589 0.00025736 -85.4007 0.36594
4.47 0.98807 5.4961e-005 3.8183 0.011987 5.8508e-005 0.001159 0.22927 0.00065927 0.22992 0.21205 0 0.032481 0.0389 0 1.2155 0.39624 0.11868 0.015104 7.7929 0.094216 0.00011823 0.7959 0.0074282 0.0082831 0.0014452 0.98618 0.99121 3.124e-006 1.2496e-005 0.1494 0.8138 0.85683 0.0014279 0.92655 0.47283 0.0019225 0.42339 1.6674 1.6654 16.0105 144.9589 0.00025691 -85.4025 0.36694
4.471 0.98807 5.496e-005 3.8183 0.011986 5.8521e-005 0.001159 0.22927 0.00065927 0.22993 0.21205 0 0.032481 0.0389 0 1.2156 0.39629 0.1187 0.015105 7.7946 0.094226 0.00011824 0.79589 0.0074289 0.0082838 0.0014447 0.98618 0.99121 3.123e-006 1.2492e-005 0.1494 0.81432 0.85712 0.0014277 0.927 0.47301 0.0019222 0.4234 1.6686 1.6666 16.0106 144.9589 0.00025646 -85.4044 0.36794
4.472 0.98807 5.496e-005 3.8183 0.011986 5.8534e-005 0.001159 0.22928 0.00065927 0.22993 0.21206 0 0.032481 0.0389 0 1.2157 0.39634 0.11871 0.015107 7.7963 0.094235 0.00011825 0.79588 0.0074296 0.0082846 0.0014443 0.98619 0.99121 3.122e-006 1.2488e-005 0.14941 0.81485 0.8574 0.0014274 0.92744 0.4732 0.0019219 0.42341 1.6698 1.6677 16.0106 144.9589 0.00025602 -85.4062 0.36894
4.473 0.98807 5.496e-005 3.8183 0.011986 5.8547e-005 0.001159 0.22928 0.00065927 0.22994 0.21206 0 0.03248 0.0389 0 1.2158 0.39638 0.11873 0.015108 7.798 0.094245 0.00011827 0.79587 0.0074302 0.0082853 0.0014438 0.9862 0.99122 3.121e-006 1.2484e-005 0.14941 0.81538 0.85769 0.0014272 0.92789 0.47338 0.0019216 0.42342 1.6709 1.6689 16.0106 144.9589 0.00025558 -85.408 0.36994
4.474 0.98807 5.496e-005 3.8183 0.011986 5.856e-005 0.001159 0.22929 0.00065927 0.22994 0.21207 0 0.03248 0.0389 0 1.2159 0.39643 0.11875 0.01511 7.7997 0.094255 0.00011828 0.79586 0.0074309 0.008286 0.0014434 0.9862 0.99122 3.12e-006 1.248e-005 0.14942 0.8159 0.85798 0.001427 0.92833 0.47356 0.0019213 0.42343 1.6721 1.6701 16.0106 144.959 0.00025514 -85.4098 0.37094
4.475 0.98807 5.496e-005 3.8183 0.011986 5.8573e-005 0.001159 0.22929 0.00065927 0.22994 0.21207 0 0.03248 0.0389 0 1.216 0.39648 0.11876 0.015112 7.8014 0.094265 0.0001183 0.79585 0.0074316 0.0082867 0.001443 0.98621 0.99122 3.119e-006 1.2476e-005 0.14942 0.81642 0.85826 0.0014268 0.92876 0.47374 0.001921 0.42345 1.6733 1.6713 16.0106 144.959 0.0002547 -85.4116 0.37194
4.476 0.98807 5.496e-005 3.8183 0.011986 5.8586e-005 0.001159 0.22929 0.00065927 0.22995 0.21207 0 0.03248 0.0389 0 1.216 0.39652 0.11878 0.015113 7.8032 0.094275 0.00011831 0.79584 0.0074322 0.0082874 0.0014426 0.98621 0.99123 3.1181e-006 1.2472e-005 0.14943 0.81695 0.85854 0.0014266 0.9292 0.47392 0.0019208 0.42346 1.6745 1.6725 16.0106 144.959 0.00025426 -85.4134 0.37294
4.477 0.98807 5.496e-005 3.8183 0.011986 5.8599e-005 0.001159 0.2293 0.00065927 0.22995 0.21208 0 0.032479 0.0389 0 1.2161 0.39657 0.11879 0.015115 7.8049 0.094285 0.00011832 0.79583 0.0074329 0.0082882 0.0014421 0.98622 0.99123 3.1171e-006 1.2468e-005 0.14943 0.81747 0.85882 0.0014263 0.92963 0.47411 0.0019205 0.42347 1.6756 1.6736 16.0106 144.959 0.00025383 -85.4151 0.37394
4.478 0.98807 5.496e-005 3.8183 0.011986 5.8612e-005 0.001159 0.2293 0.00065927 0.22996 0.21208 0 0.032479 0.0389 0 1.2162 0.39662 0.11881 0.015116 7.8066 0.094294 0.00011834 0.79582 0.0074336 0.0082889 0.0014417 0.98622 0.99123 3.1161e-006 1.2464e-005 0.14944 0.81798 0.8591 0.0014261 0.93006 0.47429 0.0019202 0.42348 1.6768 1.6748 16.0106 144.959 0.00025339 -85.4169 0.37494
4.479 0.98807 5.496e-005 3.8183 0.011986 5.8625e-005 0.001159 0.22931 0.00065927 0.22996 0.21209 0 0.032479 0.0389 0 1.2163 0.39666 0.11883 0.015118 7.8083 0.094304 0.00011835 0.79581 0.0074342 0.0082896 0.0014413 0.98623 0.99124 3.1152e-006 1.2461e-005 0.14944 0.8185 0.85938 0.0014259 0.93048 0.47447 0.0019199 0.4235 1.6779 1.676 16.0106 144.9591 0.00025296 -85.4186 0.37594
4.48 0.98807 5.496e-005 3.8183 0.011986 5.8638e-005 0.001159 0.22931 0.00065927 0.22997 0.21209 0 0.032479 0.0389 0 1.2164 0.39671 0.11884 0.015119 7.81 0.094314 0.00011837 0.7958 0.0074349 0.0082903 0.0014409 0.98623 0.99124 3.1142e-006 1.2457e-005 0.14945 0.81901 0.85966 0.0014257 0.93091 0.47465 0.0019196 0.42351 1.6791 1.6771 16.0106 144.9591 0.00025253 -85.4204 0.37694
4.481 0.98807 5.496e-005 3.8183 0.011986 5.8651e-005 0.001159 0.22932 0.00065927 0.22997 0.2121 0 0.032479 0.0389 0 1.2165 0.39676 0.11886 0.015121 7.8118 0.094324 0.00011838 0.79579 0.0074356 0.008291 0.0014405 0.98624 0.99125 3.1133e-006 1.2453e-005 0.14945 0.81953 0.85994 0.0014255 0.93133 0.47483 0.0019193 0.42352 1.6803 1.6783 16.0106 144.9591 0.00025211 -85.4221 0.37794
4.482 0.98807 5.496e-005 3.8183 0.011986 5.8664e-005 0.001159 0.22932 0.00065927 0.22998 0.2121 0 0.032478 0.0389 0 1.2166 0.3968 0.11887 0.015123 7.8135 0.094334 0.00011839 0.79578 0.0074362 0.0082917 0.0014401 0.98625 0.99125 3.1123e-006 1.2449e-005 0.14946 0.82004 0.86021 0.0014252 0.93175 0.47501 0.0019191 0.42353 1.6814 1.6795 16.0106 144.9591 0.00025168 -85.4238 0.37894
4.483 0.98808 5.496e-005 3.8183 0.011986 5.8677e-005 0.001159 0.22933 0.00065927 0.22998 0.2121 0 0.032478 0.0389 0 1.2167 0.39685 0.11889 0.015124 7.8152 0.094344 0.00011841 0.79577 0.0074369 0.0082925 0.0014396 0.98625 0.99125 3.1114e-006 1.2446e-005 0.14947 0.82055 0.86049 0.001425 0.93216 0.4752 0.0019188 0.42355 1.6826 1.6806 16.0106 144.9591 0.00025126 -85.4255 0.37994
4.484 0.98808 5.496e-005 3.8183 0.011986 5.8689e-005 0.001159 0.22933 0.00065927 0.22998 0.21211 0 0.032478 0.0389 0 1.2168 0.3969 0.1189 0.015126 7.8169 0.094353 0.00011842 0.79576 0.0074376 0.0082932 0.0014393 0.98626 0.99126 3.1105e-006 1.2442e-005 0.14947 0.82106 0.86076 0.0014248 0.93258 0.47538 0.0019185 0.42356 1.6837 1.6818 16.0106 144.9591 0.00025084 -85.4271 0.38094
4.485 0.98808 5.4959e-005 3.8183 0.011986 5.8702e-005 0.001159 0.22933 0.00065927 0.22999 0.21211 0 0.032478 0.0389 0 1.2169 0.39694 0.11892 0.015127 7.8186 0.094363 0.00011843 0.79576 0.0074382 0.0082939 0.0014389 0.98626 0.99126 3.1095e-006 1.2438e-005 0.14948 0.82156 0.86103 0.0014246 0.93299 0.47556 0.0019182 0.42357 1.6848 1.6829 16.0106 144.9592 0.00025042 -85.4288 0.38194
4.486 0.98808 5.4959e-005 3.8183 0.011986 5.8715e-005 0.001159 0.22934 0.00065927 0.22999 0.21212 0 0.032478 0.0389 0 1.217 0.39699 0.11894 0.015129 7.8204 0.094373 0.00011845 0.79575 0.0074389 0.0082946 0.0014385 0.98627 0.99126 3.1086e-006 1.2435e-005 0.14948 0.82207 0.8613 0.0014244 0.9334 0.47574 0.001918 0.42358 1.686 1.6841 16.0106 144.9592 0.00025 -85.4305 0.38294
4.487 0.98808 5.4959e-005 3.8183 0.011986 5.8728e-005 0.001159 0.22934 0.00065927 0.23 0.21212 0 0.032477 0.0389 0 1.2171 0.39704 0.11895 0.015131 7.8221 0.094383 0.00011846 0.79574 0.0074396 0.0082953 0.0014381 0.98627 0.99127 3.1077e-006 1.2431e-005 0.14949 0.82257 0.86157 0.0014242 0.9338 0.47592 0.0019177 0.4236 1.6871 1.6852 16.0106 144.9592 0.00024958 -85.4321 0.38394
4.488 0.98808 5.4959e-005 3.8183 0.011986 5.8741e-005 0.001159 0.22935 0.00065927 0.23 0.21212 0 0.032477 0.0389 0 1.2172 0.39708 0.11897 0.015132 7.8238 0.094393 0.00011848 0.79573 0.0074402 0.008296 0.0014377 0.98628 0.99127 3.1068e-006 1.2427e-005 0.14949 0.82307 0.86184 0.001424 0.93421 0.4761 0.0019174 0.42361 1.6882 1.6863 16.0106 144.9592 0.00024917 -85.4337 0.38494
4.489 0.98808 5.4959e-005 3.8183 0.011986 5.8754e-005 0.001159 0.22935 0.00065928 0.23001 0.21213 0 0.032477 0.0389 0 1.2173 0.39713 0.11898 0.015134 7.8255 0.094403 0.00011849 0.79572 0.0074409 0.0082968 0.0014373 0.98628 0.99127 3.1059e-006 1.2424e-005 0.1495 0.82357 0.86211 0.0014238 0.93461 0.47628 0.0019172 0.42362 1.6894 1.6875 16.0106 144.9592 0.00024875 -85.4354 0.38594
4.49 0.98808 5.4959e-005 3.8183 0.011986 5.8767e-005 0.001159 0.22936 0.00065928 0.23001 0.21213 0 0.032477 0.0389 0 1.2174 0.39718 0.119 0.015135 7.8273 0.094412 0.0001185 0.79571 0.0074416 0.0082975 0.0014369 0.98629 0.99128 3.1051e-006 1.242e-005 0.1495 0.82407 0.86237 0.0014236 0.935 0.47647 0.0019169 0.42363 1.6905 1.6886 16.0106 144.9593 0.00024834 -85.437 0.38694
4.491 0.98808 5.4959e-005 3.8183 0.011986 5.878e-005 0.001159 0.22936 0.00065928 0.23002 0.21214 0 0.032476 0.0389 0 1.2175 0.39722 0.11902 0.015137 7.829 0.094422 0.00011852 0.7957 0.0074422 0.0082982 0.0014365 0.98629 0.99128 3.1042e-006 1.2417e-005 0.14951 0.82457 0.86264 0.0014234 0.9354 0.47665 0.0019166 0.42365 1.6916 1.6897 16.0106 144.9593 0.00024793 -85.4386 0.38794
4.492 0.98808 5.4959e-005 3.8183 0.011986 5.8793e-005 0.001159 0.22936 0.00065928 0.23002 0.21214 0 0.032476 0.0389 0 1.2176 0.39727 0.11903 0.015139 7.8307 0.094432 0.00011853 0.79569 0.0074429 0.0082989 0.0014361 0.9863 0.99128 3.1033e-006 1.2413e-005 0.14951 0.82507 0.8629 0.0014232 0.93579 0.47683 0.0019164 0.42366 1.6927 1.6909 16.0106 144.9593 0.00024753 -85.4401 0.38894
4.493 0.98808 5.4959e-005 3.8183 0.011986 5.8806e-005 0.001159 0.22937 0.00065928 0.23002 0.21215 0 0.032476 0.0389 0 1.2177 0.39732 0.11905 0.01514 7.8324 0.094442 0.00011854 0.79568 0.0074436 0.0082996 0.0014358 0.9863 0.99129 3.1025e-006 1.241e-005 0.14952 0.82556 0.86316 0.001423 0.93618 0.47701 0.0019161 0.42367 1.6939 1.692 16.0106 144.9593 0.00024712 -85.4417 0.38994
4.494 0.98808 5.4959e-005 3.8183 0.011986 5.8819e-005 0.001159 0.22937 0.00065928 0.23003 0.21215 0 0.032476 0.0389 0 1.2178 0.39736 0.11906 0.015142 7.8342 0.094452 0.00011856 0.79567 0.0074442 0.0083003 0.0014354 0.98631 0.99129 3.1016e-006 1.2406e-005 0.14952 0.82605 0.86342 0.0014228 0.93657 0.47719 0.0019159 0.42369 1.695 1.6931 16.0106 144.9593 0.00024672 -85.4433 0.39094
4.495 0.98808 5.4959e-005 3.8183 0.011986 5.8832e-005 0.001159 0.22938 0.00065928 0.23003 0.21215 0 0.032476 0.0389 0 1.2179 0.39741 0.11908 0.015143 7.8359 0.094462 0.00011857 0.79566 0.0074449 0.0083011 0.001435 0.98631 0.99129 3.1007e-006 1.2403e-005 0.14953 0.82654 0.86368 0.0014226 0.93696 0.47737 0.0019156 0.4237 1.6961 1.6942 16.0106 144.9594 0.00024631 -85.4448 0.39194
4.496 0.98808 5.4959e-005 3.8183 0.011986 5.8845e-005 0.0011591 0.22938 0.00065928 0.23004 0.21216 0 0.032475 0.0389 0 1.218 0.39746 0.11909 0.015145 7.8376 0.094471 0.00011859 0.79565 0.0074455 0.0083018 0.0014347 0.98632 0.9913 3.0999e-006 1.24e-005 0.14953 0.82703 0.86394 0.0014224 0.93734 0.47755 0.0019154 0.42371 1.6972 1.6953 16.0106 144.9594 0.00024591 -85.4464 0.39294
4.497 0.98808 5.4959e-005 3.8183 0.011986 5.8858e-005 0.0011591 0.22939 0.00065928 0.23004 0.21216 0 0.032475 0.0389 0 1.2181 0.3975 0.11911 0.015147 7.8393 0.094481 0.0001186 0.79564 0.0074462 0.0083025 0.0014343 0.98632 0.9913 3.0991e-006 1.2396e-005 0.14954 0.82752 0.8642 0.0014222 0.93772 0.47773 0.0019151 0.42372 1.6983 1.6964 16.0106 144.9594 0.00024551 -85.4479 0.39394
4.498 0.98808 5.4959e-005 3.8183 0.011986 5.8871e-005 0.0011591 0.22939 0.00065928 0.23005 0.21217 0 0.032475 0.0389 0 1.2182 0.39755 0.11913 0.015148 7.8411 0.094491 0.00011861 0.79563 0.0074469 0.0083032 0.0014339 0.98633 0.9913 3.0982e-006 1.2393e-005 0.14955 0.82801 0.86446 0.0014221 0.9381 0.47791 0.0019149 0.42374 1.6994 1.6976 16.0106 144.9594 0.00024512 -85.4494 0.39494
4.499 0.98808 5.4958e-005 3.8183 0.011986 5.8884e-005 0.0011591 0.2294 0.00065928 0.23005 0.21217 0 0.032475 0.0389 0 1.2183 0.3976 0.11914 0.01515 7.8428 0.094501 0.00011863 0.79562 0.0074475 0.0083039 0.0014336 0.98633 0.99131 3.0974e-006 1.239e-005 0.14955 0.82849 0.86471 0.0014219 0.93848 0.47809 0.0019146 0.42375 1.7005 1.6987 16.0106 144.9594 0.00024472 -85.4509 0.39594
4.5 0.98808 5.4958e-005 3.8183 0.011986 5.8897e-005 0.0011591 0.2294 0.00065928 0.23005 0.21217 0 0.032474 0.0389 0 1.2184 0.39764 0.11916 0.015151 7.8445 0.094511 0.00011864 0.79561 0.0074482 0.0083046 0.0014332 0.98634 0.99131 3.0966e-006 1.2386e-005 0.14956 0.82898 0.86497 0.0014217 0.93885 0.47827 0.0019144 0.42376 1.7016 1.6998 16.0106 144.9594 0.00024433 -85.4524 0.39694
4.501 0.98808 5.4958e-005 3.8183 0.011986 5.891e-005 0.0011591 0.2294 0.00065928 0.23006 0.21218 0 0.032474 0.0389 0 1.2185 0.39769 0.11917 0.015153 7.8462 0.09452 0.00011866 0.7956 0.0074489 0.0083054 0.0014328 0.98634 0.99131 3.0958e-006 1.2383e-005 0.14956 0.82946 0.86522 0.0014215 0.93923 0.47845 0.0019142 0.42377 1.7027 1.7009 16.0106 144.9595 0.00024394 -85.4539 0.39794
4.502 0.98808 5.4958e-005 3.8183 0.011986 5.8923e-005 0.0011591 0.22941 0.00065928 0.23006 0.21218 0 0.032474 0.0389 0 1.2186 0.39774 0.11919 0.015154 7.848 0.09453 0.00011867 0.79559 0.0074495 0.0083061 0.0014325 0.98634 0.99131 3.095e-006 1.238e-005 0.14957 0.82994 0.86547 0.0014213 0.93959 0.47863 0.0019139 0.42379 1.7038 1.702 16.0106 144.9595 0.00024354 -85.4554 0.39894
4.503 0.98808 5.4958e-005 3.8183 0.011986 5.8936e-005 0.0011591 0.22941 0.00065928 0.23007 0.21219 0 0.032474 0.0389 0 1.2187 0.39778 0.11921 0.015156 7.8497 0.09454 0.00011868 0.79558 0.0074502 0.0083068 0.0014321 0.98635 0.99132 3.0942e-006 1.2377e-005 0.14957 0.83042 0.86573 0.0014211 0.93996 0.47882 0.0019137 0.4238 1.7049 1.703 16.0106 144.9595 0.00024316 -85.4569 0.39994
4.504 0.98808 5.4958e-005 3.8183 0.011986 5.8949e-005 0.0011591 0.22942 0.00065928 0.23007 0.21219 0 0.032474 0.0389 0 1.2188 0.39783 0.11922 0.015158 7.8514 0.09455 0.0001187 0.79557 0.0074509 0.0083075 0.0014318 0.98635 0.99132 3.0934e-006 1.2373e-005 0.14958 0.8309 0.86598 0.001421 0.94033 0.479 0.0019134 0.42381 1.7059 1.7041 16.0106 144.9595 0.00024277 -85.4583 0.40094
4.505 0.98808 5.4958e-005 3.8183 0.011986 5.8962e-005 0.0011591 0.22942 0.00065928 0.23008 0.21219 0 0.032473 0.0389 0 1.2189 0.39788 0.11924 0.015159 7.8531 0.09456 0.00011871 0.79556 0.0074515 0.0083082 0.0014315 0.98636 0.99132 3.0926e-006 1.237e-005 0.14958 0.83137 0.86622 0.0014208 0.94069 0.47918 0.0019132 0.42382 1.707 1.7052 16.0106 144.9595 0.00024238 -85.4598 0.40194
4.506 0.98808 5.4958e-005 3.8183 0.011986 5.8975e-005 0.0011591 0.22943 0.00065928 0.23008 0.2122 0 0.032473 0.0389 0 1.219 0.39792 0.11925 0.015161 7.8549 0.09457 0.00011872 0.79555 0.0074522 0.0083089 0.0014311 0.98636 0.99133 3.0918e-006 1.2367e-005 0.14959 0.83185 0.86647 0.0014206 0.94105 0.47936 0.001913 0.42384 1.7081 1.7063 16.0106 144.9596 0.000242 -85.4612 0.40294
4.507 0.98808 5.4958e-005 3.8183 0.011986 5.8988e-005 0.0011591 0.22943 0.00065928 0.23008 0.2122 0 0.032473 0.0389 0 1.2191 0.39797 0.11927 0.015162 7.8566 0.094579 0.00011874 0.79554 0.0074529 0.0083096 0.0014308 0.98637 0.99133 3.091e-006 1.2364e-005 0.14959 0.83232 0.86672 0.0014204 0.94141 0.47954 0.0019127 0.42385 1.7092 1.7074 16.0106 144.9596 0.00024162 -85.4626 0.40394
4.508 0.98808 5.4958e-005 3.8183 0.011986 5.9001e-005 0.0011591 0.22943 0.00065928 0.23009 0.21221 0 0.032473 0.0389 0 1.2192 0.39802 0.11929 0.015164 7.8583 0.094589 0.00011875 0.79553 0.0074535 0.0083104 0.0014304 0.98637 0.99133 3.0902e-006 1.2361e-005 0.1496 0.83279 0.86697 0.0014202 0.94176 0.47972 0.0019125 0.42386 1.7103 1.7085 16.0106 144.9596 0.00024124 -85.464 0.40494
4.509 0.98808 5.4958e-005 3.8183 0.011986 5.9014e-005 0.0011591 0.22944 0.00065928 0.23009 0.21221 0 0.032472 0.0389 0 1.2193 0.39806 0.1193 0.015166 7.8601 0.094599 0.00011877 0.79552 0.0074542 0.0083111 0.0014301 0.98638 0.99133 3.0895e-006 1.2358e-005 0.1496 0.83326 0.86721 0.0014201 0.94212 0.4799 0.0019123 0.42388 1.7113 1.7095 16.0106 144.9596 0.00024086 -85.4654 0.40594
4.51 0.98808 5.4958e-005 3.8183 0.011986 5.9027e-005 0.0011591 0.22944 0.00065928 0.2301 0.21221 0 0.032472 0.0389 0 1.2194 0.39811 0.11932 0.015167 7.8618 0.094609 0.00011878 0.79551 0.0074548 0.0083118 0.0014297 0.98638 0.99134 3.0887e-006 1.2355e-005 0.14961 0.83373 0.86745 0.0014199 0.94247 0.48008 0.0019121 0.42389 1.7124 1.7106 16.0106 144.9596 0.00024048 -85.4668 0.40694
4.511 0.98808 5.4958e-005 3.8183 0.011986 5.904e-005 0.0011591 0.22945 0.00065928 0.2301 0.21222 0 0.032472 0.0389 0 1.2195 0.39816 0.11933 0.015169 7.8635 0.094619 0.00011879 0.7955 0.0074555 0.0083125 0.0014294 0.98638 0.99134 3.0879e-006 1.2352e-005 0.14961 0.8342 0.8677 0.0014197 0.94282 0.48026 0.0019118 0.4239 1.7134 1.7117 16.0106 144.9597 0.0002401 -85.4682 0.40794
4.512 0.98808 5.4958e-005 3.8183 0.011986 5.9053e-005 0.0011591 0.22945 0.00065928 0.23011 0.21222 0 0.032472 0.0389 0 1.2196 0.3982 0.11935 0.01517 7.8653 0.094628 0.00011881 0.79549 0.0074562 0.0083132 0.0014291 0.98639 0.99134 3.0872e-006 1.2349e-005 0.14962 0.83466 0.86794 0.0014195 0.94317 0.48044 0.0019116 0.42391 1.7145 1.7127 16.0106 144.9597 0.00023973 -85.4696 0.40894
4.513 0.98808 5.4957e-005 3.8183 0.011986 5.9066e-005 0.0011591 0.22946 0.00065928 0.23011 0.21223 0 0.032472 0.0389 0 1.2197 0.39825 0.11936 0.015172 7.867 0.094638 0.00011882 0.79548 0.0074568 0.0083139 0.0014288 0.98639 0.99135 3.0864e-006 1.2346e-005 0.14962 0.83513 0.86818 0.0014194 0.94351 0.48062 0.0019114 0.42393 1.7156 1.7138 16.0106 144.9597 0.00023936 -85.471 0.40994
4.514 0.98808 5.4957e-005 3.8183 0.011986 5.9079e-005 0.0011591 0.22946 0.00065928 0.23011 0.21223 0 0.032471 0.0389 0 1.2198 0.3983 0.11938 0.015173 7.8687 0.094648 0.00011883 0.79547 0.0074575 0.0083147 0.0014284 0.9864 0.99135 3.0857e-006 1.2343e-005 0.14963 0.83559 0.86842 0.0014192 0.94385 0.4808 0.0019112 0.42394 1.7166 1.7149 16.0106 144.9597 0.00023898 -85.4723 0.41094
4.515 0.98808 5.4957e-005 3.8183 0.011986 5.9092e-005 0.0011591 0.22946 0.00065928 0.23012 0.21224 0 0.032471 0.0389 0 1.2199 0.39834 0.1194 0.015175 7.8704 0.094658 0.00011885 0.79546 0.0074582 0.0083154 0.0014281 0.9864 0.99135 3.085e-006 1.234e-005 0.14964 0.83605 0.86866 0.001419 0.94419 0.48098 0.0019109 0.42395 1.7177 1.7159 16.0106 144.9597 0.00023861 -85.4737 0.41194
4.516 0.98808 5.4957e-005 3.8183 0.011986 5.9105e-005 0.0011591 0.22947 0.00065928 0.23012 0.21224 0 0.032471 0.0389 0 1.22 0.39839 0.11941 0.015177 7.8722 0.094668 0.00011886 0.79545 0.0074588 0.0083161 0.0014278 0.98641 0.99135 3.0842e-006 1.2337e-005 0.14964 0.83651 0.8689 0.0014189 0.94453 0.48116 0.0019107 0.42397 1.7187 1.717 16.0106 144.9598 0.00023825 -85.475 0.41294
4.517 0.98808 5.4957e-005 3.8183 0.011986 5.9118e-005 0.0011591 0.22947 0.00065928 0.23013 0.21224 0 0.032471 0.0389 0 1.2201 0.39844 0.11943 0.015178 7.8739 0.094677 0.00011888 0.79544 0.0074595 0.0083168 0.0014275 0.98641 0.99136 3.0835e-006 1.2334e-005 0.14965 0.83697 0.86913 0.0014187 0.94487 0.48134 0.0019105 0.42398 1.7198 1.718 16.0106 144.9598 0.00023788 -85.4763 0.41394
4.518 0.98808 5.4957e-005 3.8183 0.011986 5.9131e-005 0.0011591 0.22948 0.00065928 0.23013 0.21225 0 0.032471 0.0389 0 1.2201 0.39848 0.11944 0.01518 7.8756 0.094687 0.00011889 0.79543 0.0074602 0.0083175 0.0014272 0.98641 0.99136 3.0828e-006 1.2331e-005 0.14965 0.83743 0.86937 0.0014186 0.9452 0.48152 0.0019103 0.42399 1.7208 1.7191 16.0106 144.9598 0.00023752 -85.4776 0.41494
4.519 0.98808 5.4957e-005 3.8183 0.011986 5.9144e-005 0.0011591 0.22948 0.00065928 0.23014 0.21225 0 0.03247 0.0389 0 1.2202 0.39853 0.11946 0.015181 7.8774 0.094697 0.0001189 0.79542 0.0074608 0.0083182 0.0014269 0.98642 0.99136 3.0821e-006 1.2328e-005 0.14966 0.83788 0.8696 0.0014184 0.94554 0.4817 0.0019101 0.424 1.7219 1.7201 16.0106 144.9598 0.00023715 -85.479 0.41594
4.52 0.98808 5.4957e-005 3.8183 0.011986 5.9157e-005 0.0011591 0.22949 0.00065928 0.23014 0.21226 0 0.03247 0.0389 0 1.2203 0.39858 0.11948 0.015183 7.8791 0.094707 0.00011892 0.79541 0.0074615 0.0083189 0.0014265 0.98642 0.99136 3.0814e-006 1.2325e-005 0.14966 0.83834 0.86984 0.0014182 0.94587 0.48187 0.0019099 0.42402 1.7229 1.7212 16.0106 144.9598 0.00023679 -85.4803 0.41694
4.521 0.98808 5.4957e-005 3.8183 0.011986 5.917e-005 0.0011591 0.22949 0.00065928 0.23014 0.21226 0 0.03247 0.0389 0 1.2204 0.39862 0.11949 0.015185 7.8808 0.094717 0.00011893 0.7954 0.0074621 0.0083197 0.0014262 0.98643 0.99137 3.0807e-006 1.2323e-005 0.14967 0.83879 0.87007 0.0014181 0.94619 0.48205 0.0019097 0.42403 1.7239 1.7222 16.0106 144.9598 0.00023643 -85.4815 0.41794
4.522 0.98808 5.4957e-005 3.8183 0.011986 5.9183e-005 0.0011591 0.22949 0.00065928 0.23015 0.21226 0 0.03247 0.0389 0 1.2205 0.39867 0.11951 0.015186 7.8826 0.094726 0.00011894 0.79539 0.0074628 0.0083204 0.0014259 0.98643 0.99137 3.08e-006 1.232e-005 0.14967 0.83924 0.8703 0.0014179 0.94652 0.48223 0.0019095 0.42404 1.725 1.7233 16.0106 144.9599 0.00023607 -85.4828 0.41894
4.523 0.98808 5.4957e-005 3.8183 0.011986 5.9196e-005 0.0011591 0.2295 0.00065928 0.23015 0.21227 0 0.032469 0.0389 0 1.2206 0.39872 0.11952 0.015188 7.8843 0.094736 0.00011896 0.79538 0.0074635 0.0083211 0.0014256 0.98643 0.99137 3.0793e-006 1.2317e-005 0.14968 0.83969 0.87053 0.0014177 0.94684 0.48241 0.0019092 0.42406 1.726 1.7243 16.0106 144.9599 0.00023571 -85.4841 0.41994
4.524 0.98808 5.4957e-005 3.8183 0.011986 5.9209e-005 0.0011591 0.2295 0.00065928 0.23016 0.21227 0 0.032469 0.0389 0 1.2207 0.39876 0.11954 0.015189 7.8861 0.094746 0.00011897 0.79537 0.0074641 0.0083218 0.0014253 0.98644 0.99138 3.0786e-006 1.2314e-005 0.14968 0.84014 0.87076 0.0014176 0.94717 0.48259 0.001909 0.42407 1.727 1.7253 16.0106 144.9599 0.00023536 -85.4854 0.42094
4.525 0.98808 5.4957e-005 3.8183 0.011986 5.9222e-005 0.0011591 0.22951 0.00065928 0.23016 0.21228 0 0.032469 0.0389 0 1.2208 0.39881 0.11955 0.015191 7.8878 0.094756 0.00011899 0.79536 0.0074648 0.0083225 0.0014251 0.98644 0.99138 3.0779e-006 1.2312e-005 0.14969 0.84059 0.87099 0.0014174 0.94749 0.48277 0.0019088 0.42408 1.728 1.7263 16.0106 144.9599 0.000235 -85.4866 0.42194
4.526 0.98808 5.4957e-005 3.8183 0.011986 5.9235e-005 0.0011591 0.22951 0.00065928 0.23017 0.21228 0 0.032469 0.0389 0 1.2209 0.39886 0.11957 0.015193 7.8895 0.094766 0.000119 0.79535 0.0074655 0.0083232 0.0014248 0.98645 0.99138 3.0772e-006 1.2309e-005 0.14969 0.84104 0.87122 0.0014173 0.9478 0.48295 0.0019086 0.4241 1.7291 1.7274 16.0106 144.9599 0.00023465 -85.4879 0.42294
4.527 0.98808 5.4956e-005 3.8183 0.011986 5.9248e-005 0.0011591 0.22952 0.00065928 0.23017 0.21228 0 0.032469 0.0389 0 1.221 0.3989 0.11959 0.015194 7.8913 0.094775 0.00011901 0.79534 0.0074661 0.0083239 0.0014245 0.98645 0.99138 3.0765e-006 1.2306e-005 0.1497 0.84148 0.87144 0.0014171 0.94812 0.48313 0.0019084 0.42411 1.7301 1.7284 16.0106 144.96 0.0002343 -85.4891 0.42394
4.528 0.98808 5.4956e-005 3.8183 0.011986 5.9261e-005 0.0011591 0.22952 0.00065928 0.23017 0.21229 0 0.032468 0.0389 0 1.2211 0.39895 0.1196 0.015196 7.893 0.094785 0.00011903 0.79533 0.0074668 0.0083246 0.0014242 0.98645 0.99139 3.0759e-006 1.2303e-005 0.1497 0.84192 0.87167 0.001417 0.94843 0.48331 0.0019082 0.42412 1.7311 1.7294 16.0106 144.96 0.00023395 -85.4903 0.42494
4.529 0.98808 5.4956e-005 3.8183 0.011986 5.9274e-005 0.0011591 0.22952 0.00065928 0.23018 0.21229 0 0.032468 0.0389 0 1.2212 0.399 0.11962 0.015197 7.8947 0.094795 0.00011904 0.79532 0.0074674 0.0083254 0.0014239 0.98646 0.99139 3.0752e-006 1.2301e-005 0.14971 0.84237 0.87189 0.0014168 0.94875 0.48349 0.001908 0.42413 1.7321 1.7304 16.0106 144.96 0.0002336 -85.4915 0.42594
4.53 0.98808 5.4956e-005 3.8183 0.011986 5.9287e-005 0.0011591 0.22953 0.00065928 0.23018 0.2123 0 0.032468 0.0389 0 1.2213 0.39904 0.11963 0.015199 7.8965 0.094805 0.00011905 0.79531 0.0074681 0.0083261 0.0014236 0.98646 0.99139 3.0746e-006 1.2298e-005 0.14971 0.84281 0.87212 0.0014167 0.94906 0.48367 0.0019078 0.42415 1.7331 1.7315 16.0106 144.96 0.00023325 -85.4928 0.42694
4.531 0.98808 5.4956e-005 3.8183 0.011986 5.93e-005 0.0011591 0.22953 0.00065928 0.23019 0.2123 0 0.032468 0.0389 0 1.2214 0.39909 0.11965 0.0152 7.8982 0.094814 0.00011907 0.7953 0.0074688 0.0083268 0.0014233 0.98646 0.99139 3.0739e-006 1.2296e-005 0.14972 0.84324 0.87234 0.0014165 0.94936 0.48385 0.0019076 0.42416 1.7341 1.7325 16.0106 144.96 0.00023291 -85.494 0.42794
4.532 0.98808 5.4956e-005 3.8183 0.011986 5.9313e-005 0.0011591 0.22954 0.00065928 0.23019 0.2123 0 0.032468 0.0389 0 1.2215 0.39914 0.11967 0.015202 7.8999 0.094824 0.00011908 0.79529 0.0074694 0.0083275 0.001423 0.98647 0.9914 3.0732e-006 1.2293e-005 0.14972 0.84368 0.87256 0.0014164 0.94967 0.48402 0.0019075 0.42417 1.7351 1.7335 16.0106 144.9601 0.00023256 -85.4952 0.42894
4.533 0.98808 5.4956e-005 3.8183 0.011986 5.9326e-005 0.0011591 0.22954 0.00065928 0.2302 0.21231 0 0.032467 0.0389 0 1.2216 0.39918 0.11968 0.015204 7.9017 0.094834 0.0001191 0.79529 0.0074701 0.0083282 0.0014227 0.98647 0.9914 3.0726e-006 1.229e-005 0.14973 0.84412 0.87279 0.0014162 0.94998 0.4842 0.0019073 0.42419 1.7361 1.7345 16.0106 144.9601 0.00023222 -85.4963 0.42994
4.534 0.98808 5.4956e-005 3.8183 0.011986 5.9339e-005 0.0011592 0.22954 0.00065928 0.2302 0.21231 0 0.032467 0.0389 0 1.2217 0.39923 0.1197 0.015205 7.9034 0.094844 0.00011911 0.79528 0.0074708 0.0083289 0.0014225 0.98648 0.9914 3.072e-006 1.2288e-005 0.14974 0.84455 0.87301 0.0014161 0.95028 0.48438 0.0019071 0.4242 1.7371 1.7355 16.0106 144.9601 0.00023188 -85.4975 0.43094
4.535 0.98808 5.4956e-005 3.8183 0.011985 5.9352e-005 0.0011592 0.22955 0.00065928 0.2302 0.21232 0 0.032467 0.0389 0 1.2218 0.39928 0.11971 0.015207 7.9052 0.094854 0.00011912 0.79527 0.0074714 0.0083296 0.0014222 0.98648 0.9914 3.0713e-006 1.2285e-005 0.14974 0.84499 0.87322 0.0014159 0.95058 0.48456 0.0019069 0.42421 1.7381 1.7365 16.0106 144.9601 0.00023154 -85.4987 0.43194
4.536 0.98808 5.4956e-005 3.8183 0.011985 5.9365e-005 0.0011592 0.22955 0.00065928 0.23021 0.21232 0 0.032467 0.0389 0 1.2219 0.39932 0.11973 0.015208 7.9069 0.094863 0.00011914 0.79526 0.0074721 0.0083304 0.0014219 0.98648 0.9914 3.0707e-006 1.2283e-005 0.14975 0.84542 0.87344 0.0014158 0.95088 0.48474 0.0019067 0.42423 1.7391 1.7375 16.0105 144.9601 0.0002312 -85.4999 0.43294
4.537 0.98808 5.4956e-005 3.8183 0.011985 5.9378e-005 0.0011592 0.22956 0.00065928 0.23021 0.21232 0 0.032466 0.0389 0 1.222 0.39937 0.11974 0.01521 7.9086 0.094873 0.00011915 0.79525 0.0074727 0.0083311 0.0014216 0.98649 0.99141 3.0701e-006 1.228e-005 0.14975 0.84585 0.87366 0.0014157 0.95117 0.48492 0.0019065 0.42424 1.7401 1.7385 16.0105 144.9602 0.00023086 -85.501 0.43394
4.538 0.98808 5.4956e-005 3.8183 0.011985 5.9391e-005 0.0011592 0.22956 0.00065928 0.23022 0.21233 0 0.032466 0.0389 0 1.2221 0.39942 0.11976 0.015212 7.9104 0.094883 0.00011916 0.79524 0.0074734 0.0083318 0.0014214 0.98649 0.99141 3.0694e-006 1.2278e-005 0.14976 0.84628 0.87388 0.0014155 0.95147 0.4851 0.0019063 0.42425 1.7411 1.7395 16.0105 144.9602 0.00023052 -85.5022 0.43494
4.539 0.98808 5.4956e-005 3.8183 0.011985 5.9404e-005 0.0011592 0.22957 0.00065928 0.23022 0.21233 0 0.032466 0.0389 0 1.2222 0.39946 0.11978 0.015213 7.9121 0.094893 0.00011918 0.79523 0.0074741 0.0083325 0.0014211 0.98649 0.99141 3.0688e-006 1.2275e-005 0.14976 0.84671 0.87409 0.0014154 0.95176 0.48528 0.0019061 0.42426 1.7421 1.7405 16.0105 144.9602 0.00023019 -85.5033 0.43594
4.54 0.98808 5.4955e-005 3.8183 0.011985 5.9417e-005 0.0011592 0.22957 0.00065928 0.23022 0.21234 0 0.032466 0.0389 0 1.2223 0.39951 0.11979 0.015215 7.9139 0.094903 0.00011919 0.79522 0.0074747 0.0083332 0.0014208 0.9865 0.99141 3.0682e-006 1.2273e-005 0.14977 0.84714 0.87431 0.0014152 0.95205 0.48545 0.001906 0.42428 1.7431 1.7415 16.0105 144.9602 0.00022986 -85.5044 0.43694
4.541 0.98808 5.4955e-005 3.8183 0.011985 5.943e-005 0.0011592 0.22957 0.00065928 0.23023 0.21234 0 0.032466 0.0389 0 1.2224 0.39956 0.11981 0.015216 7.9156 0.094912 0.00011921 0.79521 0.0074754 0.0083339 0.0014205 0.9865 0.99142 3.0676e-006 1.227e-005 0.14977 0.84756 0.87452 0.0014151 0.95234 0.48563 0.0019058 0.42429 1.744 1.7424 16.0105 144.9602 0.00022953 -85.5055 0.43794
4.542 0.98808 5.4955e-005 3.8183 0.011985 5.9443e-005 0.0011592 0.22958 0.00065928 0.23023 0.21234 0 0.032465 0.0389 0 1.2225 0.3996 0.11982 0.015218 7.9174 0.094922 0.00011922 0.7952 0.0074761 0.0083346 0.0014203 0.9865 0.99142 3.067e-006 1.2268e-005 0.14978 0.84799 0.87474 0.001415 0.95263 0.48581 0.0019056 0.4243 1.745 1.7434 16.0105 144.9603 0.00022919 -85.5067 0.43894
4.543 0.98808 5.4955e-005 3.8183 0.011985 5.9456e-005 0.0011592 0.22958 0.00065928 0.23024 0.21235 0 0.032465 0.0389 0 1.2226 0.39965 0.11984 0.015219 7.9191 0.094932 0.00011923 0.79519 0.0074767 0.0083353 0.00142 0.98651 0.99142 3.0664e-006 1.2266e-005 0.14978 0.84841 0.87495 0.0014148 0.95291 0.48599 0.0019054 0.42432 1.746 1.7444 16.0105 144.9603 0.00022887 -85.5078 0.43994
4.544 0.98808 5.4955e-005 3.8183 0.011985 5.9469e-005 0.0011592 0.22959 0.00065928 0.23024 0.21235 0 0.032465 0.0389 0 1.2227 0.3997 0.11985 0.015221 7.9208 0.094942 0.00011925 0.79518 0.0074774 0.0083361 0.0014198 0.98651 0.99142 3.0658e-006 1.2263e-005 0.14979 0.84883 0.87516 0.0014147 0.9532 0.48617 0.0019052 0.42433 1.747 1.7454 16.0105 144.9603 0.00022854 -85.5089 0.44094
4.545 0.98808 5.4955e-005 3.8183 0.011985 5.9482e-005 0.0011592 0.22959 0.00065928 0.23025 0.21236 0 0.032465 0.0389 0 1.2228 0.39974 0.11987 0.015223 7.9226 0.094951 0.00011926 0.79517 0.007478 0.0083368 0.0014195 0.98651 0.99142 3.0652e-006 1.2261e-005 0.14979 0.84925 0.87537 0.0014145 0.95348 0.48635 0.0019051 0.42434 1.7479 1.7464 16.0105 144.9603 0.00022821 -85.5099 0.44194
4.546 0.98808 5.4955e-005 3.8183 0.011985 5.9495e-005 0.0011592 0.22959 0.00065928 0.23025 0.21236 0 0.032465 0.0389 0 1.2229 0.39979 0.11989 0.015224 7.9243 0.094961 0.00011927 0.79516 0.0074787 0.0083375 0.0014193 0.98652 0.99143 3.0646e-006 1.2258e-005 0.1498 0.84967 0.87558 0.0014144 0.95376 0.48652 0.0019049 0.42436 1.7489 1.7473 16.0105 144.9603 0.00022789 -85.511 0.44294
4.547 0.98808 5.4955e-005 3.8183 0.011985 5.9508e-005 0.0011592 0.2296 0.00065928 0.23025 0.21236 0 0.032464 0.0389 0 1.223 0.39984 0.1199 0.015226 7.9261 0.094971 0.00011929 0.79515 0.0074794 0.0083382 0.001419 0.98652 0.99143 3.064e-006 1.2256e-005 0.1498 0.85009 0.87579 0.0014143 0.95404 0.4867 0.0019047 0.42437 1.7499 1.7483 16.0105 144.9603 0.00022756 -85.5121 0.44394
4.548 0.98808 5.4955e-005 3.8183 0.011985 5.9521e-005 0.0011592 0.2296 0.00065928 0.23026 0.21237 0 0.032464 0.0389 0 1.2231 0.39988 0.11992 0.015227 7.9278 0.094981 0.0001193 0.79514 0.00748 0.0083389 0.0014188 0.98652 0.99143 3.0635e-006 1.2254e-005 0.14981 0.8505 0.87599 0.0014141 0.95432 0.48688 0.0019045 0.42438 1.7508 1.7493 16.0105 144.9604 0.00022724 -85.5132 0.44494
4.549 0.98808 5.4955e-005 3.8183 0.011985 5.9534e-005 0.0011592 0.22961 0.00065928 0.23026 0.21237 0 0.032464 0.0389 0 1.2232 0.39993 0.11993 0.015229 7.9296 0.094991 0.00011932 0.79513 0.0074807 0.0083396 0.0014185 0.98653 0.99143 3.0629e-006 1.2252e-005 0.14981 0.85092 0.8762 0.001414 0.95459 0.48706 0.0019044 0.4244 1.7518 1.7502 16.0105 144.9604 0.00022692 -85.5142 0.44594
4.55 0.98808 5.4955e-005 3.8183 0.011985 5.9547e-005 0.0011592 0.22961 0.00065928 0.23027 0.21238 0 0.032464 0.0389 0 1.2233 0.39998 0.11995 0.01523 7.9313 0.095 0.00011933 0.79512 0.0074813 0.0083403 0.0014182 0.98653 0.99144 3.0623e-006 1.2249e-005 0.14982 0.85133 0.87641 0.0014139 0.95486 0.48724 0.0019042 0.42441 1.7528 1.7512 16.0105 144.9604 0.0002266 -85.5153 0.44694
4.551 0.98808 5.4955e-005 3.8183 0.011985 5.956e-005 0.0011592 0.22962 0.00065928 0.23027 0.21238 0 0.032464 0.0389 0 1.2234 0.40002 0.11997 0.015232 7.933 0.09501 0.00011934 0.79511 0.007482 0.008341 0.001418 0.98653 0.99144 3.0618e-006 1.2247e-005 0.14983 0.85174 0.87661 0.0014138 0.95514 0.48741 0.001904 0.42442 1.7537 1.7522 16.0105 144.9604 0.00022628 -85.5163 0.44794
4.552 0.98808 5.4955e-005 3.8183 0.011985 5.9573e-005 0.0011592 0.22962 0.00065928 0.23027 0.21238 0 0.032463 0.0389 0 1.2235 0.40007 0.11998 0.015234 7.9348 0.09502 0.00011936 0.7951 0.0074827 0.0083418 0.0014177 0.98654 0.99144 3.0612e-006 1.2245e-005 0.14983 0.85216 0.87682 0.0014136 0.95541 0.48759 0.0019039 0.42443 1.7547 1.7531 16.0105 144.9604 0.00022596 -85.5174 0.44894
4.553 0.98808 5.4955e-005 3.8183 0.011985 5.9586e-005 0.0011592 0.22962 0.00065928 0.23028 0.21239 0 0.032463 0.0389 0 1.2236 0.40012 0.12 0.015235 7.9365 0.09503 0.00011937 0.79509 0.0074833 0.0083425 0.0014175 0.98654 0.99144 3.0606e-006 1.2242e-005 0.14984 0.85257 0.87702 0.0014135 0.95567 0.48777 0.0019037 0.42445 1.7556 1.7541 16.0105 144.9605 0.00022565 -85.5184 0.44994
4.554 0.98808 5.4954e-005 3.8183 0.011985 5.9599e-005 0.0011592 0.22963 0.00065928 0.23028 0.21239 0 0.032463 0.0389 0 1.2237 0.40016 0.12001 0.015237 7.9383 0.095039 0.00011938 0.79508 0.007484 0.0083432 0.0014173 0.98654 0.99144 3.0601e-006 1.224e-005 0.14984 0.85297 0.87722 0.0014134 0.95594 0.48795 0.0019035 0.42446 1.7566 1.755 16.0104 144.9605 0.00022533 -85.5194 0.45094
4.555 0.98808 5.4954e-005 3.8183 0.011985 5.9612e-005 0.0011592 0.22963 0.00065928 0.23029 0.21239 0 0.032463 0.0389 0 1.2238 0.40021 0.12003 0.015238 7.94 0.095049 0.0001194 0.79507 0.0074846 0.0083439 0.001417 0.98655 0.99145 3.0595e-006 1.2238e-005 0.14985 0.85338 0.87743 0.0014132 0.95621 0.48812 0.0019034 0.42447 1.7575 1.756 16.0104 144.9605 0.00022502 -85.5204 0.45194
4.556 0.98808 5.4954e-005 3.8183 0.011985 5.9625e-005 0.0011592 0.22964 0.00065928 0.23029 0.2124 0 0.032463 0.0389 0 1.2239 0.40026 0.12004 0.01524 7.9418 0.095059 0.00011941 0.79506 0.0074853 0.0083446 0.0014168 0.98655 0.99145 3.059e-006 1.2236e-005 0.14985 0.85379 0.87763 0.0014131 0.95647 0.4883 0.0019032 0.42449 1.7584 1.7569 16.0104 144.9605 0.00022471 -85.5215 0.45294
4.557 0.98808 5.4954e-005 3.8183 0.011985 5.9638e-005 0.0011592 0.22964 0.00065928 0.2303 0.2124 0 0.032462 0.0389 0 1.2239 0.4003 0.12006 0.015242 7.9435 0.095069 0.00011943 0.79505 0.007486 0.0083453 0.0014166 0.98655 0.99145 3.0584e-006 1.2234e-005 0.14986 0.85419 0.87783 0.001413 0.95673 0.48848 0.001903 0.4245 1.7594 1.7579 16.0104 144.9605 0.0002244 -85.5225 0.45394
4.558 0.98808 5.4954e-005 3.8183 0.011985 5.9651e-005 0.0011592 0.22964 0.00065928 0.2303 0.21241 0 0.032462 0.0389 0 1.224 0.40035 0.12008 0.015243 7.9453 0.095078 0.00011944 0.79504 0.0074866 0.008346 0.0014163 0.98656 0.99145 3.0579e-006 1.2232e-005 0.14986 0.8546 0.87803 0.0014129 0.95699 0.48866 0.0019029 0.42451 1.7603 1.7588 16.0104 144.9606 0.00022409 -85.5235 0.45494
4.559 0.98808 5.4954e-005 3.8183 0.011985 5.9663e-005 0.0011592 0.22965 0.00065928 0.2303 0.21241 0 0.032462 0.0389 0 1.2241 0.4004 0.12009 0.015245 7.947 0.095088 0.00011945 0.79503 0.0074873 0.0083467 0.0014161 0.98656 0.99145 3.0574e-006 1.2229e-005 0.14987 0.855 0.87823 0.0014128 0.95725 0.48883 0.0019027 0.42453 1.7613 1.7597 16.0104 144.9606 0.00022378 -85.5244 0.45594
4.56 0.98808 5.4954e-005 3.8183 0.011985 5.9676e-005 0.0011592 0.22965 0.00065928 0.23031 0.21241 0 0.032462 0.0389 0 1.2242 0.40044 0.12011 0.015246 7.9488 0.095098 0.00011947 0.79502 0.0074879 0.0083474 0.0014158 0.98656 0.99146 3.0568e-006 1.2227e-005 0.14987 0.8554 0.87842 0.0014126 0.9575 0.48901 0.0019026 0.42454 1.7622 1.7607 16.0104 144.9606 0.00022347 -85.5254 0.45694
4.561 0.98808 5.4954e-005 3.8183 0.011985 5.9689e-005 0.0011592 0.22966 0.00065928 0.23031 0.21242 0 0.032461 0.0389 0 1.2243 0.40049 0.12012 0.015248 7.9505 0.095108 0.00011948 0.79501 0.0074886 0.0083482 0.0014156 0.98656 0.99146 3.0563e-006 1.2225e-005 0.14988 0.8558 0.87862 0.0014125 0.95776 0.48919 0.0019024 0.42455 1.7631 1.7616 16.0104 144.9606 0.00022317 -85.5264 0.45794
4.562 0.98808 5.4954e-005 3.8183 0.011985 5.9702e-005 0.0011592 0.22966 0.00065928 0.23032 0.21242 0 0.032461 0.0389 0 1.2244 0.40054 0.12014 0.015249 7.9523 0.095117 0.00011949 0.795 0.0074893 0.0083489 0.0014154 0.98657 0.99146 3.0558e-006 1.2223e-005 0.14988 0.8562 0.87882 0.0014124 0.95801 0.48937 0.0019022 0.42457 1.764 1.7625 16.0104 144.9606 0.00022286 -85.5274 0.45894
4.563 0.98808 5.4954e-005 3.8183 0.011985 5.9715e-005 0.0011592 0.22967 0.00065928 0.23032 0.21243 0 0.032461 0.0389 0 1.2245 0.40058 0.12016 0.015251 7.954 0.095127 0.00011951 0.79499 0.0074899 0.0083496 0.0014152 0.98657 0.99146 3.0553e-006 1.2221e-005 0.14989 0.8566 0.87901 0.0014123 0.95826 0.48954 0.0019021 0.42458 1.765 1.7635 16.0104 144.9607 0.00022256 -85.5283 0.45994
4.564 0.98808 5.4954e-005 3.8183 0.011985 5.9728e-005 0.0011592 0.22967 0.00065928 0.23032 0.21243 0 0.032461 0.0389 0 1.2246 0.40063 0.12017 0.015253 7.9558 0.095137 0.00011952 0.79498 0.0074906 0.0083503 0.0014149 0.98657 0.99146 3.0547e-006 1.2219e-005 0.14989 0.85699 0.87921 0.0014122 0.95851 0.48972 0.0019019 0.42459 1.7659 1.7644 16.0104 144.9607 0.00022226 -85.5293 0.46094
4.565 0.98808 5.4954e-005 3.8183 0.011985 5.9741e-005 0.0011592 0.22967 0.00065928 0.23033 0.21243 0 0.032461 0.0389 0 1.2247 0.40068 0.12019 0.015254 7.9575 0.095147 0.00011954 0.79497 0.0074912 0.008351 0.0014147 0.98658 0.99147 3.0542e-006 1.2217e-005 0.1499 0.85739 0.8794 0.001412 0.95876 0.4899 0.0019018 0.42461 1.7668 1.7653 16.0104 144.9607 0.00022196 -85.5302 0.46194
4.566 0.98808 5.4954e-005 3.8183 0.011985 5.9754e-005 0.0011592 0.22968 0.00065928 0.23033 0.21244 0 0.03246 0.0389 0 1.2248 0.40072 0.1202 0.015256 7.9593 0.095156 0.00011955 0.79496 0.0074919 0.0083517 0.0014145 0.98658 0.99147 3.0537e-006 1.2215e-005 0.1499 0.85778 0.87959 0.0014119 0.95901 0.49007 0.0019016 0.42462 1.7677 1.7662 16.0104 144.9607 0.00022166 -85.5312 0.46294
4.567 0.98808 5.4954e-005 3.8183 0.011985 5.9767e-005 0.0011592 0.22968 0.00065928 0.23034 0.21244 0 0.03246 0.0389 0 1.2249 0.40077 0.12022 0.015257 7.961 0.095166 0.00011956 0.79495 0.0074926 0.0083524 0.0014143 0.98658 0.99147 3.0532e-006 1.2213e-005 0.14991 0.85817 0.87979 0.0014118 0.95926 0.49025 0.0019015 0.42463 1.7686 1.7672 16.0104 144.9607 0.00022136 -85.5321 0.46394
4.568 0.98808 5.4953e-005 3.8183 0.011985 5.978e-005 0.0011592 0.22969 0.00065928 0.23034 0.21245 0 0.03246 0.0389 0 1.225 0.40082 0.12023 0.015259 7.9628 0.095176 0.00011958 0.79494 0.0074932 0.0083531 0.0014141 0.98658 0.99147 3.0527e-006 1.2211e-005 0.14991 0.85856 0.87998 0.0014117 0.9595 0.49043 0.0019013 0.42465 1.7696 1.7681 16.0103 144.9608 0.00022106 -85.533 0.46494
4.569 0.98808 5.4953e-005 3.8183 0.011985 5.9793e-005 0.0011592 0.22969 0.00065928 0.23034 0.21245 0 0.03246 0.0389 0 1.2251 0.40086 0.12025 0.015261 7.9645 0.095186 0.00011959 0.79493 0.0074939 0.0083538 0.0014138 0.98659 0.99147 3.0522e-006 1.2209e-005 0.14992 0.85895 0.88017 0.0014116 0.95974 0.4906 0.0019012 0.42466 1.7705 1.769 16.0103 144.9608 0.00022077 -85.534 0.46594
4.57 0.98808 5.4953e-005 3.8183 0.011985 5.9806e-005 0.0011592 0.22969 0.00065928 0.23035 0.21245 0 0.03246 0.0389 0 1.2252 0.40091 0.12027 0.015262 7.9663 0.095195 0.0001196 0.79492 0.0074945 0.0083545 0.0014136 0.98659 0.99147 3.0517e-006 1.2207e-005 0.14992 0.85934 0.88036 0.0014115 0.95998 0.49078 0.001901 0.42467 1.7714 1.7699 16.0103 144.9608 0.00022047 -85.5349 0.46694
4.571 0.98808 5.4953e-005 3.8183 0.011985 5.9819e-005 0.0011592 0.2297 0.00065928 0.23035 0.21246 0 0.032459 0.0389 0 1.2253 0.40096 0.12028 0.015264 7.968 0.095205 0.00011962 0.79491 0.0074952 0.0083553 0.0014134 0.98659 0.99148 3.0512e-006 1.2205e-005 0.14993 0.85973 0.88055 0.0014113 0.96022 0.49096 0.0019009 0.42469 1.7723 1.7708 16.0103 144.9608 0.00022018 -85.5358 0.46794
4.572 0.98808 5.4953e-005 3.8183 0.011985 5.9832e-005 0.0011593 0.2297 0.00065928 0.23036 0.21246 0 0.032459 0.0389 0 1.2254 0.401 0.1203 0.015265 7.9698 0.095215 0.00011963 0.7949 0.0074959 0.008356 0.0014132 0.9866 0.99148 3.0507e-006 1.2203e-005 0.14994 0.86012 0.88074 0.0014112 0.96046 0.49113 0.0019007 0.4247 1.7732 1.7717 16.0103 144.9608 0.00021989 -85.5367 0.46894
4.573 0.98808 5.4953e-005 3.8183 0.011985 5.9845e-005 0.0011593 0.22971 0.00065928 0.23036 0.21246 0 0.032459 0.0389 0 1.2255 0.40105 0.12031 0.015267 7.9715 0.095225 0.00011964 0.79489 0.0074965 0.0083567 0.001413 0.9866 0.99148 3.0503e-006 1.2201e-005 0.14994 0.8605 0.88092 0.0014111 0.9607 0.49131 0.0019006 0.42471 1.7741 1.7726 16.0103 144.9609 0.00021959 -85.5376 0.46994
4.574 0.98808 5.4953e-005 3.8183 0.011985 5.9858e-005 0.0011593 0.22971 0.00065928 0.23036 0.21247 0 0.032459 0.0389 0 1.2256 0.4011 0.12033 0.015268 7.9733 0.095234 0.00011966 0.79489 0.0074972 0.0083574 0.0014128 0.9866 0.99148 3.0498e-006 1.2199e-005 0.14995 0.86089 0.88111 0.001411 0.96093 0.49149 0.0019004 0.42472 1.775 1.7735 16.0103 144.9609 0.0002193 -85.5385 0.47094
4.575 0.98808 5.4953e-005 3.8183 0.011985 5.9871e-005 0.0011593 0.22971 0.00065928 0.23037 0.21247 0 0.032459 0.0389 0 1.2257 0.40114 0.12035 0.01527 7.975 0.095244 0.00011967 0.79488 0.0074978 0.0083581 0.0014126 0.9866 0.99148 3.0493e-006 1.2197e-005 0.14995 0.86127 0.8813 0.0014109 0.96116 0.49166 0.0019003 0.42474 1.7759 1.7744 16.0103 144.9609 0.00021902 -85.5394 0.47194
4.576 0.98808 5.4953e-005 3.8183 0.011985 5.9884e-005 0.0011593 0.22972 0.00065928 0.23037 0.21248 0 0.032458 0.0389 0 1.2258 0.40119 0.12036 0.015272 7.9768 0.095254 0.00011969 0.79487 0.0074985 0.0083588 0.0014124 0.98661 0.99149 3.0488e-006 1.2195e-005 0.14996 0.86165 0.88148 0.0014108 0.9614 0.49184 0.0019002 0.42475 1.7768 1.7753 16.0103 144.9609 0.00021873 -85.5402 0.47294
4.577 0.98808 5.4953e-005 3.8183 0.011985 5.9897e-005 0.0011593 0.22972 0.00065928 0.23038 0.21248 0 0.032458 0.0389 0 1.2259 0.40124 0.12038 0.015273 7.9785 0.095264 0.0001197 0.79486 0.0074991 0.0083595 0.0014122 0.98661 0.99149 3.0484e-006 1.2193e-005 0.14996 0.86203 0.88167 0.0014107 0.96163 0.49202 0.0019 0.42476 1.7777 1.7762 16.0103 144.9609 0.00021844 -85.5411 0.47394
4.578 0.98808 5.4953e-005 3.8183 0.011985 5.991e-005 0.0011593 0.22973 0.00065928 0.23038 0.21248 0 0.032458 0.0389 0 1.226 0.40128 0.12039 0.015275 7.9803 0.095273 0.00011971 0.79485 0.0074998 0.0083602 0.001412 0.98661 0.99149 3.0479e-006 1.2192e-005 0.14997 0.86241 0.88185 0.0014106 0.96185 0.49219 0.0018999 0.42478 1.7785 1.7771 16.0103 144.961 0.00021816 -85.542 0.47494
4.579 0.98808 5.4953e-005 3.8183 0.011985 5.9923e-005 0.0011593 0.22973 0.00065928 0.23038 0.21249 0 0.032458 0.0389 0 1.2261 0.40133 0.12041 0.015276 7.9821 0.095283 0.00011973 0.79484 0.0075005 0.0083609 0.0014117 0.98661 0.99149 3.0474e-006 1.219e-005 0.14997 0.86279 0.88203 0.0014105 0.96208 0.49237 0.0018997 0.42479 1.7794 1.778 16.0102 144.961 0.00021787 -85.5428 0.47594
4.58 0.98808 5.4953e-005 3.8183 0.011985 5.9936e-005 0.0011593 0.22973 0.00065928 0.23039 0.21249 0 0.032458 0.0389 0 1.2262 0.40137 0.12042 0.015278 7.9838 0.095293 0.00011974 0.79483 0.0075011 0.0083616 0.0014115 0.98662 0.99149 3.047e-006 1.2188e-005 0.14998 0.86317 0.88222 0.0014104 0.96231 0.49255 0.0018996 0.4248 1.7803 1.7789 16.0102 144.961 0.00021759 -85.5437 0.47694
4.581 0.98808 5.4953e-005 3.8183 0.011985 5.9949e-005 0.0011593 0.22974 0.00065928 0.23039 0.2125 0 0.032457 0.0389 0 1.2263 0.40142 0.12044 0.015279 7.9856 0.095303 0.00011975 0.79482 0.0075018 0.0083624 0.0014113 0.98662 0.99149 3.0465e-006 1.2186e-005 0.14998 0.86354 0.8824 0.0014103 0.96253 0.49272 0.0018995 0.42482 1.7812 1.7798 16.0102 144.961 0.00021731 -85.5445 0.47794
4.582 0.98808 5.4952e-005 3.8183 0.011985 5.9962e-005 0.0011593 0.22974 0.00065928 0.2304 0.2125 0 0.032457 0.0389 0 1.2264 0.40147 0.12046 0.015281 7.9873 0.095312 0.00011977 0.79481 0.0075024 0.0083631 0.0014111 0.98662 0.9915 3.0461e-006 1.2184e-005 0.14999 0.86392 0.88258 0.0014102 0.96276 0.4929 0.0018993 0.42483 1.7821 1.7807 16.0102 144.961 0.00021703 -85.5454 0.47894
4.583 0.98808 5.4952e-005 3.8183 0.011985 5.9975e-005 0.0011593 0.22975 0.00065928 0.2304 0.2125 0 0.032457 0.0389 0 1.2265 0.40151 0.12047 0.015283 7.9891 0.095322 0.00011978 0.7948 0.0075031 0.0083638 0.0014109 0.98662 0.9915 3.0456e-006 1.2182e-005 0.14999 0.86429 0.88276 0.0014101 0.96298 0.49307 0.0018992 0.42484 1.7829 1.7815 16.0102 144.9611 0.00021675 -85.5462 0.47994
4.584 0.98808 5.4952e-005 3.8183 0.011985 5.9988e-005 0.0011593 0.22975 0.00065928 0.23041 0.21251 0 0.032457 0.0389 0 1.2266 0.40156 0.12049 0.015284 7.9908 0.095332 0.0001198 0.79479 0.0075038 0.0083645 0.0014107 0.98663 0.9915 3.0452e-006 1.2181e-005 0.15 0.86466 0.88294 0.00141 0.9632 0.49325 0.0018991 0.42486 1.7838 1.7824 16.0102 144.9611 0.00021647 -85.5471 0.48094
4.585 0.98808 5.4952e-005 3.8183 0.011985 6.0001e-005 0.0011593 0.22975 0.00065928 0.23041 0.21251 0 0.032457 0.0389 0 1.2267 0.40161 0.1205 0.015286 7.9926 0.095342 0.00011981 0.79478 0.0075044 0.0083652 0.0014106 0.98663 0.9915 3.0447e-006 1.2179e-005 0.15 0.86503 0.88312 0.0014099 0.96342 0.49343 0.0018989 0.42487 1.7847 1.7833 16.0102 144.9611 0.00021619 -85.5479 0.48194
4.586 0.98808 5.4952e-005 3.8183 0.011985 6.0014e-005 0.0011593 0.22976 0.00065928 0.23041 0.21251 0 0.032456 0.0389 0 1.2268 0.40165 0.12052 0.015287 7.9943 0.095351 0.00011982 0.79477 0.0075051 0.0083659 0.0014104 0.98663 0.9915 3.0443e-006 1.2177e-005 0.15001 0.8654 0.88329 0.0014098 0.96363 0.4936 0.0018988 0.42488 1.7856 1.7842 16.0102 144.9611 0.00021591 -85.5487 0.48294
4.587 0.98808 5.4952e-005 3.8183 0.011985 6.0027e-005 0.0011593 0.22976 0.00065928 0.23042 0.21252 0 0.032456 0.0389 0 1.2269 0.4017 0.12054 0.015289 7.9961 0.095361 0.00011984 0.79476 0.0075057 0.0083666 0.0014102 0.98664 0.9915 3.0438e-006 1.2175e-005 0.15001 0.86577 0.88347 0.0014097 0.96385 0.49378 0.0018987 0.4249 1.7864 1.785 16.0102 144.9611 0.00021564 -85.5495 0.48394
4.588 0.98808 5.4952e-005 3.8183 0.011985 6.004e-005 0.0011593 0.22977 0.00065928 0.23042 0.21252 0 0.032456 0.0389 0 1.227 0.40175 0.12055 0.01529 7.9979 0.095371 0.00011985 0.79475 0.0075064 0.0083673 0.00141 0.98664 0.99151 3.0434e-006 1.2174e-005 0.15002 0.86614 0.88365 0.0014096 0.96406 0.49395 0.0018985 0.42491 1.7873 1.7859 16.0102 144.9611 0.00021536 -85.5503 0.48494
4.589 0.98808 5.4952e-005 3.8183 0.011985 6.0053e-005 0.0011593 0.22977 0.00065928 0.23043 0.21253 0 0.032456 0.0389 0 1.2271 0.40179 0.12057 0.015292 7.9996 0.095381 0.00011986 0.79474 0.007507 0.008368 0.0014098 0.98664 0.99151 3.043e-006 1.2172e-005 0.15002 0.86651 0.88382 0.0014095 0.96428 0.49413 0.0018984 0.42492 1.7882 1.7868 16.0101 144.9612 0.00021509 -85.5511 0.48594
4.59 0.98808 5.4952e-005 3.8183 0.011985 6.0066e-005 0.0011593 0.22977 0.00065928 0.23043 0.21253 0 0.032456 0.0389 0 1.2272 0.40184 0.12058 0.015294 8.0014 0.09539 0.00011988 0.79473 0.0075077 0.0083687 0.0014096 0.98664 0.99151 3.0425e-006 1.217e-005 0.15003 0.86687 0.884 0.0014094 0.96449 0.49431 0.0018983 0.42494 1.789 1.7876 16.0101 144.9612 0.00021482 -85.5519 0.48694
4.591 0.98808 5.4952e-005 3.8183 0.011985 6.0079e-005 0.0011593 0.22978 0.00065928 0.23043 0.21253 0 0.032455 0.0389 0 1.2273 0.40189 0.1206 0.015295 8.0031 0.0954 0.00011989 0.79472 0.0075084 0.0083694 0.0014094 0.98664 0.99151 3.0421e-006 1.2168e-005 0.15004 0.86723 0.88417 0.0014093 0.9647 0.49448 0.0018981 0.42495 1.7899 1.7885 16.0101 144.9612 0.00021455 -85.5527 0.48794
4.592 0.98808 5.4952e-005 3.8183 0.011985 6.0092e-005 0.0011593 0.22978 0.00065928 0.23044 0.21254 0 0.032455 0.0389 0 1.2274 0.40193 0.12061 0.015297 8.0049 0.09541 0.00011991 0.79471 0.007509 0.0083702 0.0014092 0.98665 0.99151 3.0417e-006 1.2167e-005 0.15004 0.8676 0.88435 0.0014092 0.96491 0.49466 0.001898 0.42496 1.7907 1.7894 16.0101 144.9612 0.00021428 -85.5535 0.48894
4.593 0.98808 5.4952e-005 3.8183 0.011985 6.0105e-005 0.0011593 0.22979 0.00065928 0.23044 0.21254 0 0.032455 0.0389 0 1.2275 0.40198 0.12063 0.015298 8.0067 0.095419 0.00011992 0.7947 0.0075097 0.0083709 0.001409 0.98665 0.99151 3.0413e-006 1.2165e-005 0.15005 0.86796 0.88452 0.0014091 0.96512 0.49483 0.0018979 0.42498 1.7916 1.7902 16.0101 144.9612 0.00021401 -85.5543 0.48994
4.594 0.98808 5.4952e-005 3.8183 0.011985 6.0118e-005 0.0011593 0.22979 0.00065928 0.23045 0.21255 0 0.032455 0.0389 0 1.2276 0.40203 0.12065 0.0153 8.0084 0.095429 0.00011993 0.79469 0.0075103 0.0083716 0.0014089 0.98665 0.99151 3.0408e-006 1.2163e-005 0.15005 0.86832 0.88469 0.001409 0.96532 0.49501 0.0018978 0.42499 1.7924 1.7911 16.0101 144.9613 0.00021374 -85.5551 0.49094
4.595 0.98808 5.4951e-005 3.8183 0.011985 6.0131e-005 0.0011593 0.22979 0.00065928 0.23045 0.21255 0 0.032455 0.0389 0 1.2276 0.40207 0.12066 0.015301 8.0102 0.095439 0.00011995 0.79468 0.007511 0.0083723 0.0014087 0.98665 0.99152 3.0404e-006 1.2162e-005 0.15006 0.86868 0.88486 0.0014089 0.96553 0.49518 0.0018976 0.425 1.7933 1.7919 16.0101 144.9613 0.00021347 -85.5558 0.49194
4.596 0.98808 5.4951e-005 3.8183 0.011985 6.0144e-005 0.0011593 0.2298 0.00065928 0.23045 0.21255 0 0.032454 0.0389 0 1.2277 0.40212 0.12068 0.015303 8.0119 0.095449 0.00011996 0.79467 0.0075116 0.008373 0.0014085 0.98666 0.99152 3.04e-006 1.216e-005 0.15006 0.86904 0.88504 0.0014088 0.96573 0.49536 0.0018975 0.42502 1.7941 1.7928 16.0101 144.9613 0.00021321 -85.5566 0.49294
4.597 0.98808 5.4951e-005 3.8183 0.011985 6.0157e-005 0.0011593 0.2298 0.00065928 0.23046 0.21256 0 0.032454 0.0389 0 1.2278 0.40217 0.12069 0.015305 8.0137 0.095458 0.00011997 0.79466 0.0075123 0.0083737 0.0014084 0.98666 0.99152 3.0396e-006 1.2158e-005 0.15007 0.8694 0.88521 0.0014087 0.96594 0.49553 0.0018974 0.42503 1.795 1.7936 16.0101 144.9613 0.00021294 -85.5574 0.49394
4.598 0.98808 5.4951e-005 3.8183 0.011985 6.017e-005 0.0011593 0.22981 0.00065928 0.23046 0.21256 0 0.032454 0.0389 0 1.2279 0.40221 0.12071 0.015306 8.0155 0.095468 0.00011999 0.79465 0.007513 0.0083744 0.0014082 0.98666 0.99152 3.0392e-006 1.2157e-005 0.15007 0.86975 0.88538 0.0014086 0.96614 0.49571 0.0018973 0.42504 1.7958 1.7945 16.01 144.9613 0.00021268 -85.5581 0.49494
4.599 0.98808 5.4951e-005 3.8183 0.011984 6.0183e-005 0.0011593 0.22981 0.00065928 0.23047 0.21256 0 0.032454 0.0389 0 1.228 0.40226 0.12072 0.015308 8.0172 0.095478 0.00012 0.79464 0.0075136 0.0083751 0.001408 0.98666 0.99152 3.0388e-006 1.2155e-005 0.15008 0.87011 0.88555 0.0014085 0.96634 0.49588 0.0018972 0.42506 1.7967 1.7953 16.01 144.9614 0.00021242 -85.5589 0.49594
4.6 0.98808 5.4951e-005 3.8183 0.011984 6.0196e-005 0.0011593 0.22981 0.00065928 0.23047 0.21257 0 0.032454 0.0389 0 1.2281 0.40231 0.12074 0.015309 8.019 0.095487 0.00012001 0.79463 0.0075143 0.0083758 0.0014078 0.98667 0.99152 3.0384e-006 1.2154e-005 0.15008 0.87046 0.88571 0.0014084 0.96654 0.49606 0.001897 0.42507 1.7975 1.7962 16.01 144.9614 0.00021216 -85.5596 0.49694
4.601 0.98808 5.4951e-005 3.8183 0.011984 6.0209e-005 0.0011593 0.22982 0.00065928 0.23047 0.21257 0 0.032453 0.0389 0 1.2282 0.40235 0.12076 0.015311 8.0208 0.095497 0.00012003 0.79462 0.0075149 0.0083765 0.0014076 0.98667 0.99153 3.038e-006 1.2152e-005 0.15009 0.87081 0.88588 0.0014083 0.96673 0.49623 0.0018969 0.42508 1.7983 1.797 16.01 144.9614 0.0002119 -85.5603 0.49794
4.602 0.98808 5.4951e-005 3.8183 0.011984 6.0222e-005 0.0011593 0.22982 0.00065928 0.23048 0.21258 0 0.032453 0.0389 0 1.2283 0.4024 0.12077 0.015313 8.0225 0.095507 0.00012004 0.79461 0.0075156 0.0083772 0.0014074 0.98667 0.99153 3.0376e-006 1.215e-005 0.15009 0.87117 0.88605 0.0014082 0.96693 0.49641 0.0018968 0.4251 1.7992 1.7979 16.01 144.9614 0.00021164 -85.5611 0.49894
4.603 0.98808 5.4951e-005 3.8183 0.011984 6.0235e-005 0.0011593 0.22983 0.00065928 0.23048 0.21258 0 0.032453 0.0389 0 1.2284 0.40245 0.12079 0.015314 8.0243 0.095517 0.00012006 0.7946 0.0075162 0.0083779 0.0014073 0.98667 0.99153 3.0372e-006 1.2149e-005 0.1501 0.87152 0.88621 0.0014081 0.96713 0.49658 0.0018967 0.42511 1.8 1.7987 16.01 144.9614 0.00021138 -85.5618 0.49994
4.604 0.98808 5.4951e-005 3.8183 0.011984 6.0248e-005 0.0011593 0.22983 0.00065928 0.23048 0.21258 0 0.032453 0.0389 0 1.2285 0.40249 0.1208 0.015316 8.026 0.095526 0.00012007 0.79459 0.0075169 0.0083786 0.0014071 0.98667 0.99153 3.0368e-006 1.2147e-005 0.1501 0.87187 0.88638 0.0014081 0.96732 0.49676 0.0018966 0.42512 1.8008 1.7995 16.01 144.9615 0.00021112 -85.5625 0.50094
4.605 0.98808 5.4951e-005 3.8183 0.011984 6.0261e-005 0.0011593 0.22983 0.00065928 0.23049 0.21259 0 0.032453 0.0389 0 1.2286 0.40254 0.12082 0.015317 8.0278 0.095536 0.00012008 0.79458 0.0075176 0.0083794 0.001407 0.98668 0.99153 3.0364e-006 1.2146e-005 0.15011 0.87222 0.88655 0.001408 0.96751 0.49693 0.0018964 0.42514 1.8017 1.8004 16.01 144.9615 0.00021086 -85.5632 0.50194
4.606 0.98808 5.4951e-005 3.8183 0.011984 6.0274e-005 0.0011593 0.22984 0.00065928 0.23049 0.21259 0 0.032452 0.0389 0 1.2287 0.40259 0.12084 0.015319 8.0296 0.095546 0.0001201 0.79457 0.0075182 0.0083801 0.0014068 0.98668 0.99153 3.0361e-006 1.2144e-005 0.15011 0.87256 0.88671 0.0014079 0.9677 0.49711 0.0018963 0.42515 1.8025 1.8012 16.01 144.9615 0.00021061 -85.564 0.50294
4.607 0.98808 5.4951e-005 3.8183 0.011984 6.0287e-005 0.0011593 0.22984 0.00065928 0.2305 0.21259 0 0.032452 0.0389 0 1.2288 0.40263 0.12085 0.01532 8.0313 0.095556 0.00012011 0.79456 0.0075189 0.0083808 0.0014066 0.98668 0.99153 3.0357e-006 1.2143e-005 0.15012 0.87291 0.88687 0.0014078 0.96789 0.49728 0.0018962 0.42516 1.8033 1.802 16.0099 144.9615 0.00021035 -85.5647 0.50394
4.608 0.98808 5.4951e-005 3.8183 0.011984 6.03e-005 0.0011593 0.22985 0.00065928 0.2305 0.2126 0 0.032452 0.0389 0 1.2289 0.40268 0.12087 0.015322 8.0331 0.095565 0.00012012 0.79455 0.0075195 0.0083815 0.0014065 0.98668 0.99154 3.0353e-006 1.2141e-005 0.15012 0.87326 0.88704 0.0014077 0.96808 0.49746 0.0018961 0.42518 1.8041 1.8028 16.0099 144.9615 0.0002101 -85.5654 0.50494
4.609 0.98808 5.495e-005 3.8183 0.011984 6.0313e-005 0.0011593 0.22985 0.00065928 0.2305 0.2126 0 0.032452 0.0389 0 1.229 0.40273 0.12088 0.015324 8.0349 0.095575 0.00012014 0.79455 0.0075202 0.0083822 0.0014063 0.98669 0.99154 3.0349e-006 1.214e-005 0.15013 0.8736 0.8872 0.0014076 0.96827 0.49763 0.001896 0.42519 1.805 1.8037 16.0099 144.9616 0.00020985 -85.5661 0.50594
4.61 0.98808 5.495e-005 3.8183 0.011984 6.0326e-005 0.0011594 0.22985 0.00065928 0.23051 0.21261 0 0.032452 0.0389 0 1.2291 0.40277 0.1209 0.015325 8.0366 0.095585 0.00012015 0.79454 0.0075208 0.0083829 0.0014061 0.98669 0.99154 3.0345e-006 1.2138e-005 0.15013 0.87394 0.88736 0.0014075 0.96846 0.49781 0.0018959 0.4252 1.8058 1.8045 16.0099 144.9616 0.0002096 -85.5668 0.50694
4.611 0.98808 5.495e-005 3.8183 0.011984 6.0339e-005 0.0011594 0.22986 0.00065928 0.23051 0.21261 0 0.032451 0.0389 0 1.2292 0.40282 0.12091 0.015327 8.0384 0.095594 0.00012016 0.79453 0.0075215 0.0083836 0.0014059 0.98669 0.99154 3.0342e-006 1.2137e-005 0.15014 0.87428 0.88752 0.0014074 0.96864 0.49798 0.0018958 0.42522 1.8066 1.8053 16.0099 144.9616 0.00020935 -85.5675 0.50794
4.612 0.98808 5.495e-005 3.8183 0.011984 6.0352e-005 0.0011594 0.22986 0.00065928 0.23052 0.21261 0 0.032451 0.0389 0 1.2293 0.40287 0.12093 0.015328 8.0402 0.095604 0.00012018 0.79452 0.0075222 0.0083843 0.0014058 0.98669 0.99154 3.0338e-006 1.2135e-005 0.15014 0.87463 0.88768 0.0014074 0.96883 0.49816 0.0018957 0.42523 1.8074 1.8061 16.0099 144.9616 0.0002091 -85.5681 0.50894
4.613 0.98808 5.495e-005 3.8183 0.011984 6.0365e-005 0.0011594 0.22987 0.00065928 0.23052 0.21262 0 0.032451 0.0389 0 1.2294 0.40291 0.12095 0.01533 8.0419 0.095614 0.00012019 0.79451 0.0075228 0.008385 0.0014056 0.98669 0.99154 3.0334e-006 1.2134e-005 0.15015 0.87497 0.88784 0.0014073 0.96901 0.49833 0.0018956 0.42524 1.8082 1.8069 16.0099 144.9616 0.00020885 -85.5688 0.50994
4.614 0.98808 5.495e-005 3.8183 0.011984 6.0378e-005 0.0011594 0.22987 0.00065928 0.23052 0.21262 0 0.032451 0.0389 0 1.2295 0.40296 0.12096 0.015331 8.0437 0.095623 0.00012021 0.7945 0.0075235 0.0083857 0.0014055 0.9867 0.99154 3.0331e-006 1.2132e-005 0.15016 0.8753 0.888 0.0014072 0.96919 0.4985 0.0018954 0.42526 1.809 1.8077 16.0099 144.9617 0.0002086 -85.5695 0.51094
4.615 0.98808 5.495e-005 3.8183 0.011984 6.0391e-005 0.0011594 0.22987 0.00065928 0.23053 0.21262 0 0.032451 0.0389 0 1.2296 0.40301 0.12098 0.015333 8.0455 0.095633 0.00012022 0.79449 0.0075241 0.0083864 0.0014054 0.9867 0.99154 3.0327e-006 1.2131e-005 0.15016 0.87564 0.88816 0.0014071 0.96937 0.49868 0.0018953 0.42527 1.8098 1.8086 16.0098 144.9617 0.00020835 -85.5702 0.51194
4.616 0.98808 5.495e-005 3.8183 0.011984 6.0404e-005 0.0011594 0.22988 0.00065928 0.23053 0.21263 0 0.03245 0.0389 0 1.2297 0.40305 0.12099 0.015335 8.0472 0.095643 0.00012023 0.79448 0.0075248 0.0083871 0.0014052 0.9867 0.99155 3.0324e-006 1.2129e-005 0.15017 0.87598 0.88832 0.001407 0.96955 0.49885 0.0018952 0.42528 1.8106 1.8094 16.0098 144.9617 0.00020811 -85.5708 0.51294
4.617 0.98808 5.495e-005 3.8183 0.011984 6.0417e-005 0.0011594 0.22988 0.00065928 0.23054 0.21263 0 0.03245 0.0389 0 1.2298 0.4031 0.12101 0.015336 8.049 0.095653 0.00012025 0.79447 0.0075254 0.0083878 0.001405 0.9867 0.99155 3.032e-006 1.2128e-005 0.15017 0.87632 0.88848 0.001407 0.96973 0.49903 0.0018951 0.4253 1.8114 1.8102 16.0098 144.9617 0.00020786 -85.5715 0.51394
4.618 0.98808 5.495e-005 3.8183 0.011984 6.043e-005 0.0011594 0.22989 0.00065928 0.23054 0.21264 0 0.03245 0.0389 0 1.2299 0.40315 0.12102 0.015338 8.0508 0.095662 0.00012026 0.79446 0.0075261 0.0083885 0.0014049 0.9867 0.99155 3.0317e-006 1.2127e-005 0.15018 0.87665 0.88863 0.0014069 0.96991 0.4992 0.001895 0.42531 1.8122 1.811 16.0098 144.9617 0.00020762 -85.5722 0.51494
4.619 0.98808 5.495e-005 3.8183 0.011984 6.0443e-005 0.0011594 0.22989 0.00065928 0.23054 0.21264 0 0.03245 0.0389 0 1.23 0.40319 0.12104 0.015339 8.0526 0.095672 0.00012027 0.79445 0.0075267 0.0083892 0.0014047 0.98671 0.99155 3.0313e-006 1.2125e-005 0.15018 0.87698 0.88879 0.0014068 0.97008 0.49937 0.0018949 0.42532 1.813 1.8118 16.0098 144.9618 0.00020738 -85.5728 0.51594
4.62 0.98808 5.495e-005 3.8183 0.011984 6.0455e-005 0.0011594 0.22989 0.00065928 0.23055 0.21264 0 0.03245 0.0389 0 1.2301 0.40324 0.12106 0.015341 8.0543 0.095682 0.00012029 0.79444 0.0075274 0.00839 0.0014045 0.98671 0.99155 3.031e-006 1.2124e-005 0.15019 0.87732 0.88895 0.0014067 0.97026 0.49955 0.0018948 0.42534 1.8138 1.8126 16.0098 144.9618 0.00020714 -85.5735 0.51694
4.621 0.98808 5.495e-005 3.8183 0.011984 6.0468e-005 0.0011594 0.2299 0.00065928 0.23055 0.21265 0 0.032449 0.0389 0 1.2302 0.40329 0.12107 0.015342 8.0561 0.095691 0.0001203 0.79443 0.0075281 0.0083907 0.0014043 0.98671 0.99155 3.0306e-006 1.2122e-005 0.15019 0.87765 0.8891 0.0014066 0.97043 0.49972 0.0018947 0.42535 1.8146 1.8134 16.0098 144.9618 0.0002069 -85.5741 0.51794
4.622 0.98808 5.495e-005 3.8183 0.011984 6.0481e-005 0.0011594 0.2299 0.00065928 0.23056 0.21265 0 0.032449 0.0389 0 1.2303 0.40333 0.12109 0.015344 8.0579 0.095701 0.00012032 0.79442 0.0075287 0.0083914 0.0014042 0.98671 0.99155 3.0303e-006 1.2121e-005 0.1502 0.87798 0.88925 0.0014065 0.9706 0.4999 0.0018946 0.42536 1.8154 1.8142 16.0097 144.9618 0.00020666 -85.5747 0.51894
4.623 0.98808 5.4949e-005 3.8183 0.011984 6.0494e-005 0.0011594 0.2299 0.00065928 0.23056 0.21265 0 0.032449 0.0389 0 1.2304 0.40338 0.1211 0.015346 8.0596 0.095711 0.00012033 0.79441 0.0075294 0.0083921 0.0014041 0.98671 0.99156 3.0299e-006 1.212e-005 0.1502 0.87831 0.88941 0.0014065 0.97078 0.50007 0.0018945 0.42538 1.8162 1.815 16.0097 144.9618 0.00020642 -85.5754 0.51994
4.624 0.98808 5.4949e-005 3.8183 0.011984 6.0507e-005 0.0011594 0.22991 0.00065928 0.23056 0.21266 0 0.032449 0.0389 0 1.2305 0.40343 0.12112 0.015347 8.0614 0.09572 0.00012034 0.7944 0.00753 0.0083928 0.001404 0.98672 0.99156 3.0296e-006 1.2118e-005 0.15021 0.87864 0.88956 0.0014064 0.97095 0.50024 0.0018944 0.42539 1.817 1.8158 16.0097 144.9619 0.00020618 -85.576 0.52094
4.625 0.98808 5.4949e-005 3.8183 0.011984 6.052e-005 0.0011594 0.22991 0.00065928 0.23057 0.21266 0 0.032449 0.0389 0 1.2306 0.40347 0.12114 0.015349 8.0632 0.09573 0.00012036 0.79439 0.0075307 0.0083935 0.0014038 0.98672 0.99156 3.0293e-006 1.2117e-005 0.15021 0.87896 0.88971 0.0014063 0.97112 0.50042 0.0018943 0.4254 1.8178 1.8165 16.0097 144.9619 0.00020594 -85.5766 0.52194
4.626 0.98808 5.4949e-005 3.8183 0.011984 6.0533e-005 0.0011594 0.22992 0.00065928 0.23057 0.21266 0 0.032448 0.0389 0 1.2307 0.40352 0.12115 0.01535 8.0649 0.09574 0.00012037 0.79438 0.0075313 0.0083942 0.0014037 0.98672 0.99156 3.0289e-006 1.2116e-005 0.15022 0.87929 0.88987 0.0014063 0.97128 0.50059 0.0018942 0.42542 1.8186 1.8173 16.0097 144.9619 0.00020571 -85.5773 0.52294
4.627 0.98808 5.4949e-005 3.8183 0.011984 6.0546e-005 0.0011594 0.22992 0.00065928 0.23058 0.21267 0 0.032448 0.0389 0 1.2308 0.40357 0.12117 0.015352 8.0667 0.09575 0.00012038 0.79437 0.007532 0.0083949 0.0014036 0.98672 0.99156 3.0286e-006 1.2114e-005 0.15022 0.87962 0.89002 0.0014062 0.97145 0.50076 0.0018941 0.42543 1.8193 1.8181 16.0097 144.9619 0.00020547 -85.5779 0.52394
4.628 0.98808 5.4949e-005 3.8183 0.011984 6.0559e-005 0.0011594 0.22992 0.00065928 0.23058 0.21267 0 0.032448 0.0389 0 1.2309 0.40361 0.12118 0.015353 8.0685 0.095759 0.0001204 0.79436 0.0075326 0.0083956 0.0014034 0.98672 0.99156 3.0283e-006 1.2113e-005 0.15023 0.87994 0.89017 0.0014061 0.97162 0.50094 0.001894 0.42544 1.8201 1.8189 16.0097 144.9619 0.00020524 -85.5785 0.52494
4.629 0.98808 5.4949e-005 3.8183 0.011984 6.0572e-005 0.0011594 0.22993 0.00065928 0.23058 0.21268 0 0.032448 0.0389 0 1.231 0.40366 0.1212 0.015355 8.0703 0.095769 0.00012041 0.79435 0.0075333 0.0083963 0.0014032 0.98672 0.99156 3.0279e-006 1.2112e-005 0.15023 0.88026 0.89032 0.001406 0.97178 0.50111 0.0018939 0.42546 1.8209 1.8197 16.0096 144.962 0.000205 -85.5791 0.52594
4.63 0.98808 5.4949e-005 3.8183 0.011984 6.0585e-005 0.0011594 0.22993 0.00065928 0.23059 0.21268 0 0.032448 0.0389 0 1.2311 0.40371 0.12121 0.015357 8.072 0.095779 0.00012042 0.79434 0.0075339 0.008397 0.001403 0.98673 0.99156 3.0276e-006 1.211e-005 0.15024 0.88059 0.89047 0.0014059 0.97195 0.50128 0.0018938 0.42547 1.8217 1.8205 16.0096 144.962 0.00020477 -85.5797 0.52694
4.631 0.98808 5.4949e-005 3.8183 0.011984 6.0598e-005 0.0011594 0.22994 0.00065928 0.23059 0.21268 0 0.032447 0.0389 0 1.2312 0.40375 0.12123 0.015358 8.0738 0.095788 0.00012044 0.79433 0.0075346 0.0083977 0.0014029 0.98673 0.99156 3.0273e-006 1.2109e-005 0.15024 0.88091 0.89062 0.0014058 0.97211 0.50146 0.0018937 0.42548 1.8225 1.8212 16.0096 144.962 0.00020454 -85.5803 0.52794
4.632 0.98808 5.4949e-005 3.8183 0.011984 6.0611e-005 0.0011594 0.22994 0.00065928 0.23059 0.21269 0 0.032447 0.0389 0 1.2312 0.4038 0.12125 0.01536 8.0756 0.095798 0.00012045 0.79432 0.0075353 0.0083984 0.0014028 0.98673 0.99157 3.027e-006 1.2108e-005 0.15025 0.88123 0.89077 0.0014058 0.97227 0.50163 0.0018936 0.4255 1.8232 1.822 16.0096 144.962 0.00020431 -85.5809 0.52894
4.633 0.98808 5.4949e-005 3.8183 0.011984 6.0624e-005 0.0011594 0.22994 0.00065928 0.2306 0.21269 0 0.032447 0.0389 0 1.2313 0.40385 0.12126 0.015361 8.0774 0.095808 0.00012047 0.79431 0.0075359 0.0083991 0.0014026 0.98673 0.99157 3.0267e-006 1.2107e-005 0.15025 0.88155 0.89091 0.0014057 0.97243 0.5018 0.0018935 0.42551 1.824 1.8228 16.0096 144.962 0.00020408 -85.5815 0.52994
4.634 0.98808 5.4949e-005 3.8183 0.011984 6.0637e-005 0.0011594 0.22995 0.00065928 0.2306 0.21269 0 0.032447 0.0389 0 1.2314 0.40389 0.12128 0.015363 8.0791 0.095817 0.00012048 0.7943 0.0075366 0.0083998 0.0014025 0.98673 0.99157 3.0263e-006 1.2105e-005 0.15026 0.88187 0.89106 0.0014056 0.97259 0.50198 0.0018934 0.42552 1.8248 1.8236 16.0096 144.9621 0.00020385 -85.5821 0.53094
4.635 0.98808 5.4949e-005 3.8183 0.011984 6.065e-005 0.0011594 0.22995 0.00065928 0.23061 0.2127 0 0.032447 0.0389 0 1.2315 0.40394 0.12129 0.015364 8.0809 0.095827 0.00012049 0.79429 0.0075372 0.0084005 0.0014024 0.98674 0.99157 3.026e-006 1.2104e-005 0.15026 0.88218 0.89121 0.0014056 0.97275 0.50215 0.0018933 0.42554 1.8255 1.8243 16.0096 144.9621 0.00020362 -85.5827 0.53194
4.636 0.98808 5.4949e-005 3.8183 0.011984 6.0663e-005 0.0011594 0.22996 0.00065928 0.23061 0.2127 0 0.032446 0.0389 0 1.2316 0.40399 0.12131 0.015366 8.0827 0.095837 0.00012051 0.79428 0.0075379 0.0084012 0.0014023 0.98674 0.99157 3.0257e-006 1.2103e-005 0.15027 0.8825 0.89135 0.0014055 0.97291 0.50232 0.0018932 0.42555 1.8263 1.8251 16.0095 144.9621 0.00020339 -85.5833 0.53294
4.637 0.98808 5.4948e-005 3.8183 0.011984 6.0676e-005 0.0011594 0.22996 0.00065928 0.23061 0.21271 0 0.032446 0.0389 0 1.2317 0.40403 0.12132 0.015367 8.0845 0.095846 0.00012052 0.79427 0.0075385 0.0084019 0.0014022 0.98674 0.99157 3.0254e-006 1.2102e-005 0.15028 0.88282 0.8915 0.0014054 0.97307 0.5025 0.0018931 0.42556 1.8271 1.8259 16.0095 144.9621 0.00020317 -85.5838 0.53394
4.638 0.98808 5.4948e-005 3.8183 0.011984 6.0689e-005 0.0011594 0.22996 0.00065928 0.23062 0.21271 0 0.032446 0.0389 0 1.2318 0.40408 0.12134 0.015369 8.0862 0.095856 0.00012053 0.79426 0.0075392 0.0084027 0.0014021 0.98674 0.99157 3.0251e-006 1.21e-005 0.15028 0.88313 0.89165 0.0014054 0.97322 0.50267 0.001893 0.42558 1.8278 1.8266 16.0095 144.9621 0.00020294 -85.5844 0.53494
4.639 0.98808 5.4948e-005 3.8183 0.011984 6.0702e-005 0.0011594 0.22997 0.00065928 0.23062 0.21271 0 0.032446 0.0389 0 1.2319 0.40413 0.12136 0.015371 8.088 0.095866 0.00012055 0.79425 0.0075398 0.0084034 0.0014019 0.98674 0.99157 3.0248e-006 1.2099e-005 0.15029 0.88344 0.89179 0.0014053 0.97338 0.50284 0.001893 0.42559 1.8286 1.8274 16.0095 144.9622 0.00020272 -85.585 0.53594
4.64 0.98808 5.4948e-005 3.8183 0.011984 6.0715e-005 0.0011594 0.22997 0.00065928 0.23063 0.21272 0 0.032446 0.0389 0 1.232 0.40417 0.12137 0.015372 8.0898 0.095875 0.00012056 0.79425 0.0075405 0.0084041 0.0014017 0.98674 0.99158 3.0245e-006 1.2098e-005 0.15029 0.88376 0.89193 0.0014052 0.97353 0.50302 0.0018929 0.4256 1.8293 1.8281 16.0095 144.9622 0.00020249 -85.5855 0.53694
4.641 0.98808 5.4948e-005 3.8183 0.011984 6.0728e-005 0.0011594 0.22997 0.00065928 0.23063 0.21272 0 0.032445 0.0389 0 1.2321 0.40422 0.12139 0.015374 8.0916 0.095885 0.00012057 0.79424 0.0075411 0.0084048 0.0014016 0.98675 0.99158 3.0242e-006 1.2097e-005 0.1503 0.88407 0.89208 0.0014052 0.97368 0.50319 0.0018928 0.42562 1.8301 1.8289 16.0095 144.9622 0.00020227 -85.5861 0.53794
4.642 0.98808 5.4948e-005 3.8183 0.011984 6.0741e-005 0.0011594 0.22998 0.00065928 0.23063 0.21272 0 0.032445 0.0389 0 1.2322 0.40427 0.1214 0.015375 8.0934 0.095895 0.00012059 0.79423 0.0075418 0.0084055 0.0014015 0.98675 0.99158 3.0239e-006 1.2095e-005 0.1503 0.88438 0.89222 0.0014051 0.97384 0.50336 0.0018927 0.42563 1.8308 1.8297 16.0095 144.9622 0.00020205 -85.5867 0.53894
4.643 0.98808 5.4948e-005 3.8183 0.011984 6.0754e-005 0.0011594 0.22998 0.00065928 0.23064 0.21273 0 0.032445 0.0389 0 1.2323 0.40431 0.12142 0.015377 8.0951 0.095905 0.0001206 0.79422 0.0075424 0.0084062 0.0014013 0.98675 0.99158 3.0236e-006 1.2094e-005 0.15031 0.88469 0.89236 0.001405 0.97399 0.50353 0.0018926 0.42564 1.8316 1.8304 16.0094 144.9622 0.00020183 -85.5872 0.53994
4.644 0.98808 5.4948e-005 3.8183 0.011984 6.0767e-005 0.0011594 0.22999 0.00065928 0.23064 0.21273 0 0.032445 0.0389 0 1.2324 0.40436 0.12144 0.015378 8.0969 0.095914 0.00012062 0.79421 0.0075431 0.0084069 0.0014012 0.98675 0.99158 3.0233e-006 1.2093e-005 0.15031 0.885 0.8925 0.0014049 0.97414 0.50371 0.0018925 0.42566 1.8323 1.8312 16.0094 144.9623 0.00020161 -85.5878 0.54094
4.645 0.98808 5.4948e-005 3.8183 0.011984 6.078e-005 0.0011594 0.22999 0.00065928 0.23064 0.21273 0 0.032445 0.0389 0 1.2325 0.40441 0.12145 0.01538 8.0987 0.095924 0.00012063 0.7942 0.0075438 0.0084076 0.0014011 0.98675 0.99158 3.023e-006 1.2092e-005 0.15032 0.8853 0.89265 0.0014049 0.97429 0.50388 0.0018924 0.42567 1.8331 1.8319 16.0094 144.9623 0.00020139 -85.5883 0.54194
4.646 0.98808 5.4948e-005 3.8183 0.011984 6.0793e-005 0.0011594 0.22999 0.00065928 0.23065 0.21274 0 0.032445 0.0389 0 1.2326 0.40445 0.12147 0.015382 8.1005 0.095934 0.00012064 0.79419 0.0075444 0.0084083 0.0014009 0.98675 0.99158 3.0227e-006 1.2091e-005 0.15032 0.88561 0.89279 0.0014048 0.97443 0.50405 0.0018923 0.42568 1.8338 1.8327 16.0094 144.9623 0.00020117 -85.5888 0.54294
4.647 0.98808 5.4948e-005 3.8183 0.011984 6.0806e-005 0.0011595 0.23 0.00065928 0.23065 0.21274 0 0.032444 0.0389 0 1.2327 0.4045 0.12148 0.015383 8.1022 0.095943 0.00012066 0.79418 0.0075451 0.008409 0.0014008 0.98676 0.99158 3.0224e-006 1.209e-005 0.15033 0.88592 0.89293 0.0014047 0.97458 0.50422 0.0018922 0.4257 1.8346 1.8334 16.0094 144.9623 0.00020095 -85.5894 0.54394
4.648 0.98808 5.4948e-005 3.8183 0.011984 6.0819e-005 0.0011595 0.23 0.00065928 0.23066 0.21275 0 0.032444 0.0389 0 1.2328 0.40455 0.1215 0.015385 8.104 0.095953 0.00012067 0.79417 0.0075457 0.0084097 0.0014007 0.98676 0.99158 3.0221e-006 1.2089e-005 0.15033 0.88622 0.89307 0.0014047 0.97473 0.5044 0.0018922 0.42571 1.8353 1.8342 16.0094 144.9623 0.00020073 -85.5899 0.54494
4.649 0.98808 5.4948e-005 3.8183 0.011984 6.0832e-005 0.0011595 0.23 0.00065928 0.23066 0.21275 0 0.032444 0.0389 0 1.2329 0.40459 0.12151 0.015386 8.1058 0.095963 0.00012068 0.79416 0.0075464 0.0084104 0.0014006 0.98676 0.99158 3.0219e-006 1.2087e-005 0.15034 0.88653 0.89321 0.0014046 0.97487 0.50457 0.0018921 0.42572 1.8361 1.8349 16.0093 144.9624 0.00020052 -85.5904 0.54594
4.65 0.98808 5.4947e-005 3.8183 0.011984 6.0845e-005 0.0011595 0.23001 0.00065928 0.23066 0.21275 0 0.032444 0.0389 0 1.233 0.40464 0.12153 0.015388 8.1076 0.095972 0.0001207 0.79415 0.007547 0.0084111 0.0014004 0.98676 0.99159 3.0216e-006 1.2086e-005 0.15034 0.88683 0.89334 0.0014046 0.97502 0.50474 0.001892 0.42574 1.8368 1.8356 16.0093 144.9624 0.0002003 -85.591 0.54694
4.651 0.98808 5.4947e-005 3.8183 0.011984 6.0858e-005 0.0011595 0.23001 0.00065928 0.23067 0.21276 0 0.032444 0.0389 0 1.2331 0.40469 0.12155 0.015389 8.1094 0.095982 0.00012071 0.79414 0.0075477 0.0084118 0.0014003 0.98676 0.99159 3.0213e-006 1.2085e-005 0.15035 0.88713 0.89348 0.0014045 0.97516 0.50491 0.0018919 0.42575 1.8375 1.8364 16.0093 144.9624 0.00020009 -85.5915 0.54794
4.652 0.98808 5.4947e-005 3.8183 0.011984 6.0871e-005 0.0011595 0.23002 0.00065928 0.23067 0.21276 0 0.032443 0.0389 0 1.2332 0.40473 0.12156 0.015391 8.1111 0.095992 0.00012072 0.79413 0.0075483 0.0084125 0.0014002 0.98676 0.99159 3.021e-006 1.2084e-005 0.15035 0.88743 0.89362 0.0014044 0.9753 0.50508 0.0018918 0.42576 1.8383 1.8371 16.0093 144.9624 0.00019987 -85.592 0.54894
4.653 0.98808 5.4947e-005 3.8183 0.011984 6.0884e-005 0.0011595 0.23002 0.00065928 0.23067 0.21276 0 0.032443 0.0389 0 1.2333 0.40478 0.12158 0.015393 8.1129 0.096001 0.00012074 0.79412 0.007549 0.0084132 0.0014001 0.98677 0.99159 3.0207e-006 1.2083e-005 0.15036 0.88773 0.89376 0.0014044 0.97544 0.50526 0.0018917 0.42578 1.839 1.8379 16.0093 144.9624 0.00019966 -85.5925 0.54994
4.654 0.98808 5.4947e-005 3.8183 0.011984 6.0897e-005 0.0011595 0.23002 0.00065928 0.23068 0.21277 0 0.032443 0.0389 0 1.2334 0.40483 0.12159 0.015394 8.1147 0.096011 0.00012075 0.79411 0.0075496 0.0084139 0.0014 0.98677 0.99159 3.0205e-006 1.2082e-005 0.15036 0.88803 0.89389 0.0014043 0.97558 0.50543 0.0018917 0.42579 1.8397 1.8386 16.0093 144.9625 0.00019945 -85.5931 0.55094
4.655 0.98808 5.4947e-005 3.8183 0.011984 6.091e-005 0.0011595 0.23003 0.00065928 0.23068 0.21277 0 0.032443 0.0389 0 1.2335 0.40487 0.12161 0.015396 8.1165 0.096021 0.00012077 0.7941 0.0075503 0.0084146 0.0013998 0.98677 0.99159 3.0202e-006 1.2081e-005 0.15037 0.88833 0.89403 0.0014042 0.97572 0.5056 0.0018916 0.4258 1.8405 1.8393 16.0093 144.9625 0.00019924 -85.5936 0.55194
4.656 0.98808 5.4947e-005 3.8183 0.011984 6.0923e-005 0.0011595 0.23003 0.00065928 0.23069 0.21277 0 0.032443 0.0389 0 1.2336 0.40492 0.12162 0.015397 8.1183 0.09603 0.00012078 0.79409 0.0075509 0.0084153 0.0013997 0.98677 0.99159 3.0199e-006 1.208e-005 0.15037 0.88863 0.89416 0.0014042 0.97586 0.50577 0.0018915 0.42582 1.8412 1.84 16.0092 144.9625 0.00019903 -85.5941 0.55294
4.657 0.98808 5.4947e-005 3.8183 0.011984 6.0936e-005 0.0011595 0.23004 0.00065928 0.23069 0.21278 0 0.032442 0.0389 0 1.2337 0.40497 0.12164 0.015399 8.1201 0.09604 0.00012079 0.79408 0.0075516 0.008416 0.0013996 0.98677 0.99159 3.0197e-006 1.2079e-005 0.15038 0.88892 0.8943 0.0014041 0.976 0.50594 0.0018914 0.42583 1.8419 1.8408 16.0092 144.9625 0.00019882 -85.5946 0.55394
4.658 0.98808 5.4947e-005 3.8183 0.011984 6.0949e-005 0.0011595 0.23004 0.00065928 0.23069 0.21278 0 0.032442 0.0389 0 1.2338 0.40501 0.12166 0.0154 8.1218 0.09605 0.00012081 0.79407 0.0075522 0.0084167 0.0013995 0.98677 0.99159 3.0194e-006 1.2077e-005 0.15038 0.88922 0.89443 0.001404 0.97614 0.50612 0.0018913 0.42584 1.8426 1.8415 16.0092 144.9625 0.00019861 -85.5951 0.55494
4.659 0.98808 5.4947e-005 3.8183 0.011984 6.0962e-005 0.0011595 0.23004 0.00065928 0.2307 0.21278 0 0.032442 0.0389 0 1.2339 0.40506 0.12167 0.015402 8.1236 0.096059 0.00012082 0.79406 0.0075529 0.0084174 0.0013994 0.98677 0.99159 3.0191e-006 1.2076e-005 0.15039 0.88951 0.89457 0.001404 0.97627 0.50629 0.0018912 0.42586 1.8433 1.8422 16.0092 144.9626 0.0001984 -85.5956 0.55594
4.66 0.98808 5.4947e-005 3.8183 0.011984 6.0975e-005 0.0011595 0.23005 0.00065928 0.2307 0.21279 0 0.032442 0.0389 0 1.234 0.40511 0.12169 0.015404 8.1254 0.096069 0.00012083 0.79405 0.0075535 0.0084181 0.0013993 0.98678 0.9916 3.0189e-006 1.2075e-005 0.15039 0.88981 0.8947 0.0014039 0.97641 0.50646 0.0018912 0.42587 1.8441 1.843 16.0092 144.9626 0.00019819 -85.5961 0.55694
4.661 0.98808 5.4947e-005 3.8183 0.011984 6.0988e-005 0.0011595 0.23005 0.00065928 0.23071 0.21279 0 0.032442 0.0389 0 1.2341 0.40515 0.1217 0.015405 8.1272 0.096079 0.00012085 0.79404 0.0075542 0.0084188 0.0013991 0.98678 0.9916 3.0186e-006 1.2074e-005 0.1504 0.8901 0.89483 0.0014039 0.97654 0.50663 0.0018911 0.42588 1.8448 1.8437 16.0092 144.9626 0.00019799 -85.5966 0.55794
4.662 0.98808 5.4947e-005 3.8183 0.011984 6.1001e-005 0.0011595 0.23005 0.00065928 0.23071 0.2128 0 0.032441 0.0389 0 1.2342 0.4052 0.12172 0.015407 8.129 0.096088 0.00012086 0.79403 0.0075548 0.0084195 0.001399 0.98678 0.9916 3.0183e-006 1.2073e-005 0.15041 0.89039 0.89497 0.0014038 0.97668 0.5068 0.001891 0.4259 1.8455 1.8444 16.0091 144.9626 0.00019778 -85.597 0.55894
4.663 0.98808 5.4947e-005 3.8183 0.011983 6.1014e-005 0.0011595 0.23006 0.00065928 0.23071 0.2128 0 0.032441 0.0389 0 1.2343 0.40525 0.12173 0.015408 8.1308 0.096098 0.00012087 0.79402 0.0075555 0.0084202 0.0013989 0.98678 0.9916 3.0181e-006 1.2072e-005 0.15041 0.89068 0.8951 0.0014037 0.97681 0.50697 0.0018909 0.42591 1.8462 1.8451 16.0091 144.9626 0.00019758 -85.5975 0.55994
4.664 0.98808 5.4946e-005 3.8183 0.011983 6.1027e-005 0.0011595 0.23006 0.00065928 0.23072 0.2128 0 0.032441 0.0389 0 1.2344 0.40529 0.12175 0.01541 8.1326 0.096108 0.00012089 0.79401 0.0075561 0.0084209 0.0013988 0.98678 0.9916 3.0178e-006 1.2071e-005 0.15042 0.89097 0.89523 0.0014037 0.97694 0.50715 0.0018909 0.42592 1.8469 1.8458 16.0091 144.9627 0.00019737 -85.598 0.56094
4.665 0.98808 5.4946e-005 3.8183 0.011983 6.104e-005 0.0011595 0.23007 0.00065928 0.23072 0.21281 0 0.032441 0.0389 0 1.2345 0.40534 0.12177 0.015411 8.1343 0.096117 0.0001209 0.794 0.0075568 0.0084216 0.0013987 0.98678 0.9916 3.0176e-006 1.207e-005 0.15042 0.89126 0.89536 0.0014036 0.97707 0.50732 0.0018908 0.42594 1.8476 1.8465 16.0091 144.9627 0.00019717 -85.5985 0.56194
4.666 0.98808 5.4946e-005 3.8183 0.011983 6.1053e-005 0.0011595 0.23007 0.00065928 0.23072 0.21281 0 0.032441 0.0389 0 1.2346 0.40539 0.12178 0.015413 8.1361 0.096127 0.00012092 0.79399 0.0075575 0.0084223 0.0013986 0.98678 0.9916 3.0173e-006 1.2069e-005 0.15043 0.89155 0.89549 0.0014036 0.9772 0.50749 0.0018907 0.42595 1.8483 1.8472 16.0091 144.9627 0.00019697 -85.5989 0.56294
4.667 0.98808 5.4946e-005 3.8183 0.011983 6.1066e-005 0.0011595 0.23007 0.00065928 0.23073 0.21281 0 0.032441 0.0389 0 1.2347 0.40543 0.1218 0.015414 8.1379 0.096137 0.00012093 0.79398 0.0075581 0.008423 0.0013985 0.98679 0.9916 3.0171e-006 1.2068e-005 0.15043 0.89184 0.89562 0.0014035 0.97733 0.50766 0.0018906 0.42596 1.8491 1.848 16.009 144.9627 0.00019677 -85.5994 0.56394
4.668 0.98808 5.4946e-005 3.8183 0.011983 6.1079e-005 0.0011595 0.23008 0.00065928 0.23073 0.21282 0 0.03244 0.0389 0 1.2347 0.40548 0.12181 0.015416 8.1397 0.096146 0.00012094 0.79397 0.0075588 0.0084237 0.0013984 0.98679 0.9916 3.0168e-006 1.2067e-005 0.15044 0.89212 0.89575 0.0014035 0.97746 0.50783 0.0018906 0.42598 1.8498 1.8487 16.009 144.9627 0.00019656 -85.5999 0.56494
4.669 0.98808 5.4946e-005 3.8183 0.011983 6.1092e-005 0.0011595 0.23008 0.00065928 0.23074 0.21282 0 0.03244 0.0389 0 1.2348 0.40553 0.12183 0.015418 8.1415 0.096156 0.00012096 0.79397 0.0075594 0.0084245 0.0013983 0.98679 0.9916 3.0166e-006 1.2066e-005 0.15044 0.89241 0.89588 0.0014034 0.97759 0.508 0.0018905 0.42599 1.8505 1.8494 16.009 144.9628 0.00019636 -85.6004 0.56594
4.67 0.98808 5.4946e-005 3.8183 0.011983 6.1105e-005 0.0011595 0.23008 0.00065928 0.23074 0.21282 0 0.03244 0.0389 0 1.2349 0.40557 0.12185 0.015419 8.1433 0.096165 0.00012097 0.79396 0.0075601 0.0084252 0.0013982 0.98679 0.9916 3.0163e-006 1.2065e-005 0.15045 0.89269 0.89601 0.0014033 0.97772 0.50817 0.0018904 0.426 1.8512 1.8501 16.009 144.9628 0.00019616 -85.6008 0.56694
4.671 0.98808 5.4946e-005 3.8183 0.011983 6.1118e-005 0.0011595 0.23009 0.00065928 0.23074 0.21283 0 0.03244 0.0389 0 1.235 0.40562 0.12186 0.015421 8.1451 0.096175 0.00012098 0.79395 0.0075607 0.0084259 0.001398 0.98679 0.99161 3.0161e-006 1.2064e-005 0.15045 0.89298 0.89613 0.0014033 0.97784 0.50834 0.0018903 0.42602 1.8519 1.8508 16.009 144.9628 0.00019597 -85.6013 0.56794
4.672 0.98808 5.4946e-005 3.8183 0.011983 6.1131e-005 0.0011595 0.23009 0.00065928 0.23075 0.21283 0 0.03244 0.0389 0 1.2351 0.40567 0.12188 0.015422 8.1469 0.096185 0.000121 0.79394 0.0075614 0.0084266 0.0013979 0.98679 0.99161 3.0158e-006 1.2063e-005 0.15046 0.89326 0.89626 0.0014032 0.97797 0.50852 0.0018903 0.42603 1.8526 1.8515 16.009 144.9628 0.00019577 -85.6017 0.56894
4.673 0.98808 5.4946e-005 3.8183 0.011983 6.1143e-005 0.0011595 0.2301 0.00065928 0.23075 0.21283 0 0.032439 0.0389 0 1.2352 0.40571 0.12189 0.015424 8.1486 0.096194 0.00012101 0.79393 0.007562 0.0084273 0.0013978 0.98679 0.99161 3.0156e-006 1.2062e-005 0.15046 0.89354 0.89639 0.0014032 0.97809 0.50869 0.0018902 0.42604 1.8533 1.8522 16.0089 144.9628 0.00019557 -85.6022 0.56994
4.674 0.98808 5.4946e-005 3.8183 0.011983 6.1156e-005 0.0011595 0.2301 0.00065928 0.23075 0.21284 0 0.032439 0.0389 0 1.2353 0.40576 0.12191 0.015425 8.1504 0.096204 0.00012102 0.79392 0.0075627 0.008428 0.0013977 0.9868 0.99161 3.0154e-006 1.2061e-005 0.15047 0.89382 0.89652 0.0014031 0.97821 0.50886 0.0018901 0.42606 1.854 1.8529 16.0089 144.9629 0.00019537 -85.6026 0.57094
4.675 0.98808 5.4946e-005 3.8183 0.011983 6.1169e-005 0.0011595 0.2301 0.00065928 0.23076 0.21284 0 0.032439 0.0389 0 1.2354 0.40581 0.12192 0.015427 8.1522 0.096214 0.00012104 0.79391 0.0075633 0.0084287 0.0013976 0.9868 0.99161 3.0151e-006 1.206e-005 0.15047 0.8941 0.89664 0.0014031 0.97834 0.50903 0.00189 0.42607 1.8546 1.8536 16.0089 144.9629 0.00019518 -85.6031 0.57194
4.676 0.98808 5.4946e-005 3.8183 0.011983 6.1182e-005 0.0011595 0.23011 0.00065928 0.23076 0.21285 0 0.032439 0.0389 0 1.2355 0.40585 0.12194 0.015429 8.154 0.096223 0.00012105 0.7939 0.007564 0.0084294 0.0013975 0.9868 0.99161 3.0149e-006 1.2059e-005 0.15048 0.89438 0.89677 0.001403 0.97846 0.5092 0.00189 0.42608 1.8553 1.8543 16.0089 144.9629 0.00019498 -85.6035 0.57294
4.677 0.98808 5.4946e-005 3.8183 0.011983 6.1195e-005 0.0011595 0.23011 0.00065928 0.23077 0.21285 0 0.032439 0.0389 0 1.2356 0.4059 0.12196 0.01543 8.1558 0.096233 0.00012106 0.79389 0.0075646 0.0084301 0.0013974 0.9868 0.99161 3.0147e-006 1.2059e-005 0.15048 0.89466 0.89689 0.001403 0.97858 0.50937 0.0018899 0.4261 1.856 1.855 16.0089 144.9629 0.00019479 -85.6039 0.57394
4.678 0.98808 5.4945e-005 3.8183 0.011983 6.1208e-005 0.0011595 0.23011 0.00065928 0.23077 0.21285 0 0.032438 0.0389 0 1.2357 0.40595 0.12197 0.015432 8.1576 0.096243 0.00012108 0.79388 0.0075653 0.0084308 0.0013973 0.9868 0.99161 3.0144e-006 1.2058e-005 0.15049 0.89494 0.89702 0.0014029 0.9787 0.50954 0.0018898 0.42611 1.8567 1.8557 16.0089 144.9629 0.0001946 -85.6044 0.57494
4.679 0.98808 5.4945e-005 3.8183 0.011983 6.1221e-005 0.0011595 0.23012 0.00065928 0.23077 0.21286 0 0.032438 0.0389 0 1.2358 0.40599 0.12199 0.015433 8.1594 0.096252 0.00012109 0.79387 0.0075659 0.0084315 0.0013972 0.9868 0.99161 3.0142e-006 1.2057e-005 0.15049 0.89522 0.89714 0.0014029 0.97882 0.50971 0.0018898 0.42612 1.8574 1.8563 16.0088 144.963 0.0001944 -85.6048 0.57594
4.68 0.98808 5.4945e-005 3.8183 0.011983 6.1234e-005 0.0011595 0.23012 0.00065928 0.23078 0.21286 0 0.032438 0.0389 0 1.2359 0.40604 0.122 0.015435 8.1612 0.096262 0.00012111 0.79386 0.0075666 0.0084322 0.0013971 0.9868 0.99161 3.014e-006 1.2056e-005 0.1505 0.89549 0.89726 0.0014028 0.97894 0.50988 0.0018897 0.42614 1.8581 1.857 16.0088 144.963 0.00019421 -85.6052 0.57694
4.681 0.98808 5.4945e-005 3.8183 0.011983 6.1247e-005 0.0011595 0.23013 0.00065928 0.23078 0.21286 0 0.032438 0.0389 0 1.236 0.40609 0.12202 0.015436 8.163 0.096272 0.00012112 0.79385 0.0075672 0.0084329 0.001397 0.98681 0.99161 3.0137e-006 1.2055e-005 0.1505 0.89577 0.89739 0.0014027 0.97906 0.51005 0.0018896 0.42615 1.8588 1.8577 16.0088 144.963 0.00019402 -85.6057 0.57794
4.682 0.98808 5.4945e-005 3.8183 0.011983 6.126e-005 0.0011595 0.23013 0.00065928 0.23078 0.21287 0 0.032438 0.0389 0 1.2361 0.40613 0.12203 0.015438 8.1648 0.096281 0.00012113 0.79384 0.0075679 0.0084336 0.0013969 0.98681 0.99162 3.0135e-006 1.2054e-005 0.15051 0.89604 0.89751 0.0014027 0.97918 0.51022 0.0018896 0.42616 1.8595 1.8584 16.0088 144.963 0.00019383 -85.6061 0.57894
4.683 0.98808 5.4945e-005 3.8183 0.011983 6.1273e-005 0.0011595 0.23013 0.00065928 0.23079 0.21287 0 0.032438 0.0389 0 1.2362 0.40618 0.12205 0.015439 8.1666 0.096291 0.00012115 0.79383 0.0075685 0.0084343 0.0013968 0.98681 0.99162 3.0133e-006 1.2053e-005 0.15051 0.89631 0.89763 0.0014026 0.97929 0.51039 0.0018895 0.42618 1.8601 1.8591 16.0088 144.963 0.00019364 -85.6065 0.57994
4.684 0.98808 5.4945e-005 3.8183 0.011983 6.1286e-005 0.0011596 0.23014 0.00065928 0.23079 0.21287 0 0.032437 0.0389 0 1.2363 0.40623 0.12207 0.015441 8.1683 0.0963 0.00012116 0.79382 0.0075692 0.008435 0.0013967 0.98681 0.99162 3.0131e-006 1.2052e-005 0.15052 0.89659 0.89775 0.0014026 0.97941 0.51056 0.0018894 0.42619 1.8608 1.8598 16.0087 144.9631 0.00019345 -85.6069 0.58094
4.685 0.98808 5.4945e-005 3.8183 0.011983 6.1299e-005 0.0011596 0.23014 0.00065928 0.23079 0.21288 0 0.032437 0.0389 0 1.2364 0.40627 0.12208 0.015443 8.1701 0.09631 0.00012117 0.79381 0.0075698 0.0084357 0.0013966 0.98681 0.99162 3.0128e-006 1.2051e-005 0.15052 0.89686 0.89787 0.0014025 0.97952 0.51073 0.0018894 0.4262 1.8615 1.8604 16.0087 144.9631 0.00019326 -85.6074 0.58194
4.686 0.98808 5.4945e-005 3.8183 0.011983 6.1312e-005 0.0011596 0.23014 0.00065928 0.2308 0.21288 0 0.032437 0.0389 0 1.2365 0.40632 0.1221 0.015444 8.1719 0.09632 0.00012119 0.7938 0.0075705 0.0084364 0.0013965 0.98681 0.99162 3.0126e-006 1.205e-005 0.15053 0.89713 0.898 0.0014025 0.97964 0.5109 0.0018893 0.42622 1.8622 1.8611 16.0087 144.9631 0.00019307 -85.6078 0.58294
4.687 0.98808 5.4945e-005 3.8183 0.011983 6.1325e-005 0.0011596 0.23015 0.00065928 0.2308 0.21288 0 0.032437 0.0389 0 1.2366 0.40637 0.12211 0.015446 8.1737 0.096329 0.0001212 0.79379 0.0075711 0.0084371 0.0013964 0.98681 0.99162 3.0124e-006 1.205e-005 0.15053 0.8974 0.89812 0.0014024 0.97975 0.51107 0.0018892 0.42623 1.8628 1.8618 16.0087 144.9631 0.00019288 -85.6082 0.58394
4.688 0.98808 5.4945e-005 3.8183 0.011983 6.1338e-005 0.0011596 0.23015 0.00065928 0.23081 0.21289 0 0.032437 0.0389 0 1.2367 0.40641 0.12213 0.015447 8.1755 0.096339 0.00012121 0.79378 0.0075718 0.0084378 0.0013963 0.98681 0.99162 3.0122e-006 1.2049e-005 0.15054 0.89767 0.89824 0.0014024 0.97986 0.51124 0.0018892 0.42624 1.8635 1.8625 16.0087 144.9631 0.0001927 -85.6086 0.58494
4.689 0.98808 5.4945e-005 3.8183 0.011983 6.1351e-005 0.0011596 0.23015 0.00065928 0.23081 0.21289 0 0.032436 0.0389 0 1.2368 0.40646 0.12214 0.015449 8.1773 0.096349 0.00012123 0.79377 0.0075724 0.0084385 0.0013962 0.98682 0.99162 3.012e-006 1.2048e-005 0.15054 0.89794 0.89836 0.0014023 0.97998 0.51141 0.0018891 0.42626 1.8642 1.8631 16.0086 144.9632 0.00019251 -85.609 0.58594
4.69 0.98808 5.4945e-005 3.8183 0.011983 6.1364e-005 0.0011596 0.23016 0.00065928 0.23081 0.21289 0 0.032436 0.0389 0 1.2369 0.40651 0.12216 0.01545 8.1791 0.096358 0.00012124 0.79376 0.0075731 0.0084392 0.0013962 0.98682 0.99162 3.0117e-006 1.2047e-005 0.15055 0.8982 0.89847 0.0014023 0.98009 0.51158 0.001889 0.42627 1.8648 1.8638 16.0086 144.9632 0.00019233 -85.6094 0.58694
4.691 0.98808 5.4944e-005 3.8183 0.011983 6.1377e-005 0.0011596 0.23016 0.00065928 0.23082 0.2129 0 0.032436 0.0389 0 1.237 0.40655 0.12218 0.015452 8.1809 0.096368 0.00012126 0.79375 0.0075737 0.0084399 0.0013961 0.98682 0.99162 3.0115e-006 1.2046e-005 0.15056 0.89847 0.89859 0.0014022 0.9802 0.51175 0.001889 0.42628 1.8655 1.8645 16.0086 144.9632 0.00019214 -85.6098 0.58794
4.692 0.98808 5.4944e-005 3.8183 0.011983 6.139e-005 0.0011596 0.23017 0.00065928 0.23082 0.2129 0 0.032436 0.0389 0 1.2371 0.4066 0.12219 0.015454 8.1827 0.096378 0.00012127 0.79374 0.0075744 0.0084406 0.001396 0.98682 0.99162 3.0113e-006 1.2045e-005 0.15056 0.89873 0.89871 0.0014022 0.98031 0.51192 0.0018889 0.4263 1.8662 1.8652 16.0086 144.9632 0.00019196 -85.6102 0.58894
4.693 0.98808 5.4944e-005 3.8183 0.011983 6.1403e-005 0.0011596 0.23017 0.00065928 0.23082 0.21291 0 0.032436 0.0389 0 1.2372 0.40665 0.12221 0.015455 8.1845 0.096387 0.00012128 0.79373 0.007575 0.0084413 0.0013959 0.98682 0.99162 3.0111e-006 1.2044e-005 0.15057 0.899 0.89883 0.0014021 0.98042 0.51209 0.0018888 0.42631 1.8668 1.8658 16.0086 144.9632 0.00019178 -85.6106 0.58994
4.694 0.98808 5.4944e-005 3.8183 0.011983 6.1416e-005 0.0011596 0.23017 0.00065928 0.23083 0.21291 0 0.032436 0.0389 0 1.2373 0.40669 0.12222 0.015457 8.1863 0.096397 0.0001213 0.79372 0.0075757 0.008442 0.0013958 0.98682 0.99162 3.0109e-006 1.2044e-005 0.15057 0.89926 0.89895 0.0014021 0.98053 0.51226 0.0018888 0.42632 1.8675 1.8665 16.0086 144.9633 0.00019159 -85.611 0.59094
4.695 0.98808 5.4944e-005 3.8183 0.011983 6.1429e-005 0.0011596 0.23018 0.00065928 0.23083 0.21291 0 0.032435 0.0389 0 1.2374 0.40674 0.12224 0.015458 8.1881 0.096406 0.00012131 0.79371 0.0075763 0.0084427 0.0013957 0.98682 0.99163 3.0107e-006 1.2043e-005 0.15058 0.89953 0.89906 0.001402 0.98063 0.51243 0.0018887 0.42634 1.8682 1.8671 16.0085 144.9633 0.00019141 -85.6114 0.59194
4.696 0.98808 5.4944e-005 3.8183 0.011983 6.1442e-005 0.0011596 0.23018 0.00065928 0.23084 0.21292 0 0.032435 0.0389 0 1.2375 0.40679 0.12225 0.01546 8.1899 0.096416 0.00012132 0.79371 0.007577 0.0084434 0.0013956 0.98682 0.99163 3.0105e-006 1.2042e-005 0.15058 0.89979 0.89918 0.001402 0.98074 0.5126 0.0018887 0.42635 1.8688 1.8678 16.0085 144.9633 0.00019123 -85.6117 0.59294
4.697 0.98808 5.4944e-005 3.8183 0.011983 6.1455e-005 0.0011596 0.23018 0.00065928 0.23084 0.21292 0 0.032435 0.0389 0 1.2376 0.40683 0.12227 0.015461 8.1917 0.096426 0.00012134 0.7937 0.0075776 0.0084441 0.0013955 0.98682 0.99163 3.0103e-006 1.2041e-005 0.15059 0.90005 0.8993 0.001402 0.98085 0.51277 0.0018886 0.42636 1.8695 1.8685 16.0085 144.9633 0.00019105 -85.6121 0.59394
4.698 0.98808 5.4944e-005 3.8183 0.011983 6.1468e-005 0.0011596 0.23019 0.00065928 0.23084 0.21292 0 0.032435 0.0389 0 1.2377 0.40688 0.12229 0.015463 8.1935 0.096435 0.00012135 0.79369 0.0075783 0.0084448 0.0013954 0.98683 0.99163 3.0101e-006 1.204e-005 0.15059 0.90031 0.89941 0.0014019 0.98095 0.51294 0.0018885 0.42638 1.8701 1.8691 16.0085 144.9633 0.00019087 -85.6125 0.59494
4.699 0.98808 5.4944e-005 3.8183 0.011983 6.1481e-005 0.0011596 0.23019 0.00065928 0.23085 0.21293 0 0.032435 0.0389 0 1.2378 0.40693 0.1223 0.015464 8.1953 0.096445 0.00012136 0.79368 0.0075789 0.0084455 0.0013953 0.98683 0.99163 3.0099e-006 1.2039e-005 0.1506 0.90057 0.89953 0.0014019 0.98106 0.51311 0.0018885 0.42639 1.8708 1.8698 16.0085 144.9634 0.00019069 -85.6129 0.59594
4.7 0.98808 5.4944e-005 3.8183 0.011983 6.1494e-005 0.0011596 0.23019 0.00065928 0.23085 0.21293 0 0.032434 0.0389 0 1.2379 0.40697 0.12232 0.015466 8.1971 0.096455 0.00012138 0.79367 0.0075796 0.0084462 0.0013953 0.98683 0.99163 3.0097e-006 1.2039e-005 0.1506 0.90083 0.89964 0.0014018 0.98116 0.51328 0.0018884 0.4264 1.8714 1.8704 16.0084 144.9634 0.00019051 -85.6133 0.59694
4.701 0.98808 5.4944e-005 3.8183 0.011983 6.1507e-005 0.0011596 0.2302 0.00065928 0.23085 0.21293 0 0.032434 0.0389 0 1.238 0.40702 0.12233 0.015468 8.1989 0.096464 0.00012139 0.79366 0.0075802 0.0084469 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.15061 0.90109 0.89975 0.0014018 0.98127 0.51345 0.0018884 0.42642 1.8721 1.8711 16.0084 144.9634 0.00019034 -85.6136 0.59794
4.702 0.98808 5.4944e-005 3.8183 0.011983 6.152e-005 0.0011596 0.2302 0.00065928 0.23086 0.21294 0 0.032434 0.0389 0 1.2381 0.40707 0.12235 0.015469 8.2007 0.096474 0.0001214 0.79365 0.0075809 0.0084476 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.15061 0.90135 0.89987 0.0014017 0.98137 0.51362 0.0018883 0.42643 1.8727 1.8717 16.0084 144.9634 0.00019016 -85.614 0.59894
4.703 0.98808 5.4944e-005 3.8183 0.011983 6.1533e-005 0.0011596 0.23021 0.00065928 0.23086 0.21294 0 0.032434 0.0389 0 1.2381 0.40711 0.12237 0.015471 8.2025 0.096483 0.00012142 0.79364 0.0075815 0.0084483 0.001395 0.98683 0.99163 3.0091e-006 1.2036e-005 0.15062 0.9016 0.89998 0.0014017 0.98147 0.51379 0.0018882 0.42644 1.8734 1.8724 16.0084 144.9634 0.00018998 -85.6144 0.59994
4.704 0.98808 5.4944e-005 3.8183 0.011983 6.1546e-005 0.0011596 0.23021 0.00065928 0.23086 0.21294 0 0.032434 0.0389 0 1.2382 0.40716 0.12238 0.015472 8.2043 0.096493 0.00012143 0.79363 0.0075822 0.008449 0.0013949 0.98683 0.99163 3.0089e-006 1.2036e-005 0.15062 0.90186 0.9001 0.0014016 0.98158 0.51396 0.0018882 0.42646 1.874 1.873 16.0084 144.9635 0.00018981 -85.6147 0.60094
4.705 0.98808 5.4943e-005 3.8183 0.011983 6.1559e-005 0.0011596 0.23021 0.00065928 0.23087 0.21295 0 0.032433 0.0389 0 1.2383 0.40721 0.1224 0.015474 8.2061 0.096503 0.00012145 0.79362 0.0075828 0.0084497 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.15063 0.90211 0.90021 0.0014016 0.98168 0.51413 0.0018881 0.42647 1.8747 1.8737 16.0083 144.9635 0.00018963 -85.6151 0.60194
4.706 0.98808 5.4943e-005 3.8183 0.011983 6.1572e-005 0.0011596 0.23022 0.00065928 0.23087 0.21295 0 0.032433 0.0389 0 1.2384 0.40725 0.12241 0.015475 8.2079 0.096512 0.00012146 0.79361 0.0075834 0.0084504 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.15063 0.90237 0.90032 0.0014015 0.98178 0.51429 0.0018881 0.42648 1.8753 1.8743 16.0083 144.9635 0.00018946 -85.6155 0.60294
4.707 0.98808 5.4943e-005 3.8183 0.011983 6.1585e-005 0.0011596 0.23022 0.00065928 0.23088 0.21295 0 0.032433 0.0389 0 1.2385 0.4073 0.12243 0.015477 8.2097 0.096522 0.00012147 0.7936 0.0075841 0.0084511 0.0013947 0.98684 0.99163 3.0083e-006 1.2033e-005 0.15064 0.90262 0.90043 0.0014015 0.98188 0.51446 0.001888 0.4265 1.876 1.875 16.0083 144.9635 0.00018928 -85.6158 0.60394
4.708 0.98808 5.4943e-005 3.8183 0.011983 6.1598e-005 0.0011596 0.23022 0.00065928 0.23088 0.21296 0 0.032433 0.0389 0 1.2386 0.40735 0.12244 0.015478 8.2115 0.096531 0.00012149 0.79359 0.0075847 0.0084518 0.0013946 0.98684 0.99163 3.0081e-006 1.2032e-005 0.15064 0.90288 0.90054 0.0014015 0.98198 0.51463 0.0018879 0.42651 1.8766 1.8756 16.0083 144.9635 0.00018911 -85.6162 0.60494
4.709 0.98808 5.4943e-005 3.8183 0.011983 6.1611e-005 0.0011596 0.23023 0.00065928 0.23088 0.21296 0 0.032433 0.0389 0 1.2387 0.40739 0.12246 0.01548 8.2133 0.096541 0.0001215 0.79358 0.0075854 0.0084525 0.0013945 0.98684 0.99164 3.008e-006 1.2032e-005 0.15065 0.90313 0.90065 0.0014014 0.98207 0.5148 0.0018879 0.42652 1.8772 1.8763 16.0083 144.9636 0.00018894 -85.6165 0.60594
4.71 0.98808 5.4943e-005 3.8183 0.011983 6.1624e-005 0.0011596 0.23023 0.00065928 0.23089 0.21296 0 0.032433 0.0389 0 1.2388 0.40744 0.12248 0.015482 8.2151 0.096551 0.00012151 0.79357 0.007586 0.0084532 0.0013944 0.98684 0.99164 3.0078e-006 1.2031e-005 0.15065 0.90338 0.90076 0.0014014 0.98217 0.51497 0.0018878 0.42654 1.8779 1.8769 16.0082 144.9636 0.00018877 -85.6169 0.60694
4.711 0.98808 5.4943e-005 3.8183 0.011983 6.1637e-005 0.0011596 0.23023 0.00065928 0.23089 0.21297 0 0.032432 0.0389 0 1.2389 0.40749 0.12249 0.015483 8.2169 0.09656 0.00012153 0.79356 0.0075867 0.0084539 0.0013943 0.98684 0.99164 3.0076e-006 1.203e-005 0.15066 0.90363 0.90087 0.0014013 0.98227 0.51514 0.0018878 0.42655 1.8785 1.8775 16.0082 144.9636 0.00018859 -85.6172 0.60794
4.712 0.98808 5.4943e-005 3.8183 0.011983 6.165e-005 0.0011596 0.23024 0.00065928 0.23089 0.21297 0 0.032432 0.0389 0 1.239 0.40753 0.12251 0.015485 8.2187 0.09657 0.00012154 0.79355 0.0075873 0.0084546 0.0013943 0.98684 0.99164 3.0074e-006 1.2029e-005 0.15066 0.90388 0.90098 0.0014013 0.98237 0.51531 0.0018877 0.42656 1.8791 1.8782 16.0082 144.9636 0.00018842 -85.6176 0.60894
4.713 0.98808 5.4943e-005 3.8183 0.011983 6.1663e-005 0.0011596 0.23024 0.00065928 0.2309 0.21297 0 0.032432 0.0389 0 1.2391 0.40758 0.12252 0.015486 8.2205 0.09658 0.00012155 0.79354 0.007588 0.0084553 0.0013942 0.98684 0.99164 3.0072e-006 1.2029e-005 0.15067 0.90413 0.90109 0.0014012 0.98246 0.51548 0.0018877 0.42658 1.8798 1.8788 16.0082 144.9636 0.00018825 -85.6179 0.60994
4.714 0.98808 5.4943e-005 3.8183 0.011983 6.1676e-005 0.0011596 0.23025 0.00065928 0.2309 0.21298 0 0.032432 0.0389 0 1.2392 0.40763 0.12254 0.015488 8.2223 0.096589 0.00012157 0.79353 0.0075886 0.008456 0.0013941 0.98684 0.99164 3.007e-006 1.2028e-005 0.15067 0.90438 0.9012 0.0014012 0.98256 0.51564 0.0018876 0.42659 1.8804 1.8794 16.0082 144.9637 0.00018808 -85.6182 0.61094
4.715 0.98808 5.4943e-005 3.8183 0.011983 6.1689e-005 0.0011596 0.23025 0.00065928 0.2309 0.21298 0 0.032432 0.0389 0 1.2393 0.40767 0.12255 0.015489 8.2241 0.096599 0.00012158 0.79352 0.0075893 0.0084567 0.001394 0.98684 0.99164 3.0069e-006 1.2027e-005 0.15068 0.90462 0.90131 0.0014012 0.98265 0.51581 0.0018876 0.4266 1.881 1.8801 16.0081 144.9637 0.00018792 -85.6186 0.61194
4.716 0.98808 5.4943e-005 3.8183 0.011983 6.1702e-005 0.0011596 0.23025 0.00065928 0.23091 0.21298 0 0.032431 0.0389 0 1.2394 0.40772 0.12257 0.015491 8.2259 0.096608 0.00012159 0.79351 0.0075899 0.0084574 0.0013939 0.98685 0.99164 3.0067e-006 1.2027e-005 0.15068 0.90487 0.90142 0.0014011 0.98275 0.51598 0.0018875 0.42662 1.8817 1.8807 16.0081 144.9637 0.00018775 -85.6189 0.61294
4.717 0.98808 5.4943e-005 3.8183 0.011983 6.1715e-005 0.0011596 0.23026 0.00065928 0.23091 0.21299 0 0.032431 0.0389 0 1.2395 0.40777 0.12259 0.015492 8.2277 0.096618 0.00012161 0.7935 0.0075906 0.008458 0.0013938 0.98685 0.99164 3.0065e-006 1.2026e-005 0.15069 0.90511 0.90153 0.0014011 0.98284 0.51615 0.0018874 0.42663 1.8823 1.8813 16.0081 144.9637 0.00018758 -85.6193 0.61394
4.718 0.98808 5.4943e-005 3.8183 0.011983 6.1728e-005 0.0011596 0.23026 0.00065928 0.23091 0.21299 0 0.032431 0.0389 0 1.2396 0.40781 0.1226 0.015494 8.2295 0.096628 0.00012162 0.79349 0.0075912 0.0084587 0.0013938 0.98685 0.99164 3.0063e-006 1.2025e-005 0.15069 0.90536 0.90163 0.001401 0.98293 0.51632 0.0018874 0.42664 1.8829 1.882 16.0081 144.9637 0.00018741 -85.6196 0.61494
4.719 0.98808 5.4942e-005 3.8183 0.011983 6.1741e-005 0.0011596 0.23026 0.00065928 0.23092 0.21299 0 0.032431 0.0389 0 1.2397 0.40786 0.12262 0.015496 8.2313 0.096637 0.00012164 0.79348 0.0075919 0.0084594 0.0013937 0.98685 0.99164 3.0061e-006 1.2024e-005 0.1507 0.9056 0.90174 0.001401 0.98303 0.51649 0.0018873 0.42666 1.8835 1.8826 16.0081 144.9638 0.00018725 -85.6199 0.61594
4.72 0.98808 5.4942e-005 3.8183 0.011983 6.1753e-005 0.0011596 0.23027 0.00065928 0.23092 0.213 0 0.032431 0.0389 0 1.2398 0.40791 0.12263 0.015497 8.2331 0.096647 0.00012165 0.79347 0.0075925 0.0084601 0.0013936 0.98685 0.99164 3.006e-006 1.2024e-005 0.1507 0.90585 0.90185 0.001401 0.98312 0.51666 0.0018873 0.42667 1.8842 1.8832 16.008 144.9638 0.00018708 -85.6202 0.61694
4.721 0.98808 5.4942e-005 3.8183 0.011983 6.1766e-005 0.0011597 0.23027 0.00065928 0.23093 0.213 0 0.032431 0.0389 0 1.2399 0.40795 0.12265 0.015499 8.2349 0.096656 0.00012166 0.79347 0.0075932 0.0084608 0.0013936 0.98685 0.99164 3.0058e-006 1.2023e-005 0.15071 0.90609 0.90195 0.0014009 0.98321 0.51682 0.0018872 0.42668 1.8848 1.8838 16.008 144.9638 0.00018692 -85.6206 0.61794
4.722 0.98808 5.4942e-005 3.8183 0.011983 6.1779e-005 0.0011597 0.23027 0.00065928 0.23093 0.213 0 0.03243 0.0389 0 1.24 0.408 0.12266 0.0155 8.2367 0.096666 0.00012168 0.79346 0.0075938 0.0084615 0.0013935 0.98685 0.99164 3.0056e-006 1.2022e-005 0.15072 0.90633 0.90206 0.0014009 0.9833 0.51699 0.0018872 0.4267 1.8854 1.8845 16.008 144.9638 0.00018675 -85.6209 0.61894
4.723 0.98808 5.4942e-005 3.8183 0.011983 6.1792e-005 0.0011597 0.23028 0.00065928 0.23093 0.21301 0 0.03243 0.0389 0 1.2401 0.40805 0.12268 0.015502 8.2385 0.096676 0.00012169 0.79345 0.0075945 0.0084622 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.15072 0.90657 0.90216 0.0014008 0.98339 0.51716 0.0018871 0.42671 1.886 1.8851 16.008 144.9638 0.00018659 -85.6212 0.61994
4.724 0.98808 5.4942e-005 3.8183 0.011983 6.1805e-005 0.0011597 0.23028 0.00065928 0.23094 0.21301 0 0.03243 0.0389 0 1.2402 0.40809 0.1227 0.015503 8.2404 0.096685 0.0001217 0.79344 0.0075951 0.0084629 0.0013933 0.98685 0.99165 3.0053e-006 1.2021e-005 0.15073 0.90681 0.90227 0.0014008 0.98348 0.51733 0.0018871 0.42672 1.8866 1.8857 16.0079 144.9639 0.00018642 -85.6215 0.62094
4.725 0.98808 5.4942e-005 3.8183 0.011983 6.1818e-005 0.0011597 0.23029 0.00065928 0.23094 0.21301 0 0.03243 0.0389 0 1.2403 0.40814 0.12271 0.015505 8.2422 0.096695 0.00012172 0.79343 0.0075958 0.0084636 0.0013932 0.98685 0.99165 3.0051e-006 1.202e-005 0.15073 0.90705 0.90237 0.0014008 0.98357 0.5175 0.001887 0.42674 1.8872 1.8863 16.0079 144.9639 0.00018626 -85.6219 0.62194
4.726 0.98808 5.4942e-005 3.8183 0.011983 6.1831e-005 0.0011597 0.23029 0.00065928 0.23094 0.21302 0 0.03243 0.0389 0 1.2404 0.40819 0.12273 0.015507 8.244 0.096704 0.00012173 0.79342 0.0075964 0.0084643 0.0013932 0.98685 0.99165 3.0049e-006 1.202e-005 0.15074 0.90729 0.90248 0.0014007 0.98366 0.51766 0.001887 0.42675 1.8879 1.8869 16.0079 144.9639 0.0001861 -85.6222 0.62294
4.727 0.98808 5.4942e-005 3.8183 0.011982 6.1844e-005 0.0011597 0.23029 0.00065928 0.23095 0.21302 0 0.03243 0.0389 0 1.2405 0.40823 0.12274 0.015508 8.2458 0.096714 0.00012174 0.79341 0.007597 0.008465 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.15074 0.90753 0.90258 0.0014007 0.98374 0.51783 0.0018869 0.42676 1.8885 1.8875 16.0079 144.9639 0.00018594 -85.6225 0.62394
4.728 0.98808 5.4942e-005 3.8183 0.011982 6.1857e-005 0.0011597 0.2303 0.00065928 0.23095 0.21303 0 0.032429 0.0389 0 1.2406 0.40828 0.12276 0.01551 8.2476 0.096724 0.00012176 0.7934 0.0075977 0.0084657 0.001393 0.98686 0.99165 3.0046e-006 1.2018e-005 0.15075 0.90777 0.90268 0.0014006 0.98383 0.518 0.0018869 0.42678 1.8891 1.8881 16.0079 144.964 0.00018578 -85.6228 0.62494
4.729 0.98808 5.4942e-005 3.8183 0.011982 6.187e-005 0.0011597 0.2303 0.00065928 0.23095 0.21303 0 0.032429 0.0389 0 1.2407 0.40833 0.12277 0.015511 8.2494 0.096733 0.00012177 0.79339 0.0075983 0.0084664 0.001393 0.98686 0.99165 3.0045e-006 1.2018e-005 0.15075 0.908 0.90279 0.0014006 0.98392 0.51817 0.0018868 0.42679 1.8897 1.8888 16.0078 144.964 0.00018562 -85.6231 0.62594
4.73 0.98808 5.4942e-005 3.8183 0.011982 6.1883e-005 0.0011597 0.2303 0.00065928 0.23096 0.21303 0 0.032429 0.0389 0 1.2408 0.40837 0.12279 0.015513 8.2512 0.096743 0.00012178 0.79338 0.007599 0.0084671 0.0013929 0.98686 0.99165 3.0043e-006 1.2017e-005 0.15076 0.90824 0.90289 0.0014006 0.984 0.51833 0.0018868 0.4268 1.8903 1.8894 16.0078 144.964 0.00018546 -85.6234 0.62694
4.731 0.98808 5.4942e-005 3.8183 0.011982 6.1896e-005 0.0011597 0.23031 0.00065928 0.23096 0.21304 0 0.032429 0.0389 0 1.2409 0.40842 0.12281 0.015514 8.253 0.096752 0.0001218 0.79337 0.0075996 0.0084678 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.15076 0.90848 0.90299 0.0014005 0.98409 0.5185 0.0018867 0.42682 1.8909 1.89 16.0078 144.964 0.0001853 -85.6237 0.62794
4.732 0.98808 5.4941e-005 3.8183 0.011982 6.1909e-005 0.0011597 0.23031 0.00065928 0.23096 0.21304 0 0.032429 0.0389 0 1.241 0.40847 0.12282 0.015516 8.2548 0.096762 0.00012181 0.79336 0.0076003 0.0084685 0.0013928 0.98686 0.99165 3.004e-006 1.2016e-005 0.15077 0.90871 0.90309 0.0014005 0.98417 0.51867 0.0018867 0.42683 1.8915 1.8906 16.0078 144.964 0.00018514 -85.624 0.62894
4.733 0.98808 5.4941e-005 3.8183 0.011982 6.1922e-005 0.0011597 0.23031 0.00065928 0.23097 0.21304 0 0.032428 0.0389 0 1.2411 0.40851 0.12284 0.015517 8.2566 0.096772 0.00012182 0.79335 0.0076009 0.0084692 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.15077 0.90894 0.9032 0.0014005 0.98426 0.51884 0.0018866 0.42684 1.8921 1.8912 16.0078 144.9641 0.00018498 -85.6243 0.62994
4.734 0.98808 5.4941e-005 3.8183 0.011982 6.1935e-005 0.0011597 0.23032 0.00065928 0.23097 0.21305 0 0.032428 0.0389 0 1.2412 0.40856 0.12285 0.015519 8.2584 0.096781 0.00012184 0.79334 0.0076016 0.0084699 0.0013926 0.98686 0.99165 3.0037e-006 1.2015e-005 0.15078 0.90918 0.9033 0.0014004 0.98434 0.519 0.0018866 0.42686 1.8927 1.8918 16.0077 144.9641 0.00018482 -85.6246 0.63094
4.735 0.98808 5.4941e-005 3.8183 0.011982 6.1948e-005 0.0011597 0.23032 0.00065928 0.23098 0.21305 0 0.032428 0.0389 0 1.2413 0.40861 0.12287 0.01552 8.2603 0.096791 0.00012185 0.79333 0.0076022 0.0084706 0.0013925 0.98686 0.99165 3.0035e-006 1.2014e-005 0.15078 0.90941 0.9034 0.0014004 0.98443 0.51917 0.0018865 0.42687 1.8933 1.8924 16.0077 144.9641 0.00018467 -85.6249 0.63194
4.736 0.98808 5.4941e-005 3.8183 0.011982 6.1961e-005 0.0011597 0.23032 0.00065928 0.23098 0.21305 0 0.032428 0.0389 0 1.2413 0.40865 0.12288 0.015522 8.2621 0.0968 0.00012187 0.79332 0.0076029 0.0084713 0.0013925 0.98686 0.99165 3.0033e-006 1.2013e-005 0.15079 0.90964 0.9035 0.0014003 0.98451 0.51934 0.0018865 0.42688 1.8939 1.893 16.0077 144.9641 0.00018451 -85.6252 0.63294
4.737 0.98808 5.4941e-005 3.8183 0.011982 6.1974e-005 0.0011597 0.23033 0.00065928 0.23098 0.21306 0 0.032428 0.0389 0 1.2414 0.4087 0.1229 0.015524 8.2639 0.09681 0.00012188 0.79331 0.0076035 0.008472 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.15079 0.90987 0.9036 0.0014003 0.98459 0.51951 0.0018865 0.4269 1.8945 1.8936 16.0077 144.9641 0.00018436 -85.6255 0.63394
4.738 0.98808 5.4941e-005 3.8183 0.011982 6.1987e-005 0.0011597 0.23033 0.00065928 0.23099 0.21306 0 0.032428 0.0389 0 1.2415 0.40874 0.12292 0.015525 8.2657 0.096819 0.00012189 0.7933 0.0076042 0.0084727 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.1508 0.9101 0.9037 0.0014003 0.98467 0.51967 0.0018864 0.42691 1.8951 1.8942 16.0076 144.9642 0.0001842 -85.6258 0.63494
4.739 0.98808 5.4941e-005 3.8183 0.011982 6.2e-005 0.0011597 0.23033 0.00065928 0.23099 0.21306 0 0.032427 0.0389 0 1.2416 0.40879 0.12293 0.015527 8.2675 0.096829 0.00012191 0.79329 0.0076048 0.0084734 0.0013923 0.98687 0.99165 3.0029e-006 1.2011e-005 0.1508 0.91033 0.9038 0.0014002 0.98475 0.51984 0.0018864 0.42692 1.8957 1.8948 16.0076 144.9642 0.00018405 -85.6261 0.63594
4.74 0.98808 5.4941e-005 3.8183 0.011982 6.2013e-005 0.0011597 0.23034 0.00065928 0.23099 0.21307 0 0.032427 0.0389 0 1.2417 0.40884 0.12295 0.015528 8.2693 0.096839 0.00012192 0.79328 0.0076054 0.0084741 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.15081 0.91056 0.9039 0.0014002 0.98483 0.52001 0.0018863 0.42693 1.8963 1.8954 16.0076 144.9642 0.00018389 -85.6263 0.63694
4.741 0.98808 5.4941e-005 3.8183 0.011982 6.2026e-005 0.0011597 0.23034 0.00065928 0.231 0.21307 0 0.032427 0.0389 0 1.2418 0.40888 0.12296 0.01553 8.2711 0.096848 0.00012193 0.79327 0.0076061 0.0084748 0.0013922 0.98687 0.99166 3.0026e-006 1.201e-005 0.15081 0.91079 0.90399 0.0014002 0.98492 0.52018 0.0018863 0.42695 1.8969 1.896 16.0076 144.9642 0.00018374 -85.6266 0.63794
4.742 0.98808 5.4941e-005 3.8183 0.011982 6.2039e-005 0.0011597 0.23035 0.00065928 0.231 0.21307 0 0.032427 0.0389 0 1.2419 0.40893 0.12298 0.015531 8.2729 0.096858 0.00012195 0.79326 0.0076067 0.0084755 0.0013921 0.98687 0.99166 3.0024e-006 1.201e-005 0.15082 0.91102 0.90409 0.0014001 0.98499 0.52034 0.0018862 0.42696 1.8975 1.8966 16.0076 144.9642 0.00018359 -85.6269 0.63894
4.743 0.98808 5.4941e-005 3.8183 0.011982 6.2052e-005 0.0011597 0.23035 0.00065928 0.231 0.21308 0 0.032427 0.0389 0 1.242 0.40898 0.12299 0.015533 8.2748 0.096867 0.00012196 0.79325 0.0076074 0.0084762 0.001392 0.98687 0.99166 3.0023e-006 1.2009e-005 0.15082 0.91124 0.90419 0.0014001 0.98507 0.52051 0.0018862 0.42697 1.8981 1.8972 16.0075 144.9643 0.00018343 -85.6272 0.63994
4.744 0.98808 5.4941e-005 3.8183 0.011982 6.2065e-005 0.0011597 0.23035 0.00065928 0.23101 0.21308 0 0.032427 0.0389 0 1.2421 0.40902 0.12301 0.015534 8.2766 0.096877 0.00012197 0.79325 0.007608 0.0084769 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.15083 0.91147 0.90429 0.0014001 0.98515 0.52068 0.0018861 0.42699 1.8986 1.8978 16.0075 144.9643 0.00018328 -85.6275 0.64094
4.745 0.98808 5.4941e-005 3.8183 0.011982 6.2078e-005 0.0011597 0.23036 0.00065928 0.23101 0.21308 0 0.032426 0.0389 0 1.2422 0.40907 0.12303 0.015536 8.2784 0.096887 0.00012199 0.79324 0.0076087 0.0084776 0.0013919 0.98687 0.99166 3.002e-006 1.2008e-005 0.15083 0.91169 0.90439 0.0014 0.98523 0.52084 0.0018861 0.427 1.8992 1.8983 16.0075 144.9643 0.00018313 -85.6277 0.64194
4.746 0.98808 5.494e-005 3.8183 0.011982 6.2091e-005 0.0011597 0.23036 0.00065928 0.23101 0.21309 0 0.032426 0.0389 0 1.2423 0.40912 0.12304 0.015538 8.2802 0.096896 0.000122 0.79323 0.0076093 0.0084783 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.15084 0.91192 0.90448 0.0014 0.98531 0.52101 0.001886 0.42701 1.8998 1.8989 16.0075 144.9643 0.00018298 -85.628 0.64294
4.747 0.98808 5.494e-005 3.8183 0.011982 6.2104e-005 0.0011597 0.23036 0.00065928 0.23102 0.21309 0 0.032426 0.0389 0 1.2424 0.40916 0.12306 0.015539 8.282 0.096906 0.00012201 0.79322 0.00761 0.0084789 0.0013917 0.98687 0.99166 3.0017e-006 1.2007e-005 0.15084 0.91214 0.90458 0.0014 0.98539 0.52118 0.001886 0.42703 1.9004 1.8995 16.0074 144.9643 0.00018283 -85.6283 0.64394
4.748 0.98808 5.494e-005 3.8183 0.011982 6.2117e-005 0.0011597 0.23037 0.00065928 0.23102 0.21309 0 0.032426 0.0389 0 1.2425 0.40921 0.12307 0.015541 8.2838 0.096915 0.00012203 0.79321 0.0076106 0.0084796 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.15085 0.91236 0.90467 0.0013999 0.98546 0.52134 0.001886 0.42704 1.901 1.9001 16.0074 144.9644 0.00018268 -85.6286 0.64494
4.749 0.98808 5.494e-005 3.8183 0.011982 6.213e-005 0.0011597 0.23037 0.00065928 0.23102 0.2131 0 0.032426 0.0389 0 1.2426 0.40926 0.12309 0.015542 8.2857 0.096925 0.00012204 0.7932 0.0076113 0.0084803 0.0013916 0.98687 0.99166 3.0014e-006 1.2006e-005 0.15085 0.91259 0.90477 0.0013999 0.98554 0.52151 0.0018859 0.42705 1.9016 1.9007 16.0074 144.9644 0.00018253 -85.6288 0.64594
4.75 0.98808 5.494e-005 3.8183 0.011982 6.2143e-005 0.0011597 0.23037 0.00065928 0.23103 0.2131 0 0.032425 0.0389 0 1.2427 0.4093 0.1231 0.015544 8.2875 0.096934 0.00012205 0.79319 0.0076119 0.008481 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.15086 0.91281 0.90487 0.0013999 0.98561 0.52168 0.0018859 0.42707 1.9021 1.9013 16.0074 144.9644 0.00018238 -85.6291 0.64694
4.751 0.98808 5.494e-005 3.8183 0.011982 6.2156e-005 0.0011597 0.23038 0.00065928 0.23103 0.2131 0 0.032425 0.0389 0 1.2428 0.40935 0.12312 0.015545 8.2893 0.096944 0.00012207 0.79318 0.0076125 0.0084817 0.0013915 0.98688 0.99166 3.0011e-006 1.2004e-005 0.15086 0.91303 0.90496 0.0013999 0.98569 0.52184 0.0018858 0.42708 1.9027 1.9018 16.0074 144.9644 0.00018223 -85.6294 0.64794
4.752 0.98808 5.494e-005 3.8183 0.011982 6.2169e-005 0.0011597 0.23038 0.00065928 0.23103 0.21311 0 0.032425 0.0389 0 1.2429 0.4094 0.12314 0.015547 8.2911 0.096954 0.00012208 0.79317 0.0076132 0.0084824 0.0013915 0.98688 0.99166 3.001e-006 1.2004e-005 0.15087 0.91325 0.90506 0.0013998 0.98576 0.52201 0.0018858 0.42709 1.9033 1.9024 16.0073 144.9644 0.00018209 -85.6296 0.64894
4.753 0.98808 5.494e-005 3.8183 0.011982 6.2182e-005 0.0011597 0.23038 0.00065928 0.23104 0.21311 0 0.032425 0.0389 0 1.243 0.40944 0.12315 0.015548 8.2929 0.096963 0.0001221 0.79316 0.0076138 0.0084831 0.0013914 0.98688 0.99166 3.0008e-006 1.2003e-005 0.15087 0.91347 0.90515 0.0013998 0.98584 0.52218 0.0018857 0.42711 1.9039 1.903 16.0073 144.9645 0.00018194 -85.6299 0.64994
4.754 0.98808 5.494e-005 3.8183 0.011982 6.2195e-005 0.0011597 0.23039 0.00065928 0.23104 0.21311 0 0.032425 0.0389 0 1.2431 0.40949 0.12317 0.01555 8.2947 0.096973 0.00012211 0.79315 0.0076145 0.0084838 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.15088 0.91369 0.90524 0.0013997 0.98591 0.52234 0.0018857 0.42712 1.9045 1.9036 16.0073 144.9645 0.00018179 -85.6301 0.65094
4.755 0.98808 5.494e-005 3.8183 0.011982 6.2208e-005 0.0011597 0.23039 0.00065928 0.23105 0.21312 0 0.032425 0.0389 0 1.2432 0.40954 0.12318 0.015552 8.2966 0.096982 0.00012212 0.79314 0.0076151 0.0084845 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.15088 0.91391 0.90534 0.0013997 0.98598 0.52251 0.0018857 0.42713 1.905 1.9042 16.0073 144.9645 0.00018165 -85.6304 0.65194
4.756 0.98808 5.494e-005 3.8183 0.011982 6.2221e-005 0.0011597 0.23039 0.00065928 0.23105 0.21312 0 0.032424 0.0389 0 1.2433 0.40958 0.1232 0.015553 8.2984 0.096992 0.00012214 0.79313 0.0076158 0.0084852 0.0013912 0.98688 0.99166 3.0004e-006 1.2002e-005 0.15089 0.91412 0.90543 0.0013997 0.98606 0.52267 0.0018856 0.42715 1.9056 1.9047 16.0072 144.9645 0.0001815 -85.6307 0.65294
4.757 0.98808 5.494e-005 3.8183 0.011982 6.2234e-005 0.0011598 0.2304 0.00065928 0.23105 0.21312 0 0.032424 0.0389 0 1.2434 0.40963 0.12321 0.015555 8.3002 0.097001 0.00012215 0.79312 0.0076164 0.0084859 0.0013911 0.98688 0.99166 3.0003e-006 1.2001e-005 0.15089 0.91434 0.90552 0.0013996 0.98613 0.52284 0.0018856 0.42716 1.9062 1.9053 16.0072 144.9645 0.00018136 -85.6309 0.65394
4.758 0.98808 5.494e-005 3.8183 0.011982 6.2247e-005 0.0011598 0.2304 0.00065928 0.23106 0.21313 0 0.032424 0.0389 0 1.2435 0.40968 0.12323 0.015556 8.302 0.097011 0.00012216 0.79311 0.0076171 0.0084866 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.1509 0.91456 0.90562 0.0013996 0.9862 0.52301 0.0018855 0.42717 1.9067 1.9059 16.0072 144.9646 0.00018121 -85.6312 0.65494
4.759 0.98808 5.494e-005 3.8183 0.011982 6.226e-005 0.0011598 0.2304 0.00065928 0.23106 0.21313 0 0.032424 0.0389 0 1.2436 0.40972 0.12325 0.015558 8.3038 0.09702 0.00012218 0.7931 0.0076177 0.0084873 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.15091 0.91477 0.90571 0.0013996 0.98627 0.52317 0.0018855 0.42718 1.9073 1.9064 16.0072 144.9646 0.00018107 -85.6314 0.65594
4.76 0.98808 5.4939e-005 3.8183 0.011982 6.2273e-005 0.0011598 0.23041 0.00065928 0.23106 0.21313 0 0.032424 0.0389 0 1.2437 0.40977 0.12326 0.015559 8.3057 0.09703 0.00012219 0.79309 0.0076183 0.008488 0.001391 0.98688 0.99166 2.9999e-006 1.1999e-005 0.15091 0.91499 0.9058 0.0013996 0.98634 0.52334 0.0018855 0.4272 1.9079 1.907 16.0071 144.9646 0.00018093 -85.6317 0.65694
4.761 0.98808 5.4939e-005 3.8183 0.011982 6.2286e-005 0.0011598 0.23041 0.00065928 0.23107 0.21314 0 0.032424 0.0389 0 1.2438 0.40982 0.12328 0.015561 8.3075 0.09704 0.0001222 0.79308 0.007619 0.0084887 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.15092 0.9152 0.90589 0.0013995 0.98641 0.5235 0.0018854 0.42721 1.9084 1.9076 16.0071 144.9646 0.00018078 -85.6319 0.65794
4.762 0.98808 5.4939e-005 3.8183 0.011982 6.2298e-005 0.0011598 0.23041 0.00065928 0.23107 0.21314 0 0.032423 0.0389 0 1.2439 0.40986 0.12329 0.015562 8.3093 0.097049 0.00012222 0.79307 0.0076196 0.0084894 0.0013909 0.98688 0.99167 2.9996e-006 1.1998e-005 0.15092 0.91541 0.90598 0.0013995 0.98648 0.52367 0.0018854 0.42722 1.909 1.9081 16.0071 144.9646 0.00018064 -85.6322 0.65894
4.763 0.98808 5.4939e-005 3.8183 0.011982 6.2311e-005 0.0011598 0.23042 0.00065928 0.23107 0.21314 0 0.032423 0.0389 0 1.244 0.40991 0.12331 0.015564 8.3111 0.097059 0.00012223 0.79306 0.0076203 0.0084901 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.15093 0.91563 0.90607 0.0013995 0.98655 0.52384 0.0018853 0.42724 1.9096 1.9087 16.0071 144.9647 0.0001805 -85.6324 0.65994
4.764 0.98808 5.4939e-005 3.8183 0.011982 6.2324e-005 0.0011598 0.23042 0.00065928 0.23108 0.21314 0 0.032423 0.0389 0 1.2441 0.40996 0.12332 0.015566 8.3129 0.097068 0.00012224 0.79305 0.0076209 0.0084908 0.0013907 0.98689 0.99167 2.9994e-006 1.1997e-005 0.15093 0.91584 0.90617 0.0013994 0.98662 0.524 0.0018853 0.42725 1.9101 1.9093 16.0071 144.9647 0.00018036 -85.6327 0.66094
4.765 0.98808 5.4939e-005 3.8183 0.011982 6.2337e-005 0.0011598 0.23043 0.00065928 0.23108 0.21315 0 0.032423 0.0389 0 1.2442 0.41 0.12334 0.015567 8.3148 0.097078 0.00012226 0.79304 0.0076216 0.0084914 0.0013907 0.98689 0.99167 2.9992e-006 1.1997e-005 0.15094 0.91605 0.90626 0.0013994 0.98669 0.52417 0.0018853 0.42726 1.9107 1.9098 16.007 144.9647 0.00018022 -85.6329 0.66194
4.766 0.98808 5.4939e-005 3.8183 0.011982 6.235e-005 0.0011598 0.23043 0.00065928 0.23108 0.21315 0 0.032423 0.0389 0 1.2443 0.41005 0.12336 0.015569 8.3166 0.097087 0.00012227 0.79303 0.0076222 0.0084921 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.15094 0.91626 0.90635 0.0013994 0.98676 0.52433 0.0018852 0.42728 1.9112 1.9104 16.007 144.9647 0.00018008 -85.6331 0.66294
4.767 0.98808 5.4939e-005 3.8183 0.011982 6.2363e-005 0.0011598 0.23043 0.00065928 0.23109 0.21315 0 0.032422 0.0389 0 1.2444 0.4101 0.12337 0.01557 8.3184 0.097097 0.00012228 0.79303 0.0076228 0.0084928 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.15095 0.91647 0.90644 0.0013993 0.98683 0.5245 0.0018852 0.42729 1.9118 1.911 16.007 144.9647 0.00017994 -85.6334 0.66394
4.768 0.98808 5.4939e-005 3.8183 0.011982 6.2376e-005 0.0011598 0.23044 0.00065928 0.23109 0.21316 0 0.032422 0.0389 0 1.2445 0.41014 0.12339 0.015572 8.3202 0.097107 0.0001223 0.79302 0.0076235 0.0084935 0.0013905 0.98689 0.99167 2.9989e-006 1.1995e-005 0.15095 0.91668 0.90652 0.0013993 0.98689 0.52466 0.0018851 0.4273 1.9124 1.9115 16.007 144.9648 0.0001798 -85.6336 0.66494
4.769 0.98808 5.4939e-005 3.8183 0.011982 6.2389e-005 0.0011598 0.23044 0.00065928 0.23109 0.21316 0 0.032422 0.0389 0 1.2445 0.41019 0.1234 0.015573 8.3221 0.097116 0.00012231 0.79301 0.0076241 0.0084942 0.0013905 0.98689 0.99167 2.9987e-006 1.1995e-005 0.15096 0.91689 0.90661 0.0013993 0.98696 0.52483 0.0018851 0.42732 1.9129 1.9121 16.0069 144.9648 0.00017966 -85.6338 0.66594
4.77 0.98808 5.4939e-005 3.8183 0.011982 6.2402e-005 0.0011598 0.23044 0.00065928 0.2311 0.21316 0 0.032422 0.0389 0 1.2446 0.41024 0.12342 0.015575 8.3239 0.097126 0.00012232 0.793 0.0076248 0.0084949 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.15096 0.9171 0.9067 0.0013993 0.98703 0.52499 0.0018851 0.42733 1.9135 1.9126 16.0069 144.9648 0.00017952 -85.6341 0.66694
4.771 0.98808 5.4939e-005 3.8183 0.011982 6.2415e-005 0.0011598 0.23045 0.00065928 0.2311 0.21317 0 0.032422 0.0389 0 1.2447 0.41028 0.12343 0.015576 8.3257 0.097135 0.00012234 0.79299 0.0076254 0.0084956 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.15097 0.91731 0.90679 0.0013993 0.98709 0.52516 0.001885 0.42734 1.914 1.9132 16.0069 144.9648 0.00017938 -85.6343 0.66794
4.772 0.98808 5.4939e-005 3.8183 0.011982 6.2428e-005 0.0011598 0.23045 0.00065928 0.2311 0.21317 0 0.032422 0.0389 0 1.2448 0.41033 0.12345 0.015578 8.3275 0.097145 0.00012235 0.79298 0.0076261 0.0084963 0.0013903 0.98689 0.99167 2.9984e-006 1.1993e-005 0.15097 0.91751 0.90688 0.0013992 0.98716 0.52533 0.001885 0.42736 1.9146 1.9137 16.0069 144.9648 0.00017925 -85.6345 0.66894
4.773 0.98808 5.4938e-005 3.8183 0.011982 6.2441e-005 0.0011598 0.23045 0.00065928 0.23111 0.21317 0 0.032421 0.0389 0 1.2449 0.41038 0.12347 0.015579 8.3293 0.097154 0.00012237 0.79297 0.0076267 0.008497 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.15098 0.91772 0.90697 0.0013992 0.98722 0.52549 0.001885 0.42737 1.9151 1.9143 16.0068 144.9649 0.00017911 -85.6348 0.66994
4.774 0.98808 5.4938e-005 3.8183 0.011982 6.2454e-005 0.0011598 0.23046 0.00065928 0.23111 0.21318 0 0.032421 0.0389 0 1.245 0.41042 0.12348 0.015581 8.3312 0.097164 0.00012238 0.79296 0.0076273 0.0084977 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.15098 0.91793 0.90705 0.0013992 0.98729 0.52566 0.0018849 0.42738 1.9157 1.9148 16.0068 144.9649 0.00017897 -85.635 0.67094
4.775 0.98808 5.4938e-005 3.8183 0.011982 6.2467e-005 0.0011598 0.23046 0.00065928 0.23111 0.21318 0 0.032421 0.0389 0 1.2451 0.41047 0.1235 0.015583 8.333 0.097173 0.00012239 0.79295 0.007628 0.0084984 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.15099 0.91813 0.90714 0.0013991 0.98735 0.52582 0.0018849 0.42739 1.9162 1.9154 16.0068 144.9649 0.00017884 -85.6352 0.67194
4.776 0.98808 5.4938e-005 3.8183 0.011982 6.248e-005 0.0011598 0.23046 0.00065928 0.23112 0.21318 0 0.032421 0.0389 0 1.2452 0.41052 0.12351 0.015584 8.3348 0.097183 0.00012241 0.79294 0.0076286 0.0084991 0.0013901 0.98689 0.99167 2.9979e-006 1.1992e-005 0.15099 0.91833 0.90723 0.0013991 0.98742 0.52599 0.0018849 0.42741 1.9168 1.9159 16.0068 144.9649 0.0001787 -85.6354 0.67294
4.777 0.98808 5.4938e-005 3.8183 0.011982 6.2493e-005 0.0011598 0.23047 0.00065928 0.23112 0.21319 0 0.032421 0.0389 0 1.2453 0.41056 0.12353 0.015586 8.3367 0.097192 0.00012242 0.79293 0.0076293 0.0084998 0.00139 0.9869 0.99167 2.9978e-006 1.1991e-005 0.151 0.91854 0.90731 0.0013991 0.98748 0.52615 0.0018848 0.42742 1.9173 1.9165 16.0067 144.9649 0.00017857 -85.6357 0.67394
4.778 0.98808 5.4938e-005 3.8183 0.011982 6.2506e-005 0.0011598 0.23047 0.00065928 0.23112 0.21319 0 0.032421 0.0389 0 1.2454 0.41061 0.12354 0.015587 8.3385 0.097202 0.00012243 0.79292 0.0076299 0.0085005 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.151 0.91874 0.9074 0.001399 0.98754 0.52632 0.0018848 0.42743 1.9179 1.917 16.0067 144.965 0.00017843 -85.6359 0.67494
4.779 0.98808 5.4938e-005 3.8183 0.011982 6.2519e-005 0.0011598 0.23047 0.00065928 0.23113 0.21319 0 0.03242 0.0389 0 1.2455 0.41066 0.12356 0.015589 8.3403 0.097212 0.00012245 0.79291 0.0076306 0.0085012 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.15101 0.91894 0.90749 0.001399 0.9876 0.52648 0.0018848 0.42745 1.9184 1.9176 16.0067 144.965 0.0001783 -85.6361 0.67594
4.78 0.98808 5.4938e-005 3.8183 0.011982 6.2532e-005 0.0011598 0.23048 0.00065928 0.23113 0.2132 0 0.03242 0.0389 0 1.2456 0.4107 0.12358 0.01559 8.3421 0.097221 0.00012246 0.7929 0.0076312 0.0085018 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.15101 0.91915 0.90757 0.001399 0.98767 0.52665 0.0018847 0.42746 1.9189 1.9181 16.0067 144.965 0.00017817 -85.6363 0.67694
4.781 0.98808 5.4938e-005 3.8183 0.011982 6.2545e-005 0.0011598 0.23048 0.00065928 0.23113 0.2132 0 0.03242 0.0389 0 1.2457 0.41075 0.12359 0.015592 8.344 0.097231 0.00012247 0.79289 0.0076318 0.0085025 0.0013899 0.9869 0.99167 2.9973e-006 1.1989e-005 0.15102 0.91935 0.90766 0.001399 0.98773 0.52681 0.0018847 0.42747 1.9195 1.9187 16.0066 144.965 0.00017803 -85.6365 0.67794
4.782 0.98808 5.4938e-005 3.8183 0.011982 6.2558e-005 0.0011598 0.23048 0.00065928 0.23114 0.2132 0 0.03242 0.0389 0 1.2458 0.4108 0.12361 0.015593 8.3458 0.09724 0.00012249 0.79288 0.0076325 0.0085032 0.0013898 0.9869 0.99167 2.9972e-006 1.1989e-005 0.15102 0.91955 0.90774 0.001399 0.98779 0.52698 0.0018846 0.42749 1.92 1.9192 16.0066 144.965 0.0001779 -85.6367 0.67894
4.783 0.98808 5.4938e-005 3.8183 0.011982 6.2571e-005 0.0011598 0.23049 0.00065928 0.23114 0.21321 0 0.03242 0.0389 0 1.2459 0.41084 0.12362 0.015595 8.3476 0.09725 0.0001225 0.79287 0.0076331 0.0085039 0.0013898 0.9869 0.99168 2.9971e-006 1.1988e-005 0.15103 0.91975 0.90783 0.0013989 0.98785 0.52714 0.0018846 0.4275 1.9206 1.9197 16.0066 144.9651 0.00017777 -85.637 0.67994
4.784 0.98808 5.4938e-005 3.8183 0.011982 6.2584e-005 0.0011598 0.23049 0.00065928 0.23114 0.21321 0 0.03242 0.0389 0 1.246 0.41089 0.12364 0.015596 8.3494 0.097259 0.00012251 0.79286 0.0076338 0.0085046 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.15103 0.91995 0.90791 0.0013989 0.98791 0.5273 0.0018846 0.42751 1.9211 1.9203 16.0066 144.9651 0.00017764 -85.6372 0.68094
4.785 0.98808 5.4938e-005 3.8183 0.011982 6.2597e-005 0.0011598 0.23049 0.00065928 0.23115 0.21321 0 0.032419 0.0389 0 1.2461 0.41094 0.12365 0.015598 8.3513 0.097269 0.00012253 0.79285 0.0076344 0.0085053 0.0013896 0.9869 0.99168 2.9969e-006 1.1987e-005 0.15104 0.92015 0.908 0.0013988 0.98797 0.52747 0.0018845 0.42753 1.9216 1.9208 16.0065 144.9651 0.00017751 -85.6374 0.68194
4.786 0.98808 5.4938e-005 3.8183 0.011982 6.261e-005 0.0011598 0.2305 0.00065928 0.23115 0.21322 0 0.032419 0.0389 0 1.2462 0.41098 0.12367 0.0156 8.3531 0.097278 0.00012254 0.79284 0.0076351 0.008506 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.15104 0.92034 0.90808 0.0013988 0.98803 0.52763 0.0018845 0.42754 1.9222 1.9214 16.0065 144.9651 0.00017738 -85.6376 0.68294
4.787 0.98808 5.4937e-005 3.8183 0.011982 6.2623e-005 0.0011598 0.2305 0.00065928 0.23115 0.21322 0 0.032419 0.0389 0 1.2463 0.41103 0.12369 0.015601 8.3549 0.097288 0.00012255 0.79283 0.0076357 0.0085067 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.15105 0.92054 0.90816 0.0013988 0.98809 0.5278 0.0018845 0.42755 1.9227 1.9219 16.0065 144.9651 0.00017725 -85.6378 0.68394
4.788 0.98808 5.4937e-005 3.8183 0.011982 6.2636e-005 0.0011598 0.2305 0.00065928 0.23116 0.21322 0 0.032419 0.0389 0 1.2464 0.41108 0.1237 0.015603 8.3568 0.097297 0.00012257 0.79283 0.0076363 0.0085074 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.15105 0.92074 0.90825 0.0013988 0.98815 0.52796 0.0018844 0.42756 1.9232 1.9224 16.0065 144.9652 0.00017712 -85.638 0.68494
4.789 0.98808 5.4937e-005 3.8183 0.011982 6.2649e-005 0.0011598 0.23051 0.00065928 0.23116 0.21323 0 0.032419 0.0389 0 1.2465 0.41112 0.12372 0.015604 8.3586 0.097307 0.00012258 0.79282 0.007637 0.0085081 0.0013895 0.9869 0.99168 2.9964e-006 1.1986e-005 0.15106 0.92093 0.90833 0.0013988 0.98821 0.52813 0.0018844 0.42758 1.9238 1.923 16.0064 144.9652 0.00017699 -85.6382 0.68594
4.79 0.98808 5.4937e-005 3.8183 0.011981 6.2662e-005 0.0011598 0.23051 0.00065928 0.23117 0.21323 0 0.032419 0.0389 0 1.2466 0.41117 0.12373 0.015606 8.3604 0.097316 0.00012259 0.79281 0.0076376 0.0085088 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.15106 0.92113 0.90841 0.0013988 0.98827 0.52829 0.0018844 0.42759 1.9243 1.9235 16.0064 144.9652 0.00017686 -85.6384 0.68694
4.791 0.98808 5.4937e-005 3.8183 0.011981 6.2675e-005 0.0011598 0.23051 0.00065928 0.23117 0.21323 0 0.032418 0.0389 0 1.2467 0.41122 0.12375 0.015607 8.3623 0.097326 0.00012261 0.7928 0.0076383 0.0085095 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.15107 0.92132 0.90849 0.0013987 0.98832 0.52846 0.0018843 0.4276 1.9248 1.924 16.0064 144.9652 0.00017673 -85.6386 0.68794
4.792 0.98808 5.4937e-005 3.8183 0.011981 6.2688e-005 0.0011598 0.23052 0.00065928 0.23117 0.21324 0 0.032418 0.0389 0 1.2468 0.41126 0.12376 0.015609 8.3641 0.097336 0.00012262 0.79279 0.0076389 0.0085101 0.0013894 0.9869 0.99168 2.9961e-006 1.1984e-005 0.15107 0.92152 0.90858 0.0013987 0.98838 0.52862 0.0018843 0.42762 1.9253 1.9246 16.0064 144.9653 0.0001766 -85.6388 0.68894
4.793 0.98808 5.4937e-005 3.8183 0.011981 6.2701e-005 0.0011599 0.23052 0.00065928 0.23118 0.21324 0 0.032418 0.0389 0 1.2469 0.41131 0.12378 0.01561 8.3659 0.097345 0.00012264 0.79278 0.0076395 0.0085108 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.15108 0.92171 0.90866 0.0013987 0.98844 0.52878 0.0018843 0.42763 1.9259 1.9251 16.0063 144.9653 0.00017647 -85.639 0.68994
4.794 0.98808 5.4937e-005 3.8183 0.011981 6.2714e-005 0.0011599 0.23052 0.00065928 0.23118 0.21324 0 0.032418 0.0389 0 1.247 0.41136 0.1238 0.015612 8.3678 0.097355 0.00012265 0.79277 0.0076402 0.0085115 0.0013892 0.98691 0.99168 2.9959e-006 1.1984e-005 0.15108 0.92191 0.90874 0.0013987 0.9885 0.52895 0.0018843 0.42764 1.9264 1.9256 16.0063 144.9653 0.00017635 -85.6392 0.69094
4.795 0.98808 5.4937e-005 3.8183 0.011981 6.2727e-005 0.0011599 0.23053 0.00065928 0.23118 0.21324 0 0.032418 0.0389 0 1.2471 0.4114 0.12381 0.015613 8.3696 0.097364 0.00012266 0.79276 0.0076408 0.0085122 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.15109 0.9221 0.90882 0.0013986 0.98855 0.52911 0.0018842 0.42766 1.9269 1.9261 16.0063 144.9653 0.00017622 -85.6394 0.69194
4.796 0.98808 5.4937e-005 3.8183 0.011981 6.274e-005 0.0011599 0.23053 0.00065928 0.23119 0.21325 0 0.032418 0.0389 0 1.2472 0.41145 0.12383 0.015615 8.3714 0.097374 0.00012268 0.79275 0.0076415 0.0085129 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.15109 0.92229 0.9089 0.0013986 0.98861 0.52928 0.0018842 0.42767 1.9274 1.9267 16.0063 144.9653 0.0001761 -85.6396 0.69294
4.797 0.98808 5.4937e-005 3.8183 0.011981 6.2753e-005 0.0011599 0.23053 0.00065928 0.23119 0.21325 0 0.032417 0.0389 0 1.2473 0.4115 0.12384 0.015617 8.3733 0.097383 0.00012269 0.79274 0.0076421 0.0085136 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.1511 0.92248 0.90898 0.0013986 0.98866 0.52944 0.0018842 0.42768 1.928 1.9272 16.0062 144.9654 0.00017597 -85.6398 0.69394
4.798 0.98808 5.4937e-005 3.8183 0.011981 6.2766e-005 0.0011599 0.23054 0.00065928 0.23119 0.21325 0 0.032417 0.0389 0 1.2474 0.41154 0.12386 0.015618 8.3751 0.097393 0.0001227 0.79273 0.0076428 0.0085143 0.001389 0.98691 0.99168 2.9955e-006 1.1982e-005 0.1511 0.92267 0.90906 0.0013985 0.98872 0.5296 0.0018841 0.42769 1.9285 1.9277 16.0062 144.9654 0.00017584 -85.64 0.69494
4.799 0.98808 5.4937e-005 3.8183 0.011981 6.2779e-005 0.0011599 0.23054 0.00065928 0.2312 0.21326 0 0.032417 0.0389 0 1.2475 0.41159 0.12387 0.01562 8.3769 0.097402 0.00012272 0.79272 0.0076434 0.008515 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.15111 0.92286 0.90914 0.0013985 0.98877 0.52977 0.0018841 0.42771 1.929 1.9282 16.0062 144.9654 0.00017572 -85.6402 0.69594
4.8 0.98808 5.4937e-005 3.8183 0.011981 6.2792e-005 0.0011599 0.23054 0.00065928 0.2312 0.21326 0 0.032417 0.0389 0 1.2475 0.41164 0.12389 0.015621 8.3788 0.097412 0.00012273 0.79271 0.007644 0.0085157 0.001389 0.98691 0.99168 2.9953e-006 1.1981e-005 0.15111 0.92305 0.90922 0.0013985 0.98883 0.52993 0.0018841 0.42772 1.9295 1.9287 16.0062 144.9654 0.0001756 -85.6404 0.69694
4.801 0.98808 5.4936e-005 3.8183 0.011981 6.2805e-005 0.0011599 0.23055 0.00065928 0.2312 0.21326 0 0.032417 0.0389 0 1.2476 0.41168 0.12391 0.015623 8.3806 0.097421 0.00012274 0.7927 0.0076447 0.0085164 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.15112 0.92324 0.9093 0.0013985 0.98888 0.53009 0.001884 0.42773 1.93 1.9293 16.0061 144.9654 0.00017547 -85.6406 0.69794
4.802 0.98808 5.4936e-005 3.8183 0.011981 6.2817e-005 0.0011599 0.23055 0.00065928 0.23121 0.21327 0 0.032417 0.0389 0 1.2477 0.41173 0.12392 0.015624 8.3824 0.097431 0.00012276 0.79269 0.0076453 0.0085171 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.15112 0.92343 0.90938 0.0013985 0.98894 0.53026 0.001884 0.42775 1.9306 1.9298 16.0061 144.9655 0.00017535 -85.6407 0.69894
4.803 0.98808 5.4936e-005 3.8183 0.011981 6.283e-005 0.0011599 0.23055 0.00065928 0.23121 0.21327 0 0.032416 0.0389 0 1.2478 0.41178 0.12394 0.015626 8.3843 0.09744 0.00012277 0.79268 0.007646 0.0085178 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.15113 0.92362 0.90946 0.0013984 0.98899 0.53042 0.001884 0.42776 1.9311 1.9303 16.0061 144.9655 0.00017523 -85.6409 0.69994
4.804 0.98808 5.4936e-005 3.8183 0.011981 6.2843e-005 0.0011599 0.23056 0.00065928 0.23121 0.21327 0 0.032416 0.0389 0 1.2479 0.41182 0.12395 0.015627 8.3861 0.09745 0.00012278 0.79267 0.0076466 0.0085184 0.0013888 0.98691 0.99168 2.9949e-006 1.1979e-005 0.15113 0.9238 0.90954 0.0013984 0.98904 0.53059 0.0018839 0.42777 1.9316 1.9308 16.0061 144.9655 0.0001751 -85.6411 0.70094
4.805 0.98808 5.4936e-005 3.8183 0.011981 6.2856e-005 0.0011599 0.23056 0.00065928 0.23122 0.21328 0 0.032416 0.0389 0 1.248 0.41187 0.12397 0.015629 8.3879 0.097459 0.0001228 0.79266 0.0076472 0.0085191 0.0013887 0.98691 0.99168 2.9948e-006 1.1979e-005 0.15114 0.92399 0.90962 0.0013984 0.9891 0.53075 0.0018839 0.42779 1.9321 1.9313 16.006 144.9655 0.00017498 -85.6413 0.70194
4.806 0.98808 5.4936e-005 3.8183 0.011981 6.2869e-005 0.0011599 0.23056 0.00065928 0.23122 0.21328 0 0.032416 0.0389 0 1.2481 0.41192 0.12398 0.01563 8.3898 0.097469 0.00012281 0.79265 0.0076479 0.0085198 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.15114 0.92418 0.90969 0.0013984 0.98915 0.53091 0.0018839 0.4278 1.9326 1.9318 16.006 144.9655 0.00017486 -85.6415 0.70294
4.807 0.98808 5.4936e-005 3.8183 0.011981 6.2882e-005 0.0011599 0.23057 0.00065928 0.23122 0.21328 0 0.032416 0.0389 0 1.2482 0.41196 0.124 0.015632 8.3916 0.097478 0.00012282 0.79264 0.0076485 0.0085205 0.0013886 0.98691 0.99168 2.9946e-006 1.1978e-005 0.15115 0.92436 0.90977 0.0013983 0.9892 0.53108 0.0018839 0.42781 1.9331 1.9324 16.006 144.9656 0.00017474 -85.6417 0.70394
4.808 0.98808 5.4936e-005 3.8183 0.011981 6.2895e-005 0.0011599 0.23057 0.00065928 0.23123 0.21329 0 0.032416 0.0389 0 1.2483 0.41201 0.12402 0.015634 8.3934 0.097488 0.00012284 0.79263 0.0076492 0.0085212 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.15115 0.92455 0.90985 0.0013983 0.98925 0.53124 0.0018838 0.42782 1.9336 1.9329 16.006 144.9656 0.00017462 -85.6418 0.70494
4.809 0.98808 5.4936e-005 3.8183 0.011981 6.2908e-005 0.0011599 0.23057 0.00065928 0.23123 0.21329 0 0.032415 0.0389 0 1.2484 0.41206 0.12403 0.015635 8.3953 0.097497 0.00012285 0.79263 0.0076498 0.0085219 0.0013886 0.98691 0.99168 2.9944e-006 1.1978e-005 0.15116 0.92473 0.90993 0.0013983 0.98931 0.5314 0.0018838 0.42784 1.9341 1.9334 16.0059 144.9656 0.0001745 -85.642 0.70594
4.81 0.98808 5.4936e-005 3.8183 0.011981 6.2921e-005 0.0011599 0.23058 0.00065929 0.23123 0.21329 0 0.032415 0.0389 0 1.2485 0.4121 0.12405 0.015637 8.3971 0.097507 0.00012286 0.79262 0.0076504 0.0085226 0.0013885 0.98691 0.99169 2.9943e-006 1.1977e-005 0.15117 0.92492 0.91 0.0013983 0.98936 0.53156 0.0018838 0.42785 1.9346 1.9339 16.0059 144.9656 0.00017438 -85.6422 0.70694
4.811 0.98808 5.4936e-005 3.8183 0.011981 6.2934e-005 0.0011599 0.23058 0.00065929 0.23124 0.2133 0 0.032415 0.0389 0 1.2486 0.41215 0.12406 0.015638 8.399 0.097516 0.00012288 0.79261 0.0076511 0.0085233 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.15117 0.9251 0.91008 0.0013983 0.98941 0.53173 0.0018837 0.42786 1.9351 1.9344 16.0059 144.9656 0.00017426 -85.6424 0.70794
4.812 0.98808 5.4936e-005 3.8183 0.011981 6.2947e-005 0.0011599 0.23058 0.00065929 0.23124 0.2133 0 0.032415 0.0389 0 1.2487 0.4122 0.12408 0.01564 8.4008 0.097526 0.00012289 0.7926 0.0076517 0.008524 0.0013885 0.98692 0.99169 2.9941e-006 1.1976e-005 0.15118 0.92528 0.91016 0.0013982 0.98946 0.53189 0.0018837 0.42788 1.9357 1.9349 16.0059 144.9657 0.00017414 -85.6425 0.70894
4.813 0.98808 5.4936e-005 3.8183 0.011981 6.296e-005 0.0011599 0.23059 0.00065929 0.23124 0.2133 0 0.032415 0.0389 0 1.2488 0.41224 0.12409 0.015641 8.4026 0.097535 0.0001229 0.79259 0.0076524 0.0085247 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.15118 0.92546 0.91023 0.0013982 0.98951 0.53205 0.0018837 0.42789 1.9362 1.9354 16.0058 144.9657 0.00017402 -85.6427 0.70994
4.814 0.98808 5.4935e-005 3.8183 0.011981 6.2973e-005 0.0011599 0.23059 0.00065929 0.23125 0.2133 0 0.032415 0.0389 0 1.2489 0.41229 0.12411 0.015643 8.4045 0.097545 0.00012292 0.79258 0.007653 0.0085253 0.0013884 0.98692 0.99169 2.9939e-006 1.1976e-005 0.15119 0.92565 0.91031 0.0013982 0.98956 0.53222 0.0018837 0.4279 1.9367 1.9359 16.0058 144.9657 0.0001739 -85.6429 0.71094
4.815 0.98808 5.4935e-005 3.8183 0.011981 6.2986e-005 0.0011599 0.23059 0.00065929 0.23125 0.21331 0 0.032414 0.0389 0 1.249 0.41234 0.12413 0.015644 8.4063 0.097554 0.00012293 0.79257 0.0076536 0.008526 0.0013883 0.98692 0.99169 2.9939e-006 1.1975e-005 0.15119 0.92583 0.91038 0.0013982 0.98961 0.53238 0.0018836 0.42791 1.9372 1.9364 16.0058 144.9657 0.00017378 -85.6431 0.71194
4.816 0.98808 5.4935e-005 3.8183 0.011981 6.2999e-005 0.0011599 0.2306 0.00065929 0.23125 0.21331 0 0.032414 0.0389 0 1.2491 0.41238 0.12414 0.015646 8.4082 0.097564 0.00012294 0.79256 0.0076543 0.0085267 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.1512 0.92601 0.91046 0.0013981 0.98966 0.53254 0.0018836 0.42793 1.9377 1.9369 16.0058 144.9657 0.00017367 -85.6432 0.71294
4.817 0.98808 5.4935e-005 3.8183 0.011981 6.3012e-005 0.0011599 0.2306 0.00065929 0.23126 0.21331 0 0.032414 0.0389 0 1.2492 0.41243 0.12416 0.015647 8.41 0.097574 0.00012296 0.79255 0.0076549 0.0085274 0.0013882 0.98692 0.99169 2.9937e-006 1.1975e-005 0.1512 0.92619 0.91053 0.0013981 0.98971 0.53271 0.0018836 0.42794 1.9382 1.9374 16.0057 144.9658 0.00017355 -85.6434 0.71394
4.818 0.98808 5.4935e-005 3.8183 0.011981 6.3025e-005 0.0011599 0.2306 0.00065929 0.23126 0.21332 0 0.032414 0.0389 0 1.2493 0.41248 0.12417 0.015649 8.4118 0.097583 0.00012297 0.79254 0.0076556 0.0085281 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.15121 0.92637 0.91061 0.0013981 0.98975 0.53287 0.0018836 0.42795 1.9387 1.9379 16.0057 144.9658 0.00017343 -85.6436 0.71494
4.819 0.98808 5.4935e-005 3.8183 0.011981 6.3038e-005 0.0011599 0.23061 0.00065929 0.23126 0.21332 0 0.032414 0.0389 0 1.2494 0.41252 0.12419 0.015651 8.4137 0.097593 0.00012299 0.79253 0.0076562 0.0085288 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.15121 0.92654 0.91068 0.0013981 0.9898 0.53303 0.0018835 0.42797 1.9392 1.9384 16.0057 144.9658 0.00017332 -85.6437 0.71594
4.82 0.98808 5.4935e-005 3.8183 0.011981 6.3051e-005 0.0011599 0.23061 0.00065929 0.23126 0.21332 0 0.032414 0.0389 0 1.2495 0.41257 0.1242 0.015652 8.4155 0.097602 0.000123 0.79252 0.0076568 0.0085295 0.0013881 0.98692 0.99169 2.9934e-006 1.1974e-005 0.15122 0.92672 0.91076 0.0013981 0.98985 0.53319 0.0018835 0.42798 1.9397 1.9389 16.0057 144.9658 0.0001732 -85.6439 0.71694
4.821 0.98808 5.4935e-005 3.8183 0.011981 6.3064e-005 0.0011599 0.23061 0.00065929 0.23127 0.21333 0 0.032413 0.0389 0 1.2496 0.41262 0.12422 0.015654 8.4174 0.097612 0.00012301 0.79251 0.0076575 0.0085302 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.15122 0.9269 0.91083 0.0013981 0.9899 0.53336 0.0018835 0.42799 1.9402 1.9394 16.0056 144.9658 0.00017308 -85.6441 0.71794
4.822 0.98808 5.4935e-005 3.8183 0.011981 6.3077e-005 0.0011599 0.23062 0.00065929 0.23127 0.21333 0 0.032413 0.0389 0 1.2497 0.41266 0.12424 0.015655 8.4192 0.097621 0.00012303 0.7925 0.0076581 0.0085309 0.0013881 0.98692 0.99169 2.9932e-006 1.1973e-005 0.15123 0.92708 0.9109 0.001398 0.98995 0.53352 0.0018834 0.42801 1.9406 1.9399 16.0056 144.9659 0.00017297 -85.6442 0.71894
4.823 0.98808 5.4935e-005 3.8183 0.011981 6.309e-005 0.0011599 0.23062 0.00065929 0.23127 0.21333 0 0.032413 0.0389 0 1.2498 0.41271 0.12425 0.015657 8.421 0.097631 0.00012304 0.79249 0.0076587 0.0085315 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.15123 0.92725 0.91098 0.001398 0.98999 0.53368 0.0018834 0.42802 1.9411 1.9404 16.0056 144.9659 0.00017286 -85.6444 0.71994
4.824 0.98808 5.4935e-005 3.8183 0.011981 6.3103e-005 0.0011599 0.23062 0.00065929 0.23128 0.21334 0 0.032413 0.0389 0 1.2499 0.41276 0.12427 0.015658 8.4229 0.09764 0.00012305 0.79248 0.0076594 0.0085322 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.15124 0.92743 0.91105 0.001398 0.99004 0.53384 0.0018834 0.42803 1.9416 1.9409 16.0056 144.9659 0.00017274 -85.6445 0.72094
4.825 0.98808 5.4935e-005 3.8183 0.011981 6.3116e-005 0.0011599 0.23063 0.00065929 0.23128 0.21334 0 0.032413 0.0389 0 1.25 0.4128 0.12428 0.01566 8.4247 0.09765 0.00012307 0.79247 0.00766 0.0085329 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.15124 0.9276 0.91112 0.001398 0.99009 0.53401 0.0018834 0.42804 1.9421 1.9414 16.0055 144.9659 0.00017263 -85.6447 0.72194
4.826 0.98808 5.4935e-005 3.8183 0.011981 6.3129e-005 0.0011599 0.23063 0.00065929 0.23128 0.21334 0 0.032413 0.0389 0 1.2501 0.41285 0.1243 0.015661 8.4266 0.097659 0.00012308 0.79246 0.0076607 0.0085336 0.0013879 0.98692 0.99169 2.9929e-006 1.1972e-005 0.15125 0.92778 0.9112 0.0013979 0.99013 0.53417 0.0018833 0.42806 1.9426 1.9419 16.0055 144.9659 0.00017251 -85.6449 0.72294
4.827 0.98808 5.4935e-005 3.8183 0.011981 6.3142e-005 0.0011599 0.23063 0.00065929 0.23129 0.21335 0 0.032412 0.0389 0 1.2502 0.4129 0.12431 0.015663 8.4284 0.097669 0.00012309 0.79245 0.0076613 0.0085343 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.15125 0.92795 0.91127 0.0013979 0.99018 0.53433 0.0018833 0.42807 1.9431 1.9424 16.0055 144.966 0.0001724 -85.645 0.72394
4.828 0.98808 5.4934e-005 3.8183 0.011981 6.3155e-005 0.0011599 0.23064 0.00065929 0.23129 0.21335 0 0.032412 0.0389 0 1.2503 0.41294 0.12433 0.015664 8.4303 0.097678 0.00012311 0.79245 0.0076619 0.008535 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.15126 0.92813 0.91134 0.0013979 0.99022 0.53449 0.0018833 0.42808 1.9436 1.9429 16.0054 144.966 0.00017229 -85.6452 0.72494
4.829 0.98808 5.4934e-005 3.8183 0.011981 6.3168e-005 0.00116 0.23064 0.00065929 0.23129 0.21335 0 0.032412 0.0389 0 1.2504 0.41299 0.12435 0.015666 8.4321 0.097688 0.00012312 0.79244 0.0076626 0.0085357 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.15126 0.9283 0.91141 0.0013979 0.99027 0.53465 0.0018833 0.4281 1.9441 1.9434 16.0054 144.966 0.00017218 -85.6453 0.72594
4.83 0.98808 5.4934e-005 3.8183 0.011981 6.3181e-005 0.00116 0.23064 0.00065929 0.2313 0.21335 0 0.032412 0.0389 0 1.2505 0.41304 0.12436 0.015667 8.434 0.097697 0.00012313 0.79243 0.0076632 0.0085364 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.15127 0.92847 0.91149 0.0013979 0.99031 0.53482 0.0018832 0.42811 1.9446 1.9438 16.0054 144.966 0.00017206 -85.6455 0.72694
4.831 0.98808 5.4934e-005 3.8183 0.011981 6.3194e-005 0.00116 0.23065 0.00065929 0.2313 0.21336 0 0.032412 0.0389 0 1.2505 0.41308 0.12438 0.015669 8.4358 0.097706 0.00012315 0.79242 0.0076639 0.008537 0.0013878 0.98692 0.99169 2.9925e-006 1.197e-005 0.15127 0.92865 0.91156 0.0013979 0.99036 0.53498 0.0018832 0.42812 1.945 1.9443 16.0054 144.966 0.00017195 -85.6456 0.72794
4.832 0.98808 5.4934e-005 3.8183 0.011981 6.3207e-005 0.00116 0.23065 0.00065929 0.2313 0.21336 0 0.032412 0.0389 0 1.2506 0.41313 0.12439 0.015671 8.4376 0.097716 0.00012316 0.79241 0.0076645 0.0085377 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.15128 0.92882 0.91163 0.0013978 0.9904 0.53514 0.0018832 0.42813 1.9455 1.9448 16.0053 144.9661 0.00017184 -85.6458 0.72894
4.833 0.98808 5.4934e-005 3.8183 0.011981 6.322e-005 0.00116 0.23065 0.00065929 0.23131 0.21336 0 0.032411 0.0389 0 1.2507 0.41318 0.12441 0.015672 8.4395 0.097725 0.00012317 0.7924 0.0076651 0.0085384 0.0013877 0.98693 0.99169 2.9923e-006 1.1969e-005 0.15128 0.92899 0.9117 0.0013978 0.99045 0.5353 0.0018832 0.42815 1.946 1.9453 16.0053 144.9661 0.00017173 -85.6459 0.72994
4.834 0.98808 5.4934e-005 3.8183 0.011981 6.3233e-005 0.00116 0.23066 0.00065929 0.23131 0.21337 0 0.032411 0.0389 0 1.2508 0.41322 0.12442 0.015674 8.4413 0.097735 0.00012319 0.79239 0.0076658 0.0085391 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.15129 0.92916 0.91177 0.0013978 0.99049 0.53546 0.0018832 0.42816 1.9465 1.9458 16.0053 144.9661 0.00017162 -85.6461 0.73094
4.835 0.98808 5.4934e-005 3.8183 0.011981 6.3246e-005 0.00116 0.23066 0.00065929 0.23131 0.21337 0 0.032411 0.0389 0 1.2509 0.41327 0.12444 0.015675 8.4432 0.097744 0.0001232 0.79238 0.0076664 0.0085398 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.15129 0.92933 0.91184 0.0013978 0.99053 0.53563 0.0018831 0.42817 1.947 1.9463 16.0053 144.9661 0.00017151 -85.6462 0.73194
4.836 0.98808 5.4934e-005 3.8183 0.011981 6.3259e-005 0.00116 0.23066 0.00065929 0.23132 0.21337 0 0.032411 0.0389 0 1.251 0.41332 0.12445 0.015677 8.445 0.097754 0.00012321 0.79237 0.007667 0.0085405 0.0013875 0.98693 0.99169 2.9921e-006 1.1968e-005 0.1513 0.9295 0.91191 0.0013977 0.99058 0.53579 0.0018831 0.42819 1.9475 1.9467 16.0052 144.9661 0.0001714 -85.6464 0.73294
4.837 0.98808 5.4934e-005 3.8183 0.011981 6.3272e-005 0.00116 0.23067 0.00065929 0.23132 0.21338 0 0.032411 0.0389 0 1.2511 0.41336 0.12447 0.015678 8.4469 0.097763 0.00012323 0.79236 0.0076677 0.0085412 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.1513 0.92967 0.91198 0.0013977 0.99062 0.53595 0.0018831 0.4282 1.9479 1.9472 16.0052 144.9662 0.00017129 -85.6465 0.73394
4.838 0.98808 5.4934e-005 3.8183 0.011981 6.3285e-005 0.00116 0.23067 0.00065929 0.23132 0.21338 0 0.032411 0.0389 0 1.2512 0.41341 0.12449 0.01568 8.4487 0.097773 0.00012324 0.79235 0.0076683 0.0085419 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.15131 0.92983 0.91205 0.0013977 0.99066 0.53611 0.0018831 0.42821 1.9484 1.9477 16.0052 144.9662 0.00017118 -85.6467 0.73494
4.839 0.98808 5.4934e-005 3.8183 0.011981 6.3297e-005 0.00116 0.23067 0.00065929 0.23133 0.21338 0 0.03241 0.0389 0 1.2513 0.41346 0.1245 0.015681 8.4506 0.097782 0.00012325 0.79234 0.007669 0.0085426 0.0013875 0.98693 0.99169 2.9919e-006 1.1967e-005 0.15131 0.93 0.91212 0.0013977 0.9907 0.53627 0.001883 0.42822 1.9489 1.9482 16.0052 144.9662 0.00017108 -85.6468 0.73594
4.84 0.98808 5.4934e-005 3.8183 0.011981 6.331e-005 0.00116 0.23068 0.00065929 0.23133 0.21339 0 0.03241 0.0389 0 1.2514 0.4135 0.12452 0.015683 8.4524 0.097792 0.00012327 0.79233 0.0076696 0.0085432 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.15132 0.93017 0.91219 0.0013977 0.99075 0.53643 0.001883 0.42824 1.9494 1.9487 16.0051 144.9662 0.00017097 -85.647 0.73694
4.841 0.98808 5.4934e-005 3.8183 0.011981 6.3323e-005 0.00116 0.23068 0.00065929 0.23133 0.21339 0 0.03241 0.0389 0 1.2515 0.41355 0.12453 0.015684 8.4543 0.097801 0.00012328 0.79232 0.0076702 0.0085439 0.0013874 0.98693 0.99169 2.9917e-006 1.1967e-005 0.15132 0.93034 0.91226 0.0013977 0.99079 0.53659 0.001883 0.42825 1.9498 1.9491 16.0051 144.9663 0.00017086 -85.6471 0.73794
4.842 0.98808 5.4933e-005 3.8183 0.011981 6.3336e-005 0.00116 0.23068 0.00065929 0.23134 0.21339 0 0.03241 0.0389 0 1.2516 0.41359 0.12455 0.015686 8.4561 0.097811 0.00012329 0.79231 0.0076709 0.0085446 0.0013874 0.98693 0.9917 2.9916e-006 1.1966e-005 0.15133 0.9305 0.91233 0.0013977 0.99083 0.53676 0.001883 0.42826 1.9503 1.9496 16.0051 144.9663 0.00017075 -85.6473 0.73894
4.843 0.98808 5.4933e-005 3.8183 0.011981 6.3349e-005 0.00116 0.23068 0.00065929 0.23134 0.21339 0 0.03241 0.0389 0 1.2517 0.41364 0.12456 0.015687 8.458 0.09782 0.00012331 0.7923 0.0076715 0.0085453 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.15133 0.93067 0.91239 0.0013976 0.99087 0.53692 0.0018829 0.42827 1.9508 1.9501 16.005 144.9663 0.00017065 -85.6474 0.73994
4.844 0.98808 5.4933e-005 3.8183 0.011981 6.3362e-005 0.00116 0.23069 0.00065929 0.23134 0.2134 0 0.03241 0.0389 0 1.2518 0.41369 0.12458 0.015689 8.4598 0.09783 0.00012332 0.79229 0.0076721 0.008546 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.15134 0.93083 0.91246 0.0013976 0.99091 0.53708 0.0018829 0.42829 1.9513 1.9506 16.005 144.9663 0.00017054 -85.6475 0.74094
4.845 0.98808 5.4933e-005 3.8183 0.011981 6.3375e-005 0.00116 0.23069 0.00065929 0.23135 0.2134 0 0.032409 0.0389 0 1.2519 0.41373 0.1246 0.015691 8.4617 0.097839 0.00012333 0.79228 0.0076728 0.0085467 0.0013872 0.98693 0.9917 2.9914e-006 1.1966e-005 0.15134 0.931 0.91253 0.0013976 0.99095 0.53724 0.0018829 0.4283 1.9517 1.951 16.005 144.9663 0.00017043 -85.6477 0.74194
4.846 0.98808 5.4933e-005 3.8183 0.011981 6.3388e-005 0.00116 0.23069 0.00065929 0.23135 0.2134 0 0.032409 0.0389 0 1.252 0.41378 0.12461 0.015692 8.4635 0.097849 0.00012335 0.79227 0.0076734 0.0085474 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.15135 0.93116 0.9126 0.0013976 0.99099 0.5374 0.0018829 0.42831 1.9522 1.9515 16.005 144.9664 0.00017033 -85.6478 0.74294
4.847 0.98808 5.4933e-005 3.8183 0.011981 6.3401e-005 0.00116 0.2307 0.00065929 0.23135 0.21341 0 0.032409 0.0389 0 1.2521 0.41383 0.12463 0.015694 8.4654 0.097858 0.00012336 0.79227 0.0076741 0.008548 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.15135 0.93133 0.91267 0.0013975 0.99103 0.53756 0.0018829 0.42833 1.9527 1.952 16.0049 144.9664 0.00017022 -85.6479 0.74394
4.848 0.98808 5.4933e-005 3.8183 0.011981 6.3414e-005 0.00116 0.2307 0.00065929 0.23136 0.21341 0 0.032409 0.0389 0 1.2522 0.41387 0.12464 0.015695 8.4672 0.097868 0.00012337 0.79226 0.0076747 0.0085487 0.0013871 0.98693 0.9917 2.9912e-006 1.1965e-005 0.15136 0.93149 0.91273 0.0013975 0.99107 0.53772 0.0018828 0.42834 1.9531 1.9524 16.0049 144.9664 0.00017012 -85.6481 0.74494
4.849 0.98808 5.4933e-005 3.8183 0.011981 6.3427e-005 0.00116 0.2307 0.00065929 0.23136 0.21341 0 0.032409 0.0389 0 1.2523 0.41392 0.12466 0.015697 8.4691 0.097877 0.00012339 0.79225 0.0076753 0.0085494 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.15136 0.93165 0.9128 0.0013975 0.99111 0.53788 0.0018828 0.42835 1.9536 1.9529 16.0049 144.9664 0.00017001 -85.6482 0.74594
4.85 0.98808 5.4933e-005 3.8183 0.011981 6.344e-005 0.00116 0.23071 0.00065929 0.23136 0.21342 0 0.032409 0.0389 0 1.2524 0.41397 0.12467 0.015698 8.4709 0.097887 0.0001234 0.79224 0.007676 0.0085501 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.15137 0.93181 0.91287 0.0013975 0.99115 0.53805 0.0018828 0.42836 1.9541 1.9534 16.0049 144.9664 0.00016991 -85.6484 0.74694
4.851 0.98808 5.4933e-005 3.8183 0.011981 6.3453e-005 0.00116 0.23071 0.00065929 0.23137 0.21342 0 0.032409 0.0389 0 1.2525 0.41401 0.12469 0.0157 8.4728 0.097896 0.00012341 0.79223 0.0076766 0.0085508 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.15137 0.93198 0.91293 0.0013975 0.99119 0.53821 0.0018828 0.42838 1.9545 1.9539 16.0048 144.9665 0.0001698 -85.6485 0.74794
4.852 0.98808 5.4933e-005 3.8183 0.011981 6.3466e-005 0.00116 0.23071 0.00065929 0.23137 0.21342 0 0.032408 0.0389 0 1.2526 0.41406 0.12471 0.015701 8.4746 0.097906 0.00012343 0.79222 0.0076772 0.0085515 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.15138 0.93214 0.913 0.0013975 0.99123 0.53837 0.0018827 0.42839 1.955 1.9543 16.0048 144.9665 0.0001697 -85.6486 0.74894
4.853 0.98808 5.4933e-005 3.8183 0.011981 6.3479e-005 0.00116 0.23072 0.00065929 0.23137 0.21343 0 0.032408 0.0389 0 1.2527 0.41411 0.12472 0.015703 8.4765 0.097915 0.00012344 0.79221 0.0076779 0.0085522 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.15138 0.9323 0.91307 0.0013975 0.99127 0.53853 0.0018827 0.4284 1.9555 1.9548 16.0048 144.9665 0.0001696 -85.6488 0.74994
4.854 0.98808 5.4933e-005 3.8183 0.01198 6.3492e-005 0.00116 0.23072 0.00065929 0.23137 0.21343 0 0.032408 0.0389 0 1.2528 0.41415 0.12474 0.015704 8.4783 0.097925 0.00012346 0.7922 0.0076785 0.0085529 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.15139 0.93246 0.91313 0.0013974 0.99131 0.53869 0.0018827 0.42842 1.9559 1.9552 16.0047 144.9665 0.00016949 -85.6489 0.75094
4.855 0.98808 5.4932e-005 3.8183 0.01198 6.3505e-005 0.00116 0.23072 0.00065929 0.23138 0.21343 0 0.032408 0.0389 0 1.2529 0.4142 0.12475 0.015706 8.4802 0.097934 0.00012347 0.79219 0.0076791 0.0085535 0.0013869 0.98693 0.9917 2.9907e-006 1.1963e-005 0.15139 0.93262 0.9132 0.0013974 0.99135 0.53885 0.0018827 0.42843 1.9564 1.9557 16.0047 144.9665 0.00016939 -85.649 0.75194
4.856 0.98808 5.4932e-005 3.8183 0.01198 6.3518e-005 0.00116 0.23073 0.00065929 0.23138 0.21343 0 0.032408 0.0389 0 1.253 0.41425 0.12477 0.015707 8.4821 0.097943 0.00012348 0.79218 0.0076798 0.0085542 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.1514 0.93278 0.91326 0.0013974 0.99138 0.53901 0.0018827 0.42844 1.9569 1.9562 16.0047 144.9666 0.00016929 -85.6491 0.75294
4.857 0.98808 5.4932e-005 3.8183 0.01198 6.3531e-005 0.00116 0.23073 0.00065929 0.23138 0.21344 0 0.032408 0.0389 0 1.2531 0.41429 0.12478 0.015709 8.4839 0.097953 0.0001235 0.79217 0.0076804 0.0085549 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.1514 0.93294 0.91333 0.0013974 0.99142 0.53917 0.0018826 0.42845 1.9573 1.9566 16.0047 144.9666 0.00016919 -85.6493 0.75394
4.858 0.98808 5.4932e-005 3.8183 0.01198 6.3544e-005 0.00116 0.23073 0.00065929 0.23139 0.21344 0 0.032407 0.0389 0 1.2532 0.41434 0.1248 0.015711 8.4858 0.097962 0.00012351 0.79216 0.0076811 0.0085556 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.15141 0.93309 0.91339 0.0013974 0.99146 0.53933 0.0018826 0.42847 1.9578 1.9571 16.0046 144.9666 0.00016909 -85.6494 0.75494
4.859 0.98808 5.4932e-005 3.8183 0.01198 6.3557e-005 0.00116 0.23074 0.00065929 0.23139 0.21344 0 0.032407 0.0389 0 1.2533 0.41439 0.12482 0.015712 8.4876 0.097972 0.00012352 0.79215 0.0076817 0.0085563 0.0013868 0.98694 0.9917 2.9904e-006 1.1962e-005 0.15141 0.93325 0.91346 0.0013974 0.9915 0.53949 0.0018826 0.42848 1.9582 1.9576 16.0046 144.9666 0.00016898 -85.6495 0.75594
4.86 0.98808 5.4932e-005 3.8183 0.01198 6.357e-005 0.00116 0.23074 0.00065929 0.23139 0.21345 0 0.032407 0.0389 0 1.2534 0.41443 0.12483 0.015714 8.4895 0.097981 0.00012354 0.79214 0.0076823 0.008557 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.15142 0.93341 0.91352 0.0013974 0.99153 0.53965 0.0018826 0.42849 1.9587 1.958 16.0046 144.9666 0.00016888 -85.6496 0.75694
4.861 0.98808 5.4932e-005 3.8183 0.01198 6.3583e-005 0.00116 0.23074 0.00065929 0.2314 0.21345 0 0.032407 0.0389 0 1.2534 0.41448 0.12485 0.015715 8.4913 0.097991 0.00012355 0.79213 0.007683 0.0085577 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.15142 0.93356 0.91359 0.0013974 0.99157 0.53981 0.0018826 0.4285 1.9591 1.9585 16.0045 144.9667 0.00016878 -85.6498 0.75794
4.862 0.98808 5.4932e-005 3.8183 0.01198 6.3596e-005 0.00116 0.23075 0.00065929 0.2314 0.21345 0 0.032407 0.0389 0 1.2535 0.41453 0.12486 0.015717 8.4932 0.098 0.00012356 0.79212 0.0076836 0.0085583 0.0013868 0.98694 0.9917 2.9902e-006 1.1961e-005 0.15143 0.93372 0.91365 0.0013973 0.99161 0.53997 0.0018825 0.42852 1.9596 1.9589 16.0045 144.9667 0.00016868 -85.6499 0.75894
4.863 0.98808 5.4932e-005 3.8183 0.01198 6.3609e-005 0.00116 0.23075 0.00065929 0.2314 0.21346 0 0.032407 0.0389 0 1.2536 0.41457 0.12488 0.015718 8.495 0.09801 0.00012358 0.79211 0.0076842 0.008559 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.15143 0.93388 0.91372 0.0013973 0.99164 0.54013 0.0018825 0.42853 1.96 1.9594 16.0045 144.9667 0.00016858 -85.65 0.75994
4.864 0.98808 5.4932e-005 3.8183 0.01198 6.3622e-005 0.00116 0.23075 0.00065929 0.23141 0.21346 0 0.032406 0.0389 0 1.2537 0.41462 0.12489 0.01572 8.4969 0.098019 0.00012359 0.7921 0.0076849 0.0085597 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.15144 0.93403 0.91378 0.0013973 0.99168 0.54029 0.0018825 0.42854 1.9605 1.9598 16.0045 144.9667 0.00016848 -85.6501 0.76094
4.865 0.98808 5.4932e-005 3.8183 0.01198 6.3635e-005 0.0011601 0.23076 0.00065929 0.23141 0.21346 0 0.032406 0.0389 0 1.2538 0.41467 0.12491 0.015721 8.4988 0.098029 0.0001236 0.79209 0.0076855 0.0085604 0.0013867 0.98694 0.9917 2.99e-006 1.196e-005 0.15144 0.93419 0.91384 0.0013973 0.99171 0.54045 0.0018825 0.42856 1.961 1.9603 16.0044 144.9667 0.00016838 -85.6503 0.76194
4.866 0.98808 5.4932e-005 3.8183 0.01198 6.3648e-005 0.0011601 0.23076 0.00065929 0.23141 0.21346 0 0.032406 0.0389 0 1.2539 0.41471 0.12492 0.015723 8.5006 0.098038 0.00012362 0.79209 0.0076861 0.0085611 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.15145 0.93434 0.91391 0.0013973 0.99175 0.54061 0.0018825 0.42857 1.9614 1.9607 16.0044 144.9668 0.00016829 -85.6504 0.76294
4.867 0.98808 5.4932e-005 3.8183 0.01198 6.3661e-005 0.0011601 0.23076 0.00065929 0.23142 0.21347 0 0.032406 0.0389 0 1.254 0.41476 0.12494 0.015724 8.5025 0.098048 0.00012363 0.79208 0.0076868 0.0085618 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.15145 0.93449 0.91397 0.0013972 0.99179 0.54077 0.0018824 0.42858 1.9619 1.9612 16.0044 144.9668 0.00016819 -85.6505 0.76394
4.868 0.98808 5.4932e-005 3.8183 0.01198 6.3674e-005 0.0011601 0.23076 0.00065929 0.23142 0.21347 0 0.032406 0.0389 0 1.2541 0.41481 0.12496 0.015726 8.5043 0.098057 0.00012364 0.79207 0.0076874 0.0085624 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.15146 0.93465 0.91403 0.0013972 0.99182 0.54093 0.0018824 0.42859 1.9623 1.9616 16.0044 144.9668 0.00016809 -85.6506 0.76494
4.869 0.98808 5.4931e-005 3.8183 0.01198 6.3687e-005 0.0011601 0.23077 0.00065929 0.23142 0.21347 0 0.032406 0.0389 0 1.2542 0.41485 0.12497 0.015727 8.5062 0.098066 0.00012366 0.79206 0.007688 0.0085631 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.15146 0.9348 0.91409 0.0013972 0.99185 0.54109 0.0018824 0.42861 1.9628 1.9621 16.0043 144.9668 0.00016799 -85.6507 0.76594
4.87 0.98808 5.4931e-005 3.8183 0.01198 6.37e-005 0.0011601 0.23077 0.00065929 0.23143 0.21348 0 0.032405 0.0389 0 1.2543 0.4149 0.12499 0.015729 8.5081 0.098076 0.00012367 0.79205 0.0076887 0.0085638 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.15147 0.93495 0.91416 0.0013972 0.99189 0.54125 0.0018824 0.42862 1.9632 1.9625 16.0043 144.9668 0.00016789 -85.6509 0.76694
4.871 0.98808 5.4931e-005 3.8183 0.01198 6.3713e-005 0.0011601 0.23077 0.00065929 0.23143 0.21348 0 0.032405 0.0389 0 1.2544 0.41495 0.125 0.015731 8.5099 0.098085 0.00012368 0.79204 0.0076893 0.0085645 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.15147 0.9351 0.91422 0.0013972 0.99192 0.54141 0.0018824 0.42863 1.9636 1.963 16.0043 144.9669 0.0001678 -85.651 0.76794
4.872 0.98808 5.4931e-005 3.8183 0.01198 6.3726e-005 0.0011601 0.23078 0.00065929 0.23143 0.21348 0 0.032405 0.0389 0 1.2545 0.41499 0.12502 0.015732 8.5118 0.098095 0.0001237 0.79203 0.0076899 0.0085652 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.15148 0.93526 0.91428 0.0013972 0.99196 0.54157 0.0018824 0.42864 1.9641 1.9634 16.0042 144.9669 0.0001677 -85.6511 0.76894
4.873 0.98808 5.4931e-005 3.8183 0.01198 6.3739e-005 0.0011601 0.23078 0.00065929 0.23143 0.21349 0 0.032405 0.0389 0 1.2546 0.41504 0.12503 0.015734 8.5136 0.098104 0.00012371 0.79202 0.0076906 0.0085659 0.0013865 0.98694 0.9917 2.9895e-006 1.1958e-005 0.15148 0.93541 0.91434 0.0013972 0.99199 0.54173 0.0018823 0.42866 1.9645 1.9639 16.0042 144.9669 0.0001676 -85.6512 0.76994
4.874 0.98808 5.4931e-005 3.8183 0.01198 6.3751e-005 0.0011601 0.23078 0.00065929 0.23144 0.21349 0 0.032405 0.0389 0 1.2547 0.41509 0.12505 0.015735 8.5155 0.098114 0.00012372 0.79201 0.0076912 0.0085666 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.15149 0.93556 0.9144 0.0013972 0.99203 0.54189 0.0018823 0.42867 1.965 1.9643 16.0042 144.9669 0.00016751 -85.6513 0.77094
4.875 0.98808 5.4931e-005 3.8183 0.01198 6.3764e-005 0.0011601 0.23079 0.00065929 0.23144 0.21349 0 0.032405 0.0389 0 1.2548 0.41513 0.12507 0.015737 8.5174 0.098123 0.00012374 0.792 0.0076918 0.0085672 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.15149 0.93571 0.91446 0.0013971 0.99206 0.54205 0.0018823 0.42868 1.9654 1.9648 16.0042 144.9669 0.00016741 -85.6514 0.77194
4.876 0.98808 5.4931e-005 3.8183 0.01198 6.3777e-005 0.0011601 0.23079 0.00065929 0.23144 0.21349 0 0.032405 0.0389 0 1.2549 0.41518 0.12508 0.015738 8.5192 0.098133 0.00012375 0.79199 0.0076925 0.0085679 0.0013863 0.98694 0.9917 2.9894e-006 1.1957e-005 0.1515 0.93586 0.91453 0.0013971 0.99209 0.54221 0.0018823 0.42869 1.9659 1.9652 16.0041 144.967 0.00016732 -85.6515 0.77294
4.877 0.98808 5.4931e-005 3.8183 0.01198 6.379e-005 0.0011601 0.23079 0.00065929 0.23145 0.2135 0 0.032404 0.0389 0 1.255 0.41523 0.1251 0.01574 8.5211 0.098142 0.00012376 0.79198 0.0076931 0.0085686 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.1515 0.93601 0.91459 0.0013971 0.99213 0.54237 0.0018823 0.42871 1.9663 1.9657 16.0041 144.967 0.00016722 -85.6516 0.77394
4.878 0.98808 5.4931e-005 3.8183 0.01198 6.3803e-005 0.0011601 0.2308 0.00065929 0.23145 0.2135 0 0.032404 0.0389 0 1.2551 0.41527 0.12511 0.015741 8.5229 0.098152 0.00012378 0.79197 0.0076938 0.0085693 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.15151 0.93615 0.91465 0.0013971 0.99216 0.54253 0.0018822 0.42872 1.9668 1.9661 16.0041 144.967 0.00016713 -85.6518 0.77494
4.879 0.98808 5.4931e-005 3.8183 0.01198 6.3816e-005 0.0011601 0.2308 0.00065929 0.23145 0.2135 0 0.032404 0.0389 0 1.2552 0.41532 0.12513 0.015743 8.5248 0.098161 0.00012379 0.79196 0.0076944 0.00857 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.15151 0.9363 0.91471 0.0013971 0.99219 0.54269 0.0018822 0.42873 1.9672 1.9665 16.004 144.967 0.00016703 -85.6519 0.77594
4.88 0.98808 5.4931e-005 3.8183 0.01198 6.3829e-005 0.0011601 0.2308 0.00065929 0.23146 0.21351 0 0.032404 0.0389 0 1.2553 0.41537 0.12514 0.015744 8.5267 0.09817 0.0001238 0.79195 0.007695 0.0085707 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.15152 0.93645 0.91477 0.0013971 0.99222 0.54285 0.0018822 0.42875 1.9676 1.967 16.004 144.967 0.00016694 -85.652 0.77694
4.881 0.98808 5.4931e-005 3.8183 0.01198 6.3842e-005 0.0011601 0.23081 0.00065929 0.23146 0.21351 0 0.032404 0.0389 0 1.2554 0.41541 0.12516 0.015746 8.5285 0.09818 0.00012382 0.79194 0.0076957 0.0085713 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.15152 0.9366 0.91483 0.0013971 0.99226 0.54301 0.0018822 0.42876 1.9681 1.9674 16.004 144.9671 0.00016684 -85.6521 0.77794
4.882 0.98808 5.493e-005 3.8183 0.01198 6.3855e-005 0.0011601 0.23081 0.00065929 0.23146 0.21351 0 0.032404 0.0389 0 1.2555 0.41546 0.12518 0.015747 8.5304 0.098189 0.00012383 0.79193 0.0076963 0.008572 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.15153 0.93674 0.91489 0.0013971 0.99229 0.54317 0.0018822 0.42877 1.9685 1.9679 16.004 144.9671 0.00016675 -85.6522 0.77894
4.883 0.98808 5.493e-005 3.8183 0.01198 6.3868e-005 0.0011601 0.23081 0.00065929 0.23147 0.21351 0 0.032403 0.0389 0 1.2556 0.41551 0.12519 0.015749 8.5323 0.098199 0.00012384 0.79193 0.0076969 0.0085727 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.15153 0.93689 0.91495 0.001397 0.99232 0.54332 0.0018822 0.42878 1.9689 1.9683 16.0039 144.9671 0.00016666 -85.6523 0.77994
4.884 0.98808 5.493e-005 3.8183 0.01198 6.3881e-005 0.0011601 0.23081 0.00065929 0.23147 0.21352 0 0.032403 0.0389 0 1.2557 0.41555 0.12521 0.01575 8.5341 0.098208 0.00012386 0.79192 0.0076976 0.0085734 0.0013862 0.98695 0.9917 2.9889e-006 1.1956e-005 0.15154 0.93704 0.91501 0.001397 0.99235 0.54348 0.0018821 0.4288 1.9694 1.9687 16.0039 144.9671 0.00016657 -85.6524 0.78094
4.885 0.98808 5.493e-005 3.8183 0.01198 6.3894e-005 0.0011601 0.23082 0.00065929 0.23147 0.21352 0 0.032403 0.0389 0 1.2558 0.4156 0.12522 0.015752 8.536 0.098218 0.00012387 0.79191 0.0076982 0.0085741 0.0013861 0.98695 0.99171 2.9889e-006 1.1955e-005 0.15154 0.93718 0.91507 0.001397 0.99238 0.54364 0.0018821 0.42881 1.9698 1.9692 16.0039 144.9672 0.00016647 -85.6525 0.78194
4.886 0.98808 5.493e-005 3.8183 0.01198 6.3907e-005 0.0011601 0.23082 0.00065929 0.23148 0.21352 0 0.032403 0.0389 0 1.2559 0.41565 0.12524 0.015754 8.5379 0.098227 0.00012388 0.7919 0.0076988 0.0085748 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.15155 0.93733 0.91512 0.001397 0.99241 0.5438 0.0018821 0.42882 1.9702 1.9696 16.0038 144.9672 0.00016638 -85.6526 0.78294
4.887 0.98808 5.493e-005 3.8183 0.01198 6.392e-005 0.0011601 0.23082 0.00065929 0.23148 0.21353 0 0.032403 0.0389 0 1.256 0.41569 0.12525 0.015755 8.5397 0.098237 0.0001239 0.79189 0.0076995 0.0085754 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.15155 0.93747 0.91518 0.001397 0.99244 0.54396 0.0018821 0.42883 1.9707 1.97 16.0038 144.9672 0.00016629 -85.6527 0.78394
4.888 0.98808 5.493e-005 3.8183 0.01198 6.3933e-005 0.0011601 0.23083 0.00065929 0.23148 0.21353 0 0.032403 0.0389 0 1.2561 0.41574 0.12527 0.015757 8.5416 0.098246 0.00012391 0.79188 0.0077001 0.0085761 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.15156 0.93761 0.91524 0.001397 0.99248 0.54412 0.0018821 0.42885 1.9711 1.9705 16.0038 144.9672 0.0001662 -85.6528 0.78494
4.889 0.98808 5.493e-005 3.8183 0.01198 6.3946e-005 0.0011601 0.23083 0.00065929 0.23148 0.21353 0 0.032403 0.0389 0 1.2562 0.41579 0.12529 0.015758 8.5435 0.098255 0.00012392 0.79187 0.0077007 0.0085768 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.15156 0.93776 0.9153 0.001397 0.99251 0.54428 0.0018821 0.42886 1.9715 1.9709 16.0038 144.9672 0.00016611 -85.6529 0.78594
4.89 0.98808 5.493e-005 3.8183 0.01198 6.3959e-005 0.0011601 0.23083 0.00065929 0.23149 0.21354 0 0.032402 0.0389 0 1.2563 0.41583 0.1253 0.01576 8.5453 0.098265 0.00012394 0.79186 0.0077014 0.0085775 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.15157 0.9379 0.91536 0.001397 0.99254 0.54444 0.001882 0.42887 1.972 1.9713 16.0037 144.9673 0.00016601 -85.653 0.78694
4.891 0.98808 5.493e-005 3.8183 0.01198 6.3972e-005 0.0011601 0.23084 0.00065929 0.23149 0.21354 0 0.032402 0.0389 0 1.2563 0.41588 0.12532 0.015761 8.5472 0.098274 0.00012395 0.79185 0.007702 0.0085782 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.15157 0.93804 0.91542 0.001397 0.99257 0.54459 0.001882 0.42888 1.9724 1.9718 16.0037 144.9673 0.00016592 -85.6531 0.78794
4.892 0.98808 5.493e-005 3.8183 0.01198 6.3985e-005 0.0011601 0.23084 0.00065929 0.23149 0.21354 0 0.032402 0.0389 0 1.2564 0.41593 0.12533 0.015763 8.5491 0.098284 0.00012396 0.79184 0.0077026 0.0085789 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.15158 0.93819 0.91547 0.0013969 0.9926 0.54475 0.001882 0.4289 1.9728 1.9722 16.0037 144.9673 0.00016583 -85.6532 0.78894
4.893 0.98808 5.493e-005 3.8183 0.01198 6.3998e-005 0.0011601 0.23084 0.00065929 0.2315 0.21354 0 0.032402 0.0389 0 1.2565 0.41597 0.12535 0.015764 8.5509 0.098293 0.00012398 0.79183 0.0077033 0.0085795 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.15158 0.93833 0.91553 0.0013969 0.99263 0.54491 0.001882 0.42891 1.9733 1.9726 16.0036 144.9673 0.00016574 -85.6533 0.78994
4.894 0.98808 5.493e-005 3.8183 0.01198 6.4011e-005 0.0011601 0.23085 0.00065929 0.2315 0.21355 0 0.032402 0.0389 0 1.2566 0.41602 0.12536 0.015766 8.5528 0.098303 0.00012399 0.79182 0.0077039 0.0085802 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.15159 0.93847 0.91559 0.0013969 0.99266 0.54507 0.001882 0.42892 1.9737 1.9731 16.0036 144.9673 0.00016565 -85.6534 0.79094
4.895 0.98808 5.493e-005 3.8183 0.01198 6.4024e-005 0.0011601 0.23085 0.00065929 0.2315 0.21355 0 0.032402 0.0389 0 1.2567 0.41607 0.12538 0.015767 8.5547 0.098312 0.000124 0.79181 0.0077045 0.0085809 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15159 0.93861 0.91565 0.0013969 0.99269 0.54523 0.001882 0.42893 1.9741 1.9735 16.0036 144.9674 0.00016556 -85.6535 0.79194
4.896 0.98808 5.4929e-005 3.8183 0.01198 6.4037e-005 0.0011601 0.23085 0.00065929 0.23151 0.21355 0 0.032401 0.0389 0 1.2568 0.41611 0.12539 0.015769 8.5565 0.098321 0.00012402 0.7918 0.0077052 0.0085816 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.1516 0.93875 0.9157 0.0013969 0.99271 0.54539 0.0018819 0.42895 1.9745 1.9739 16.0036 144.9674 0.00016548 -85.6536 0.79294
4.897 0.98808 5.4929e-005 3.8183 0.01198 6.405e-005 0.0011601 0.23085 0.00065929 0.23151 0.21356 0 0.032401 0.0389 0 1.2569 0.41616 0.12541 0.01577 8.5584 0.098331 0.00012403 0.79179 0.0077058 0.0085823 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.1516 0.93889 0.91576 0.0013968 0.99274 0.54555 0.0018819 0.42896 1.975 1.9743 16.0035 144.9674 0.00016539 -85.6537 0.79394
4.898 0.98808 5.4929e-005 3.8183 0.01198 6.4063e-005 0.0011601 0.23086 0.00065929 0.23151 0.21356 0 0.032401 0.0389 0 1.257 0.41621 0.12543 0.015772 8.5603 0.09834 0.00012404 0.79178 0.0077064 0.0085829 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.15161 0.93903 0.91582 0.0013968 0.99277 0.5457 0.0018819 0.42897 1.9754 1.9748 16.0035 144.9674 0.0001653 -85.6538 0.79494
4.899 0.98808 5.4929e-005 3.8183 0.01198 6.4076e-005 0.0011601 0.23086 0.00065929 0.23152 0.21356 0 0.032401 0.0389 0 1.2571 0.41625 0.12544 0.015773 8.5621 0.09835 0.00012406 0.79177 0.0077071 0.0085836 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.15161 0.93917 0.91587 0.0013968 0.9928 0.54586 0.0018819 0.42898 1.9758 1.9752 16.0035 144.9674 0.00016521 -85.6539 0.79594
4.9 0.98808 5.4929e-005 3.8183 0.01198 6.4089e-005 0.0011602 0.23086 0.00065929 0.23152 0.21356 0 0.032401 0.0389 0 1.2572 0.4163 0.12546 0.015775 8.564 0.098359 0.00012407 0.79176 0.0077077 0.0085843 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.15162 0.93931 0.91593 0.0013968 0.99283 0.54602 0.0018819 0.429 1.9762 1.9756 16.0034 144.9675 0.00016512 -85.654 0.79694
4.901 0.98808 5.4929e-005 3.8183 0.01198 6.4102e-005 0.0011602 0.23087 0.00065929 0.23152 0.21357 0 0.032401 0.0389 0 1.2573 0.41635 0.12547 0.015776 8.5659 0.098369 0.00012408 0.79176 0.0077083 0.008585 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.15162 0.93945 0.91599 0.0013968 0.99286 0.54618 0.0018819 0.42901 1.9766 1.976 16.0034 144.9675 0.00016503 -85.6541 0.79794
4.902 0.98808 5.4929e-005 3.8183 0.01198 6.4115e-005 0.0011602 0.23087 0.00065929 0.23152 0.21357 0 0.032401 0.0389 0 1.2574 0.41639 0.12549 0.015778 8.5677 0.098378 0.0001241 0.79175 0.007709 0.0085857 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.15163 0.93958 0.91604 0.0013968 0.99289 0.54634 0.0018819 0.42902 1.9771 1.9765 16.0034 144.9675 0.00016495 -85.6542 0.79894
4.903 0.98808 5.4929e-005 3.8183 0.01198 6.4128e-005 0.0011602 0.23087 0.00065929 0.23153 0.21357 0 0.0324 0.0389 0 1.2575 0.41644 0.1255 0.01578 8.5696 0.098387 0.00012411 0.79174 0.0077096 0.0085864 0.0013858 0.98695 0.99171 2.9879e-006 1.1952e-005 0.15163 0.93972 0.9161 0.0013968 0.99291 0.54649 0.0018818 0.42903 1.9775 1.9769 16.0033 144.9675 0.00016486 -85.6543 0.79994
4.904 0.98808 5.4929e-005 3.8183 0.01198 6.4141e-005 0.0011602 0.23088 0.00065929 0.23153 0.21358 0 0.0324 0.0389 0 1.2576 0.41649 0.12552 0.015781 8.5715 0.098397 0.00012412 0.79173 0.0077102 0.008587 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.15164 0.93986 0.91615 0.0013968 0.99294 0.54665 0.0018818 0.42905 1.9779 1.9773 16.0033 144.9675 0.00016477 -85.6544 0.80094
4.905 0.98808 5.4929e-005 3.8183 0.01198 6.4154e-005 0.0011602 0.23088 0.00065929 0.23153 0.21358 0 0.0324 0.0389 0 1.2577 0.41653 0.12554 0.015783 8.5734 0.098406 0.00012414 0.79172 0.0077108 0.0085877 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.15164 0.93999 0.91621 0.0013968 0.99297 0.54681 0.0018818 0.42906 1.9783 1.9777 16.0033 144.9676 0.00016469 -85.6545 0.80194
4.906 0.98808 5.4929e-005 3.8183 0.01198 6.4167e-005 0.0011602 0.23088 0.00065929 0.23154 0.21358 0 0.0324 0.0389 0 1.2578 0.41658 0.12555 0.015784 8.5752 0.098416 0.00012415 0.79171 0.0077115 0.0085884 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.15165 0.94013 0.91626 0.0013968 0.993 0.54697 0.0018818 0.42907 1.9787 1.9781 16.0033 144.9676 0.0001646 -85.6545 0.80294
4.907 0.98808 5.4929e-005 3.8183 0.01198 6.4179e-005 0.0011602 0.23089 0.00065929 0.23154 0.21358 0 0.0324 0.0389 0 1.2579 0.41663 0.12557 0.015786 8.5771 0.098425 0.00012416 0.7917 0.0077121 0.0085891 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.15165 0.94027 0.91632 0.0013968 0.99302 0.54713 0.0018818 0.42908 1.9792 1.9786 16.0032 144.9676 0.00016452 -85.6546 0.80394
4.908 0.98808 5.4929e-005 3.8183 0.01198 6.4192e-005 0.0011602 0.23089 0.00065929 0.23154 0.21359 0 0.0324 0.0389 0 1.258 0.41667 0.12558 0.015787 8.579 0.098434 0.00012418 0.79169 0.0077127 0.0085898 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.15166 0.9404 0.91637 0.0013967 0.99305 0.54728 0.0018818 0.4291 1.9796 1.979 16.0032 144.9676 0.00016443 -85.6547 0.80494
4.909 0.98808 5.4928e-005 3.8183 0.01198 6.4205e-005 0.0011602 0.23089 0.00065929 0.23155 0.21359 0 0.032399 0.0389 0 1.2581 0.41672 0.1256 0.015789 8.5808 0.098444 0.00012419 0.79168 0.0077134 0.0085904 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.15166 0.94054 0.91643 0.0013967 0.99308 0.54744 0.0018818 0.42911 1.98 1.9794 16.0032 144.9676 0.00016434 -85.6548 0.80594
4.91 0.98808 5.4928e-005 3.8183 0.01198 6.4218e-005 0.0011602 0.23089 0.00065929 0.23155 0.21359 0 0.032399 0.0389 0 1.2582 0.41677 0.12561 0.01579 8.5827 0.098453 0.0001242 0.79167 0.007714 0.0085911 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.15167 0.94067 0.91648 0.0013967 0.9931 0.5476 0.0018817 0.42912 1.9804 1.9798 16.0031 144.9677 0.00016426 -85.6549 0.80694
4.911 0.98808 5.4928e-005 3.8183 0.01198 6.4231e-005 0.0011602 0.2309 0.00065929 0.23155 0.2136 0 0.032399 0.0389 0 1.2583 0.41681 0.12563 0.015792 8.5846 0.098463 0.00012422 0.79166 0.0077146 0.0085918 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.15167 0.9408 0.91654 0.0013967 0.99313 0.54776 0.0018817 0.42913 1.9808 1.9802 16.0031 144.9677 0.00016417 -85.655 0.80794
4.912 0.98808 5.4928e-005 3.8183 0.01198 6.4244e-005 0.0011602 0.2309 0.00065929 0.23155 0.2136 0 0.032399 0.0389 0 1.2584 0.41686 0.12564 0.015793 8.5865 0.098472 0.00012423 0.79165 0.0077153 0.0085925 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.15168 0.94094 0.91659 0.0013967 0.99316 0.54791 0.0018817 0.42915 1.9812 1.9806 16.0031 144.9677 0.00016409 -85.6551 0.80894
4.913 0.98808 5.4928e-005 3.8183 0.01198 6.4257e-005 0.0011602 0.2309 0.00065929 0.23156 0.2136 0 0.032399 0.0389 0 1.2585 0.41691 0.12566 0.015795 8.5883 0.098482 0.00012424 0.79164 0.0077159 0.0085932 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.15168 0.94107 0.91664 0.0013967 0.99318 0.54807 0.0018817 0.42916 1.9816 1.981 16.0031 144.9677 0.00016401 -85.6552 0.80994
4.914 0.98808 5.4928e-005 3.8183 0.01198 6.427e-005 0.0011602 0.23091 0.00065929 0.23156 0.21361 0 0.032399 0.0389 0 1.2586 0.41695 0.12568 0.015796 8.5902 0.098491 0.00012426 0.79163 0.0077165 0.0085939 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.15169 0.9412 0.9167 0.0013967 0.99321 0.54823 0.0018817 0.42917 1.982 1.9815 16.003 144.9677 0.00016392 -85.6552 0.81094
4.915 0.98808 5.4928e-005 3.8183 0.01198 6.4283e-005 0.0011602 0.23091 0.00065929 0.23156 0.21361 0 0.032399 0.0389 0 1.2587 0.417 0.12569 0.015798 8.5921 0.0985 0.00012427 0.79162 0.0077172 0.0085945 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.15169 0.94134 0.91675 0.0013967 0.99323 0.54839 0.0018817 0.42918 1.9825 1.9819 16.003 144.9678 0.00016384 -85.6553 0.81194
4.916 0.98808 5.4928e-005 3.8183 0.01198 6.4296e-005 0.0011602 0.23091 0.00065929 0.23157 0.21361 0 0.032398 0.0389 0 1.2588 0.41704 0.12571 0.015799 8.594 0.09851 0.00012428 0.79161 0.0077178 0.0085952 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.1517 0.94147 0.9168 0.0013966 0.99326 0.54854 0.0018817 0.4292 1.9829 1.9823 16.003 144.9678 0.00016376 -85.6554 0.81294
4.917 0.98808 5.4928e-005 3.8183 0.011979 6.4309e-005 0.0011602 0.23092 0.00065929 0.23157 0.21361 0 0.032398 0.0389 0 1.2589 0.41709 0.12572 0.015801 8.5958 0.098519 0.0001243 0.79161 0.0077184 0.0085959 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.1517 0.9416 0.91686 0.0013966 0.99329 0.5487 0.0018816 0.42921 1.9833 1.9827 16.0029 144.9678 0.00016367 -85.6555 0.81394
4.918 0.98808 5.4928e-005 3.8183 0.011979 6.4322e-005 0.0011602 0.23092 0.00065929 0.23157 0.21362 0 0.032398 0.0389 0 1.259 0.41714 0.12574 0.015802 8.5977 0.098529 0.00012431 0.7916 0.0077191 0.0085966 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.15171 0.94173 0.91691 0.0013966 0.99331 0.54886 0.0018816 0.42922 1.9837 1.9831 16.0029 144.9678 0.00016359 -85.6556 0.81494
4.919 0.98808 5.4928e-005 3.8183 0.011979 6.4335e-005 0.0011602 0.23092 0.00065929 0.23158 0.21362 0 0.032398 0.0389 0 1.259 0.41718 0.12575 0.015804 8.5996 0.098538 0.00012432 0.79159 0.0077197 0.0085973 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.15171 0.94186 0.91696 0.0013966 0.99334 0.54901 0.0018816 0.42923 1.9841 1.9835 16.0029 144.9678 0.00016351 -85.6557 0.81594
4.92 0.98808 5.4928e-005 3.8183 0.011979 6.4348e-005 0.0011602 0.23092 0.00065929 0.23158 0.21362 0 0.032398 0.0389 0 1.2591 0.41723 0.12577 0.015806 8.6015 0.098547 0.00012434 0.79158 0.0077203 0.0085979 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15172 0.94199 0.91701 0.0013966 0.99336 0.54917 0.0018816 0.42925 1.9845 1.9839 16.0028 144.9679 0.00016343 -85.6557 0.81694
4.921 0.98808 5.4928e-005 3.8183 0.011979 6.4361e-005 0.0011602 0.23093 0.00065929 0.23158 0.21363 0 0.032398 0.0389 0 1.2592 0.41728 0.12579 0.015807 8.6034 0.098557 0.00012435 0.79157 0.0077209 0.0085986 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15172 0.94212 0.91707 0.0013966 0.99339 0.54933 0.0018816 0.42926 1.9849 1.9843 16.0028 144.9679 0.00016334 -85.6558 0.81794
4.922 0.98808 5.4928e-005 3.8183 0.011979 6.4374e-005 0.0011602 0.23093 0.00065929 0.23159 0.21363 0 0.032397 0.0389 0 1.2593 0.41732 0.1258 0.015809 8.6052 0.098566 0.00012436 0.79156 0.0077216 0.0085993 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15173 0.94225 0.91712 0.0013966 0.99341 0.54949 0.0018816 0.42927 1.9853 1.9847 16.0028 144.9679 0.00016326 -85.6559 0.81894
4.923 0.98808 5.4927e-005 3.8183 0.011979 6.4387e-005 0.0011602 0.23093 0.00065929 0.23159 0.21363 0 0.032397 0.0389 0 1.2594 0.41737 0.12582 0.01581 8.6071 0.098576 0.00012438 0.79155 0.0077222 0.0086 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.15173 0.94238 0.91717 0.0013966 0.99344 0.54964 0.0018816 0.42928 1.9857 1.9851 16.0028 144.9679 0.00016318 -85.656 0.81994
4.924 0.98808 5.4927e-005 3.8183 0.011979 6.44e-005 0.0011602 0.23094 0.00065929 0.23159 0.21363 0 0.032397 0.0389 0 1.2595 0.41742 0.12583 0.015812 8.609 0.098585 0.00012439 0.79154 0.0077228 0.0086007 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.15174 0.94251 0.91722 0.0013966 0.99346 0.5498 0.0018816 0.4293 1.9861 1.9855 16.0027 144.968 0.0001631 -85.6561 0.82094
4.925 0.98808 5.4927e-005 3.8183 0.011979 6.4413e-005 0.0011602 0.23094 0.00065929 0.23159 0.21364 0 0.032397 0.0389 0 1.2596 0.41746 0.12585 0.015813 8.6109 0.098594 0.0001244 0.79153 0.0077235 0.0086013 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.15174 0.94264 0.91727 0.0013966 0.99348 0.54996 0.0018815 0.42931 1.9865 1.9859 16.0027 144.968 0.00016302 -85.6561 0.82194
4.926 0.98808 5.4927e-005 3.8183 0.011979 6.4426e-005 0.0011602 0.23094 0.00065929 0.2316 0.21364 0 0.032397 0.0389 0 1.2597 0.41751 0.12586 0.015815 8.6128 0.098604 0.00012442 0.79152 0.0077241 0.008602 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.15175 0.94276 0.91733 0.0013965 0.99351 0.55011 0.0018815 0.42932 1.9869 1.9863 16.0027 144.968 0.00016294 -85.6562 0.82294
4.927 0.98808 5.4927e-005 3.8183 0.011979 6.4439e-005 0.0011602 0.23095 0.00065929 0.2316 0.21364 0 0.032397 0.0389 0 1.2598 0.41756 0.12588 0.015816 8.6146 0.098613 0.00012443 0.79151 0.0077247 0.0086027 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.15175 0.94289 0.91738 0.0013965 0.99353 0.55027 0.0018815 0.42933 1.9873 1.9867 16.0026 144.968 0.00016286 -85.6563 0.82394
4.928 0.98808 5.4927e-005 3.8183 0.011979 6.4452e-005 0.0011602 0.23095 0.00065929 0.2316 0.21364 0 0.032397 0.0389 0 1.2599 0.4176 0.12589 0.015818 8.6165 0.098623 0.00012444 0.7915 0.0077254 0.0086034 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.15176 0.94302 0.91743 0.0013965 0.99356 0.55043 0.0018815 0.42935 1.9877 1.9871 16.0026 144.968 0.00016278 -85.6564 0.82494
4.929 0.98808 5.4927e-005 3.8183 0.011979 6.4465e-005 0.0011602 0.23095 0.00065929 0.23161 0.21365 0 0.032396 0.0389 0 1.26 0.41765 0.12591 0.015819 8.6184 0.098632 0.00012446 0.79149 0.007726 0.0086041 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.15176 0.94315 0.91748 0.0013965 0.99358 0.55058 0.0018815 0.42936 1.9881 1.9875 16.0026 144.9681 0.0001627 -85.6565 0.82594
4.93 0.98808 5.4927e-005 3.8183 0.011979 6.4478e-005 0.0011602 0.23095 0.00065929 0.23161 0.21365 0 0.032396 0.0389 0 1.2601 0.4177 0.12593 0.015821 8.6203 0.098641 0.00012447 0.79148 0.0077266 0.0086047 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.15177 0.94327 0.91753 0.0013965 0.9936 0.55074 0.0018815 0.42937 1.9885 1.9879 16.0025 144.9681 0.00016262 -85.6565 0.82694
4.931 0.98808 5.4927e-005 3.8183 0.011979 6.4491e-005 0.0011602 0.23096 0.00065929 0.23161 0.21365 0 0.032396 0.0389 0 1.2602 0.41774 0.12594 0.015822 8.6222 0.098651 0.00012448 0.79147 0.0077272 0.0086054 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.15177 0.9434 0.91758 0.0013965 0.99363 0.5509 0.0018815 0.42938 1.9889 1.9883 16.0025 144.9681 0.00016254 -85.6566 0.82794
4.932 0.98808 5.4927e-005 3.8183 0.011979 6.4504e-005 0.0011602 0.23096 0.00065929 0.23161 0.21366 0 0.032396 0.0389 0 1.2603 0.41779 0.12596 0.015824 8.624 0.09866 0.0001245 0.79146 0.0077279 0.0086061 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.15178 0.94352 0.91763 0.0013965 0.99365 0.55105 0.0018815 0.4294 1.9893 1.9887 16.0025 144.9681 0.00016246 -85.6567 0.82894
4.933 0.98808 5.4927e-005 3.8183 0.011979 6.4517e-005 0.0011602 0.23096 0.00065929 0.23162 0.21366 0 0.032396 0.0389 0 1.2604 0.41784 0.12597 0.015825 8.6259 0.09867 0.00012451 0.79145 0.0077285 0.0086068 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.15178 0.94365 0.91768 0.0013965 0.99367 0.55121 0.0018814 0.42941 1.9897 1.9891 16.0025 144.9681 0.00016238 -85.6568 0.82994
4.934 0.98808 5.4927e-005 3.8183 0.011979 6.453e-005 0.0011602 0.23097 0.00065929 0.23162 0.21366 0 0.032396 0.0389 0 1.2605 0.41788 0.12599 0.015827 8.6278 0.098679 0.00012452 0.79145 0.0077291 0.0086074 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.15179 0.94377 0.91773 0.0013965 0.99369 0.55136 0.0018814 0.42942 1.9901 1.9895 16.0024 144.9682 0.0001623 -85.6568 0.83094
4.935 0.98808 5.4927e-005 3.8183 0.011979 6.4543e-005 0.0011603 0.23097 0.00065929 0.23162 0.21366 0 0.032396 0.0389 0 1.2606 0.41793 0.126 0.015828 8.6297 0.098688 0.00012454 0.79144 0.0077298 0.0086081 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.15179 0.9439 0.91778 0.0013965 0.99372 0.55152 0.0018814 0.42943 1.9905 1.9899 16.0024 144.9682 0.00016223 -85.6569 0.83194
4.936 0.98808 5.4927e-005 3.8183 0.011979 6.4556e-005 0.0011603 0.23097 0.00065929 0.23163 0.21367 0 0.032395 0.0389 0 1.2607 0.41798 0.12602 0.01583 8.6316 0.098698 0.00012455 0.79143 0.0077304 0.0086088 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.1518 0.94402 0.91783 0.0013965 0.99374 0.55168 0.0018814 0.42944 1.9909 1.9903 16.0024 144.9682 0.00016215 -85.657 0.83294
4.937 0.98808 5.4926e-005 3.8183 0.011979 6.4569e-005 0.0011603 0.23098 0.00065929 0.23163 0.21367 0 0.032395 0.0389 0 1.2608 0.41802 0.12604 0.015831 8.6334 0.098707 0.00012456 0.79142 0.007731 0.0086095 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.1518 0.94414 0.91788 0.0013964 0.99376 0.55183 0.0018814 0.42946 1.9913 1.9907 16.0023 144.9682 0.00016207 -85.657 0.83394
4.938 0.98808 5.4926e-005 3.8183 0.011979 6.4582e-005 0.0011603 0.23098 0.00065929 0.23163 0.21367 0 0.032395 0.0389 0 1.2609 0.41807 0.12605 0.015833 8.6353 0.098716 0.00012458 0.79141 0.0077317 0.0086102 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.15181 0.94427 0.91793 0.0013964 0.99378 0.55199 0.0018814 0.42947 1.9917 1.9911 16.0023 144.9682 0.00016199 -85.6571 0.83494
4.939 0.98808 5.4926e-005 3.8183 0.011979 6.4594e-005 0.0011603 0.23098 0.00065929 0.23164 0.21368 0 0.032395 0.0389 0 1.261 0.41812 0.12607 0.015834 8.6372 0.098726 0.00012459 0.7914 0.0077323 0.0086108 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.15181 0.94439 0.91798 0.0013964 0.99381 0.55215 0.0018814 0.42948 1.9921 1.9915 16.0023 144.9683 0.00016192 -85.6572 0.83594
4.94 0.98808 5.4926e-005 3.8183 0.011979 6.4607e-005 0.0011603 0.23098 0.00065929 0.23164 0.21368 0 0.032395 0.0389 0 1.2611 0.41816 0.12608 0.015836 8.6391 0.098735 0.0001246 0.79139 0.0077329 0.0086115 0.0013851 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15182 0.94451 0.91803 0.0013964 0.99383 0.5523 0.0018814 0.42949 1.9925 1.9919 16.0022 144.9683 0.00016184 -85.6573 0.83694
4.941 0.98808 5.4926e-005 3.8183 0.011979 6.462e-005 0.0011603 0.23099 0.00065929 0.23164 0.21368 0 0.032395 0.0389 0 1.2612 0.41821 0.1261 0.015838 8.641 0.098745 0.00012462 0.79138 0.0077335 0.0086122 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15182 0.94463 0.91808 0.0013964 0.99385 0.55246 0.0018814 0.42951 1.9929 1.9923 16.0022 144.9683 0.00016176 -85.6573 0.83794
4.942 0.98808 5.4926e-005 3.8183 0.011979 6.4633e-005 0.0011603 0.23099 0.00065929 0.23164 0.21368 0 0.032395 0.0389 0 1.2613 0.41826 0.12611 0.015839 8.6429 0.098754 0.00012463 0.79137 0.0077342 0.0086129 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15183 0.94476 0.91813 0.0013964 0.99387 0.55261 0.0018813 0.42952 1.9932 1.9927 16.0022 144.9683 0.00016169 -85.6574 0.83894
4.943 0.98808 5.4926e-005 3.8183 0.011979 6.4646e-005 0.0011603 0.23099 0.00065929 0.23165 0.21369 0 0.032394 0.0389 0 1.2614 0.4183 0.12613 0.015841 8.6448 0.098763 0.00012464 0.79136 0.0077348 0.0086136 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.15183 0.94488 0.91817 0.0013964 0.99389 0.55277 0.0018813 0.42953 1.9936 1.9931 16.0021 144.9683 0.00016161 -85.6575 0.83994
4.944 0.98808 5.4926e-005 3.8183 0.011979 6.4659e-005 0.0011603 0.231 0.00065929 0.23165 0.21369 0 0.032394 0.0389 0 1.2615 0.41835 0.12614 0.015842 8.6466 0.098773 0.00012466 0.79135 0.0077354 0.0086142 0.001385 0.98696 0.99171 2.9862e-006 1.1945e-005 0.15184 0.945 0.91822 0.0013964 0.99391 0.55292 0.0018813 0.42954 1.994 1.9935 16.0021 144.9684 0.00016153 -85.6575 0.84094
4.945 0.98808 5.4926e-005 3.8183 0.011979 6.4672e-005 0.0011603 0.231 0.00065929 0.23165 0.21369 0 0.032394 0.0389 0 1.2616 0.4184 0.12616 0.015844 8.6485 0.098782 0.00012467 0.79134 0.0077361 0.0086149 0.0013849 0.98696 0.99172 2.9862e-006 1.1945e-005 0.15184 0.94512 0.91827 0.0013964 0.99394 0.55308 0.0018813 0.42956 1.9944 1.9938 16.0021 144.9684 0.00016146 -85.6576 0.84194
4.946 0.98808 5.4926e-005 3.8183 0.011979 6.4685e-005 0.0011603 0.231 0.00065929 0.23166 0.2137 0 0.032394 0.0389 0 1.2617 0.41844 0.12618 0.015845 8.6504 0.098792 0.00012468 0.79133 0.0077367 0.0086156 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.15185 0.94524 0.91832 0.0013964 0.99396 0.55324 0.0018813 0.42957 1.9948 1.9942 16.0021 144.9684 0.00016138 -85.6577 0.84294
4.947 0.98808 5.4926e-005 3.8183 0.011979 6.4698e-005 0.0011603 0.231 0.00065929 0.23166 0.2137 0 0.032394 0.0389 0 1.2617 0.41849 0.12619 0.015847 8.6523 0.098801 0.0001247 0.79132 0.0077373 0.0086163 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.15185 0.94536 0.91837 0.0013964 0.99398 0.55339 0.0018813 0.42958 1.9952 1.9946 16.002 144.9684 0.00016131 -85.6577 0.84394
4.948 0.98808 5.4926e-005 3.8183 0.011979 6.4711e-005 0.0011603 0.23101 0.00065929 0.23166 0.2137 0 0.032394 0.0389 0 1.2618 0.41854 0.12621 0.015848 8.6542 0.09881 0.00012471 0.79131 0.0077379 0.0086169 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.15186 0.94548 0.91841 0.0013964 0.994 0.55355 0.0018813 0.42959 1.9956 1.995 16.002 144.9684 0.00016123 -85.6578 0.84494
4.949 0.98808 5.4926e-005 3.8183 0.011979 6.4724e-005 0.0011603 0.23101 0.00065929 0.23167 0.2137 0 0.032393 0.0389 0 1.2619 0.41858 0.12622 0.01585 8.6561 0.09882 0.00012472 0.79131 0.0077386 0.0086176 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.15186 0.9456 0.91846 0.0013964 0.99402 0.5537 0.0018813 0.4296 1.996 1.9954 16.002 144.9685 0.00016116 -85.6579 0.84594
4.95 0.98808 5.4925e-005 3.8183 0.011979 6.4737e-005 0.0011603 0.23101 0.00065929 0.23167 0.21371 0 0.032393 0.0389 0 1.262 0.41863 0.12624 0.015851 8.658 0.098829 0.00012474 0.7913 0.0077392 0.0086183 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.15187 0.94572 0.91851 0.0013964 0.99404 0.55386 0.0018813 0.42962 1.9963 1.9958 16.0019 144.9685 0.00016109 -85.6579 0.84694
4.951 0.98808 5.4925e-005 3.8183 0.011979 6.475e-005 0.0011603 0.23102 0.00065929 0.23167 0.21371 0 0.032393 0.0389 0 1.2621 0.41868 0.12625 0.015853 8.6599 0.098838 0.00012475 0.79129 0.0077398 0.008619 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.15187 0.94583 0.91856 0.0013964 0.99406 0.55401 0.0018812 0.42963 1.9967 1.9962 16.0019 144.9685 0.00016101 -85.658 0.84794
4.952 0.98808 5.4925e-005 3.8183 0.011979 6.4763e-005 0.0011603 0.23102 0.00065929 0.23167 0.21371 0 0.032393 0.0389 0 1.2622 0.41872 0.12627 0.015854 8.6617 0.098848 0.00012476 0.79128 0.0077405 0.0086197 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.15188 0.94595 0.9186 0.0013963 0.99408 0.55417 0.0018812 0.42964 1.9971 1.9966 16.0019 144.9685 0.00016094 -85.6581 0.84894
4.953 0.98808 5.4925e-005 3.8183 0.011979 6.4776e-005 0.0011603 0.23102 0.00065929 0.23168 0.21372 0 0.032393 0.0389 0 1.2623 0.41877 0.12629 0.015856 8.6636 0.098857 0.00012478 0.79127 0.0077411 0.0086203 0.0013849 0.98696 0.99172 2.9859e-006 1.1943e-005 0.15188 0.94607 0.91865 0.0013963 0.9941 0.55432 0.0018812 0.42965 1.9975 1.9969 16.0018 144.9685 0.00016086 -85.6581 0.84994
4.954 0.98808 5.4925e-005 3.8183 0.011979 6.4789e-005 0.0011603 0.23103 0.00065929 0.23168 0.21372 0 0.032393 0.0389 0 1.2624 0.41882 0.1263 0.015857 8.6655 0.098867 0.00012479 0.79126 0.0077417 0.008621 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.15189 0.94619 0.9187 0.0013963 0.99412 0.55448 0.0018812 0.42967 1.9979 1.9973 16.0018 144.9686 0.00016079 -85.6582 0.85094
4.955 0.98808 5.4925e-005 3.8183 0.011979 6.4802e-005 0.0011603 0.23103 0.00065929 0.23168 0.21372 0 0.032393 0.0389 0 1.2625 0.41886 0.12632 0.015859 8.6674 0.098876 0.0001248 0.79125 0.0077423 0.0086217 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.15189 0.9463 0.91874 0.0013963 0.99414 0.55463 0.0018812 0.42968 1.9983 1.9977 16.0018 144.9686 0.00016072 -85.6583 0.85194
4.956 0.98808 5.4925e-005 3.8183 0.011979 6.4815e-005 0.0011603 0.23103 0.00065929 0.23169 0.21372 0 0.032392 0.0389 0 1.2626 0.41891 0.12633 0.01586 8.6693 0.098885 0.00012482 0.79124 0.007743 0.0086224 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.1519 0.94642 0.91879 0.0013963 0.99416 0.55479 0.0018812 0.42969 1.9986 1.9981 16.0017 144.9686 0.00016064 -85.6583 0.85294
4.957 0.98808 5.4925e-005 3.8183 0.011979 6.4828e-005 0.0011603 0.23103 0.00065929 0.23169 0.21373 0 0.032392 0.0389 0 1.2627 0.41896 0.12635 0.015862 8.6712 0.098895 0.00012483 0.79123 0.0077436 0.008623 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.1519 0.94654 0.91884 0.0013963 0.99418 0.55494 0.0018812 0.4297 1.999 1.9985 16.0017 144.9686 0.00016057 -85.6584 0.85394
4.958 0.98808 5.4925e-005 3.8183 0.011979 6.4841e-005 0.0011603 0.23104 0.00065929 0.23169 0.21373 0 0.032392 0.0389 0 1.2628 0.419 0.12636 0.015863 8.6731 0.098904 0.00012484 0.79122 0.0077442 0.0086237 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15191 0.94665 0.91888 0.0013963 0.9942 0.5551 0.0018812 0.42972 1.9994 1.9988 16.0017 144.9686 0.0001605 -85.6584 0.85494
4.959 0.98808 5.4925e-005 3.8183 0.011979 6.4854e-005 0.0011603 0.23104 0.00065929 0.23169 0.21373 0 0.032392 0.0389 0 1.2629 0.41905 0.12638 0.015865 8.675 0.098913 0.00012486 0.79121 0.0077449 0.0086244 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15191 0.94677 0.91893 0.0013963 0.99422 0.55525 0.0018812 0.42973 1.9998 1.9992 16.0017 144.9687 0.00016043 -85.6585 0.85594
4.96 0.98808 5.4925e-005 3.8183 0.011979 6.4867e-005 0.0011603 0.23104 0.00065929 0.2317 0.21373 0 0.032392 0.0389 0 1.263 0.4191 0.12639 0.015866 8.6769 0.098923 0.00012487 0.7912 0.0077455 0.0086251 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15192 0.94688 0.91897 0.0013963 0.99424 0.55541 0.0018812 0.42974 2.0001 1.9996 16.0016 144.9687 0.00016036 -85.6586 0.85694
4.961 0.98808 5.4925e-005 3.8183 0.011979 6.488e-005 0.0011603 0.23105 0.00065929 0.2317 0.21374 0 0.032392 0.0389 0 1.2631 0.41914 0.12641 0.015868 8.6788 0.098932 0.00012488 0.79119 0.0077461 0.0086257 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.15192 0.947 0.91902 0.0013963 0.99426 0.55556 0.0018811 0.42975 2.0005 2 16.0016 144.9687 0.00016028 -85.6586 0.85794
4.962 0.98808 5.4925e-005 3.8183 0.011979 6.4893e-005 0.0011603 0.23105 0.00065929 0.2317 0.21374 0 0.032392 0.0389 0 1.2632 0.41919 0.12643 0.01587 8.6806 0.098941 0.0001249 0.79118 0.0077467 0.0086264 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.15193 0.94711 0.91907 0.0013962 0.99428 0.55572 0.0018811 0.42976 2.0009 2.0004 16.0016 144.9687 0.00016021 -85.6587 0.85894
4.963 0.98808 5.4925e-005 3.8183 0.011979 6.4906e-005 0.0011603 0.23105 0.00065929 0.23171 0.21374 0 0.032391 0.0389 0 1.2633 0.41924 0.12644 0.015871 8.6825 0.098951 0.00012491 0.79117 0.0077474 0.0086271 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.15193 0.94722 0.91911 0.0013962 0.99429 0.55587 0.0018811 0.42978 2.0013 2.0007 16.0015 144.9688 0.00016014 -85.6587 0.85994
4.964 0.98808 5.4924e-005 3.8183 0.011979 6.4919e-005 0.0011603 0.23105 0.00065929 0.23171 0.21375 0 0.032391 0.0389 0 1.2634 0.41928 0.12646 0.015873 8.6844 0.09896 0.00012492 0.79116 0.007748 0.0086278 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.15194 0.94734 0.91916 0.0013962 0.99431 0.55603 0.0018811 0.42979 2.0016 2.0011 16.0015 144.9688 0.00016007 -85.6588 0.86094
4.965 0.98808 5.4924e-005 3.8183 0.011979 6.4932e-005 0.0011603 0.23106 0.00065929 0.23171 0.21375 0 0.032391 0.0389 0 1.2635 0.41933 0.12647 0.015874 8.6863 0.09897 0.00012494 0.79116 0.0077486 0.0086284 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.15194 0.94745 0.9192 0.0013962 0.99433 0.55618 0.0018811 0.4298 2.002 2.0015 16.0015 144.9688 0.00016 -85.6589 0.86194
4.966 0.98808 5.4924e-005 3.8183 0.011979 6.4945e-005 0.0011603 0.23106 0.00065929 0.23171 0.21375 0 0.032391 0.0389 0 1.2636 0.41938 0.12649 0.015876 8.6882 0.098979 0.00012495 0.79115 0.0077492 0.0086291 0.0013846 0.98696 0.99172 2.9855e-006 1.1942e-005 0.15195 0.94756 0.91925 0.0013962 0.99435 0.55634 0.0018811 0.42981 2.0024 2.0019 16.0014 144.9688 0.00015993 -85.6589 0.86294
4.967 0.98808 5.4924e-005 3.8183 0.011979 6.4958e-005 0.0011603 0.23106 0.00065929 0.23172 0.21375 0 0.032391 0.0389 0 1.2637 0.41942 0.1265 0.015877 8.6901 0.098988 0.00012496 0.79114 0.0077499 0.0086298 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.15195 0.94768 0.91929 0.0013962 0.99437 0.55649 0.0018811 0.42983 2.0028 2.0022 16.0014 144.9688 0.00015986 -85.659 0.86394
4.968 0.98808 5.4924e-005 3.8183 0.011979 6.4971e-005 0.0011603 0.23107 0.00065929 0.23172 0.21376 0 0.032391 0.0389 0 1.2638 0.41947 0.12652 0.015879 8.692 0.098998 0.00012498 0.79113 0.0077505 0.0086305 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.15196 0.94779 0.91934 0.0013962 0.99439 0.55665 0.0018811 0.42984 2.0031 2.0026 16.0014 144.9689 0.00015979 -85.659 0.86494
4.969 0.98808 5.4924e-005 3.8183 0.011979 6.4983e-005 0.0011604 0.23107 0.00065929 0.23172 0.21376 0 0.032391 0.0389 0 1.2639 0.41952 0.12654 0.01588 8.6939 0.099007 0.00012499 0.79112 0.0077511 0.0086312 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.15196 0.9479 0.91938 0.0013962 0.99441 0.5568 0.0018811 0.42985 2.0035 2.003 16.0013 144.9689 0.00015972 -85.6591 0.86594
4.97 0.98808 5.4924e-005 3.8183 0.011979 6.4996e-005 0.0011604 0.23107 0.00065929 0.23173 0.21376 0 0.03239 0.0389 0 1.264 0.41956 0.12655 0.015882 8.6958 0.099016 0.000125 0.79111 0.0077517 0.0086318 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15197 0.94801 0.91943 0.0013962 0.99442 0.55696 0.0018811 0.42986 2.0039 2.0033 16.0013 144.9689 0.00015965 -85.6592 0.86694
4.971 0.98808 5.4924e-005 3.8183 0.011979 6.5009e-005 0.0011604 0.23107 0.00065929 0.23173 0.21376 0 0.03239 0.0389 0 1.2641 0.41961 0.12657 0.015883 8.6977 0.099026 0.00012502 0.7911 0.0077524 0.0086325 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15197 0.94812 0.91947 0.0013962 0.99444 0.55711 0.0018811 0.42987 2.0043 2.0037 16.0013 144.9689 0.00015958 -85.6592 0.86794
4.972 0.98808 5.4924e-005 3.8183 0.011979 6.5022e-005 0.0011604 0.23108 0.00065929 0.23173 0.21377 0 0.03239 0.0389 0 1.2642 0.41965 0.12658 0.015885 8.6996 0.099035 0.00012503 0.79109 0.007753 0.0086332 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15198 0.94823 0.91951 0.0013962 0.99446 0.55726 0.001881 0.42989 2.0046 2.0041 16.0013 144.9689 0.00015951 -85.6593 0.86894
4.973 0.98808 5.4924e-005 3.8183 0.011979 6.5035e-005 0.0011604 0.23108 0.00065929 0.23173 0.21377 0 0.03239 0.0389 0 1.2643 0.4197 0.1266 0.015886 8.7015 0.099044 0.00012504 0.79108 0.0077536 0.0086339 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15198 0.94834 0.91956 0.0013962 0.99448 0.55742 0.001881 0.4299 2.005 2.0045 16.0012 144.969 0.00015944 -85.6593 0.86994
4.974 0.98808 5.4924e-005 3.8183 0.011979 6.5048e-005 0.0011604 0.23108 0.00065929 0.23174 0.21377 0 0.03239 0.0389 0 1.2644 0.41975 0.12661 0.015888 8.7034 0.099054 0.00012506 0.79107 0.0077543 0.0086345 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.15199 0.94845 0.9196 0.0013962 0.99449 0.55757 0.001881 0.42991 2.0054 2.0048 16.0012 144.969 0.00015938 -85.6594 0.87094
4.975 0.98808 5.4924e-005 3.8183 0.011979 6.5061e-005 0.0011604 0.23109 0.00065929 0.23174 0.21378 0 0.03239 0.0389 0 1.2644 0.41979 0.12663 0.015889 8.7053 0.099063 0.00012507 0.79106 0.0077549 0.0086352 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.15199 0.94856 0.91964 0.0013962 0.99451 0.55773 0.001881 0.42992 2.0057 2.0052 16.0012 144.969 0.00015931 -85.6594 0.87194
4.976 0.98808 5.4924e-005 3.8183 0.011979 6.5074e-005 0.0011604 0.23109 0.00065929 0.23174 0.21378 0 0.03239 0.0389 0 1.2645 0.41984 0.12664 0.015891 8.7072 0.099072 0.00012508 0.79105 0.0077555 0.0086359 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.152 0.94867 0.91969 0.0013962 0.99453 0.55788 0.001881 0.42993 2.0061 2.0056 16.0011 144.969 0.00015924 -85.6595 0.87294
4.977 0.98808 5.4923e-005 3.8183 0.011979 6.5087e-005 0.0011604 0.23109 0.00065929 0.23175 0.21378 0 0.032389 0.0389 0 1.2646 0.41989 0.12666 0.015892 8.7091 0.099082 0.0001251 0.79104 0.0077561 0.0086366 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.152 0.94878 0.91973 0.0013961 0.99455 0.55803 0.001881 0.42995 2.0065 2.0059 16.0011 144.969 0.00015917 -85.6595 0.87394
4.978 0.98808 5.4923e-005 3.8183 0.011979 6.51e-005 0.0011604 0.23109 0.00065929 0.23175 0.21378 0 0.032389 0.0389 0 1.2647 0.41993 0.12668 0.015894 8.711 0.099091 0.00012511 0.79103 0.0077568 0.0086372 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.15201 0.94889 0.91977 0.0013961 0.99456 0.55819 0.001881 0.42996 2.0068 2.0063 16.0011 144.9691 0.0001591 -85.6596 0.87494
4.979 0.98808 5.4923e-005 3.8183 0.011979 6.5113e-005 0.0011604 0.2311 0.00065929 0.23175 0.21379 0 0.032389 0.0389 0 1.2648 0.41998 0.12669 0.015895 8.7129 0.099101 0.00012512 0.79102 0.0077574 0.0086379 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.15201 0.949 0.91982 0.0013961 0.99458 0.55834 0.001881 0.42997 2.0072 2.0067 16.001 144.9691 0.00015904 -85.6596 0.87594
4.98 0.98808 5.4923e-005 3.8183 0.011978 6.5126e-005 0.0011604 0.2311 0.00065929 0.23175 0.21379 0 0.032389 0.0389 0 1.2649 0.42003 0.12671 0.015897 8.7148 0.09911 0.00012514 0.79102 0.007758 0.0086386 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.15202 0.94911 0.91986 0.0013961 0.9946 0.5585 0.001881 0.42998 2.0076 2.007 16.001 144.9691 0.00015897 -85.6597 0.87694
4.981 0.98808 5.4923e-005 3.8183 0.011978 6.5139e-005 0.0011604 0.2311 0.00065929 0.23176 0.21379 0 0.032389 0.0389 0 1.265 0.42007 0.12672 0.015898 8.7167 0.099119 0.00012515 0.79101 0.0077586 0.0086393 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.15202 0.94921 0.9199 0.0013961 0.99461 0.55865 0.001881 0.43 2.0079 2.0074 16.001 144.9691 0.0001589 -85.6597 0.87794
4.982 0.98808 5.4923e-005 3.8183 0.011978 6.5152e-005 0.0011604 0.23111 0.00065929 0.23176 0.21379 0 0.032389 0.0389 0 1.2651 0.42012 0.12674 0.0159 8.7186 0.099129 0.00012516 0.791 0.0077593 0.0086399 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.15203 0.94932 0.91995 0.0013961 0.99463 0.5588 0.001881 0.43001 2.0083 2.0078 16.0009 144.9691 0.00015884 -85.6598 0.87894
4.983 0.98808 5.4923e-005 3.8183 0.011978 6.5165e-005 0.0011604 0.23111 0.00065929 0.23176 0.2138 0 0.032389 0.0389 0 1.2652 0.42017 0.12675 0.015901 8.7205 0.099138 0.00012518 0.79099 0.0077599 0.0086406 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.15203 0.94943 0.91999 0.0013961 0.99465 0.55896 0.001881 0.43002 2.0086 2.0081 16.0009 144.9692 0.00015877 -85.6598 0.87994
4.984 0.98808 5.4923e-005 3.8183 0.011978 6.5178e-005 0.0011604 0.23111 0.00065929 0.23177 0.2138 0 0.032388 0.0389 0 1.2653 0.42021 0.12677 0.015903 8.7224 0.099147 0.00012519 0.79098 0.0077605 0.0086413 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.15204 0.94953 0.92003 0.0013961 0.99466 0.55911 0.0018809 0.43003 2.009 2.0085 16.0009 144.9692 0.0001587 -85.6599 0.88094
4.985 0.98808 5.4923e-005 3.8183 0.011978 6.5191e-005 0.0011604 0.23111 0.00065929 0.23177 0.2138 0 0.032388 0.0389 0 1.2654 0.42026 0.12678 0.015904 8.7243 0.099157 0.0001252 0.79097 0.0077611 0.008642 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.15204 0.94964 0.92007 0.0013961 0.99468 0.55926 0.0018809 0.43004 2.0094 2.0088 16.0008 144.9692 0.00015864 -85.6599 0.88194
4.986 0.98808 5.4923e-005 3.8183 0.011978 6.5204e-005 0.0011604 0.23112 0.00065929 0.23177 0.21381 0 0.032388 0.0389 0 1.2655 0.42031 0.1268 0.015906 8.7262 0.099166 0.00012522 0.79096 0.0077618 0.0086426 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.15205 0.94975 0.92011 0.0013961 0.9947 0.55942 0.0018809 0.43006 2.0097 2.0092 16.0008 144.9692 0.00015857 -85.66 0.88294
4.987 0.98808 5.4923e-005 3.8183 0.011978 6.5217e-005 0.0011604 0.23112 0.00065929 0.23177 0.21381 0 0.032388 0.0389 0 1.2656 0.42035 0.12682 0.015907 8.7281 0.099175 0.00012523 0.79095 0.0077624 0.0086433 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.15205 0.94985 0.92016 0.0013961 0.99471 0.55957 0.0018809 0.43007 2.0101 2.0096 16.0008 144.9692 0.0001585 -85.66 0.88394
4.988 0.98808 5.4923e-005 3.8183 0.011978 6.523e-005 0.0011604 0.23112 0.00065929 0.23178 0.21381 0 0.032388 0.0389 0 1.2657 0.4204 0.12683 0.015909 8.73 0.099185 0.00012524 0.79094 0.007763 0.008644 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.15206 0.94996 0.9202 0.0013961 0.99473 0.55972 0.0018809 0.43008 2.0104 2.0099 16.0007 144.9693 0.00015844 -85.6601 0.88494
4.989 0.98808 5.4923e-005 3.8183 0.011978 6.5243e-005 0.0011604 0.23113 0.00065929 0.23178 0.21381 0 0.032388 0.0389 0 1.2658 0.42045 0.12685 0.015911 8.7319 0.099194 0.00012526 0.79093 0.0077636 0.0086446 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.15206 0.95006 0.92024 0.0013961 0.99474 0.55988 0.0018809 0.43009 2.0108 2.0103 16.0007 144.9693 0.00015837 -85.6601 0.88594
4.99 0.98808 5.4923e-005 3.8183 0.011978 6.5256e-005 0.0011604 0.23113 0.00065929 0.23178 0.21382 0 0.032388 0.0389 0 1.2659 0.42049 0.12686 0.015912 8.7338 0.099203 0.00012527 0.79092 0.0077643 0.0086453 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.15207 0.95017 0.92028 0.0013961 0.99476 0.56003 0.0018809 0.4301 2.0112 2.0107 16.0007 144.9693 0.00015831 -85.6602 0.88694
4.991 0.98808 5.4922e-005 3.8183 0.011978 6.5269e-005 0.0011604 0.23113 0.00065929 0.23179 0.21382 0 0.032387 0.0389 0 1.266 0.42054 0.12688 0.015914 8.7357 0.099213 0.00012528 0.79091 0.0077649 0.008646 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.15207 0.95027 0.92032 0.0013961 0.99478 0.56018 0.0018809 0.43012 2.0115 2.011 16.0007 144.9693 0.00015824 -85.6602 0.88794
4.992 0.98808 5.4922e-005 3.8183 0.011978 6.5282e-005 0.0011604 0.23113 0.00065929 0.23179 0.21382 0 0.032387 0.0389 0 1.2661 0.42059 0.12689 0.015915 8.7376 0.099222 0.0001253 0.7909 0.0077655 0.0086467 0.0013844 0.98697 0.99172 2.9847e-006 1.1939e-005 0.15208 0.95038 0.92036 0.0013961 0.99479 0.56034 0.0018809 0.43013 2.0119 2.0114 16.0006 144.9693 0.00015818 -85.6603 0.88894
4.993 0.98808 5.4922e-005 3.8183 0.011978 6.5295e-005 0.0011604 0.23114 0.00065929 0.23179 0.21382 0 0.032387 0.0389 0 1.2662 0.42063 0.12691 0.015917 8.7395 0.099231 0.00012531 0.79089 0.0077661 0.0086473 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.15208 0.95048 0.9204 0.0013961 0.99481 0.56049 0.0018809 0.43014 2.0122 2.0117 16.0006 144.9694 0.00015812 -85.6603 0.88994
4.994 0.98808 5.4922e-005 3.8183 0.011978 6.5308e-005 0.0011604 0.23114 0.00065929 0.23179 0.21383 0 0.032387 0.0389 0 1.2663 0.42068 0.12693 0.015918 8.7414 0.099241 0.00012532 0.79088 0.0077668 0.008648 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.15209 0.95058 0.92045 0.001396 0.99482 0.56064 0.0018809 0.43015 2.0126 2.0121 16.0006 144.9694 0.00015805 -85.6604 0.89094
4.995 0.98808 5.4922e-005 3.8183 0.011978 6.5321e-005 0.0011604 0.23114 0.00065929 0.2318 0.21383 0 0.032387 0.0389 0 1.2664 0.42073 0.12694 0.01592 8.7433 0.09925 0.00012534 0.79088 0.0077674 0.0086487 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.15209 0.95069 0.92049 0.001396 0.99484 0.5608 0.0018809 0.43016 2.0129 2.0124 16.0005 144.9694 0.00015799 -85.6604 0.89194
4.996 0.98808 5.4922e-005 3.8183 0.011978 6.5334e-005 0.0011604 0.23115 0.00065929 0.2318 0.21383 0 0.032387 0.0389 0 1.2665 0.42077 0.12696 0.015921 8.7452 0.099259 0.00012535 0.79087 0.007768 0.0086494 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.1521 0.95079 0.92053 0.001396 0.99485 0.56095 0.0018809 0.43018 2.0133 2.0128 16.0005 144.9694 0.00015792 -85.6605 0.89294
4.997 0.98808 5.4922e-005 3.8183 0.011978 6.5347e-005 0.0011604 0.23115 0.00065929 0.2318 0.21383 0 0.032387 0.0389 0 1.2666 0.42082 0.12697 0.015923 8.7471 0.099269 0.00012536 0.79086 0.0077686 0.00865 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.1521 0.95089 0.92057 0.001396 0.99487 0.5611 0.0018808 0.43019 2.0137 2.0131 16.0005 144.9694 0.00015786 -85.6605 0.89394
4.998 0.98808 5.4922e-005 3.8183 0.011978 6.5359e-005 0.0011604 0.23115 0.00065929 0.23181 0.21384 0 0.032386 0.0389 0 1.2667 0.42087 0.12699 0.015924 8.749 0.099278 0.00012538 0.79085 0.0077693 0.0086507 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.15211 0.95099 0.92061 0.001396 0.99488 0.56126 0.0018808 0.4302 2.014 2.0135 16.0004 144.9695 0.0001578 -85.6606 0.89494
4.999 0.98808 5.4922e-005 3.8183 0.011978 6.5372e-005 0.0011604 0.23115 0.00065929 0.23181 0.21384 0 0.032386 0.0389 0 1.2668 0.42091 0.127 0.015926 8.7509 0.099287 0.00012539 0.79084 0.0077699 0.0086514 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.15211 0.95109 0.92065 0.001396 0.9949 0.56141 0.0018808 0.43021 2.0144 2.0139 16.0004 144.9695 0.00015773 -85.6606 0.89594
5 0.98808 5.4922e-005 3.8183 0.011978 6.5385e-005 0.0011604 0.23116 0.00065929 0.23181 0.21384 0 0.032386 0.0389 0 1.2669 0.42096 0.12702 0.015927 8.7528 0.099297 0.0001254 0.79083 0.0077705 0.0086521 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15212 0.9512 0.92069 0.001396 0.99491 0.56156 0.0018808 0.43022 2.0147 2.0142 16.0004 144.9695 0.00015767 -85.6607 0.89694
5.001 0.98808 5.4922e-005 3.8183 0.011978 6.5398e-005 0.0011604 0.23116 0.00065929 0.23181 0.21385 0 0.032386 0.0389 0 1.267 0.42101 0.12703 0.015929 8.7547 0.099306 0.00012541 0.79082 0.0077711 0.0086527 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15212 0.9513 0.92073 0.001396 0.99493 0.56171 0.0018808 0.43024 2.0151 2.0146 16.0003 144.9695 0.00015761 -85.6607 0.89794
5.002 0.98808 5.4922e-005 3.8183 0.011978 6.5411e-005 0.0011604 0.23116 0.00065929 0.23182 0.21385 0 0.032386 0.0389 0 1.267 0.42105 0.12705 0.01593 8.7566 0.099315 0.00012543 0.79081 0.0077718 0.0086534 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15213 0.9514 0.92077 0.001396 0.99494 0.56187 0.0018808 0.43025 2.0154 2.0149 16.0003 144.9696 0.00015755 -85.6607 0.89894
5.003 0.98808 5.4922e-005 3.8183 0.011978 6.5424e-005 0.0011605 0.23116 0.00065929 0.23182 0.21385 0 0.032386 0.0389 0 1.2671 0.4211 0.12707 0.015932 8.7585 0.099325 0.00012544 0.7908 0.0077724 0.0086541 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15213 0.9515 0.92081 0.001396 0.99496 0.56202 0.0018808 0.43026 2.0158 2.0153 16.0003 144.9696 0.00015748 -85.6608 0.89994
5.004 0.98808 5.4921e-005 3.8183 0.011978 6.5437e-005 0.0011605 0.23117 0.00065929 0.23182 0.21385 0 0.032386 0.0389 0 1.2672 0.42115 0.12708 0.015933 8.7604 0.099334 0.00012545 0.79079 0.007773 0.0086547 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15214 0.9516 0.92085 0.001396 0.99497 0.56217 0.0018808 0.43027 2.0161 2.0156 16.0002 144.9696 0.00015742 -85.6608 0.90094
5.005 0.98808 5.4921e-005 3.8183 0.011978 6.545e-005 0.0011605 0.23117 0.00065929 0.23183 0.21386 0 0.032385 0.0389 0 1.2673 0.42119 0.1271 0.015935 8.7623 0.099343 0.00012547 0.79078 0.0077736 0.0086554 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.15214 0.9517 0.92089 0.001396 0.99498 0.56232 0.0018808 0.43028 2.0165 2.016 16.0002 144.9696 0.00015736 -85.6609 0.90194
5.006 0.98808 5.4921e-005 3.8183 0.011978 6.5463e-005 0.0011605 0.23117 0.00065929 0.23183 0.21386 0 0.032385 0.0389 0 1.2674 0.42124 0.12711 0.015936 8.7643 0.099352 0.00012548 0.79077 0.0077742 0.0086561 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.15215 0.9518 0.92093 0.001396 0.995 0.56248 0.0018808 0.4303 2.0168 2.0163 16.0002 144.9696 0.0001573 -85.6609 0.90294
5.007 0.98808 5.4921e-005 3.8183 0.011978 6.5476e-005 0.0011605 0.23118 0.00065929 0.23183 0.21386 0 0.032385 0.0389 0 1.2675 0.42129 0.12713 0.015938 8.7662 0.099362 0.00012549 0.79076 0.0077749 0.0086568 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.15215 0.9519 0.92097 0.001396 0.99501 0.56263 0.0018808 0.43031 2.0172 2.0167 16.0001 144.9697 0.00015724 -85.661 0.90394
5.008 0.98808 5.4921e-005 3.8183 0.011978 6.5489e-005 0.0011605 0.23118 0.00065929 0.23183 0.21386 0 0.032385 0.0389 0 1.2676 0.42133 0.12714 0.015939 8.7681 0.099371 0.00012551 0.79075 0.0077755 0.0086574 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.15216 0.952 0.921 0.001396 0.99503 0.56278 0.0018808 0.43032 2.0175 2.017 16.0001 144.9697 0.00015718 -85.661 0.90494
5.009 0.98808 5.4921e-005 3.8183 0.011978 6.5502e-005 0.0011605 0.23118 0.00065929 0.23184 0.21387 0 0.032385 0.0389 0 1.2677 0.42138 0.12716 0.015941 8.77 0.09938 0.00012552 0.79075 0.0077761 0.0086581 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15216 0.95209 0.92104 0.001396 0.99504 0.56293 0.0018808 0.43033 2.0179 2.0174 16.0001 144.9697 0.00015711 -85.661 0.90594
5.01 0.98808 5.4921e-005 3.8183 0.011978 6.5515e-005 0.0011605 0.23118 0.00065929 0.23184 0.21387 0 0.032385 0.0389 0 1.2678 0.42143 0.12717 0.015942 8.7719 0.09939 0.00012553 0.79074 0.0077767 0.0086588 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15217 0.95219 0.92108 0.001396 0.99506 0.56309 0.0018808 0.43034 2.0182 2.0177 16 144.9697 0.00015705 -85.6611 0.90694
5.011 0.98808 5.4921e-005 3.8183 0.011978 6.5528e-005 0.0011605 0.23119 0.00065929 0.23184 0.21387 0 0.032385 0.0389 0 1.2679 0.42147 0.12719 0.015944 8.7738 0.099399 0.00012555 0.79073 0.0077774 0.0086595 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15217 0.95229 0.92112 0.001396 0.99507 0.56324 0.0018807 0.43036 2.0186 2.0181 16 144.9697 0.00015699 -85.6611 0.90794
5.012 0.98808 5.4921e-005 3.8183 0.011978 6.5541e-005 0.0011605 0.23119 0.00065929 0.23184 0.21387 0 0.032384 0.0389 0 1.268 0.42152 0.12721 0.015945 8.7757 0.099408 0.00012556 0.79072 0.007778 0.0086601 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15218 0.95239 0.92116 0.001396 0.99508 0.56339 0.0018807 0.43037 2.0189 2.0184 16 144.9698 0.00015693 -85.6612 0.90894
5.013 0.98808 5.4921e-005 3.8183 0.011978 6.5554e-005 0.0011605 0.23119 0.00065929 0.23185 0.21388 0 0.032384 0.0389 0 1.2681 0.42157 0.12722 0.015947 8.7776 0.099418 0.00012557 0.79071 0.0077786 0.0086608 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15218 0.95249 0.9212 0.001396 0.9951 0.56354 0.0018807 0.43038 2.0192 2.0187 15.9999 144.9698 0.00015687 -85.6612 0.90994
5.014 0.98808 5.4921e-005 3.8183 0.011978 6.5567e-005 0.0011605 0.2312 0.00065929 0.23185 0.21388 0 0.032384 0.0389 0 1.2682 0.42161 0.12724 0.015948 8.7795 0.099427 0.00012559 0.7907 0.0077792 0.0086615 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.15219 0.95258 0.92124 0.001396 0.99511 0.56369 0.0018807 0.43039 2.0196 2.0191 15.9999 144.9698 0.00015681 -85.6612 0.91094
5.015 0.98808 5.4921e-005 3.8183 0.011978 6.558e-005 0.0011605 0.2312 0.00065929 0.23185 0.21388 0 0.032384 0.0389 0 1.2683 0.42166 0.12725 0.01595 8.7814 0.099436 0.0001256 0.79069 0.0077799 0.0086621 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.15219 0.95268 0.92127 0.0013959 0.99512 0.56385 0.0018807 0.4304 2.0199 2.0194 15.9999 144.9698 0.00015675 -85.6613 0.91194
5.016 0.98808 5.4921e-005 3.8183 0.011978 6.5593e-005 0.0011605 0.2312 0.00065929 0.23186 0.21388 0 0.032384 0.0389 0 1.2684 0.42171 0.12727 0.015951 8.7834 0.099446 0.00012561 0.79068 0.0077805 0.0086628 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.1522 0.95278 0.92131 0.0013959 0.99514 0.564 0.0018807 0.43042 2.0203 2.0198 15.9998 144.9698 0.00015669 -85.6613 0.91294
5.017 0.98808 5.4921e-005 3.8183 0.011978 6.5606e-005 0.0011605 0.2312 0.00065929 0.23186 0.21389 0 0.032384 0.0389 0 1.2685 0.42175 0.12728 0.015953 8.7853 0.099455 0.00012563 0.79067 0.0077811 0.0086635 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.1522 0.95287 0.92135 0.0013959 0.99515 0.56415 0.0018807 0.43043 2.0206 2.0201 15.9998 144.9699 0.00015663 -85.6614 0.91394
5.018 0.98808 5.492e-005 3.8183 0.011978 6.5619e-005 0.0011605 0.23121 0.00065929 0.23186 0.21389 0 0.032384 0.0389 0 1.2686 0.4218 0.1273 0.015954 8.7872 0.099464 0.00012564 0.79066 0.0077817 0.0086642 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.15221 0.95297 0.92139 0.0013959 0.99516 0.5643 0.0018807 0.43044 2.021 2.0205 15.9998 144.9699 0.00015657 -85.6614 0.91494
5.019 0.98808 5.492e-005 3.8183 0.011978 6.5632e-005 0.0011605 0.23121 0.00065929 0.23186 0.21389 0 0.032384 0.0389 0 1.2687 0.42185 0.12731 0.015956 8.7891 0.099474 0.00012565 0.79065 0.0077823 0.0086648 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15221 0.95306 0.92143 0.0013959 0.99518 0.56445 0.0018807 0.43045 2.0213 2.0208 15.9998 144.9699 0.00015652 -85.6614 0.91594
5.02 0.98808 5.492e-005 3.8183 0.011978 6.5645e-005 0.0011605 0.23121 0.00065929 0.23187 0.2139 0 0.032383 0.0389 0 1.2688 0.42189 0.12733 0.015957 8.791 0.099483 0.00012567 0.79064 0.007783 0.0086655 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15222 0.95316 0.92146 0.0013959 0.99519 0.5646 0.0018807 0.43046 2.0216 2.0211 15.9997 144.9699 0.00015646 -85.6615 0.91694
5.021 0.98808 5.492e-005 3.8183 0.011978 6.5658e-005 0.0011605 0.23121 0.00065929 0.23187 0.2139 0 0.032383 0.0389 0 1.2689 0.42194 0.12735 0.015959 8.7929 0.099492 0.00012568 0.79063 0.0077836 0.0086662 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15222 0.95325 0.9215 0.0013959 0.9952 0.56476 0.0018807 0.43048 2.022 2.0215 15.9997 144.9699 0.0001564 -85.6615 0.91794
5.022 0.98808 5.492e-005 3.8183 0.011978 6.5671e-005 0.0011605 0.23122 0.00065929 0.23187 0.2139 0 0.032383 0.0389 0 1.269 0.42198 0.12736 0.015961 8.7948 0.099501 0.00012569 0.79062 0.0077842 0.0086668 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15223 0.95335 0.92154 0.0013959 0.99521 0.56491 0.0018807 0.43049 2.0223 2.0218 15.9997 144.97 0.00015634 -85.6616 0.91894
5.023 0.98808 5.492e-005 3.8183 0.011978 6.5684e-005 0.0011605 0.23122 0.00065929 0.23187 0.2139 0 0.032383 0.0389 0 1.2691 0.42203 0.12738 0.015962 8.7967 0.099511 0.00012571 0.79061 0.0077848 0.0086675 0.001384 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15223 0.95344 0.92158 0.0013959 0.99523 0.56506 0.0018807 0.4305 2.0227 2.0222 15.9996 144.97 0.00015628 -85.6616 0.91994
5.024 0.98808 5.492e-005 3.8183 0.011978 6.5697e-005 0.0011605 0.23122 0.00065929 0.23188 0.21391 0 0.032383 0.0389 0 1.2692 0.42208 0.12739 0.015964 8.7987 0.09952 0.00012572 0.79061 0.0077855 0.0086682 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.15224 0.95354 0.92161 0.0013959 0.99524 0.56521 0.0018807 0.43051 2.023 2.0225 15.9996 144.97 0.00015622 -85.6616 0.92094
5.025 0.98808 5.492e-005 3.8183 0.011978 6.571e-005 0.0011605 0.23123 0.00065929 0.23188 0.21391 0 0.032383 0.0389 0 1.2693 0.42212 0.12741 0.015965 8.8006 0.099529 0.00012573 0.7906 0.0077861 0.0086689 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.15224 0.95363 0.92165 0.0013959 0.99525 0.56536 0.0018807 0.43052 2.0233 2.0228 15.9996 144.97 0.00015617 -85.6617 0.92194
5.026 0.98808 5.492e-005 3.8183 0.011978 6.5722e-005 0.0011605 0.23123 0.00065929 0.23188 0.21391 0 0.032383 0.0389 0 1.2694 0.42217 0.12742 0.015967 8.8025 0.099539 0.00012575 0.79059 0.0077867 0.0086695 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.15225 0.95372 0.92169 0.0013959 0.99527 0.56551 0.0018807 0.43054 2.0237 2.0232 15.9995 144.97 0.00015611 -85.6617 0.92294
5.027 0.98808 5.492e-005 3.8183 0.011978 6.5735e-005 0.0011605 0.23123 0.00065929 0.23189 0.21391 0 0.032382 0.0389 0 1.2695 0.42222 0.12744 0.015968 8.8044 0.099548 0.00012576 0.79058 0.0077873 0.0086702 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.15225 0.95382 0.92172 0.0013959 0.99528 0.56566 0.0018806 0.43055 2.024 2.0235 15.9995 144.9701 0.00015605 -85.6617 0.92394
5.028 0.98808 5.492e-005 3.8183 0.011978 6.5748e-005 0.0011605 0.23123 0.00065929 0.23189 0.21392 0 0.032382 0.0389 0 1.2695 0.42226 0.12746 0.01597 8.8063 0.099557 0.00012577 0.79057 0.0077879 0.0086709 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.15226 0.95391 0.92176 0.0013959 0.99529 0.56582 0.0018806 0.43056 2.0243 2.0239 15.9995 144.9701 0.00015599 -85.6618 0.92494
5.029 0.98808 5.492e-005 3.8183 0.011978 6.5761e-005 0.0011605 0.23124 0.00065929 0.23189 0.21392 0 0.032382 0.0389 0 1.2696 0.42231 0.12747 0.015971 8.8082 0.099567 0.00012579 0.79056 0.0077886 0.0086715 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.15226 0.954 0.9218 0.0013959 0.9953 0.56597 0.0018806 0.43057 2.0247 2.0242 15.9994 144.9701 0.00015594 -85.6618 0.92594
5.03 0.98808 5.492e-005 3.8183 0.011978 6.5774e-005 0.0011605 0.23124 0.00065929 0.23189 0.21392 0 0.032382 0.0389 0 1.2697 0.42236 0.12749 0.015973 8.8101 0.099576 0.0001258 0.79055 0.0077892 0.0086722 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.15227 0.95409 0.92183 0.0013959 0.99531 0.56612 0.0018806 0.43058 2.025 2.0245 15.9994 144.9701 0.00015588 -85.6618 0.92694
5.031 0.98808 5.4919e-005 3.8183 0.011978 6.5787e-005 0.0011605 0.23124 0.00065929 0.2319 0.21392 0 0.032382 0.0389 0 1.2698 0.4224 0.1275 0.015974 8.8121 0.099585 0.00012581 0.79054 0.0077898 0.0086729 0.001384 0.98697 0.99172 2.9839e-006 1.1936e-005 0.15227 0.95419 0.92187 0.0013959 0.99533 0.56627 0.0018806 0.4306 2.0253 2.0249 15.9994 144.9701 0.00015582 -85.6619 0.92794
5.032 0.98808 5.4919e-005 3.8183 0.011978 6.58e-005 0.0011605 0.23124 0.00065929 0.2319 0.21393 0 0.032382 0.0389 0 1.2699 0.42245 0.12752 0.015976 8.814 0.099594 0.00012583 0.79053 0.0077904 0.0086735 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.15228 0.95428 0.9219 0.0013959 0.99534 0.56642 0.0018806 0.43061 2.0257 2.0252 15.9993 144.9702 0.00015577 -85.6619 0.92894
5.033 0.98808 5.4919e-005 3.8183 0.011978 6.5813e-005 0.0011605 0.23125 0.00065929 0.2319 0.21393 0 0.032382 0.0389 0 1.27 0.4225 0.12753 0.015977 8.8159 0.099604 0.00012584 0.79052 0.0077911 0.0086742 0.001384 0.98697 0.99172 2.9839e-006 1.1935e-005 0.15228 0.95437 0.92194 0.0013959 0.99535 0.56657 0.0018806 0.43062 2.026 2.0255 15.9993 144.9702 0.00015571 -85.6619 0.92994
5.034 0.98808 5.4919e-005 3.8183 0.011978 6.5826e-005 0.0011605 0.23125 0.00065929 0.23191 0.21393 0 0.032381 0.0389 0 1.2701 0.42254 0.12755 0.015979 8.8178 0.099613 0.00012585 0.79051 0.0077917 0.0086749 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.15229 0.95446 0.92198 0.0013959 0.99536 0.56672 0.0018806 0.43063 2.0263 2.0259 15.9993 144.9702 0.00015565 -85.662 0.93094
5.035 0.98808 5.4919e-005 3.8183 0.011978 6.5839e-005 0.0011605 0.23125 0.00065929 0.23191 0.21393 0 0.032381 0.0389 0 1.2702 0.42259 0.12756 0.01598 8.8197 0.099622 0.00012586 0.7905 0.0077923 0.0086756 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.15229 0.95455 0.92201 0.0013958 0.99537 0.56687 0.0018806 0.43064 2.0267 2.0262 15.9992 144.9702 0.0001556 -85.662 0.93194
5.036 0.98808 5.4919e-005 3.8183 0.011978 6.5852e-005 0.0011605 0.23126 0.00065929 0.23191 0.21394 0 0.032381 0.0389 0 1.2703 0.42264 0.12758 0.015982 8.8217 0.099632 0.00012588 0.79049 0.0077929 0.0086762 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.1523 0.95464 0.92205 0.0013958 0.99539 0.56702 0.0018806 0.43065 2.027 2.0265 15.9992 144.9703 0.00015554 -85.6621 0.93294
5.037 0.98808 5.4919e-005 3.8183 0.011978 6.5865e-005 0.0011606 0.23126 0.00065929 0.23191 0.21394 0 0.032381 0.0389 0 1.2704 0.42268 0.1276 0.015983 8.8236 0.099641 0.00012589 0.79048 0.0077935 0.0086769 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.1523 0.95473 0.92208 0.0013958 0.9954 0.56717 0.0018806 0.43067 2.0273 2.0269 15.9992 144.9703 0.00015549 -85.6621 0.93394
5.038 0.98808 5.4919e-005 3.8183 0.011978 6.5878e-005 0.0011606 0.23126 0.00065929 0.23192 0.21394 0 0.032381 0.0389 0 1.2705 0.42273 0.12761 0.015985 8.8255 0.09965 0.0001259 0.79048 0.0077942 0.0086776 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.15231 0.95482 0.92212 0.0013958 0.99541 0.56733 0.0018806 0.43068 2.0277 2.0272 15.9991 144.9703 0.00015543 -85.6621 0.93494
5.039 0.98808 5.4919e-005 3.8183 0.011978 6.5891e-005 0.0011606 0.23126 0.00065929 0.23192 0.21394 0 0.032381 0.0389 0 1.2706 0.42278 0.12763 0.015986 8.8274 0.099659 0.00012592 0.79047 0.0077948 0.0086782 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.15231 0.95491 0.92215 0.0013958 0.99542 0.56748 0.0018806 0.43069 2.028 2.0275 15.9991 144.9703 0.00015537 -85.6621 0.93594
5.04 0.98808 5.4919e-005 3.8183 0.011978 6.5904e-005 0.0011606 0.23127 0.00065929 0.23192 0.21395 0 0.032381 0.0389 0 1.2707 0.42282 0.12764 0.015988 8.8293 0.099669 0.00012593 0.79046 0.0077954 0.0086789 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15232 0.955 0.92219 0.0013958 0.99543 0.56763 0.0018806 0.4307 2.0283 2.0279 15.9991 144.9703 0.00015532 -85.6622 0.93694
5.041 0.98808 5.4919e-005 3.8183 0.011978 6.5917e-005 0.0011606 0.23127 0.00065929 0.23192 0.21395 0 0.03238 0.0389 0 1.2708 0.42287 0.12766 0.015989 8.8313 0.099678 0.00012594 0.79045 0.007796 0.0086796 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15232 0.95509 0.92222 0.0013958 0.99544 0.56778 0.0018806 0.43071 2.0287 2.0282 15.999 144.9704 0.00015526 -85.6622 0.93794
5.042 0.98808 5.4919e-005 3.8183 0.011978 6.593e-005 0.0011606 0.23127 0.00065929 0.23193 0.21395 0 0.03238 0.0389 0 1.2709 0.42292 0.12767 0.015991 8.8332 0.099687 0.00012596 0.79044 0.0077966 0.0086802 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15232 0.95518 0.92226 0.0013958 0.99545 0.56793 0.0018806 0.43073 2.029 2.0285 15.999 144.9704 0.00015521 -85.6622 0.93894
5.043 0.98808 5.4919e-005 3.8183 0.011977 6.5943e-005 0.0011606 0.23127 0.00065929 0.23193 0.21395 0 0.03238 0.0389 0 1.271 0.42296 0.12769 0.015992 8.8351 0.099697 0.00012597 0.79043 0.0077973 0.0086809 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15233 0.95527 0.92229 0.0013958 0.99547 0.56808 0.0018806 0.43074 2.0293 2.0289 15.999 144.9704 0.00015516 -85.6623 0.93994
5.044 0.98808 5.4919e-005 3.8183 0.011977 6.5956e-005 0.0011606 0.23128 0.00065929 0.23193 0.21396 0 0.03238 0.0389 0 1.2711 0.42301 0.1277 0.015994 8.837 0.099706 0.00012598 0.79042 0.0077979 0.0086816 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15233 0.95536 0.92233 0.0013958 0.99548 0.56823 0.0018806 0.43075 2.0297 2.0292 15.9989 144.9704 0.0001551 -85.6623 0.94094
5.045 0.98808 5.4918e-005 3.8183 0.011977 6.5969e-005 0.0011606 0.23128 0.00065929 0.23193 0.21396 0 0.03238 0.0389 0 1.2712 0.42306 0.12772 0.015995 8.8389 0.099715 0.000126 0.79041 0.0077985 0.0086822 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15234 0.95544 0.92236 0.0013958 0.99549 0.56838 0.0018806 0.43076 2.03 2.0295 15.9989 144.9704 0.00015505 -85.6623 0.94194
5.046 0.98808 5.4918e-005 3.8183 0.011977 6.5982e-005 0.0011606 0.23128 0.00065929 0.23194 0.21396 0 0.03238 0.0389 0 1.2713 0.4231 0.12774 0.015997 8.8409 0.099724 0.00012601 0.7904 0.0077991 0.0086829 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.15234 0.95553 0.9224 0.0013958 0.9955 0.56853 0.0018805 0.43077 2.0303 2.0298 15.9989 144.9705 0.00015499 -85.6624 0.94294
5.047 0.98808 5.4918e-005 3.8183 0.011977 6.5995e-005 0.0011606 0.23129 0.00065929 0.23194 0.21397 0 0.03238 0.0389 0 1.2714 0.42315 0.12775 0.015998 8.8428 0.099734 0.00012602 0.79039 0.0077997 0.0086836 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.15235 0.95562 0.92243 0.0013958 0.99551 0.56868 0.0018805 0.43078 2.0306 2.0302 15.9988 144.9705 0.00015494 -85.6624 0.94394
5.048 0.98808 5.4918e-005 3.8183 0.011977 6.6008e-005 0.0011606 0.23129 0.00065929 0.23194 0.21397 0 0.03238 0.0389 0 1.2715 0.4232 0.12777 0.016 8.8447 0.099743 0.00012604 0.79038 0.0078004 0.0086843 0.0013838 0.98697 0.99172 2.9836e-006 1.1934e-005 0.15235 0.95571 0.92247 0.0013958 0.99552 0.56883 0.0018805 0.4308 2.031 2.0305 15.9988 144.9705 0.00015489 -85.6624 0.94494
5.049 0.98808 5.4918e-005 3.8183 0.011977 6.6021e-005 0.0011606 0.23129 0.00065929 0.23195 0.21397 0 0.032379 0.0389 0 1.2716 0.42324 0.12778 0.016001 8.8466 0.099752 0.00012605 0.79037 0.007801 0.0086849 0.0013838 0.98698 0.99172 2.9836e-006 1.1934e-005 0.15236 0.95579 0.9225 0.0013958 0.99553 0.56898 0.0018805 0.43081 2.0313 2.0308 15.9988 144.9705 0.00015483 -85.6625 0.94594
5.05 0.98808 5.4918e-005 3.8183 0.011977 6.6034e-005 0.0011606 0.23129 0.00065929 0.23195 0.21397 0 0.032379 0.0389 0 1.2717 0.42329 0.1278 0.016003 8.8486 0.099762 0.00012606 0.79036 0.0078016 0.0086856 0.0013839 0.98698 0.99172 2.9836e-006 1.1934e-005 0.15236 0.95588 0.92253 0.0013958 0.99554 0.56913 0.0018805 0.43082 2.0316 2.0311 15.9987 144.9705 0.00015478 -85.6625 0.94694
5.051 0.98808 5.4918e-005 3.8183 0.011977 6.6047e-005 0.0011606 0.2313 0.00065929 0.23195 0.21398 0 0.032379 0.0389 0 1.2718 0.42334 0.12781 0.016004 8.8505 0.099771 0.00012608 0.79036 0.0078022 0.0086863 0.0013839 0.98698 0.99172 2.9836e-006 1.1934e-005 0.15237 0.95597 0.92257 0.0013958 0.99555 0.56928 0.0018805 0.43083 2.0319 2.0315 15.9987 144.9706 0.00015473 -85.6625 0.94794
5.052 0.98808 5.4918e-005 3.8183 0.011977 6.606e-005 0.0011606 0.2313 0.00065929 0.23195 0.21398 0 0.032379 0.0389 0 1.2719 0.42338 0.12783 0.016006 8.8524 0.09978 0.00012609 0.79035 0.0078028 0.0086869 0.0013838 0.98698 0.99172 2.9836e-006 1.1934e-005 0.15237 0.95605 0.9226 0.0013958 0.99556 0.56943 0.0018805 0.43084 2.0323 2.0318 15.9987 144.9706 0.00015467 -85.6625 0.94894
5.053 0.98808 5.4918e-005 3.8183 0.011977 6.6072e-005 0.0011606 0.2313 0.00065929 0.23196 0.21398 0 0.032379 0.0389 0 1.272 0.42343 0.12784 0.016007 8.8543 0.099789 0.0001261 0.79034 0.0078035 0.0086876 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.15238 0.95614 0.92263 0.0013958 0.99557 0.56958 0.0018805 0.43085 2.0326 2.0321 15.9986 144.9706 0.00015462 -85.6626 0.94994
5.054 0.98808 5.4918e-005 3.8183 0.011977 6.6085e-005 0.0011606 0.2313 0.00065929 0.23196 0.21398 0 0.032379 0.0389 0 1.272 0.42348 0.12786 0.016009 8.8562 0.099799 0.00012612 0.79033 0.0078041 0.0086883 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.15238 0.95623 0.92267 0.0013958 0.99558 0.56973 0.0018805 0.43087 2.0329 2.0324 15.9986 144.9706 0.00015457 -85.6626 0.95094
5.055 0.98808 5.4918e-005 3.8183 0.011977 6.6098e-005 0.0011606 0.23131 0.00065929 0.23196 0.21399 0 0.032379 0.0389 0 1.2721 0.42352 0.12788 0.01601 8.8582 0.099808 0.00012613 0.79032 0.0078047 0.0086889 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.15239 0.95631 0.9227 0.0013958 0.99559 0.56988 0.0018805 0.43088 2.0332 2.0328 15.9986 144.9706 0.00015451 -85.6626 0.95194
5.056 0.98808 5.4918e-005 3.8183 0.011977 6.6111e-005 0.0011606 0.23131 0.00065929 0.23196 0.21399 0 0.032378 0.0389 0 1.2722 0.42357 0.12789 0.016012 8.8601 0.099817 0.00012614 0.79031 0.0078053 0.0086896 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.15239 0.9564 0.92273 0.0013958 0.9956 0.57003 0.0018805 0.43089 2.0335 2.0331 15.9985 144.9707 0.00015446 -85.6627 0.95294
5.057 0.98808 5.4918e-005 3.8183 0.011977 6.6124e-005 0.0011606 0.23131 0.00065929 0.23197 0.21399 0 0.032378 0.0389 0 1.2723 0.42362 0.12791 0.016013 8.862 0.099826 0.00012616 0.7903 0.0078059 0.0086903 0.0013838 0.98698 0.99172 2.9835e-006 1.1934e-005 0.1524 0.95648 0.92277 0.0013958 0.99561 0.57018 0.0018805 0.4309 2.0339 2.0334 15.9985 144.9707 0.00015441 -85.6627 0.95394
5.058 0.98808 5.4917e-005 3.8183 0.011977 6.6137e-005 0.0011606 0.23131 0.00065929 0.23197 0.21399 0 0.032378 0.0389 0 1.2724 0.42366 0.12792 0.016015 8.864 0.099836 0.00012617 0.79029 0.0078066 0.0086909 0.0013838 0.98698 0.99173 2.9835e-006 1.1934e-005 0.1524 0.95657 0.9228 0.0013958 0.99562 0.57033 0.0018805 0.43091 2.0342 2.0337 15.9985 144.9707 0.00015436 -85.6627 0.95494
5.059 0.98808 5.4917e-005 3.8183 0.011977 6.615e-005 0.0011606 0.23132 0.00065929 0.23197 0.214 0 0.032378 0.0389 0 1.2725 0.42371 0.12794 0.016016 8.8659 0.099845 0.00012618 0.79028 0.0078072 0.0086916 0.0013838 0.98698 0.99173 2.9834e-006 1.1934e-005 0.15241 0.95665 0.92283 0.0013958 0.99563 0.57048 0.0018805 0.43093 2.0345 2.0341 15.9984 144.9707 0.00015431 -85.6627 0.95594
5.06 0.98808 5.4917e-005 3.8183 0.011977 6.6163e-005 0.0011606 0.23132 0.00065929 0.23197 0.214 0 0.032378 0.0389 0 1.2726 0.42376 0.12795 0.016018 8.8678 0.099854 0.00012619 0.79027 0.0078078 0.0086923 0.0013838 0.98698 0.99173 2.9834e-006 1.1934e-005 0.15241 0.95673 0.92287 0.0013958 0.99564 0.57063 0.0018805 0.43094 2.0348 2.0344 15.9984 144.9707 0.00015425 -85.6628 0.95694
5.061 0.98808 5.4917e-005 3.8183 0.011977 6.6176e-005 0.0011606 0.23132 0.00065929 0.23198 0.214 0 0.032378 0.0389 0 1.2727 0.4238 0.12797 0.016019 8.8697 0.099864 0.00012621 0.79026 0.0078084 0.0086929 0.0013838 0.98698 0.99173 2.9834e-006 1.1934e-005 0.15242 0.95682 0.9229 0.0013958 0.99565 0.57078 0.0018805 0.43095 2.0351 2.0347 15.9984 144.9708 0.0001542 -85.6628 0.95794
5.062 0.98808 5.4917e-005 3.8183 0.011977 6.6189e-005 0.0011606 0.23133 0.00065929 0.23198 0.214 0 0.032378 0.0389 0 1.2728 0.42385 0.12798 0.016021 8.8717 0.099873 0.00012622 0.79025 0.007809 0.0086936 0.0013838 0.98698 0.99173 2.9834e-006 1.1934e-005 0.15242 0.9569 0.92293 0.0013958 0.99566 0.57093 0.0018805 0.43096 2.0355 2.035 15.9983 144.9708 0.00015415 -85.6628 0.95894
5.063 0.98808 5.4917e-005 3.8183 0.011977 6.6202e-005 0.0011606 0.23133 0.00065929 0.23198 0.21401 0 0.032378 0.0389 0 1.2729 0.42389 0.128 0.016022 8.8736 0.099882 0.00012623 0.79024 0.0078096 0.0086943 0.0013838 0.98698 0.99173 2.9834e-006 1.1933e-005 0.15243 0.95698 0.92296 0.0013958 0.99567 0.57108 0.0018805 0.43097 2.0358 2.0353 15.9983 144.9708 0.0001541 -85.6629 0.95994
5.064 0.98808 5.4917e-005 3.8183 0.011977 6.6215e-005 0.0011606 0.23133 0.00065929 0.23199 0.21401 0 0.032377 0.0389 0 1.273 0.42394 0.12802 0.016024 8.8755 0.099891 0.00012625 0.79023 0.0078103 0.0086949 0.0013838 0.98698 0.99173 2.9834e-006 1.1933e-005 0.15243 0.95707 0.923 0.0013958 0.99568 0.57123 0.0018805 0.43098 2.0361 2.0356 15.9983 144.9708 0.00015405 -85.6629 0.96094
5.065 0.98808 5.4917e-005 3.8183 0.011977 6.6228e-005 0.0011606 0.23133 0.00065929 0.23199 0.21401 0 0.032377 0.0389 0 1.2731 0.42399 0.12803 0.016025 8.8774 0.099901 0.00012626 0.79023 0.0078109 0.0086956 0.0013837 0.98698 0.99173 2.9834e-006 1.1933e-005 0.15244 0.95715 0.92303 0.0013957 0.99569 0.57138 0.0018805 0.431 2.0364 2.036 15.9982 144.9708 0.000154 -85.6629 0.96194
5.066 0.98808 5.4917e-005 3.8183 0.011977 6.6241e-005 0.0011606 0.23134 0.00065929 0.23199 0.21401 0 0.032377 0.0389 0 1.2732 0.42403 0.12805 0.016027 8.8794 0.09991 0.00012627 0.79022 0.0078115 0.0086963 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15244 0.95723 0.92306 0.0013957 0.9957 0.57152 0.0018805 0.43101 2.0367 2.0363 15.9982 144.9709 0.00015395 -85.6629 0.96294
5.067 0.98808 5.4917e-005 3.8183 0.011977 6.6254e-005 0.0011606 0.23134 0.00065929 0.23199 0.21402 0 0.032377 0.0389 0 1.2733 0.42408 0.12806 0.016028 8.8813 0.099919 0.00012629 0.79021 0.0078121 0.0086969 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15245 0.95731 0.92309 0.0013957 0.99571 0.57167 0.0018805 0.43102 2.0371 2.0366 15.9982 144.9709 0.0001539 -85.663 0.96394
5.068 0.98808 5.4917e-005 3.8183 0.011977 6.6267e-005 0.0011606 0.23134 0.00065929 0.232 0.21402 0 0.032377 0.0389 0 1.2734 0.42413 0.12808 0.01603 8.8832 0.099928 0.0001263 0.7902 0.0078127 0.0086976 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15245 0.9574 0.92313 0.0013957 0.99572 0.57182 0.0018804 0.43103 2.0374 2.0369 15.9981 144.9709 0.00015385 -85.663 0.96494
5.069 0.98808 5.4917e-005 3.8183 0.011977 6.628e-005 0.0011606 0.23134 0.00065929 0.232 0.21402 0 0.032377 0.0389 0 1.2735 0.42417 0.12809 0.016031 8.8852 0.099938 0.00012631 0.79019 0.0078134 0.0086983 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15246 0.95748 0.92316 0.0013957 0.99573 0.57197 0.0018804 0.43104 2.0377 2.0372 15.9981 144.9709 0.0001538 -85.663 0.96594
5.07 0.98808 5.4917e-005 3.8183 0.011977 6.6293e-005 0.0011606 0.23135 0.00065929 0.232 0.21402 0 0.032377 0.0389 0 1.2736 0.42422 0.12811 0.016033 8.8871 0.099947 0.00012633 0.79018 0.007814 0.0086989 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15246 0.95756 0.92319 0.0013957 0.99574 0.57212 0.0018804 0.43105 2.038 2.0376 15.9981 144.971 0.00015375 -85.663 0.96694
5.071 0.98808 5.4917e-005 3.8183 0.011977 6.6306e-005 0.0011607 0.23135 0.00065929 0.232 0.21403 0 0.032376 0.0389 0 1.2737 0.42427 0.12812 0.016034 8.889 0.099956 0.00012634 0.79017 0.0078146 0.0086996 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15247 0.95764 0.92322 0.0013957 0.99575 0.57227 0.0018804 0.43107 2.0383 2.0379 15.998 144.971 0.0001537 -85.6631 0.96794
5.072 0.98808 5.4916e-005 3.8183 0.011977 6.6319e-005 0.0011607 0.23135 0.00065929 0.23201 0.21403 0 0.032376 0.0389 0 1.2738 0.42431 0.12814 0.016036 8.891 0.099965 0.00012635 0.79016 0.0078152 0.0087003 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15247 0.95772 0.92325 0.0013957 0.99576 0.57242 0.0018804 0.43108 2.0386 2.0382 15.998 144.971 0.00015365 -85.6631 0.96894
5.073 0.98808 5.4916e-005 3.8183 0.011977 6.6332e-005 0.0011607 0.23135 0.00065929 0.23201 0.21403 0 0.032376 0.0389 0 1.2739 0.42436 0.12816 0.016037 8.8929 0.099975 0.00012637 0.79015 0.0078158 0.0087009 0.0013837 0.98698 0.99173 2.9833e-006 1.1933e-005 0.15248 0.9578 0.92328 0.0013957 0.99577 0.57257 0.0018804 0.43109 2.0389 2.0385 15.998 144.971 0.0001536 -85.6631 0.96994
5.074 0.98808 5.4916e-005 3.8183 0.011977 6.6345e-005 0.0011607 0.23136 0.00065929 0.23201 0.21403 0 0.032376 0.0389 0 1.274 0.42441 0.12817 0.016039 8.8948 0.099984 0.00012638 0.79014 0.0078164 0.0087016 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.15248 0.95788 0.92332 0.0013957 0.99578 0.57272 0.0018804 0.4311 2.0393 2.0388 15.9979 144.971 0.00015355 -85.6631 0.97094
5.075 0.98808 5.4916e-005 3.8183 0.011977 6.6358e-005 0.0011607 0.23136 0.00065929 0.23201 0.21404 0 0.032376 0.0389 0 1.2741 0.42445 0.12819 0.01604 8.8968 0.099993 0.00012639 0.79013 0.0078171 0.0087023 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.15249 0.95796 0.92335 0.0013957 0.99579 0.57287 0.0018804 0.43111 2.0396 2.0391 15.9979 144.9711 0.0001535 -85.6632 0.97194
5.076 0.98808 5.4916e-005 3.8183 0.011977 6.6371e-005 0.0011607 0.23136 0.00065929 0.23202 0.21404 0 0.032376 0.0389 0 1.2742 0.4245 0.1282 0.016042 8.8987 0.1 0.00012641 0.79012 0.0078177 0.0087029 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.15249 0.95804 0.92338 0.0013957 0.9958 0.57301 0.0018804 0.43112 2.0399 2.0394 15.9979 144.9711 0.00015345 -85.6632 0.97294
5.077 0.98808 5.4916e-005 3.8183 0.011977 6.6384e-005 0.0011607 0.23136 0.00065929 0.23202 0.21404 0 0.032376 0.0389 0 1.2743 0.42455 0.12822 0.016043 8.9006 0.10001 0.00012642 0.79011 0.0078183 0.0087036 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.1525 0.95812 0.92341 0.0013957 0.99581 0.57316 0.0018804 0.43114 2.0402 2.0397 15.9978 144.9711 0.0001534 -85.6632 0.97394
5.078 0.98808 5.4916e-005 3.8183 0.011977 6.6397e-005 0.0011607 0.23137 0.00065929 0.23202 0.21404 0 0.032376 0.0389 0 1.2744 0.42459 0.12823 0.016045 8.9026 0.10002 0.00012643 0.79011 0.0078189 0.0087043 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.1525 0.9582 0.92344 0.0013957 0.99581 0.57331 0.0018804 0.43115 2.0405 2.0401 15.9978 144.9711 0.00015335 -85.6632 0.97494
5.079 0.98808 5.4916e-005 3.8183 0.011977 6.6409e-005 0.0011607 0.23137 0.00065929 0.23202 0.21405 0 0.032375 0.0389 0 1.2744 0.42464 0.12825 0.016046 8.9045 0.10003 0.00012644 0.7901 0.0078195 0.0087049 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.15251 0.95828 0.92347 0.0013957 0.99582 0.57346 0.0018804 0.43116 2.0408 2.0404 15.9978 144.9711 0.00015331 -85.6632 0.97594
5.08 0.98808 5.4916e-005 3.8183 0.011977 6.6422e-005 0.0011607 0.23137 0.00065929 0.23203 0.21405 0 0.032375 0.0389 0 1.2745 0.42469 0.12826 0.016048 8.9064 0.10004 0.00012646 0.79009 0.0078202 0.0087056 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.15251 0.95836 0.9235 0.0013957 0.99583 0.57361 0.0018804 0.43117 2.0411 2.0407 15.9977 144.9712 0.00015326 -85.6633 0.97694
5.081 0.98808 5.4916e-005 3.8183 0.011977 6.6435e-005 0.0011607 0.23138 0.00065929 0.23203 0.21405 0 0.032375 0.0389 0 1.2746 0.42473 0.12828 0.016049 8.9084 0.10005 0.00012647 0.79008 0.0078208 0.0087063 0.0013837 0.98698 0.99173 2.9832e-006 1.1933e-005 0.15252 0.95844 0.92353 0.0013957 0.99584 0.57376 0.0018804 0.43118 2.0414 2.041 15.9977 144.9712 0.00015321 -85.6633 0.97794
5.082 0.98808 5.4916e-005 3.8183 0.011977 6.6448e-005 0.0011607 0.23138 0.00065929 0.23203 0.21405 0 0.032375 0.0389 0 1.2747 0.42478 0.1283 0.016051 8.9103 0.10006 0.00012648 0.79007 0.0078214 0.0087069 0.0013837 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15252 0.95852 0.92356 0.0013957 0.99585 0.57391 0.0018804 0.43119 2.0417 2.0413 15.9977 144.9712 0.00015316 -85.6633 0.97894
5.083 0.98808 5.4916e-005 3.8183 0.011977 6.6461e-005 0.0011607 0.23138 0.00065929 0.23204 0.21406 0 0.032375 0.0389 0 1.2748 0.42483 0.12831 0.016052 8.9122 0.10007 0.0001265 0.79006 0.007822 0.0087076 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15253 0.9586 0.92359 0.0013957 0.99586 0.57405 0.0018804 0.4312 2.042 2.0416 15.9976 144.9712 0.00015311 -85.6633 0.97994
5.084 0.98808 5.4916e-005 3.8183 0.011977 6.6474e-005 0.0011607 0.23138 0.00065929 0.23204 0.21406 0 0.032375 0.0389 0 1.2749 0.42487 0.12833 0.016054 8.9142 0.10008 0.00012651 0.79005 0.0078226 0.0087083 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15253 0.95867 0.92362 0.0013957 0.99587 0.5742 0.0018804 0.43122 2.0424 2.0419 15.9976 144.9712 0.00015307 -85.6634 0.98094
5.085 0.98808 5.4915e-005 3.8183 0.011977 6.6487e-005 0.0011607 0.23139 0.00065929 0.23204 0.21406 0 0.032375 0.0389 0 1.275 0.42492 0.12834 0.016055 8.9161 0.10009 0.00012652 0.79004 0.0078232 0.0087089 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15254 0.95875 0.92365 0.0013957 0.99587 0.57435 0.0018804 0.43123 2.0427 2.0422 15.9976 144.9713 0.00015302 -85.6634 0.98194
5.086 0.98808 5.4915e-005 3.8183 0.011977 6.65e-005 0.0011607 0.23139 0.00065929 0.23204 0.21406 0 0.032375 0.0389 0 1.2751 0.42497 0.12836 0.016057 8.918 0.10009 0.00012654 0.79003 0.0078239 0.0087096 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15254 0.95883 0.92369 0.0013957 0.99588 0.5745 0.0018804 0.43124 2.043 2.0425 15.9975 144.9713 0.00015297 -85.6634 0.98294
5.087 0.98808 5.4915e-005 3.8183 0.011977 6.6513e-005 0.0011607 0.23139 0.00065929 0.23205 0.21407 0 0.032374 0.0389 0 1.2752 0.42501 0.12837 0.016058 8.92 0.1001 0.00012655 0.79002 0.0078245 0.0087103 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15255 0.95891 0.92372 0.0013957 0.99589 0.57465 0.0018804 0.43125 2.0433 2.0428 15.9975 144.9713 0.00015292 -85.6634 0.98394
5.088 0.98808 5.4915e-005 3.8183 0.011977 6.6526e-005 0.0011607 0.23139 0.00065929 0.23205 0.21407 0 0.032374 0.0389 0 1.2753 0.42506 0.12839 0.01606 8.9219 0.10011 0.00012656 0.79001 0.0078251 0.0087109 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15255 0.95898 0.92375 0.0013957 0.9959 0.5748 0.0018804 0.43126 2.0436 2.0432 15.9975 144.9713 0.00015288 -85.6634 0.98494
5.089 0.98808 5.4915e-005 3.8183 0.011977 6.6539e-005 0.0011607 0.2314 0.00065929 0.23205 0.21407 0 0.032374 0.0389 0 1.2754 0.42511 0.1284 0.016061 8.9238 0.10012 0.00012658 0.79 0.0078257 0.0087116 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15256 0.95906 0.92378 0.0013957 0.99591 0.57494 0.0018804 0.43127 2.0439 2.0435 15.9974 144.9713 0.00015283 -85.6635 0.98594
5.09 0.98808 5.4915e-005 3.8183 0.011977 6.6552e-005 0.0011607 0.2314 0.00065929 0.23205 0.21407 0 0.032374 0.0389 0 1.2755 0.42515 0.12842 0.016063 8.9258 0.10013 0.00012659 0.78999 0.0078263 0.0087123 0.0013836 0.98698 0.99173 2.9831e-006 1.1932e-005 0.15256 0.95914 0.9238 0.0013957 0.99592 0.57509 0.0018804 0.43129 2.0442 2.0438 15.9974 144.9714 0.00015278 -85.6635 0.98694
5.091 0.98808 5.4915e-005 3.8183 0.011977 6.6565e-005 0.0011607 0.2314 0.00065929 0.23206 0.21408 0 0.032374 0.0389 0 1.2756 0.4252 0.12843 0.016065 8.9277 0.10014 0.0001266 0.78999 0.0078269 0.0087129 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15256 0.95921 0.92383 0.0013957 0.99592 0.57524 0.0018804 0.4313 2.0445 2.0441 15.9974 144.9714 0.00015274 -85.6635 0.98794
5.092 0.98808 5.4915e-005 3.8183 0.011977 6.6578e-005 0.0011607 0.2314 0.00065929 0.23206 0.21408 0 0.032374 0.0389 0 1.2757 0.42525 0.12845 0.016066 8.9297 0.10015 0.00012662 0.78998 0.0078276 0.0087136 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15257 0.95929 0.92386 0.0013957 0.99593 0.57539 0.0018804 0.43131 2.0448 2.0444 15.9973 144.9714 0.00015269 -85.6635 0.98894
5.093 0.98808 5.4915e-005 3.8183 0.011977 6.6591e-005 0.0011607 0.23141 0.00065929 0.23206 0.21408 0 0.032374 0.0389 0 1.2758 0.42529 0.12847 0.016068 8.9316 0.10016 0.00012663 0.78997 0.0078282 0.0087142 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15257 0.95936 0.92389 0.0013957 0.99594 0.57553 0.0018804 0.43132 2.0451 2.0447 15.9973 144.9714 0.00015264 -85.6635 0.98994
5.094 0.98808 5.4915e-005 3.8183 0.011977 6.6604e-005 0.0011607 0.23141 0.00065929 0.23206 0.21408 0 0.032373 0.0389 0 1.2759 0.42534 0.12848 0.016069 8.9335 0.10017 0.00012664 0.78996 0.0078288 0.0087149 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15258 0.95944 0.92392 0.0013957 0.99595 0.57568 0.0018804 0.43133 2.0454 2.045 15.9973 144.9714 0.0001526 -85.6636 0.99094
5.095 0.98808 5.4915e-005 3.8183 0.011977 6.6617e-005 0.0011607 0.23141 0.00065929 0.23207 0.21408 0 0.032373 0.0389 0 1.276 0.42539 0.1285 0.016071 8.9355 0.10018 0.00012666 0.78995 0.0078294 0.0087156 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15258 0.95951 0.92395 0.0013956 0.99596 0.57583 0.0018804 0.43134 2.0457 2.0453 15.9972 144.9715 0.00015255 -85.6636 0.99194
5.096 0.98808 5.4915e-005 3.8183 0.011977 6.663e-005 0.0011607 0.23141 0.00065929 0.23207 0.21409 0 0.032373 0.0389 0 1.2761 0.42543 0.12851 0.016072 8.9374 0.10019 0.00012667 0.78994 0.00783 0.0087162 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15259 0.95959 0.92398 0.0013956 0.99596 0.57598 0.0018804 0.43135 2.046 2.0456 15.9972 144.9715 0.00015251 -85.6636 0.99294
5.097 0.98808 5.4915e-005 3.8183 0.011977 6.6643e-005 0.0011607 0.23142 0.00065929 0.23207 0.21409 0 0.032373 0.0389 0 1.2762 0.42548 0.12853 0.016074 8.9394 0.1002 0.00012668 0.78993 0.0078306 0.0087169 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15259 0.95966 0.92401 0.0013957 0.99597 0.57613 0.0018803 0.43137 2.0463 2.0459 15.9972 144.9715 0.00015246 -85.6636 0.99394
5.098 0.98808 5.4915e-005 3.8183 0.011977 6.6656e-005 0.0011607 0.23142 0.00065929 0.23207 0.21409 0 0.032373 0.0389 0 1.2763 0.42553 0.12854 0.016075 8.9413 0.10021 0.00012669 0.78992 0.0078312 0.0087176 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.1526 0.95974 0.92404 0.0013957 0.99598 0.57627 0.0018803 0.43138 2.0466 2.0462 15.9971 144.9715 0.00015241 -85.6636 0.99494
5.099 0.98808 5.4914e-005 3.8183 0.011977 6.6669e-005 0.0011607 0.23142 0.00065929 0.23208 0.21409 0 0.032373 0.0389 0 1.2764 0.42557 0.12856 0.016077 8.9432 0.10021 0.00012671 0.78991 0.0078319 0.0087182 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.1526 0.95981 0.92407 0.0013956 0.99599 0.57642 0.0018803 0.43139 2.0469 2.0465 15.9971 144.9715 0.00015237 -85.6637 0.99594
5.1 0.98808 5.4914e-005 3.8183 0.011977 6.6682e-005 0.0011607 0.23142 0.00065929 0.23208 0.2141 0 0.032373 0.0389 0 1.2765 0.42562 0.12857 0.016078 8.9452 0.10022 0.00012672 0.7899 0.0078325 0.0087189 0.0013836 0.98698 0.99173 2.983e-006 1.1932e-005 0.15261 0.95989 0.9241 0.0013956 0.996 0.57657 0.0018803 0.4314 2.0472 2.0468 15.9971 144.9716 0.00015232 -85.6626 0.99694
5.101 0.98808 5.4914e-005 3.8183 0.011977 6.6695e-005 0.0011607 0.23143 0.00065929 0.23208 0.2141 0 0.032373 0.0389 0 1.2766 0.42566 0.12859 0.01608 8.9471 0.10023 0.00012673 0.78989 0.0078331 0.0087196 0.006473 0.98323 0.99099 1.4518e-005 5.3335e-005 0.15261 0.95991 0.92413 0.0027731 0.99599 0.5767 0.0023955 0.43136 2.0475 2.0471 15.997 144.9716 0.00015229 -76.1611 0.99794
5.102 0.98808 5.4914e-005 3.8183 0.011977 6.6708e-005 0.0011607 0.23143 0.00065929 0.23208 0.2141 0 0.032372 0.0389 0 1.2767 0.42571 0.12861 0.016081 8.9491 0.10024 0.00012675 0.78988 0.0078337 0.0087202 0.026219 0.97171 0.98767 6.5971e-005 0.00022947 0.15262 0.95971 0.92415 0.0053006 0.99594 0.57681 0.0033362 0.43124 2.0478 2.0474 15.9969 144.9715 0.00015227 -67.1471 0.99894
5.103 0.98808 5.4914e-005 3.8183 0.011977 6.6721e-005 0.0011607 0.23143 0.00065929 0.23209 0.2141 0 0.032372 0.0389 0 1.2768 0.42576 0.12862 0.016083 8.951 0.10025 0.00012676 0.78987 0.0078343 0.0087209 0.094871 0.94722 0.97733 0.00028439 0.00091309 0.15262 0.95897 0.92418 0.0092474 0.99567 0.5769 0.004425 0.43108 2.0481 2.0477 15.9968 144.9715 0.00015228 -58.0155 0.99994
5.104 0.98808 5.4914e-005 3.8183 0.011977 6.6733e-005 0.0011607 0.23143 0.00065929 0.23209 0.21411 0 0.032372 0.0389 0 1.2768 0.4258 0.12864 0.016084 8.9529 0.10026 0.00012677 0.78987 0.0078349 0.0087215 0.48802 0.85635 0.93874 0.0021791 0.0054754 0.15263 0.95696 0.9242 0.015752 0.99157 0.57693 0.0056239 0.43089 2.0484 2.048 15.9976 144.9715 0.00015232 -37.2183 0.15609
5.105 0.98808 5.4914e-005 3.8183 0.011977 6.6746e-005 0.0011608 0.23144 0.00065929 0.23209 0.21411 0 0.032372 0.0389 0 1.2769 0.42585 0.12865 0.016086 8.9549 0.10027 0.00012679 0.78986 0.0078356 0.0087222 0.99962 0.0021695 0.71212 0.94071 0.99631 0.15263 0.92357 0.92119 0.33431 0.96415 0.56426 0.044314 0.43068 1.9996 0.95043 16.0015 144.9712 0.00024115 24.693 0.0019407
5.106 0.98808 5.4914e-005 3.8183 0.011976 6.6759e-005 0.0011608 0.23144 0.00065929 0.23209 0.21411 0 0.032372 0.0389 0 1.277 0.4259 0.12867 0.016087 8.9568 0.10028 0.0001268 0.78985 0.0078362 0.0087229 0.99945 1.345e-006 0.5282 0.99773 0.99949 0.15264 0.88358 0.90309 0.61722 0.93699 0.54848 0.098389 0.43048 1.8039 0.59501 16.0011 144.9698 0.00035337 20.6743 0.0029407
5.107 0.98808 5.4914e-005 3.8183 0.011976 6.6772e-005 0.0011608 0.23144 0.00065929 0.2321 0.21411 0 0.032372 0.0389 0 1.2771 0.42594 0.12868 0.016089 8.9588 0.10029 0.00012681 0.78984 0.0078368 0.0087235 0.99905 4.2851e-010 0.3921 0.99571 0.99878 0.15264 0.84588 0.87968 0.74014 0.9106 0.53334 0.13977 0.43027 1.6191 0.57379 16.0007 144.9681 0.00042513 15.46 0.0039407
5.108 0.98808 5.4914e-005 3.8183 0.011976 6.6785e-005 0.0011608 0.23144 0.00065929 0.2321 0.21412 0 0.032372 0.0389 0 1.2772 0.42599 0.1287 0.01609 8.9607 0.1003 0.00012683 0.78983 0.0078374 0.0087242 0.99859 -7.962e-011 0.29139 0.99197 0.9977 0.15265 0.81093 0.85358 0.79383 0.88496 0.51897 0.17212 0.43007 1.4654 0.61481 16.0004 144.9663 0.00047915 11.8864 0.0049407
5.109 0.98808 5.4914e-005 3.8183 0.011976 6.6798e-005 0.0011608 0.23145 0.00065929 0.2321 0.21412 0 0.032372 0.0389 0 1.2773 0.42604 0.12871 0.016092 8.9627 0.10031 0.00012684 0.78982 0.007838 0.0087249 0.99817 2.6301e-011 0.21677 0.98756 0.99645 0.15265 0.77861 0.82603 0.81692 0.86004 0.5054 0.19909 0.42986 1.3434 0.67564 16.0001 144.9645 0.00052087 9.5232 0.0059407
5.11 0.98808 5.4914e-005 3.8183 0.011976 6.6811e-005 0.0011608 0.23145 0.00065929 0.2321 0.21412 0 0.032371 0.0389 0 1.2774 0.42608 0.12873 0.016093 8.9646 0.10032 0.00012685 0.78981 0.0078386 0.0087255 0.99779 -1.0275e-010 0.1614 0.98281 0.99512 0.15266 0.74861 0.79791 0.82484 0.83583 0.49257 0.22248 0.42966 1.2499 0.74091 15.9998 144.9628 0.00055297 7.7683 0.0069407
5.111 0.98808 5.4914e-005 3.8183 0.011976 6.6824e-005 0.0011608 0.23145 0.00065929 0.23211 0.21412 0 0.032371 0.0389 0 1.2775 0.42613 0.12875 0.016095 8.9666 0.10033 0.00012687 0.7898 0.0078392 0.0087262 0.99741 2.8709e-011 0.12028 0.9777 0.99368 0.15266 0.72068 0.76984 0.82441 0.8123 0.48045 0.24319 0.42945 1.1804 0.80267 15.9995 144.9611 0.00057752 6.3062 0.0079407
5.112 0.98808 5.4913e-005 3.8183 0.011976 6.6837e-005 0.0011608 0.23146 0.00065929 0.23211 0.21413 0 0.032371 0.0389 0 1.2776 0.42618 0.12876 0.016096 8.9685 0.10033 0.00012688 0.78979 0.0078399 0.0087269 0.997 1.1645e-011 0.089717 0.97208 0.99207 0.15267 0.69464 0.74226 0.81898 0.78944 0.46901 0.26168 0.42925 1.1304 0.85664 15.9992 144.9595 0.00059634 4.9873 0.0089407
5.113 0.98808 5.4913e-005 3.8183 0.011976 6.685e-005 0.0011608 0.23146 0.00065929 0.23211 0.21413 0 0.032371 0.0389 0 1.2777 0.42622 0.12878 0.016098 8.9704 0.10034 0.00012689 0.78978 0.0078405 0.0087275 0.99656 -2.9935e-011 0.066978 0.96575 0.9902 0.15267 0.67037 0.7155 0.81029 0.76722 0.45823 0.27825 0.42904 1.0955 0.90105 15.9989 144.958 0.00061094 3.7351 0.0099407
5.114 0.98808 5.4913e-005 3.8183 0.011976 6.6863e-005 0.0011608 0.23146 0.00065929 0.23211 0.21413 0 0.032371 0.0389 0 1.2778 0.42627 0.12879 0.016099 8.9724 0.10035 0.00012691 0.78977 0.0078411 0.0087282 0.99607 2.4874e-011 0.050052 0.95848 0.988 0.15268 0.64776 0.68978 0.7993 0.74564 0.44812 0.29311 0.42884 1.072 0.93596 15.9986 144.9566 0.00062249 2.5054 0.010941
5.115 0.98808 5.4913e-005 3.8183 0.011976 6.6876e-005 0.0011608 0.23146 0.00065929 0.23212 0.21413 0 0.032371 0.0389 0 1.2779 0.42632 0.12881 0.016101 8.9743 0.10036 0.00012692 0.78976 0.0078417 0.0087288 0.99549 -4.6297e-011 0.037445 0.94999 0.98536 0.15268 0.62674 0.66527 0.7865 0.72466 0.43869 0.30639 0.42863 1.0567 0.96249 15.9983 144.9552 0.00063187 1.2679 0.011941
5.116 0.98808 5.4913e-005 3.8183 0.011976 6.6889e-005 0.0011608 0.23147 0.00065929 0.23212 0.21414 0 0.032371 0.0389 0 1.278 0.42636 0.12882 0.016102 8.9763 0.10037 0.00012693 0.78976 0.0078423 0.0087295 0.99482 8.7226e-011 0.028048 0.93994 0.9821 0.15269 0.60726 0.64209 0.77214 0.70429 0.42993 0.31819 0.42843 1.0473 0.98221 15.998 144.954 0.00063966 -0.0026911 0.012941
5.117 0.98808 5.4913e-005 3.8183 0.011976 6.6902e-005 0.0011608 0.23147 0.00065929 0.23212 0.21414 0 0.032371 0.0389 0 1.2781 0.42641 0.12884 0.016104 8.9782 0.10038 0.00012694 0.78975 0.0078429 0.0087302 0.994 2.6201e-011 0.021041 0.92789 0.9781 0.15269 0.58928 0.62035 0.75629 0.68449 0.42188 0.3286 0.42823 1.0418 0.99673 15.9978 144.9528 0.00064629 -1.3318 0.013941
5.118 0.98808 5.4913e-005 3.8183 0.011976 6.6915e-005 0.0011608 0.23147 0.00065929 0.23212 0.21414 0 0.03237 0.0389 0 1.2782 0.42646 0.12885 0.016105 8.9802 0.10039 0.00012696 0.78974 0.0078435 0.0087308 0.99298 8.5574e-011 0.015812 0.91325 0.97301 0.1527 0.57277 0.60014 0.7389 0.66526 0.41456 0.33766 0.42802 1.0392 1.0074 15.9975 144.9517 0.000652 -2.7491 0.014941
5.119 0.98808 5.4913e-005 3.8183 0.011976 6.6928e-005 0.0011608 0.23147 0.00065929 0.23213 0.21414 0 0.03237 0.0389 0 1.2783 0.4265 0.12887 0.016107 8.9821 0.1004 0.00012697 0.78973 0.0078442 0.0087315 0.99168 4.7763e-010 0.011908 0.89522 0.96648 0.1527 0.55772 0.58157 0.71981 0.64659 0.40798 0.34542 0.42782 1.0383 1.0155 15.9973 144.9506 0.00065694 -4.2931 0.015941
5.12 0.98809 5.4913e-005 3.8183 0.011976 6.6941e-005 0.0011608 0.23148 0.00065929 0.23213 0.21415 0 0.03237 0.0389 0 1.2784 0.42655 0.12889 0.016108 8.9841 0.10041 0.00012698 0.78972 0.0078448 0.0087322 0.98992 4.5991e-010 0.0089924 0.87266 0.9578 0.15271 0.54415 0.56475 0.69877 0.62846 0.4022 0.35188 0.42762 1.0387 1.0216 15.997 144.9497 0.00066119 -6.0163 0.016941
5.121 0.98809 5.4913e-005 3.8183 0.011976 6.6954e-005 0.0011608 0.23148 0.00065929 0.23213 0.21415 0 0.03237 0.0389 0 1.2785 0.4266 0.1289 0.01611 8.986 0.10042 0.000127 0.78971 0.0078454 0.0087328 0.98745 5.6129e-011 0.0068149 0.84388 0.94604 0.15271 0.53209 0.54983 0.67542 0.61087 0.39724 0.35704 0.42741 1.0398 1.0265 15.9968 144.9488 0.00066477 -7.993 0.017941
5.122 0.98809 5.4913e-005 3.8183 0.011976 6.6967e-005 0.0011608 0.23148 0.00065929 0.23213 0.21415 0 0.03237 0.0389 0 1.2786 0.42664 0.12892 0.016111 8.988 0.10043 0.00012701 0.7897 0.007846 0.0087335 0.98372 -3.5432e-012 0.0051904 0.80645 0.92955 0.15272 0.52161 0.53696 0.64931 0.59381 0.39314 0.36087 0.42721 1.0414 1.0306 15.9966 144.948 0.00066765 -10.3292 0.018941
5.123 0.98809 5.4913e-005 3.8183 0.011976 6.698e-005 0.0011608 0.23148 0.00065929 0.23214 0.21415 0 0.03237 0.0389 0 1.2787 0.42669 0.12893 0.016112 8.9899 0.10044 0.00012702 0.78969 0.0078466 0.0087341 0.97766 -1.602e-012 0.0039816 0.75669 0.90571 0.15272 0.51277 0.52633 0.61996 0.5773 0.38993 0.36335 0.42701 1.0434 1.0341 15.9963 144.9472 0.00066978 -13.1712 0.019941
5.124 0.98809 5.4913e-005 3.8183 0.011976 6.6993e-005 0.0011608 0.23149 0.00065929 0.23214 0.21415 0 0.03237 0.0389 0 1.2788 0.42674 0.12895 0.016114 8.9919 0.10045 0.00012704 0.78968 0.0078472 0.0087348 0.96689 4.9523e-013 0.0030884 0.6894 0.87012 0.15273 0.50563 0.5181 0.58696 0.56137 0.38758 0.36446 0.4268 1.0456 1.0373 15.9961 144.9466 0.00067103 -16.7028 0.020941
5.125 0.98809 5.4913e-005 3.8183 0.011976 6.7006e-005 0.0011608 0.23149 0.00065929 0.23214 0.21416 0 0.03237 0.0389 0 1.2789 0.42678 0.12896 0.016115 8.9938 0.10045 0.00012705 0.78967 0.0078478 0.0087355 0.946 -2.2414e-013 0.0024382 0.59782 0.81582 0.15273 0.50015 0.51234 0.55025 0.54616 0.38602 0.36426 0.4266 1.0479 1.0403 15.996 144.9461 0.00067132 -21.0933 0.021941
5.126 0.98809 5.4912e-005 3.8183 0.011976 6.7019e-005 0.0011608 0.23149 0.00065929 0.23214 0.21416 0 0.032369 0.0389 0 1.279 0.42683 0.12898 0.016117 8.9958 0.10046 0.00012706 0.78966 0.0078485 0.0087361 0.90361 8.1271e-014 0.0019785 0.47637 0.73308 0.15274 0.49616 0.50883 0.51002 0.53198 0.38509 0.36287 0.4264 1.0503 1.0432 15.9958 144.9456 0.00067062 -26.3322 0.022941
5.127 0.98809 5.4912e-005 3.8183 0.011976 6.7032e-005 0.0011608 0.23149 0.00065929 0.23215 0.21416 0 0.032369 0.0389 0 1.2791 0.42688 0.12899 0.016118 8.9977 0.10047 0.00012708 0.78965 0.0078491 0.0087368 0.82264 7.0868e-014 0.0016674 0.32972 0.61335 0.15274 0.49331 0.50697 0.46587 0.5196 0.3846 0.36044 0.4262 1.0528 1.0459 15.9957 144.9452 0.00066915 -31.9922 0.023941
5.128 0.98809 5.4912e-005 3.8183 0.011976 6.7045e-005 0.0011608 0.2315 0.00065929 0.23215 0.21416 0 0.032369 0.0389 0 1.2791 0.42692 0.12901 0.01612 8.9997 0.10048 0.00012709 0.78964 0.0078497 0.0087374 0.6974 1.5513e-014 0.0014643 0.18484 0.46085 0.15274 0.49122 0.50602 0.41589 0.5104 0.38438 0.3569 0.426 1.0553 1.0485 15.9956 144.9449 0.00066727 -37.327 0.024941
5.129 0.98809 5.4912e-005 3.8183 0.011976 6.7057e-005 0.0011608 0.2315 0.00065929 0.23215 0.21417 0 0.032369 0.0389 0 1.2792 0.42697 0.12902 0.016121 9.0016 0.10049 0.0001271 0.78964 0.0078503 0.0087381 0.55179 0.00017701 0.0013833 0.07934 0.30118 0.15275 0.48965 0.50566 0.35832 0.50548 0.38432 0.35195 0.4258 1.0578 1.0512 15.9955 144.9447 0.00066525 -41.8788 0.025941
5.13 0.98809 5.4912e-005 3.8183 0.011976 6.707e-005 0.0011608 0.2315 0.00065929 0.23215 0.21417 0 0.032369 0.0389 0 1.2793 0.42702 0.12904 0.016123 9.0036 0.1005 0.00012711 0.78963 0.0078509 0.0087388 0.41896 0.00076827 0.0015651 0.025826 0.1679 0.15275 0.4885 0.50612 0.29418 0.5043 0.38436 0.34521 0.4256 1.0603 1.0537 15.9954 144.9445 0.00066318 -45.6269 0.026941
5.131 0.98809 5.4912e-005 3.8183 0.011976 6.7083e-005 0.0011608 0.2315 0.00065929 0.23216 0.21417 0 0.032369 0.0389 0 1.2794 0.42706 0.12906 0.016124 9.0055 0.10051 0.00012713 0.78962 0.0078515 0.0087394 0.3159 0.0017351 0.002025 0.007088 0.079704 0.15276 0.48768 0.50762 0.22809 0.50518 0.38444 0.3364 0.42541 1.0629 1.0563 15.9954 144.9443 0.00066106 -48.6788 0.027941
5.132 0.98809 5.4912e-005 3.8183 0.011976 6.7096e-005 0.0011608 0.23151 0.00065929 0.23216 0.21417 0 0.032369 0.0389 0 1.2795 0.42711 0.12907 0.016126 9.0075 0.10052 0.00012714 0.78961 0.0078521 0.0087401 0.2425 0.0031847 0.0027853 0.0022863 0.033103 0.15276 0.48716 0.50995 0.1666 0.50684 0.38456 0.32543 0.42522 1.0654 1.0589 15.9953 144.9442 0.00065892 -51.1543 0.028941
5.133 0.98809 5.4912e-005 3.8183 0.011976 6.7109e-005 0.0011608 0.23151 0.00065929 0.23216 0.21418 0 0.032369 0.0389 0 1.2796 0.42716 0.12909 0.016127 9.0094 0.10053 0.00012715 0.7896 0.0078527 0.0087407 0.19143 0.0051948 0.0038548 0.001156 0.013006 0.15277 0.48689 0.51274 0.11526 0.50868 0.38469 0.31243 0.42503 1.0679 1.0614 15.9953 144.9442 0.00065676 -53.1781 0.029941
5.134 0.98809 5.4912e-005 3.8183 0.011976 6.7122e-005 0.0011608 0.23151 0.00065929 0.23216 0.21418 0 0.032368 0.0389 0 1.2797 0.4272 0.1291 0.016129 9.0114 0.10054 0.00012717 0.78959 0.0078534 0.0087414 0.15523 0.0078211 0.0052337 0.00077966 0.0055984 0.15277 0.48683 0.51571 0.076639 0.51051 0.38483 0.29763 0.42485 1.0704 1.064 15.9953 144.9441 0.00065458 -54.8703 0.030941
5.135 0.98809 5.4912e-005 3.8183 0.011976 6.7135e-005 0.0011608 0.23151 0.00065929 0.23217 0.21418 0 0.032368 0.0389 0 1.2798 0.42725 0.12912 0.01613 9.0133 0.10055 0.00012718 0.78958 0.007854 0.0087421 0.12853 0.011112 0.0069214 0.00058268 0.0030361 0.15278 0.48694 0.51872 0.050172 0.51227 0.38498 0.28131 0.42467 1.073 1.0665 15.9953 144.9441 0.0006524 -56.3336 0.031941
5.136 0.98809 5.4912e-005 3.8183 0.011976 6.7148e-005 0.0011608 0.23152 0.00065929 0.23217 0.21418 0 0.032368 0.0389 0 1.2799 0.42729 0.12913 0.016132 9.0153 0.10056 0.00012719 0.78957 0.0078546 0.0087427 0.10794 0.015122 0.0089218 0.00045397 0.0020526 0.15278 0.4872 0.52172 0.033417 0.51393 0.38512 0.26377 0.42449 1.0755 1.0691 15.9953 144.944 0.0006502 -57.6465 0.032941
5.137 0.98809 5.4912e-005 3.8183 0.011976 6.7161e-005 0.0011608 0.23152 0.00065929 0.23217 0.21419 0 0.032368 0.0389 0 1.28 0.42734 0.12915 0.016133 9.0172 0.10056 0.00012721 0.78956 0.0078552 0.0087434 0.091464 0.019923 0.011246 0.00036194 0.0015585 0.15279 0.48759 0.52469 0.023437 0.5155 0.38527 0.24529 0.42431 1.078 1.0716 15.9953 144.944 0.000648 -58.8623 0.033941
5.138 0.98809 5.4912e-005 3.8183 0.011976 6.7174e-005 0.0011609 0.23152 0.00065929 0.23217 0.21419 0 0.032368 0.0389 0 1.2801 0.42739 0.12916 0.016135 9.0192 0.10057 0.00012722 0.78955 0.0078558 0.0087441 0.07792 0.025606 0.013913 0.00029253 0.0012388 0.15279 0.4881 0.52764 0.017687 0.51699 0.38543 0.22613 0.42414 1.0805 1.0741 15.9953 144.944 0.00064579 -60.0145 0.034941
5.139 0.98809 5.4911e-005 3.8183 0.011976 6.7187e-005 0.0011609 0.23152 0.00065929 0.23218 0.21419 0 0.032368 0.0389 0 1.2802 0.42743 0.12918 0.016136 9.0212 0.10058 0.00012723 0.78954 0.0078564 0.0087447 0.066608 0.032281 0.016946 0.00023927 0.0010032 0.1528 0.48871 0.53057 0.014342 0.51841 0.38558 0.20653 0.42397 1.083 1.0767 15.9954 144.944 0.00064358 -61.122 0.035941
5.14 0.98809 5.4911e-005 3.8183 0.011976 6.72e-005 0.0011609 0.23153 0.00065929 0.23218 0.21419 0 0.032368 0.0389 0 1.2803 0.42748 0.1292 0.016138 9.0231 0.10059 0.00012725 0.78953 0.007857 0.0087454 0.057078 0.040074 0.020374 0.00019697 0.00082089 0.1528 0.48942 0.53346 0.012267 0.51977 0.38573 0.18676 0.4238 1.0855 1.0792 15.9954 144.9439 0.00064137 -62.195 0.036941
5.141 0.98809 5.4911e-005 3.8183 0.011976 6.7213e-005 0.0011609 0.23153 0.00065929 0.23218 0.2142 0 0.032368 0.0389 0 1.2804 0.42753 0.12921 0.016139 9.0251 0.1006 0.00012726 0.78953 0.0078576 0.008746 0.049015 0.049123 0.024228 0.00016306 0.00067651 0.15281 0.49022 0.53632 0.010835 0.52107 0.38588 0.1671 0.42364 1.0881 1.0817 15.9954 144.9439 0.00063915 -63.2388 0.037941
5.142 0.98809 5.4911e-005 3.8183 0.011976 6.7226e-005 0.0011609 0.23153 0.00065929 0.23218 0.2142 0 0.032367 0.0389 0 1.2805 0.42757 0.12923 0.016141 9.027 0.10061 0.00012727 0.78952 0.0078583 0.0087467 0.042177 0.059578 0.028543 0.00013578 0.00056093 0.15281 0.49109 0.53916 0.0097365 0.52233 0.38604 0.14781 0.42348 1.0906 1.0843 15.9954 144.9439 0.00063693 -64.2559 0.038941
5.143 0.98809 5.4911e-005 3.8183 0.011976 6.7239e-005 0.0011609 0.23153 0.00065929 0.23219 0.2142 0 0.032367 0.0389 0 1.2806 0.42762 0.12924 0.016142 9.029 0.10062 0.00012729 0.78951 0.0078589 0.0087474 0.03637 0.071591 0.033357 0.00011355 0.00046762 0.15282 0.49203 0.54196 0.0088285 0.52355 0.38619 0.12918 0.42333 1.0931 1.0868 15.9955 144.9439 0.00063472 -65.2478 0.039941
5.144 0.98809 5.4911e-005 3.8183 0.011976 6.7252e-005 0.0011609 0.23153 0.00065929 0.23219 0.2142 0 0.032367 0.0389 0 1.2807 0.42767 0.12926 0.016144 9.0309 0.10063 0.0001273 0.7895 0.0078595 0.008748 0.031434 0.085318 0.038709 9.5469e-005 0.00039186 0.15282 0.49303 0.54473 0.0080472 0.52474 0.38635 0.11146 0.42318 1.0956 1.0893 15.9955 144.9438 0.00063249 -66.2152 0.040941
5.145 0.98809 5.4911e-005 3.8183 0.011976 6.7265e-005 0.0011609 0.23154 0.00065929 0.23219 0.2142 0 0.032367 0.0389 0 1.2808 0.42771 0.12927 0.016145 9.0329 0.10064 0.00012731 0.78949 0.0078601 0.0087487 0.027232 0.10091 0.044645 8.0564e-005 0.00032999 0.15283 0.49409 0.54748 0.0073629 0.52591 0.3865 0.094905 0.42303 1.0981 1.0918 15.9956 144.9438 0.00063027 -67.1583 0.041941
5.146 0.98809 5.4911e-005 3.8183 0.011976 6.7278e-005 0.0011609 0.23154 0.00065929 0.23219 0.21421 0 0.032367 0.0389 0 1.2809 0.42776 0.12929 0.016147 9.0349 0.10065 0.00012732 0.78948 0.0078607 0.0087493 0.023653 0.11852 0.051214 6.8347e-005 0.00027924 0.15283 0.4952 0.55019 0.0067579 0.52707 0.38666 0.079703 0.42289 1.1006 1.0943 15.9956 144.9438 0.00062805 -68.0772 0.042941
5.147 0.98809 5.4911e-005 3.8183 0.011976 6.7291e-005 0.0011609 0.23154 0.00065929 0.2322 0.21421 0 0.032367 0.0389 0 1.281 0.42781 0.1293 0.016148 9.0368 0.10066 0.00012734 0.78947 0.0078613 0.00875 0.020603 0.13827 0.058467 5.8244e-005 0.00023743 0.15284 0.49635 0.55288 0.0062207 0.52822 0.38681 0.066009 0.42275 1.1031 1.0969 15.9957 144.9437 0.00062583 -68.9716 0.043941
5.148 0.98809 5.4911e-005 3.8183 0.011976 6.7304e-005 0.0011609 0.23154 0.00065929 0.2322 0.21421 0 0.032367 0.0389 0 1.2811 0.42785 0.12932 0.01615 9.0388 0.10067 0.00012735 0.78946 0.0078619 0.0087507 0.017998 0.16028 0.066465 4.9845e-005 0.00020286 0.15284 0.49754 0.55554 0.0057424 0.52937 0.38697 0.053916 0.42262 1.1056 1.0994 15.9957 144.9437 0.00062361 -69.8411 0.044941
5.149 0.98809 5.4911e-005 3.8183 0.011976 6.7317e-005 0.0011609 0.23155 0.00065929 0.2322 0.21421 0 0.032367 0.0389 0 1.2812 0.4279 0.12934 0.016151 9.0407 0.10068 0.00012736 0.78945 0.0078625 0.0087513 0.015774 0.1846 0.075269 4.2871e-005 0.00017418 0.15285 0.49877 0.55817 0.0053154 0.53053 0.38713 0.043459 0.4225 1.1081 1.1019 15.9958 144.9437 0.00062139 -70.6848 0.045941
5.15 0.98809 5.4911e-005 3.8183 0.011976 6.733e-005 0.0011609 0.23155 0.00065929 0.2322 0.21422 0 0.032366 0.0389 0 1.2813 0.42795 0.12935 0.016153 9.0427 0.10068 0.00012738 0.78944 0.0078631 0.008752 0.013874 0.21129 0.084949 3.7047e-005 0.0001503 0.15285 0.50002 0.56077 0.0049337 0.53169 0.38728 0.034609 0.42238 1.1105 1.1044 15.9959 144.9436 0.00061917 -71.502 0.046941
5.151 0.98809 5.4911e-005 3.8183 0.011976 6.7343e-005 0.0011609 0.23155 0.00065929 0.23221 0.21422 0 0.032366 0.0389 0 1.2814 0.42799 0.12937 0.016154 9.0446 0.10069 0.00012739 0.78943 0.0078638 0.0087526 0.012247 0.24032 0.095574 3.2176e-005 0.00013036 0.15286 0.5013 0.56335 0.0045922 0.53287 0.38744 0.027287 0.42226 1.113 1.1069 15.9959 144.9436 0.00061696 -72.2915 0.047941
5.152 0.98809 5.4911e-005 3.8183 0.011976 6.7356e-005 0.0011609 0.23155 0.00065929 0.23221 0.21422 0 0.032366 0.0389 0 1.2814 0.42804 0.12938 0.016156 9.0466 0.1007 0.0001274 0.78942 0.0078644 0.0087533 0.010855 0.27161 0.10721 2.8092e-005 0.00011367 0.15286 0.5026 0.5659 0.0042865 0.53407 0.3876 0.021366 0.42215 1.1155 1.1094 15.996 144.9436 0.00061474 -73.0522 0.048941
5.153 0.98809 5.491e-005 3.8183 0.011976 6.7368e-005 0.0011609 0.23156 0.00065929 0.23221 0.21422 0 0.032366 0.0389 0 1.2815 0.42809 0.1294 0.016157 9.0486 0.10071 0.00012742 0.78942 0.007865 0.0087539 0.0096626 0.30502 0.11993 2.4658e-005 9.9671e-005 0.15287 0.50392 0.56842 0.0040126 0.53529 0.38777 0.016685 0.42205 1.118 1.1119 15.9961 144.9436 0.00061253 -73.783 0.049941
5.154 0.98809 5.491e-005 3.8183 0.011976 6.7381e-005 0.0011609 0.23156 0.00065929 0.23221 0.21423 0 0.032366 0.0389 0 1.2816 0.42813 0.12941 0.016159 9.0505 0.10072 0.00012743 0.78941 0.0078656 0.0087546 0.0086401 0.34035 0.13379 2.1766e-005 8.7892e-005 0.15287 0.50525 0.57091 0.0037674 0.53654 0.38793 0.013069 0.42195 1.1205 1.1144 15.9962 144.9435 0.00061033 -74.4827 0.050941
5.155 0.98809 5.491e-005 3.8183 0.011976 6.7394e-005 0.0011609 0.23156 0.00065929 0.23222 0.21423 0 0.032366 0.0389 0 1.2817 0.42818 0.12943 0.01616 9.0525 0.10073 0.00012744 0.7894 0.0078662 0.0087553 0.0077628 0.3773 0.14882 1.9324e-005 7.7959e-005 0.15288 0.5066 0.57338 0.0035478 0.53782 0.38809 0.010334 0.42186 1.1229 1.1169 15.9963 144.9435 0.00060813 -75.1502 0.051941
5.156 0.98809 5.491e-005 3.8183 0.011976 6.7407e-005 0.0011609 0.23156 0.00065929 0.23222 0.21423 0 0.032366 0.0389 0 1.2818 0.42823 0.12944 0.016162 9.0544 0.10074 0.00012746 0.78939 0.0078668 0.0087559 0.0070092 0.41552 0.16504 1.7258e-005 6.9565e-005 0.15288 0.50796 0.57583 0.0033512 0.53914 0.38826 0.0083063 0.42177 1.1254 1.1194 15.9963 144.9435 0.00060593 -75.7849 0.052941
5.157 0.98809 5.491e-005 3.8183 0.011976 6.742e-005 0.0011609 0.23157 0.00065929 0.23222 0.21423 0 0.032366 0.0389 0 1.2819 0.42827 0.12946 0.016163 9.0564 0.10075 0.00012747 0.78938 0.0078674 0.0087566 0.0063615 0.45463 0.18245 1.5505e-005 6.2453e-005 0.15289 0.50932 0.57824 0.0031754 0.54049 0.38843 0.0068273 0.42169 1.1279 1.1219 15.9964 144.9435 0.00060374 -76.386 0.053941
5.158 0.98809 5.491e-005 3.8183 0.011976 6.7433e-005 0.0011609 0.23157 0.00065929 0.23222 0.21423 0 0.032365 0.0389 0 1.282 0.42832 0.12947 0.016165 9.0584 0.10076 0.00012748 0.78937 0.007868 0.0087572 0.0058038 0.49416 0.201 1.4015e-005 5.6413e-005 0.15289 0.5107 0.58064 0.0030182 0.54188 0.38859 0.0057614 0.42161 1.1304 1.1244 15.9965 144.9434 0.00060155 -76.9531 0.054941
5.159 0.98809 5.491e-005 3.8183 0.011976 6.7446e-005 0.0011609 0.23157 0.00065929 0.23223 0.21424 0 0.032365 0.0389 0 1.2821 0.42837 0.12949 0.016166 9.0603 0.10077 0.00012749 0.78936 0.0078686 0.0087579 0.0053229 0.53367 0.22064 1.2746e-005 5.127e-005 0.15289 0.51208 0.58301 0.0028776 0.54332 0.38877 0.004998 0.42154 1.1328 1.1268 15.9966 144.9434 0.00059937 -77.4863 0.055941
5.16 0.98809 5.491e-005 3.8183 0.011976 6.7459e-005 0.0011609 0.23157 0.00065929 0.23223 0.21424 0 0.032365 0.0389 0 1.2822 0.42841 0.12951 0.016168 9.0623 0.10078 0.00012751 0.78935 0.0078693 0.0087586 0.004908 0.57267 0.24126 1.1661e-005 4.6881e-005 0.1529 0.51347 0.58535 0.002752 0.54479 0.38894 0.0044502 0.42147 1.1353 1.1293 15.9967 144.9434 0.00059719 -77.9858 0.056941
5.161 0.98809 5.491e-005 3.8183 0.011976 6.7472e-005 0.0011609 0.23158 0.00065929 0.23223 0.21424 0 0.032365 0.0389 0 1.2823 0.42846 0.12952 0.016169 9.0643 0.10079 0.00012752 0.78934 0.0078699 0.0087592 0.0045492 0.61072 0.26276 1.0733e-005 4.3126e-005 0.1529 0.51486 0.58767 0.0026399 0.54631 0.38911 0.0040529 0.4214 1.1377 1.1318 15.9968 144.9434 0.00059502 -78.452 0.057941
5.162 0.98809 5.491e-005 3.8183 0.011976 6.7485e-005 0.0011609 0.23158 0.00065929 0.23223 0.21424 0 0.032365 0.0389 0 1.2824 0.42851 0.12954 0.016171 9.0662 0.10079 0.00012753 0.78933 0.0078705 0.0087599 0.0042384 0.64741 0.28499 9.9354e-006 3.9903e-005 0.15291 0.51625 0.58997 0.0025397 0.54787 0.38929 0.0037594 0.42135 1.1402 1.1343 15.9969 144.9433 0.00059286 -78.8858 0.058941
5.163 0.98809 5.491e-005 3.8183 0.011976 6.7498e-005 0.0011609 0.23158 0.00065929 0.23224 0.21425 0 0.032365 0.0389 0 1.2825 0.42855 0.12955 0.016172 9.0682 0.1008 0.00012755 0.78932 0.0078711 0.0087605 0.0039688 0.68237 0.3078 9.249e-006 3.7131e-005 0.15291 0.51765 0.59224 0.0024503 0.54947 0.38946 0.0035368 0.42129 1.1427 1.1367 15.997 144.9433 0.00059071 -79.2881 0.059941
5.164 0.98809 5.491e-005 3.8183 0.011976 6.7511e-005 0.0011609 0.23158 0.00065929 0.23224 0.21425 0 0.032365 0.0389 0 1.2826 0.4286 0.12957 0.016174 9.0701 0.10081 0.00012756 0.78931 0.0078717 0.0087612 0.0037344 0.71531 0.33105 8.6565e-006 3.4739e-005 0.15292 0.51905 0.59449 0.0023705 0.55111 0.38964 0.0033629 0.42124 1.1451 1.1392 15.9971 144.9433 0.00058856 -79.6601 0.060941
5.165 0.98809 5.491e-005 3.8183 0.011976 6.7524e-005 0.0011609 0.23159 0.00065929 0.23224 0.21425 0 0.032365 0.0389 0 1.2827 0.42865 0.12958 0.016175 9.0721 0.10082 0.00012757 0.78931 0.0078723 0.0087618 0.0035302 0.74601 0.35459 8.1438e-006 3.2671e-005 0.15292 0.52045 0.59672 0.0022992 0.55279 0.38982 0.003223 0.42119 1.1475 1.1417 15.9972 144.9433 0.00058643 -80.0034 0.061941
5.166 0.98809 5.4909e-005 3.8183 0.011976 6.7537e-005 0.0011609 0.23159 0.00065929 0.23224 0.21425 0 0.032365 0.0389 0 1.2828 0.42869 0.1296 0.016177 9.0741 0.10083 0.00012759 0.7893 0.0078729 0.0087625 0.0033519 0.77432 0.37825 7.6989e-006 3.0876e-005 0.15293 0.52184 0.59893 0.0022355 0.55451 0.39 0.0031072 0.42115 1.15 1.1441 15.9973 144.9433 0.0005843 -80.3192 0.062941
5.167 0.98809 5.4909e-005 3.8183 0.011976 6.755e-005 0.0011609 0.23159 0.00065929 0.23225 0.21426 0 0.032364 0.0389 0 1.2829 0.42874 0.12961 0.016178 9.076 0.10084 0.0001276 0.78929 0.0078735 0.0087632 0.0031961 0.80018 0.40192 7.3119e-006 2.9316e-005 0.15293 0.52324 0.60111 0.0021786 0.55626 0.39019 0.0030093 0.42111 1.1524 1.1466 15.9974 144.9433 0.00058218 -80.6092 0.063941
5.168 0.98809 5.4909e-005 3.8183 0.011975 6.7563e-005 0.0011609 0.23159 0.00065929 0.23225 0.21426 0 0.032364 0.0389 0 1.283 0.42878 0.12963 0.01618 9.078 0.10085 0.00012761 0.78928 0.0078741 0.0087638 0.0030594 0.82356 0.42546 6.9743e-006 2.7956e-005 0.15294 0.52464 0.60327 0.0021278 0.55805 0.39037 0.0029253 0.42107 1.1549 1.149 15.9975 144.9433 0.00058007 -80.8751 0.064941
5.169 0.98809 5.4909e-005 3.8183 0.011975 6.7576e-005 0.0011609 0.2316 0.00065929 0.23225 0.21426 0 0.032364 0.0389 0 1.2831 0.42883 0.12965 0.016181 9.08 0.10086 0.00012763 0.78927 0.0078747 0.0087645 0.0029393 0.84453 0.44875 6.679e-006 2.6767e-005 0.15294 0.52603 0.60541 0.0020823 0.55987 0.39055 0.0028522 0.42104 1.1573 1.1515 15.9976 144.9432 0.00057797 -81.1183 0.065941
5.17 0.98809 5.4909e-005 3.8183 0.011975 6.7589e-005 0.0011609 0.2316 0.00065929 0.23225 0.21426 0 0.032364 0.0389 0 1.2832 0.42888 0.12966 0.016183 9.0819 0.10087 0.00012764 0.78926 0.0078754 0.0087651 0.0028337 0.86317 0.4717 6.4202e-006 2.5724e-005 0.15295 0.52742 0.60753 0.0020417 0.56172 0.39074 0.002788 0.421 1.1597 1.154 15.9977 144.9432 0.00057588 -81.3407 0.066941
5.171 0.98809 5.4909e-005 3.8183 0.011975 6.7602e-005 0.001161 0.2316 0.00065929 0.23226 0.21426 0 0.032364 0.0389 0 1.2833 0.42892 0.12968 0.016184 9.0839 0.10088 0.00012765 0.78925 0.007876 0.0087658 0.0027406 0.87962 0.49422 6.1927e-006 2.4808e-005 0.15295 0.52882 0.60963 0.0020052 0.56359 0.39093 0.0027314 0.42097 1.1622 1.1564 15.9978 144.9432 0.0005738 -81.5436 0.067941
5.172 0.98809 5.4909e-005 3.8183 0.011975 6.7615e-005 0.001161 0.2316 0.00065929 0.23226 0.21427 0 0.032364 0.0389 0 1.2834 0.42897 0.12969 0.016186 9.0859 0.10089 0.00012766 0.78924 0.0078766 0.0087664 0.0026582 0.89403 0.51624 5.9922e-006 2.4002e-005 0.15296 0.5302 0.61171 0.0019726 0.56549 0.39111 0.0026812 0.42094 1.1646 1.1588 15.9979 144.9432 0.00057173 -81.7287 0.068941
5.173 0.98809 5.4909e-005 3.8183 0.011975 6.7628e-005 0.001161 0.23161 0.00065929 0.23226 0.21427 0 0.032364 0.0389 0 1.2835 0.42902 0.12971 0.016187 9.0878 0.1009 0.00012768 0.78923 0.0078772 0.0087671 0.0025849 0.90657 0.53769 5.8152e-006 2.3289e-005 0.15296 0.53159 0.61377 0.0019433 0.56741 0.3913 0.0026367 0.42092 1.167 1.1613 15.9981 144.9432 0.00056967 -81.8974 0.069941
5.174 0.98809 5.4909e-005 3.8183 0.011975 6.7641e-005 0.001161 0.23161 0.00065929 0.23226 0.21427 0 0.032364 0.0389 0 1.2836 0.42906 0.12972 0.016189 9.0898 0.1009 0.00012769 0.78922 0.0078778 0.0087678 0.0025199 0.91743 0.55854 5.6585e-006 2.2659e-005 0.15297 0.53297 0.61581 0.001917 0.56935 0.39149 0.002597 0.42089 1.1694 1.1637 15.9982 144.9432 0.00056762 -82.0512 0.070941
5.175 0.98809 5.4909e-005 3.8183 0.011975 6.7654e-005 0.001161 0.23161 0.00065929 0.23226 0.21427 0 0.032363 0.0389 0 1.2837 0.42911 0.12974 0.01619 9.0918 0.10091 0.0001277 0.78921 0.0078784 0.0087684 0.0024626 0.92677 0.57875 5.5194e-006 2.2099e-005 0.15297 0.53435 0.61783 0.0018934 0.5713 0.39168 0.0025616 0.42087 1.1718 1.1662 15.9983 144.9432 0.00056558 -82.1913 0.071941
5.176 0.98809 5.4909e-005 3.8183 0.011975 6.7666e-005 0.001161 0.23161 0.00065929 0.23227 0.21428 0 0.032363 0.0389 0 1.2837 0.42916 0.12975 0.016192 9.0937 0.10092 0.00012772 0.78921 0.007879 0.0087691 0.0024113 0.93478 0.59828 5.3956e-006 2.1601e-005 0.15298 0.53573 0.61983 0.0018721 0.57328 0.39187 0.0025298 0.42085 1.1743 1.1686 15.9984 144.9432 0.00056355 -82.3189 0.072941
5.177 0.98809 5.4909e-005 3.8183 0.011975 6.7679e-005 0.001161 0.23161 0.00065929 0.23227 0.21428 0 0.032363 0.0389 0 1.2838 0.4292 0.12977 0.016193 9.0957 0.10093 0.00012773 0.7892 0.0078796 0.0087697 0.0023654 0.94161 0.61713 5.2852e-006 2.1158e-005 0.15298 0.53711 0.62181 0.0018529 0.57526 0.39206 0.0025014 0.42083 1.1767 1.171 15.9985 144.9432 0.00056153 -82.4352 0.073941
5.178 0.98809 5.4909e-005 3.8183 0.011975 6.7692e-005 0.001161 0.23162 0.00065929 0.23227 0.21428 0 0.032363 0.0389 0 1.2839 0.42925 0.12978 0.016195 9.0977 0.10094 0.00012774 0.78919 0.0078802 0.0087704 0.0023242 0.94743 0.63528 5.1865e-006 2.0761e-005 0.15299 0.53848 0.62377 0.0018356 0.57726 0.39226 0.0024758 0.42081 1.1791 1.1734 15.9986 144.9432 0.00055952 -82.5413 0.074941
5.179 0.98809 5.4908e-005 3.8183 0.011975 6.7705e-005 0.001161 0.23162 0.00065929 0.23227 0.21428 0 0.032363 0.0389 0 1.284 0.4293 0.1298 0.016196 9.0996 0.10095 0.00012776 0.78918 0.0078808 0.008771 0.0022873 0.95235 0.65272 5.0981e-006 2.0406e-005 0.15299 0.53985 0.62571 0.00182 0.57926 0.39245 0.0024529 0.42079 1.1815 1.1759 15.9987 144.9432 0.00055752 -82.6381 0.075941
5.18 0.98809 5.4908e-005 3.8183 0.011975 6.7718e-005 0.001161 0.23162 0.00065929 0.23228 0.21428 0 0.032363 0.0389 0 1.2841 0.42934 0.12982 0.016198 9.1016 0.10096 0.00012777 0.78917 0.0078814 0.0087717 0.0022541 0.95652 0.66945 5.0186e-006 2.0086e-005 0.153 0.54121 0.62763 0.0018058 0.58128 0.39264 0.0024321 0.42077 1.1839 1.1783 15.9988 144.9432 0.00055554 -82.7266 0.076941
5.181 0.98809 5.4908e-005 3.8183 0.011975 6.7731e-005 0.001161 0.23162 0.00065929 0.23228 0.21429 0 0.032363 0.0389 0 1.2842 0.42939 0.12983 0.016199 9.1036 0.10097 0.00012778 0.78916 0.0078821 0.0087724 0.0022241 0.96003 0.68549 4.947e-006 1.9799e-005 0.153 0.54257 0.62954 0.0017929 0.5833 0.39283 0.0024134 0.42076 1.1863 1.1807 15.9989 144.9432 0.00055356 -82.8075 0.077941
5.182 0.98809 5.4908e-005 3.8183 0.011975 6.7744e-005 0.001161 0.23163 0.00065929 0.23228 0.21429 0 0.032363 0.0389 0 1.2843 0.42944 0.12985 0.016201 9.1056 0.10098 0.0001278 0.78915 0.0078827 0.008773 0.0021969 0.963 0.70085 4.8824e-006 1.9539e-005 0.15301 0.54393 0.63143 0.0017812 0.58533 0.39303 0.0023965 0.42074 1.1886 1.1831 15.999 144.9432 0.0005516 -82.8816 0.078941
5.183 0.98809 5.4908e-005 3.8183 0.011975 6.7757e-005 0.001161 0.23163 0.00065929 0.23228 0.21429 0 0.032362 0.0389 0 1.2844 0.42948 0.12986 0.016202 9.1075 0.10099 0.00012781 0.78914 0.0078833 0.0087737 0.0021724 0.96549 0.71553 4.8238e-006 1.9304e-005 0.15301 0.54528 0.6333 0.0017706 0.58735 0.39322 0.0023811 0.42073 1.191 1.1855 15.9991 144.9432 0.00054964 -82.9495 0.079941
5.184 0.98809 5.4908e-005 3.8183 0.011975 6.777e-005 0.001161 0.23163 0.00065929 0.23229 0.21429 0 0.032362 0.0389 0 1.2845 0.42953 0.12988 0.016204 9.1095 0.101 0.00012782 0.78913 0.0078839 0.0087743 0.0021501 0.9676 0.72955 4.7706e-006 1.909e-005 0.15302 0.54664 0.63515 0.0017608 0.58939 0.39341 0.0023671 0.42071 1.1934 1.1879 15.9992 144.9432 0.0005477 -83.0119 0.080941
5.185 0.98809 5.4908e-005 3.8183 0.011975 6.7783e-005 0.001161 0.23163 0.00065929 0.23229 0.2143 0 0.032362 0.0389 0 1.2846 0.42958 0.12989 0.016205 9.1115 0.101 0.00012783 0.78912 0.0078845 0.008775 0.0021297 0.96937 0.74293 4.7222e-006 1.8896e-005 0.15302 0.54798 0.63698 0.0017519 0.59142 0.39361 0.0023543 0.4207 1.1958 1.1903 15.9993 144.9432 0.00054577 -83.0694 0.081941
5.186 0.98809 5.4908e-005 3.8183 0.011975 6.7796e-005 0.001161 0.23164 0.00065929 0.23229 0.2143 0 0.032362 0.0389 0 1.2847 0.42962 0.12991 0.016207 9.1134 0.10101 0.00012785 0.78911 0.0078851 0.0087756 0.002111 0.97086 0.75568 4.678e-006 1.8718e-005 0.15303 0.54933 0.6388 0.0017437 0.59345 0.3938 0.0023427 0.42069 1.1982 1.1927 15.9994 144.9432 0.00054384 -83.1224 0.082941
5.187 0.98809 5.4908e-005 3.8183 0.011975 6.7809e-005 0.001161 0.23164 0.00065929 0.23229 0.2143 0 0.032362 0.0389 0 1.2848 0.42967 0.12992 0.016208 9.1154 0.10102 0.00012786 0.7891 0.0078857 0.0087763 0.0020942 0.97212 0.76784 4.6375e-006 1.8556e-005 0.15303 0.55066 0.6406 0.0017362 0.59549 0.394 0.002332 0.42068 1.2006 1.1951 15.9995 144.9432 0.00054193 -83.1715 0.083941
5.188 0.98809 5.4908e-005 3.8183 0.011975 6.7822e-005 0.001161 0.23164 0.00065929 0.2323 0.2143 0 0.032362 0.0389 0 1.2849 0.42972 0.12994 0.01621 9.1174 0.10103 0.00012787 0.7891 0.0078863 0.008777 0.0020783 0.97318 0.77941 4.6002e-006 1.8406e-005 0.15303 0.552 0.64239 0.0017293 0.59752 0.39419 0.0023221 0.42067 1.2029 1.1975 15.9996 144.9432 0.00054003 -83.2169 0.084941
5.189 0.98809 5.4908e-005 3.8183 0.011975 6.7835e-005 0.001161 0.23164 0.00065929 0.2323 0.21431 0 0.032362 0.0389 0 1.285 0.42976 0.12995 0.016211 9.1194 0.10104 0.00012789 0.78909 0.0078869 0.0087776 0.0020634 0.97408 0.79042 4.5658e-006 1.8268e-005 0.15304 0.55333 0.64416 0.0017228 0.59955 0.39439 0.0023131 0.42066 1.2053 1.1999 15.9997 144.9432 0.00053814 -83.2591 0.085941
5.19 0.98809 5.4908e-005 3.8183 0.011975 6.7848e-005 0.001161 0.23165 0.00065929 0.2323 0.21431 0 0.032362 0.0389 0 1.2851 0.42981 0.12997 0.016212 9.1213 0.10105 0.0001279 0.78908 0.0078875 0.0087783 0.0020501 0.97484 0.80089 4.5341e-006 1.8141e-005 0.15304 0.55466 0.64591 0.0017169 0.60158 0.39459 0.0023047 0.42065 1.2077 1.2022 15.9998 144.9432 0.00053626 -83.2985 0.086941
5.191 0.98809 5.4908e-005 3.8183 0.011975 6.7861e-005 0.001161 0.23165 0.00065929 0.2323 0.21431 0 0.032362 0.0389 0 1.2852 0.42986 0.12999 0.016214 9.1233 0.10106 0.00012791 0.78907 0.0078881 0.0087789 0.002038 0.97549 0.81084 4.5047e-006 1.8023e-005 0.15305 0.55598 0.64764 0.0017113 0.60361 0.39478 0.0022969 0.42064 1.21 1.2046 15.9999 144.9432 0.00053439 -83.3352 0.087941
5.192 0.98809 5.4908e-005 3.8183 0.011975 6.7874e-005 0.001161 0.23165 0.00065929 0.23231 0.21431 0 0.032361 0.0389 0 1.2853 0.4299 0.13 0.016215 9.1253 0.10107 0.00012793 0.78906 0.0078887 0.0087796 0.0020264 0.97605 0.82029 4.4773e-006 1.7913e-005 0.15305 0.5573 0.64936 0.0017062 0.60563 0.39498 0.0022897 0.42063 1.2124 1.207 16 144.9432 0.00053253 -83.3696 0.088941
5.193 0.98809 5.4907e-005 3.8183 0.011975 6.7887e-005 0.001161 0.23165 0.00065929 0.23231 0.21431 0 0.032361 0.0389 0 1.2854 0.42995 0.13002 0.016217 9.1273 0.10108 0.00012794 0.78905 0.0078894 0.0087802 0.0020155 0.97653 0.82927 4.4516e-006 1.781e-005 0.15306 0.55862 0.65107 0.0017013 0.60765 0.39517 0.002283 0.42062 1.2147 1.2094 16.0001 144.9432 0.00053068 -83.402 0.089941
5.194 0.98809 5.4907e-005 3.8183 0.011975 6.79e-005 0.001161 0.23166 0.00065929 0.23231 0.21432 0 0.032361 0.0389 0 1.2855 0.43 0.13003 0.016218 9.1292 0.10109 0.00012795 0.78904 0.00789 0.0087809 0.0020053 0.97694 0.8378 4.4277e-006 1.7714e-005 0.15306 0.55993 0.65276 0.0016968 0.60967 0.39537 0.0022767 0.42061 1.2171 1.2117 16.0002 144.9432 0.00052885 -83.4324 0.090941
5.195 0.98809 5.4907e-005 3.8183 0.011975 6.7913e-005 0.001161 0.23166 0.00065929 0.23231 0.21432 0 0.032361 0.0389 0 1.2856 0.43004 0.13005 0.01622 9.1312 0.1011 0.00012796 0.78903 0.0078906 0.0087815 0.0019957 0.9773 0.84589 4.4051e-006 1.7624e-005 0.15307 0.56124 0.65443 0.0016925 0.61168 0.39556 0.0022707 0.4206 1.2194 1.2141 16.0003 144.9432 0.00052702 -83.4612 0.091941
5.196 0.98809 5.4907e-005 3.8183 0.011975 6.7926e-005 0.001161 0.23166 0.00065929 0.23231 0.21432 0 0.032361 0.0389 0 1.2857 0.43009 0.13006 0.016221 9.1332 0.10111 0.00012798 0.78902 0.0078912 0.0087822 0.0019868 0.97761 0.85356 4.3839e-006 1.7538e-005 0.15307 0.56255 0.65609 0.0016884 0.61368 0.39576 0.0022652 0.42059 1.2218 1.2165 16.0004 144.9432 0.0005252 -83.4885 0.092941
5.197 0.98809 5.4907e-005 3.8183 0.011975 6.7939e-005 0.001161 0.23166 0.00065929 0.23232 0.21432 0 0.032361 0.0389 0 1.2858 0.43013 0.13008 0.016223 9.1352 0.10111 0.00012799 0.78901 0.0078918 0.0087828 0.0019783 0.97789 0.86084 4.3638e-006 1.7458e-005 0.15308 0.56385 0.65773 0.0016846 0.61568 0.39596 0.0022599 0.42058 1.2241 1.2188 16.0005 144.9433 0.00052339 -83.5144 0.093941
5.198 0.98809 5.4907e-005 3.8183 0.011975 6.7952e-005 0.001161 0.23166 0.00065929 0.23232 0.21433 0 0.032361 0.0389 0 1.2859 0.43018 0.13009 0.016224 9.1371 0.10112 0.000128 0.789 0.0078924 0.0087835 0.0019702 0.97813 0.86774 4.3447e-006 1.7381e-005 0.15308 0.56514 0.65936 0.0016809 0.61768 0.39615 0.0022549 0.42058 1.2264 1.2212 16.0006 144.9433 0.0005216 -83.5391 0.094941
5.199 0.98809 5.4907e-005 3.8183 0.011975 6.7964e-005 0.001161 0.23167 0.00065929 0.23232 0.21433 0 0.032361 0.0389 0 1.2859 0.43023 0.13011 0.016226 9.1391 0.10113 0.00012802 0.789 0.007893 0.0087842 0.0019625 0.97835 0.87428 4.3266e-006 1.7309e-005 0.15309 0.56644 0.66098 0.0016774 0.61967 0.39635 0.0022502 0.42057 1.2288 1.2235 16.0007 144.9433 0.00051981 -83.5627 0.095941
5.2 0.98809 5.4907e-005 3.8183 0.011975 6.7977e-005 0.001161 0.23167 0.00065929 0.23232 0.21433 0 0.03236 0.0389 0 1.286 0.43027 0.13012 0.016227 9.1411 0.10114 0.00012803 0.78899 0.0078936 0.0087848 0.0019551 0.97854 0.88048 4.3093e-006 1.7239e-005 0.15309 0.56773 0.66258 0.0016741 0.62165 0.39655 0.0022457 0.42056 1.2311 1.2259 16.0008 144.9433 0.00051803 -83.5853 0.096941
5.201 0.98809 5.4907e-005 3.8183 0.011975 6.799e-005 0.001161 0.23167 0.00065929 0.23233 0.21433 0 0.03236 0.0389 0 1.2861 0.43032 0.13014 0.016229 9.1431 0.10115 0.00012804 0.78898 0.0078942 0.0087855 0.0019481 0.97872 0.88636 4.2927e-006 1.7173e-005 0.1531 0.56901 0.66416 0.0016709 0.62363 0.39674 0.0022414 0.42055 1.2334 1.2282 16.0009 144.9433 0.00051626 -83.607 0.097941
5.202 0.98809 5.4907e-005 3.8183 0.011975 6.8003e-005 0.001161 0.23167 0.00065929 0.23233 0.21433 0 0.03236 0.0389 0 1.2862 0.43037 0.13016 0.01623 9.145 0.10116 0.00012806 0.78897 0.0078948 0.0087861 0.0019414 0.97888 0.89192 4.2769e-006 1.711e-005 0.1531 0.57029 0.66574 0.0016679 0.6256 0.39694 0.0022372 0.42055 1.2357 1.2305 16.001 144.9433 0.00051451 -83.6279 0.098941
5.203 0.98809 5.4907e-005 3.8183 0.011975 6.8016e-005 0.001161 0.23168 0.00065929 0.23233 0.21434 0 0.03236 0.0389 0 1.2863 0.43041 0.13017 0.016232 9.147 0.10117 0.00012807 0.78896 0.0078954 0.0087868 0.0019349 0.97903 0.89719 4.2616e-006 1.7048e-005 0.15311 0.57157 0.6673 0.0016649 0.62757 0.39714 0.0022332 0.42054 1.2381 1.2329 16.0011 144.9433 0.00051276 -83.6481 0.099941
5.204 0.98809 5.4907e-005 3.8183 0.011975 6.8029e-005 0.0011611 0.23168 0.00065929 0.23233 0.21434 0 0.03236 0.0389 0 1.2864 0.43046 0.13019 0.016233 9.149 0.10118 0.00012808 0.78895 0.007896 0.0087874 0.0019286 0.97916 0.90218 4.2469e-006 1.699e-005 0.15311 0.57285 0.66884 0.0016621 0.62952 0.39733 0.0022294 0.42054 1.2404 1.2352 16.0012 144.9433 0.00051102 -83.6676 0.10094
5.205 0.98809 5.4907e-005 3.8183 0.011975 6.8042e-005 0.0011611 0.23168 0.00065929 0.23234 0.21434 0 0.03236 0.0389 0 1.2865 0.43051 0.1302 0.016235 9.151 0.10119 0.0001281 0.78894 0.0078966 0.0087881 0.0019226 0.97928 0.90691 4.2327e-006 1.6933e-005 0.15312 0.57412 0.67037 0.0016593 0.63148 0.39753 0.0022257 0.42053 1.2427 1.2375 16.0013 144.9433 0.00050929 -83.6865 0.10194
5.206 0.98809 5.4906e-005 3.8183 0.011975 6.8055e-005 0.0011611 0.23168 0.00065929 0.23234 0.21434 0 0.03236 0.0389 0 1.2866 0.43055 0.13022 0.016236 9.1529 0.1012 0.00012811 0.78893 0.0078972 0.0087887 0.0019168 0.9794 0.91138 4.219e-006 1.6878e-005 0.15312 0.57538 0.67189 0.0016566 0.63342 0.39773 0.0022222 0.42052 1.245 1.2398 16.0014 144.9433 0.00050757 -83.7049 0.10294
5.207 0.98809 5.4906e-005 3.8183 0.011975 6.8068e-005 0.0011611 0.23169 0.00065929 0.23234 0.21435 0 0.03236 0.0389 0 1.2867 0.4306 0.13023 0.016238 9.1549 0.10121 0.00012812 0.78892 0.0078978 0.0087894 0.0019111 0.97951 0.91562 4.2057e-006 1.6824e-005 0.15313 0.57665 0.6734 0.001654 0.63536 0.39793 0.0022187 0.42052 1.2473 1.2422 16.0015 144.9433 0.00050587 -83.7227 0.10394
5.208 0.98809 5.4906e-005 3.8183 0.011975 6.8081e-005 0.0011611 0.23169 0.00065929 0.23234 0.21435 0 0.03236 0.0389 0 1.2868 0.43065 0.13025 0.016239 9.1569 0.10121 0.00012813 0.78891 0.0078985 0.00879 0.0019056 0.97961 0.91963 4.1927e-006 1.6773e-005 0.15313 0.5779 0.67489 0.0016515 0.63729 0.39812 0.0022154 0.42051 1.2496 1.2445 16.0016 144.9433 0.00050417 -83.7401 0.10494
5.209 0.98809 5.4906e-005 3.8183 0.011975 6.8094e-005 0.0011611 0.23169 0.00065929 0.23235 0.21435 0 0.032359 0.0389 0 1.2869 0.43069 0.13026 0.016241 9.1589 0.10122 0.00012815 0.7889 0.0078991 0.0087907 0.0019002 0.97971 0.92342 4.1801e-006 1.6722e-005 0.15314 0.57916 0.67637 0.0016491 0.63921 0.39832 0.0022121 0.42051 1.2519 1.2468 16.0017 144.9433 0.00050248 -83.7571 0.10594
5.21 0.98809 5.4906e-005 3.8183 0.011975 6.8107e-005 0.0011611 0.23169 0.00065929 0.23235 0.21435 0 0.032359 0.0389 0 1.287 0.43074 0.13028 0.016242 9.1609 0.10123 0.00012816 0.7889 0.0078997 0.0087914 0.001895 0.9798 0.92701 4.1679e-006 1.6673e-005 0.15314 0.58041 0.67784 0.0016467 0.64113 0.39852 0.0022089 0.4205 1.2542 1.2491 16.0018 144.9433 0.00050079 -83.7737 0.10694
5.211 0.98809 5.4906e-005 3.8183 0.011975 6.812e-005 0.0011611 0.23169 0.00065929 0.23235 0.21435 0 0.032359 0.0389 0 1.2871 0.43079 0.1303 0.016244 9.1628 0.10124 0.00012817 0.78889 0.0079003 0.008792 0.0018899 0.97989 0.93041 4.1559e-006 1.6625e-005 0.15315 0.58166 0.67929 0.0016443 0.64304 0.39871 0.0022058 0.4205 1.2565 1.2514 16.0018 144.9433 0.00049912 -83.7899 0.10794
5.212 0.98809 5.4906e-005 3.8183 0.011975 6.8133e-005 0.0011611 0.2317 0.00065929 0.23235 0.21436 0 0.032359 0.0389 0 1.2872 0.43083 0.13031 0.016245 9.1648 0.10125 0.00012819 0.78888 0.0079009 0.0087927 0.0018849 0.97997 0.93362 4.1442e-006 1.6578e-005 0.15315 0.5829 0.68073 0.001642 0.64494 0.39891 0.0022028 0.42049 1.2587 1.2537 16.0019 144.9433 0.00049746 -83.8058 0.10894
5.213 0.98809 5.4906e-005 3.8183 0.011975 6.8146e-005 0.0011611 0.2317 0.00065929 0.23235 0.21436 0 0.032359 0.0389 0 1.2873 0.43088 0.13033 0.016247 9.1668 0.10126 0.0001282 0.78887 0.0079015 0.0087933 0.00188 0.98005 0.93666 4.1327e-006 1.6532e-005 0.15315 0.58414 0.68216 0.0016398 0.64684 0.39911 0.0021998 0.42049 1.261 1.256 16.002 144.9433 0.00049581 -83.8214 0.10994
5.214 0.98809 5.4906e-005 3.8183 0.011975 6.8159e-005 0.0011611 0.2317 0.00065929 0.23236 0.21436 0 0.032359 0.0389 0 1.2874 0.43093 0.13034 0.016248 9.1688 0.10127 0.00012821 0.78886 0.0079021 0.008794 0.0018752 0.98013 0.93954 4.1216e-006 1.6488e-005 0.15316 0.58538 0.68358 0.0016376 0.64873 0.39931 0.0021969 0.42049 1.2633 1.2583 16.0021 144.9434 0.00049416 -83.8368 0.11094
5.215 0.98809 5.4906e-005 3.8183 0.011975 6.8172e-005 0.0011611 0.2317 0.00065929 0.23236 0.21436 0 0.032359 0.0389 0 1.2875 0.43097 0.13036 0.01625 9.1708 0.10128 0.00012823 0.78885 0.0079027 0.0087946 0.0018706 0.98021 0.94225 4.1106e-006 1.6444e-005 0.15316 0.58661 0.68498 0.0016354 0.65061 0.3995 0.0021941 0.42048 1.2656 1.2606 16.0022 144.9434 0.00049253 -83.8519 0.11194
5.216 0.98809 5.4906e-005 3.8183 0.011975 6.8185e-005 0.0011611 0.23171 0.00065929 0.23236 0.21437 0 0.032359 0.0389 0 1.2876 0.43102 0.13037 0.016251 9.1728 0.10129 0.00012824 0.78884 0.0079033 0.0087953 0.001866 0.98028 0.94483 4.0998e-006 1.6401e-005 0.15317 0.58784 0.68638 0.0016333 0.65248 0.3997 0.0021912 0.42048 1.2678 1.2629 16.0023 144.9434 0.0004909 -83.8667 0.11294
5.217 0.98809 5.4906e-005 3.8183 0.011975 6.8198e-005 0.0011611 0.23171 0.00065929 0.23236 0.21437 0 0.032358 0.0389 0 1.2877 0.43107 0.13039 0.016253 9.1747 0.1013 0.00012825 0.78883 0.0079039 0.0087959 0.0018615 0.98036 0.94726 4.0892e-006 1.6358e-005 0.15317 0.58906 0.68776 0.0016312 0.65434 0.3999 0.0021885 0.42047 1.2701 1.2651 16.0024 144.9434 0.00048929 -83.8813 0.11394
5.218 0.98809 5.4906e-005 3.8183 0.011975 6.8211e-005 0.0011611 0.23171 0.00065929 0.23237 0.21437 0 0.032358 0.0389 0 1.2878 0.43111 0.1304 0.016254 9.1767 0.10131 0.00012826 0.78882 0.0079045 0.0087966 0.001857 0.98043 0.94956 4.0788e-006 1.6317e-005 0.15318 0.59029 0.68913 0.0016292 0.6562 0.40009 0.0021858 0.42047 1.2724 1.2674 16.0025 144.9434 0.00048768 -83.8957 0.11494
5.219 0.98809 5.4906e-005 3.8183 0.011975 6.8224e-005 0.0011611 0.23171 0.00065929 0.23237 0.21437 0 0.032358 0.0389 0 1.2879 0.43116 0.13042 0.016256 9.1787 0.10132 0.00012828 0.78881 0.0079051 0.0087972 0.0018527 0.98049 0.95174 4.0686e-006 1.6276e-005 0.15318 0.5915 0.69049 0.0016271 0.65805 0.40029 0.0021831 0.42047 1.2746 1.2697 16.0025 144.9434 0.00048608 -83.9099 0.11594
5.22 0.98809 5.4905e-005 3.8183 0.011975 6.8237e-005 0.0011611 0.23172 0.00065929 0.23237 0.21437 0 0.032358 0.0389 0 1.288 0.43121 0.13043 0.016257 9.1807 0.10132 0.00012829 0.7888 0.0079057 0.0087979 0.0018483 0.98056 0.95379 4.0585e-006 1.6235e-005 0.15319 0.59272 0.69184 0.0016251 0.6599 0.40049 0.0021805 0.42047 1.2769 1.272 16.0026 144.9434 0.00048449 -83.9239 0.11694
5.221 0.98809 5.4905e-005 3.8183 0.011975 6.8249e-005 0.0011611 0.23172 0.00065929 0.23237 0.21438 0 0.032358 0.0389 0 1.2881 0.43125 0.13045 0.016259 9.1827 0.10133 0.0001283 0.78879 0.0079063 0.0087985 0.0018441 0.98062 0.95574 4.0486e-006 1.6196e-005 0.15319 0.59393 0.69318 0.0016232 0.66173 0.40069 0.0021779 0.42046 1.2791 1.2742 16.0027 144.9434 0.00048291 -83.9377 0.11794
5.222 0.98809 5.4905e-005 3.8183 0.011975 6.8262e-005 0.0011611 0.23172 0.00065929 0.23238 0.21438 0 0.032358 0.0389 0 1.2881 0.4313 0.13047 0.01626 9.1847 0.10134 0.00012832 0.78879 0.0079069 0.0087992 0.0018399 0.98069 0.95758 4.0388e-006 1.6156e-005 0.1532 0.59513 0.6945 0.0016212 0.66356 0.40088 0.0021754 0.42046 1.2814 1.2765 16.0028 144.9434 0.00048134 -83.9514 0.11894
5.223 0.98809 5.4905e-005 3.8183 0.011975 6.8275e-005 0.0011611 0.23172 0.00065929 0.23238 0.21438 0 0.032358 0.0389 0 1.2882 0.43134 0.13048 0.016262 9.1866 0.10135 0.00012833 0.78878 0.0079075 0.0087998 0.0018358 0.98075 0.95931 4.0292e-006 1.6118e-005 0.1532 0.59634 0.69582 0.0016193 0.66538 0.40108 0.0021729 0.42046 1.2836 1.2787 16.0029 144.9434 0.00047977 -83.9649 0.11994
5.224 0.98809 5.4905e-005 3.8183 0.011975 6.8288e-005 0.0011611 0.23172 0.00065929 0.23238 0.21438 0 0.032358 0.0389 0 1.2883 0.43139 0.1305 0.016263 9.1886 0.10136 0.00012834 0.78877 0.0079081 0.0088005 0.0018317 0.98081 0.96096 4.0197e-006 1.608e-005 0.15321 0.59753 0.69712 0.0016174 0.6672 0.40128 0.0021704 0.42045 1.2858 1.281 16.003 144.9434 0.00047822 -83.9782 0.12094
5.225 0.98809 5.4905e-005 3.8183 0.011975 6.8301e-005 0.0011611 0.23173 0.00065929 0.23238 0.21438 0 0.032358 0.0389 0 1.2884 0.43144 0.13051 0.016264 9.1906 0.10137 0.00012836 0.78876 0.0079087 0.0088011 0.0018277 0.98087 0.96251 4.0103e-006 1.6042e-005 0.15321 0.59873 0.69842 0.0016156 0.669 0.40148 0.002168 0.42045 1.2881 1.2832 16.003 144.9434 0.00047667 -83.9914 0.12194
5.226 0.98809 5.4905e-005 3.8183 0.011975 6.8314e-005 0.0011611 0.23173 0.00065929 0.23238 0.21439 0 0.032357 0.0389 0 1.2885 0.43148 0.13053 0.016266 9.1926 0.10138 0.00012837 0.78875 0.0079094 0.0088018 0.0018238 0.98093 0.96398 4.0011e-006 1.6005e-005 0.15322 0.59992 0.6997 0.0016137 0.6708 0.40167 0.0021655 0.42045 1.2903 1.2855 16.0031 144.9434 0.00047513 -84.0044 0.12294
5.227 0.98809 5.4905e-005 3.8183 0.011975 6.8327e-005 0.0011611 0.23173 0.00065929 0.23239 0.21439 0 0.032357 0.0389 0 1.2886 0.43153 0.13054 0.016267 9.1946 0.10139 0.00012838 0.78874 0.00791 0.0088025 0.0018199 0.98099 0.96537 3.992e-006 1.5969e-005 0.15322 0.60111 0.70097 0.0016119 0.67259 0.40187 0.0021632 0.42045 1.2925 1.2877 16.0032 144.9435 0.0004736 -84.0173 0.12394
5.228 0.98809 5.4905e-005 3.8183 0.011975 6.834e-005 0.0011611 0.23173 0.00065929 0.23239 0.21439 0 0.032357 0.0389 0 1.2887 0.43158 0.13056 0.016269 9.1966 0.1014 0.00012839 0.78873 0.0079106 0.0088031 0.001816 0.98104 0.96668 3.983e-006 1.5933e-005 0.15323 0.60229 0.70224 0.0016101 0.67438 0.40207 0.0021608 0.42045 1.2947 1.29 16.0033 144.9435 0.00047208 -84.0301 0.12494
5.229 0.98809 5.4905e-005 3.8183 0.011975 6.8353e-005 0.0011611 0.23174 0.00065929 0.23239 0.21439 0 0.032357 0.0389 0 1.2888 0.43162 0.13057 0.01627 9.1986 0.10141 0.00012841 0.78872 0.0079112 0.0088038 0.0018122 0.9811 0.96792 3.9741e-006 1.5897e-005 0.15323 0.60348 0.70349 0.0016083 0.67615 0.40227 0.0021585 0.42044 1.2969 1.2922 16.0034 144.9435 0.00047056 -84.0427 0.12594
5.23 0.98809 5.4905e-005 3.8183 0.011975 6.8366e-005 0.0011611 0.23174 0.00065929 0.23239 0.2144 0 0.032357 0.0389 0 1.2889 0.43167 0.13059 0.016272 9.2005 0.10142 0.00012842 0.78871 0.0079118 0.0088044 0.0018085 0.98115 0.96909 3.9653e-006 1.5862e-005 0.15324 0.60465 0.70473 0.0016066 0.67792 0.40246 0.0021562 0.42044 1.2992 1.2944 16.0035 144.9435 0.00046906 -84.0552 0.12694
5.231 0.98809 5.4905e-005 3.8183 0.011974 6.8379e-005 0.0011611 0.23174 0.00065929 0.2324 0.2144 0 0.032357 0.0389 0 1.289 0.43172 0.1306 0.016273 9.2025 0.10142 0.00012843 0.7887 0.0079124 0.0088051 0.0018047 0.98121 0.9702 3.9566e-006 1.5827e-005 0.15324 0.60583 0.70596 0.0016048 0.67968 0.40266 0.0021539 0.42044 1.3014 1.2966 16.0035 144.9435 0.00046756 -84.0676 0.12794
5.232 0.98809 5.4905e-005 3.8183 0.011974 6.8392e-005 0.0011611 0.23174 0.00065929 0.2324 0.2144 0 0.032357 0.0389 0 1.2891 0.43176 0.13062 0.016275 9.2045 0.10143 0.00012845 0.78869 0.007913 0.0088057 0.0018011 0.98126 0.97124 3.948e-006 1.5793e-005 0.15325 0.607 0.70719 0.0016031 0.68144 0.40286 0.0021516 0.42044 1.3036 1.2989 16.0036 144.9435 0.00046607 -84.0798 0.12894
5.233 0.98809 5.4904e-005 3.8183 0.011974 6.8405e-005 0.0011611 0.23175 0.00065929 0.2324 0.2144 0 0.032357 0.0389 0 1.2892 0.43181 0.13064 0.016276 9.2065 0.10144 0.00012846 0.78869 0.0079136 0.0088064 0.0017974 0.98132 0.97223 3.9395e-006 1.5759e-005 0.15325 0.60816 0.7084 0.0016014 0.68318 0.40306 0.0021494 0.42044 1.3058 1.3011 16.0037 144.9435 0.00046459 -84.092 0.12994
5.234 0.98809 5.4904e-005 3.8183 0.011974 6.8418e-005 0.0011611 0.23175 0.00065929 0.2324 0.2144 0 0.032357 0.0389 0 1.2893 0.43186 0.13065 0.016278 9.2085 0.10145 0.00012847 0.78868 0.0079142 0.008807 0.0017938 0.98137 0.97317 3.9311e-006 1.5726e-005 0.15326 0.60933 0.7096 0.0015997 0.68492 0.40326 0.0021472 0.42044 1.308 1.3033 16.0038 144.9435 0.00046312 -84.104 0.13094
5.235 0.98809 5.4904e-005 3.8183 0.011974 6.8431e-005 0.0011611 0.23175 0.00065929 0.2324 0.21441 0 0.032356 0.0389 0 1.2894 0.4319 0.13067 0.016279 9.2105 0.10146 0.00012849 0.78867 0.0079148 0.0088077 0.0017903 0.98142 0.97405 3.9228e-006 1.5692e-005 0.15326 0.61049 0.7108 0.0015981 0.68665 0.40345 0.002145 0.42044 1.3102 1.3055 16.0038 144.9435 0.00046165 -84.116 0.13194
5.236 0.98809 5.4904e-005 3.8183 0.011974 6.8444e-005 0.0011611 0.23175 0.00065929 0.23241 0.21441 0 0.032356 0.0389 0 1.2895 0.43195 0.13068 0.016281 9.2125 0.10147 0.0001285 0.78866 0.0079154 0.0088083 0.0017868 0.98147 0.97489 3.9146e-006 1.566e-005 0.15326 0.61164 0.71198 0.0015964 0.68838 0.40365 0.0021428 0.42044 1.3123 1.3077 16.0039 144.9435 0.00046019 -84.1278 0.13294
5.237 0.98809 5.4904e-005 3.8183 0.011974 6.8457e-005 0.0011612 0.23175 0.00065929 0.23241 0.21441 0 0.032356 0.0389 0 1.2896 0.432 0.1307 0.016282 9.2145 0.10148 0.00012851 0.78865 0.007916 0.008809 0.0017833 0.98152 0.97568 3.9065e-006 1.5627e-005 0.15327 0.61279 0.71316 0.0015948 0.69009 0.40385 0.0021407 0.42043 1.3145 1.3099 16.004 144.9435 0.00045874 -84.1395 0.13394
5.238 0.98809 5.4904e-005 3.8183 0.011974 6.847e-005 0.0011612 0.23176 0.00065929 0.23241 0.21441 0 0.032356 0.0389 0 1.2897 0.43204 0.13071 0.016284 9.2165 0.10149 0.00012852 0.78864 0.0079166 0.0088096 0.0017799 0.98157 0.97642 3.8985e-006 1.5595e-005 0.15327 0.61394 0.71433 0.0015931 0.6918 0.40405 0.0021386 0.42043 1.3167 1.3121 16.0041 144.9435 0.0004573 -84.1511 0.13494
5.239 0.98809 5.4904e-005 3.8183 0.011974 6.8483e-005 0.0011612 0.23176 0.00065929 0.23241 0.21441 0 0.032356 0.0389 0 1.2898 0.43209 0.13073 0.016285 9.2184 0.1015 0.00012854 0.78863 0.0079172 0.0088103 0.0017765 0.98162 0.97713 3.8906e-006 1.5563e-005 0.15328 0.61509 0.71548 0.0015915 0.6935 0.40424 0.0021365 0.42043 1.3189 1.3143 16.0042 144.9436 0.00045587 -84.1626 0.13594
5.24 0.98809 5.4904e-005 3.8183 0.011974 6.8496e-005 0.0011612 0.23176 0.00065929 0.23242 0.21442 0 0.032356 0.0389 0 1.2899 0.43214 0.13074 0.016287 9.2204 0.10151 0.00012855 0.78862 0.0079178 0.0088109 0.0017731 0.98167 0.9778 3.8827e-006 1.5532e-005 0.15328 0.61623 0.71663 0.0015899 0.6952 0.40444 0.0021344 0.42043 1.3211 1.3165 16.0042 144.9436 0.00045444 -84.1741 0.13694
5.241 0.98809 5.4904e-005 3.8183 0.011974 6.8509e-005 0.0011612 0.23176 0.00065929 0.23242 0.21442 0 0.032356 0.0389 0 1.29 0.43218 0.13076 0.016288 9.2224 0.10152 0.00012856 0.78861 0.0079184 0.0088116 0.0017698 0.98172 0.97843 3.8749e-006 1.5501e-005 0.15329 0.61737 0.71777 0.0015884 0.69688 0.40464 0.0021324 0.42043 1.3232 1.3187 16.0043 144.9436 0.00045302 -84.1854 0.13794
5.242 0.98809 5.4904e-005 3.8183 0.011974 6.8522e-005 0.0011612 0.23177 0.00065929 0.23242 0.21442 0 0.032356 0.0389 0 1.2901 0.43223 0.13077 0.01629 9.2244 0.10152 0.00012858 0.7886 0.007919 0.0088122 0.0017665 0.98177 0.97902 3.8673e-006 1.547e-005 0.15329 0.6185 0.7189 0.0015868 0.69856 0.40484 0.0021303 0.42043 1.3254 1.3208 16.0044 144.9436 0.00045161 -84.1966 0.13894
5.243 0.98809 5.4904e-005 3.8183 0.011974 6.8534e-005 0.0011612 0.23177 0.00065929 0.23242 0.21442 0 0.032356 0.0389 0 1.2902 0.43228 0.13079 0.016291 9.2264 0.10153 0.00012859 0.7886 0.0079196 0.0088129 0.0017632 0.98181 0.97959 3.8596e-006 1.5439e-005 0.1533 0.61964 0.72003 0.0015853 0.70023 0.40503 0.0021283 0.42043 1.3275 1.323 16.0045 144.9436 0.00045021 -84.2077 0.13994
5.244 0.98809 5.4904e-005 3.8183 0.011974 6.8547e-005 0.0011612 0.23177 0.00065929 0.23242 0.21443 0 0.032355 0.0389 0 1.2902 0.43232 0.13081 0.016293 9.2284 0.10154 0.0001286 0.78859 0.0079202 0.0088135 0.00176 0.98186 0.98012 3.8521e-006 1.5409e-005 0.1533 0.62076 0.72114 0.0015837 0.70189 0.40523 0.0021263 0.42043 1.3297 1.3252 16.0045 144.9436 0.00044881 -84.2188 0.14094
5.245 0.98809 5.4904e-005 3.8183 0.011974 6.856e-005 0.0011612 0.23177 0.00065929 0.23243 0.21443 0 0.032355 0.0389 0 1.2903 0.43237 0.13082 0.016294 9.2304 0.10155 0.00012862 0.78858 0.0079208 0.0088142 0.0017568 0.9819 0.98063 3.8447e-006 1.538e-005 0.15331 0.62189 0.72224 0.0015822 0.70355 0.40543 0.0021243 0.42043 1.3318 1.3273 16.0046 144.9436 0.00044742 -84.2297 0.14194
5.246 0.98809 5.4904e-005 3.8183 0.011974 6.8573e-005 0.0011612 0.23177 0.00065929 0.23243 0.21443 0 0.032355 0.0389 0 1.2904 0.43242 0.13084 0.016296 9.2324 0.10156 0.00012863 0.78857 0.0079214 0.0088148 0.0017536 0.98195 0.9811 3.8373e-006 1.535e-005 0.15331 0.62301 0.72334 0.0015807 0.7052 0.40563 0.0021223 0.42043 1.334 1.3295 16.0047 144.9436 0.00044604 -84.2405 0.14294
5.247 0.98809 5.4903e-005 3.8183 0.011974 6.8586e-005 0.0011612 0.23178 0.00065929 0.23243 0.21443 0 0.032355 0.0389 0 1.2905 0.43246 0.13085 0.016297 9.2344 0.10157 0.00012864 0.78856 0.007922 0.0088155 0.0017505 0.98199 0.98155 3.83e-006 1.5321e-005 0.15332 0.62413 0.72443 0.0015792 0.70684 0.40583 0.0021204 0.42043 1.3361 1.3317 16.0047 144.9436 0.00044467 -84.2513 0.14394
5.248 0.98809 5.4903e-005 3.8183 0.011974 6.8599e-005 0.0011612 0.23178 0.00065929 0.23243 0.21443 0 0.032355 0.0389 0 1.2906 0.43251 0.13087 0.016299 9.2364 0.10158 0.00012865 0.78855 0.0079226 0.0088161 0.0017474 0.98204 0.98198 3.8228e-006 1.5292e-005 0.15332 0.62524 0.72551 0.0015778 0.70847 0.40602 0.0021185 0.42044 1.3383 1.3338 16.0048 144.9436 0.0004433 -84.262 0.14494
5.249 0.98809 5.4903e-005 3.8183 0.011974 6.8612e-005 0.0011612 0.23178 0.00065929 0.23244 0.21444 0 0.032355 0.0389 0 1.2907 0.43255 0.13088 0.0163 9.2384 0.10159 0.00012867 0.78854 0.0079232 0.0088168 0.0017443 0.98208 0.98238 3.8156e-006 1.5263e-005 0.15333 0.62635 0.72658 0.0015763 0.7101 0.40622 0.0021166 0.42044 1.3404 1.336 16.0049 144.9437 0.00044194 -84.2726 0.14594
5.25 0.98809 5.4903e-005 3.8183 0.011974 6.8625e-005 0.0011612 0.23178 0.00065929 0.23244 0.21444 0 0.032355 0.0389 0 1.2908 0.4326 0.1309 0.016301 9.2404 0.1016 0.00012868 0.78853 0.0079238 0.0088174 0.0017413 0.98213 0.98277 3.8085e-006 1.5235e-005 0.15333 0.62746 0.72765 0.0015749 0.71172 0.40642 0.0021147 0.42044 1.3425 1.3381 16.005 144.9437 0.00044059 -84.283 0.14694
5.251 0.98809 5.4903e-005 3.8183 0.011974 6.8638e-005 0.0011612 0.23179 0.00065929 0.23244 0.21444 0 0.032355 0.0389 0 1.2909 0.43265 0.13091 0.016303 9.2424 0.10161 0.00012869 0.78852 0.0079244 0.0088181 0.0017383 0.98217 0.98313 3.8015e-006 1.5207e-005 0.15334 0.62856 0.7287 0.0015734 0.71333 0.40662 0.0021128 0.42044 1.3447 1.3402 16.005 144.9437 0.00043925 -84.2934 0.14794
5.252 0.98809 5.4903e-005 3.8183 0.011974 6.8651e-005 0.0011612 0.23179 0.00065929 0.23244 0.21444 0 0.032355 0.0389 0 1.291 0.43269 0.13093 0.016304 9.2444 0.10162 0.00012871 0.78851 0.007925 0.0088187 0.0017353 0.98221 0.98347 3.7946e-006 1.5179e-005 0.15334 0.62967 0.72975 0.001572 0.71493 0.40681 0.0021109 0.42044 1.3468 1.3424 16.0051 144.9437 0.00043791 -84.3038 0.14894
5.253 0.98809 5.4903e-005 3.8183 0.011974 6.8664e-005 0.0011612 0.23179 0.00065929 0.23245 0.21444 0 0.032354 0.0389 0 1.2911 0.43274 0.13094 0.016306 9.2463 0.10162 0.00012872 0.7885 0.0079256 0.0088194 0.0017323 0.98225 0.98379 3.7877e-006 1.5152e-005 0.15335 0.63076 0.73079 0.0015706 0.71653 0.40701 0.0021091 0.42044 1.3489 1.3445 16.0052 144.9437 0.00043658 -84.314 0.14994
5.254 0.98809 5.4903e-005 3.8183 0.011974 6.8677e-005 0.0011612 0.23179 0.00065929 0.23245 0.21445 0 0.032354 0.0389 0 1.2912 0.43279 0.13096 0.016307 9.2483 0.10163 0.00012873 0.7885 0.0079263 0.00882 0.0017294 0.9823 0.9841 3.7809e-006 1.5124e-005 0.15335 0.63186 0.73183 0.0015692 0.71812 0.40721 0.0021073 0.42044 1.351 1.3466 16.0052 144.9437 0.00043525 -84.3242 0.15094
5.255 0.98809 5.4903e-005 3.8183 0.011974 6.869e-005 0.0011612 0.23179 0.00065929 0.23245 0.21445 0 0.032354 0.0389 0 1.2913 0.43283 0.13098 0.016309 9.2503 0.10164 0.00012874 0.78849 0.0079269 0.0088207 0.0017265 0.98234 0.98439 3.7742e-006 1.5098e-005 0.15336 0.63295 0.73285 0.0015678 0.7197 0.40741 0.0021055 0.42044 1.3531 1.3488 16.0053 144.9437 0.00043394 -84.3342 0.15194
5.256 0.98809 5.4903e-005 3.8183 0.011974 6.8703e-005 0.0011612 0.2318 0.00065929 0.23245 0.21445 0 0.032354 0.0389 0 1.2914 0.43288 0.13099 0.01631 9.2523 0.10165 0.00012876 0.78848 0.0079275 0.0088213 0.0017236 0.98238 0.98466 3.7675e-006 1.5071e-005 0.15336 0.63404 0.73387 0.0015664 0.72128 0.4076 0.0021037 0.42045 1.3552 1.3509 16.0054 144.9437 0.00043263 -84.3442 0.15294
5.257 0.98809 5.4903e-005 3.8183 0.011974 6.8716e-005 0.0011612 0.2318 0.00065929 0.23245 0.21445 0 0.032354 0.0389 0 1.2915 0.43293 0.13101 0.016312 9.2543 0.10166 0.00012877 0.78847 0.0079281 0.008822 0.0017208 0.98242 0.98492 3.7609e-006 1.5044e-005 0.15336 0.63512 0.73488 0.0015651 0.72284 0.4078 0.0021019 0.42045 1.3573 1.353 16.0054 144.9437 0.00043133 -84.3541 0.15394
5.258 0.98809 5.4903e-005 3.8183 0.011974 6.8729e-005 0.0011612 0.2318 0.00065929 0.23246 0.21446 0 0.032354 0.0389 0 1.2916 0.43297 0.13102 0.016313 9.2563 0.10167 0.00012878 0.78846 0.0079287 0.0088226 0.001718 0.98246 0.98517 3.7544e-006 1.5018e-005 0.15337 0.6362 0.73588 0.0015637 0.7244 0.408 0.0021001 0.42045 1.3594 1.3551 16.0055 144.9437 0.00043003 -84.364 0.15494
5.259 0.98809 5.4903e-005 3.8183 0.011974 6.8742e-005 0.0011612 0.2318 0.00065929 0.23246 0.21446 0 0.032354 0.0389 0 1.2917 0.43302 0.13104 0.016315 9.2583 0.10168 0.0001288 0.78845 0.0079293 0.0088233 0.0017152 0.9825 0.9854 3.7479e-006 1.4992e-005 0.15337 0.63728 0.73688 0.0015624 0.72596 0.4082 0.0020984 0.42045 1.3615 1.3572 16.0056 144.9438 0.00042874 -84.3737 0.15594
5.26 0.98809 5.4902e-005 3.8183 0.011974 6.8755e-005 0.0011612 0.23181 0.00065929 0.23246 0.21446 0 0.032354 0.0389 0 1.2918 0.43307 0.13105 0.016316 9.2603 0.10169 0.00012881 0.78844 0.0079299 0.0088239 0.0017125 0.98254 0.98562 3.7415e-006 1.4967e-005 0.15338 0.63835 0.73787 0.0015611 0.7275 0.4084 0.0020967 0.42045 1.3636 1.3593 16.0056 144.9438 0.00042746 -84.3834 0.15694
5.261 0.98809 5.4902e-005 3.8183 0.011974 6.8768e-005 0.0011612 0.23181 0.00065929 0.23246 0.21446 0 0.032354 0.0389 0 1.2919 0.43311 0.13107 0.016318 9.2623 0.1017 0.00012882 0.78843 0.0079305 0.0088246 0.0017097 0.98257 0.98583 3.7351e-006 1.4941e-005 0.15338 0.63942 0.73885 0.0015598 0.72904 0.40859 0.002095 0.42046 1.3657 1.3614 16.0057 144.9438 0.00042618 -84.393 0.15794
5.262 0.98809 5.4902e-005 3.8183 0.011974 6.8781e-005 0.0011612 0.23181 0.00065929 0.23247 0.21446 0 0.032353 0.0389 0 1.292 0.43316 0.13108 0.016319 9.2643 0.10171 0.00012884 0.78842 0.0079311 0.0088252 0.001707 0.98261 0.98603 3.7289e-006 1.4916e-005 0.15339 0.64049 0.73982 0.0015585 0.73057 0.40879 0.0020933 0.42046 1.3678 1.3635 16.0058 144.9438 0.00042491 -84.4025 0.15894
5.263 0.98809 5.4902e-005 3.8183 0.011974 6.8794e-005 0.0011612 0.23181 0.00065929 0.23247 0.21447 0 0.032353 0.0389 0 1.2921 0.43321 0.1311 0.016321 9.2663 0.10171 0.00012885 0.78841 0.0079317 0.0088259 0.0017044 0.98265 0.98622 3.7226e-006 1.4891e-005 0.15339 0.64155 0.74079 0.0015572 0.73209 0.40899 0.0020916 0.42046 1.3698 1.3656 16.0058 144.9438 0.00042365 -84.412 0.15994
5.264 0.98809 5.4902e-005 3.8183 0.011974 6.8806e-005 0.0011612 0.23181 0.00065929 0.23247 0.21447 0 0.032353 0.0389 0 1.2922 0.43325 0.13111 0.016322 9.2683 0.10172 0.00012886 0.7884 0.0079323 0.0088265 0.0017017 0.98269 0.98639 3.7165e-006 1.4867e-005 0.1534 0.64262 0.74175 0.0015559 0.73361 0.40919 0.0020899 0.42046 1.3719 1.3677 16.0059 144.9438 0.0004224 -84.4213 0.16094
5.265 0.98809 5.4902e-005 3.8183 0.011974 6.8819e-005 0.0011612 0.23182 0.00065929 0.23247 0.21447 0 0.032353 0.0389 0 1.2923 0.4333 0.13113 0.016324 9.2703 0.10173 0.00012887 0.7884 0.0079329 0.0088272 0.0016991 0.98272 0.98656 3.7104e-006 1.4842e-005 0.1534 0.64367 0.7427 0.0015546 0.73512 0.40938 0.0020883 0.42047 1.374 1.3698 16.006 144.9438 0.00042115 -84.4306 0.16194
5.266 0.98809 5.4902e-005 3.8183 0.011974 6.8832e-005 0.0011612 0.23182 0.0006593 0.23247 0.21447 0 0.032353 0.0389 0 1.2924 0.43335 0.13114 0.016325 9.2723 0.10174 0.00012889 0.78839 0.0079335 0.0088278 0.0016965 0.98276 0.98672 3.7043e-006 1.4818e-005 0.15341 0.64473 0.74365 0.0015534 0.73662 0.40958 0.0020866 0.42047 1.376 1.3718 16.006 144.9438 0.0004199 -84.4398 0.16294
5.267 0.98809 5.4902e-005 3.8183 0.011974 6.8845e-005 0.0011612 0.23182 0.0006593 0.23248 0.21447 0 0.032353 0.0389 0 1.2924 0.43339 0.13116 0.016327 9.2743 0.10175 0.0001289 0.78838 0.0079341 0.0088285 0.0016939 0.9828 0.98688 3.6983e-006 1.4794e-005 0.15341 0.64578 0.74459 0.0015522 0.73811 0.40978 0.002085 0.42047 1.3781 1.3739 16.0061 144.9438 0.00041867 -84.449 0.16394
5.268 0.98809 5.4902e-005 3.8183 0.011974 6.8858e-005 0.0011612 0.23182 0.0006593 0.23248 0.21448 0 0.032353 0.0389 0 1.2925 0.43344 0.13118 0.016328 9.2763 0.10176 0.00012891 0.78837 0.0079347 0.0088291 0.0016913 0.98283 0.98702 3.6924e-006 1.477e-005 0.15342 0.64683 0.74552 0.0015509 0.7396 0.40998 0.0020834 0.42047 1.3801 1.376 16.0061 144.9439 0.00041744 -84.4581 0.16494
5.269 0.98809 5.4902e-005 3.8183 0.011974 6.8871e-005 0.0011613 0.23183 0.0006593 0.23248 0.21448 0 0.032353 0.0389 0 1.2926 0.43349 0.13119 0.01633 9.2783 0.10177 0.00012893 0.78836 0.0079353 0.0088298 0.0016888 0.98287 0.98716 3.6865e-006 1.4747e-005 0.15342 0.64787 0.74645 0.0015497 0.74108 0.41017 0.0020818 0.42048 1.3822 1.378 16.0062 144.9439 0.00041621 -84.4671 0.16594
5.27 0.98809 5.4902e-005 3.8183 0.011974 6.8884e-005 0.0011613 0.23183 0.0006593 0.23248 0.21448 0 0.032353 0.0389 0 1.2927 0.43353 0.13121 0.016331 9.2803 0.10178 0.00012894 0.78835 0.0079359 0.0088304 0.0016863 0.9829 0.98729 3.6807e-006 1.4723e-005 0.15343 0.64891 0.74737 0.0015485 0.74255 0.41037 0.0020802 0.42048 1.3842 1.3801 16.0063 144.9439 0.000415 -84.476 0.16694
5.271 0.98809 5.4902e-005 3.8183 0.011974 6.8897e-005 0.0011613 0.23183 0.0006593 0.23248 0.21448 0 0.032352 0.0389 0 1.2928 0.43358 0.13122 0.016333 9.2823 0.10179 0.00012895 0.78834 0.0079365 0.0088311 0.0016838 0.98294 0.98741 3.6749e-006 1.47e-005 0.15343 0.64995 0.74829 0.0015473 0.74402 0.41057 0.0020786 0.42048 1.3863 1.3822 16.0063 144.9439 0.00041379 -84.4848 0.16794
5.272 0.98809 5.4902e-005 3.8183 0.011974 6.891e-005 0.0011613 0.23183 0.0006593 0.23249 0.21448 0 0.032352 0.0389 0 1.2929 0.43362 0.13124 0.016334 9.2843 0.1018 0.00012897 0.78833 0.0079371 0.0088317 0.0016814 0.98297 0.98753 3.6692e-006 1.4677e-005 0.15344 0.65099 0.74919 0.0015461 0.74548 0.41077 0.0020771 0.42049 1.3883 1.3842 16.0064 144.9439 0.00041258 -84.4936 0.16894
5.273 0.98809 5.4901e-005 3.8183 0.011974 6.8923e-005 0.0011613 0.23183 0.0006593 0.23249 0.21449 0 0.032352 0.0389 0 1.293 0.43367 0.13125 0.016335 9.2863 0.10181 0.00012898 0.78832 0.0079377 0.0088324 0.0016789 0.98301 0.98764 3.6635e-006 1.4655e-005 0.15344 0.65202 0.7501 0.0015449 0.74693 0.41097 0.0020755 0.42049 1.3903 1.3862 16.0065 144.9439 0.00041138 -84.5024 0.16994
5.274 0.98809 5.4901e-005 3.8183 0.011974 6.8936e-005 0.0011613 0.23184 0.0006593 0.23249 0.21449 0 0.032352 0.0389 0 1.2931 0.43372 0.13127 0.016337 9.2883 0.10181 0.00012899 0.78831 0.0079383 0.008833 0.0016765 0.98304 0.98775 3.6579e-006 1.4632e-005 0.15345 0.65305 0.75099 0.0015438 0.74838 0.41116 0.002074 0.42049 1.3924 1.3883 16.0065 144.9439 0.00041019 -84.511 0.17094
5.275 0.98809 5.4901e-005 3.8183 0.011974 6.8949e-005 0.0011613 0.23184 0.0006593 0.23249 0.21449 0 0.032352 0.0389 0 1.2932 0.43376 0.13128 0.016338 9.2903 0.10182 0.000129 0.78831 0.0079389 0.0088336 0.0016741 0.98308 0.98785 3.6524e-006 1.461e-005 0.15345 0.65407 0.75188 0.0015426 0.74981 0.41136 0.0020725 0.4205 1.3944 1.3903 16.0066 144.9439 0.00040901 -84.5196 0.17194
5.276 0.98809 5.4901e-005 3.8183 0.011974 6.8962e-005 0.0011613 0.23184 0.0006593 0.2325 0.21449 0 0.032352 0.0389 0 1.2933 0.43381 0.1313 0.01634 9.2923 0.10183 0.00012902 0.7883 0.0079395 0.0088343 0.0016717 0.98311 0.98795 3.6469e-006 1.4588e-005 0.15345 0.6551 0.75276 0.0015414 0.75124 0.41156 0.002071 0.4205 1.3964 1.3924 16.0066 144.9439 0.00040783 -84.5281 0.17294
5.277 0.98809 5.4901e-005 3.8183 0.011974 6.8975e-005 0.0011613 0.23184 0.0006593 0.2325 0.2145 0 0.032352 0.0389 0 1.2934 0.43386 0.13131 0.016341 9.2943 0.10184 0.00012903 0.78829 0.0079401 0.0088349 0.0016694 0.98314 0.98804 3.6414e-006 1.4566e-005 0.15346 0.65612 0.75364 0.0015403 0.75267 0.41176 0.0020695 0.4205 1.3984 1.3944 16.0067 144.944 0.00040665 -84.5366 0.17394
5.278 0.98809 5.4901e-005 3.8183 0.011974 6.8988e-005 0.0011613 0.23185 0.0006593 0.2325 0.2145 0 0.032352 0.0389 0 1.2935 0.4339 0.13133 0.016343 9.2963 0.10185 0.00012904 0.78828 0.0079407 0.0088356 0.0016671 0.98317 0.98813 3.636e-006 1.4545e-005 0.15346 0.65713 0.75451 0.0015392 0.75408 0.41195 0.002068 0.42051 1.4004 1.3964 16.0067 144.944 0.00040549 -84.5449 0.17494
5.279 0.98809 5.4901e-005 3.8183 0.011974 6.9001e-005 0.0011613 0.23185 0.0006593 0.2325 0.2145 0 0.032352 0.0389 0 1.2936 0.43395 0.13135 0.016344 9.2983 0.10186 0.00012906 0.78827 0.0079413 0.0088362 0.0016648 0.98321 0.98821 3.6307e-006 1.4523e-005 0.15347 0.65815 0.75537 0.0015381 0.75549 0.41215 0.0020666 0.42051 1.4024 1.3984 16.0068 144.944 0.00040433 -84.5533 0.17594
5.28 0.98809 5.4901e-005 3.8183 0.011974 6.9014e-005 0.0011613 0.23185 0.0006593 0.2325 0.2145 0 0.032351 0.0389 0 1.2937 0.434 0.13136 0.016346 9.3004 0.10187 0.00012907 0.78826 0.0079419 0.0088369 0.0016625 0.98324 0.98829 3.6254e-006 1.4502e-005 0.15347 0.65916 0.75623 0.001537 0.7569 0.41235 0.0020651 0.42052 1.4044 1.4004 16.0069 144.944 0.00040317 -84.5615 0.17694
5.281 0.98809 5.4901e-005 3.8183 0.011974 6.9027e-005 0.0011613 0.23185 0.0006593 0.23251 0.2145 0 0.032351 0.0389 0 1.2938 0.43404 0.13138 0.016347 9.3024 0.10188 0.00012908 0.78825 0.0079425 0.0088375 0.0016603 0.98327 0.98837 3.6202e-006 1.4481e-005 0.15348 0.66016 0.75709 0.0015359 0.75829 0.41255 0.0020637 0.42052 1.4064 1.4025 16.0069 144.944 0.00040202 -84.5697 0.17794
5.282 0.98809 5.4901e-005 3.8183 0.011974 6.904e-005 0.0011613 0.23185 0.0006593 0.23251 0.21451 0 0.032351 0.0389 0 1.2939 0.43409 0.13139 0.016349 9.3044 0.10189 0.00012909 0.78824 0.0079431 0.0088382 0.0016581 0.9833 0.98844 3.615e-006 1.446e-005 0.15348 0.66117 0.75793 0.0015348 0.75968 0.41274 0.0020622 0.42052 1.4084 1.4045 16.007 144.944 0.00040088 -84.5778 0.17894
5.283 0.98809 5.4901e-005 3.8183 0.011974 6.9053e-005 0.0011613 0.23186 0.0006593 0.23251 0.21451 0 0.032351 0.0389 0 1.294 0.43414 0.13141 0.01635 9.3064 0.1019 0.00012911 0.78823 0.0079437 0.0088388 0.0016558 0.98333 0.98851 3.6098e-006 1.444e-005 0.15349 0.66217 0.75877 0.0015337 0.76106 0.41294 0.0020608 0.42053 1.4104 1.4065 16.007 144.944 0.00039974 -84.5859 0.17994
5.284 0.98809 5.4901e-005 3.8183 0.011974 6.9066e-005 0.0011613 0.23186 0.0006593 0.23251 0.21451 0 0.032351 0.0389 0 1.2941 0.43418 0.13142 0.016352 9.3084 0.10191 0.00012912 0.78822 0.0079443 0.0088395 0.0016535 0.98336 0.98858 3.6047e-006 1.4419e-005 0.15349 0.66317 0.75961 0.0015326 0.76244 0.41314 0.0020594 0.42053 1.4124 1.4085 16.0071 144.944 0.00039861 -84.5939 0.18094
5.285 0.98809 5.4901e-005 3.8183 0.011974 6.9078e-005 0.0011613 0.23186 0.0006593 0.23252 0.21451 0 0.032351 0.0389 0 1.2942 0.43423 0.13144 0.016353 9.3104 0.10191 0.00012913 0.78821 0.0079449 0.0088401 0.0016512 0.98339 0.98864 3.5996e-006 1.4399e-005 0.1535 0.66416 0.76044 0.0015315 0.7638 0.41334 0.002058 0.42054 1.4144 1.4105 16.0071 144.9441 0.00039748 -84.6018 0.18194
5.286 0.98809 5.4901e-005 3.8183 0.011974 6.9091e-005 0.0011613 0.23186 0.0006593 0.23252 0.21451 0 0.032351 0.0389 0 1.2943 0.43428 0.13145 0.016355 9.3124 0.10192 0.00012915 0.78821 0.0079455 0.0088408 0.001649 0.98342 0.9887 3.5946e-006 1.4379e-005 0.1535 0.66515 0.76127 0.0015304 0.76516 0.41353 0.0020567 0.42054 1.4164 1.4124 16.0072 144.9441 0.00039636 -84.6097 0.18294
5.287 0.98809 5.49e-005 3.8183 0.011974 6.9104e-005 0.0011613 0.23187 0.0006593 0.23252 0.21452 0 0.032351 0.0389 0 1.2944 0.43432 0.13147 0.016356 9.3144 0.10193 0.00012916 0.7882 0.0079461 0.0088414 0.0016468 0.98345 0.98876 3.5896e-006 1.4359e-005 0.15351 0.66614 0.76208 0.0015294 0.76652 0.41373 0.0020553 0.42055 1.4183 1.4144 16.0073 144.9441 0.00039525 -84.6175 0.18394
5.288 0.98809 5.49e-005 3.8183 0.011974 6.9117e-005 0.0011613 0.23187 0.0006593 0.23252 0.21452 0 0.032351 0.0389 0 1.2944 0.43437 0.13148 0.016358 9.3164 0.10194 0.00012917 0.78819 0.0079467 0.0088421 0.0016447 0.98348 0.98882 3.5847e-006 1.4339e-005 0.15351 0.66713 0.7629 0.0015284 0.76787 0.41393 0.0020539 0.42055 1.4203 1.4164 16.0073 144.9441 0.00039414 -84.6252 0.18494
5.289 0.98809 5.49e-005 3.8183 0.011974 6.913e-005 0.0011613 0.23187 0.0006593 0.23252 0.21452 0 0.03235 0.0389 0 1.2945 0.43442 0.1315 0.016359 9.3184 0.10195 0.00012919 0.78818 0.0079473 0.0088427 0.0016426 0.98351 0.98887 3.5798e-006 1.432e-005 0.15352 0.66811 0.76371 0.0015273 0.76921 0.41413 0.0020526 0.42056 1.4222 1.4184 16.0074 144.9441 0.00039303 -84.6329 0.18594
5.29 0.98809 5.49e-005 3.8183 0.011974 6.9143e-005 0.0011613 0.23187 0.0006593 0.23253 0.21452 0 0.03235 0.0389 0 1.2946 0.43446 0.13152 0.016361 9.3204 0.10196 0.0001292 0.78817 0.0079479 0.0088433 0.0016406 0.98354 0.98892 3.575e-006 1.4301e-005 0.15352 0.66909 0.76451 0.0015263 0.77054 0.41432 0.0020513 0.42056 1.4242 1.4204 16.0074 144.9441 0.00039194 -84.6405 0.18694
5.291 0.98809 5.49e-005 3.8183 0.011974 6.9156e-005 0.0011613 0.23187 0.0006593 0.23253 0.21452 0 0.03235 0.0389 0 1.2947 0.43451 0.13153 0.016362 9.3224 0.10197 0.00012921 0.78816 0.0079485 0.008844 0.0016386 0.98357 0.98897 3.5702e-006 1.4281e-005 0.15353 0.67007 0.76531 0.0015253 0.77187 0.41452 0.0020499 0.42057 1.4262 1.4223 16.0075 144.9441 0.00039084 -84.6481 0.18794
5.292 0.98809 5.49e-005 3.8183 0.011974 6.9169e-005 0.0011613 0.23188 0.0006593 0.23253 0.21453 0 0.03235 0.0389 0 1.2948 0.43456 0.13155 0.016363 9.3244 0.10198 0.00012922 0.78815 0.0079491 0.0088446 0.0016366 0.9836 0.98902 3.5655e-006 1.4263e-005 0.15353 0.67104 0.7661 0.0015243 0.77319 0.41472 0.0020486 0.42057 1.4281 1.4243 16.0075 144.9441 0.00038976 -84.6556 0.18894
5.293 0.98809 5.49e-005 3.8183 0.011973 6.9182e-005 0.0011613 0.23188 0.0006593 0.23253 0.21453 0 0.03235 0.0389 0 1.2949 0.4346 0.13156 0.016365 9.3264 0.10199 0.00012924 0.78814 0.0079497 0.0088453 0.0016346 0.98362 0.98906 3.5608e-006 1.4244e-005 0.15354 0.67201 0.76689 0.0015233 0.7745 0.41491 0.0020473 0.42058 1.4301 1.4262 16.0076 144.9442 0.00038868 -84.6631 0.18994
5.294 0.98809 5.49e-005 3.8183 0.011973 6.9195e-005 0.0011613 0.23188 0.0006593 0.23253 0.21453 0 0.03235 0.0389 0 1.295 0.43465 0.13158 0.016366 9.3285 0.102 0.00012925 0.78813 0.0079503 0.0088459 0.0016327 0.98365 0.98911 3.5562e-006 1.4225e-005 0.15354 0.67298 0.76767 0.0015224 0.77581 0.41511 0.002046 0.42058 1.432 1.4282 16.0076 144.9442 0.0003876 -84.6705 0.19094
5.295 0.98809 5.49e-005 3.8183 0.011973 6.9208e-005 0.0011613 0.23188 0.0006593 0.23254 0.21453 0 0.03235 0.0389 0 1.2951 0.43469 0.13159 0.016368 9.3305 0.102 0.00012926 0.78812 0.0079509 0.0088466 0.0016307 0.98368 0.98915 3.5516e-006 1.4207e-005 0.15354 0.67394 0.76845 0.0015214 0.77711 0.41531 0.0020448 0.42059 1.4339 1.4301 16.0077 144.9442 0.00038653 -84.6778 0.19194
5.296 0.98809 5.49e-005 3.8183 0.011973 6.9221e-005 0.0011613 0.23188 0.0006593 0.23254 0.21453 0 0.03235 0.0389 0 1.2952 0.43474 0.13161 0.016369 9.3325 0.10201 0.00012928 0.78812 0.0079515 0.0088472 0.0016287 0.98371 0.98919 3.547e-006 1.4188e-005 0.15355 0.6749 0.76922 0.0015204 0.7784 0.41551 0.0020435 0.42059 1.4359 1.4321 16.0077 144.9442 0.00038547 -84.6851 0.19294
5.297 0.98809 5.49e-005 3.8183 0.011973 6.9234e-005 0.0011613 0.23189 0.0006593 0.23254 0.21454 0 0.03235 0.0389 0 1.2953 0.43479 0.13162 0.016371 9.3345 0.10202 0.00012929 0.78811 0.0079521 0.0088479 0.0016268 0.98373 0.98923 3.5425e-006 1.417e-005 0.15355 0.67586 0.76999 0.0015195 0.77969 0.4157 0.0020422 0.4206 1.4378 1.434 16.0078 144.9442 0.00038441 -84.6923 0.19394
5.298 0.98809 5.49e-005 3.8183 0.011973 6.9247e-005 0.0011613 0.23189 0.0006593 0.23254 0.21454 0 0.032349 0.0389 0 1.2954 0.43483 0.13164 0.016372 9.3365 0.10203 0.0001293 0.7881 0.0079527 0.0088485 0.0016248 0.98376 0.98927 3.538e-006 1.4152e-005 0.15356 0.67682 0.77075 0.0015185 0.78097 0.4159 0.002041 0.4206 1.4397 1.436 16.0078 144.9442 0.00038335 -84.6995 0.19494
5.299 0.98809 5.49e-005 3.8183 0.011973 6.926e-005 0.0011613 0.23189 0.0006593 0.23255 0.21454 0 0.032349 0.0389 0 1.2955 0.43488 0.13165 0.016374 9.3385 0.10204 0.00012931 0.78809 0.0079533 0.0088492 0.0016229 0.98379 0.9893 3.5335e-006 1.4135e-005 0.15356 0.67777 0.77151 0.0015176 0.78224 0.4161 0.0020398 0.42061 1.4416 1.4379 16.0079 144.9442 0.00038231 -84.7066 0.19594
5.3 0.98809 5.4899e-005 3.8183 0.011973 6.9273e-005 0.0011613 0.23189 0.0006593 0.23255 0.21454 0 0.032349 0.0389 0 1.2956 0.43493 0.13167 0.016375 9.3405 0.10205 0.00012933 0.78808 0.0079539 0.0088498 0.0016209 0.98381 0.98934 3.5291e-006 1.4117e-005 0.15357 0.67872 0.77226 0.0015166 0.78351 0.4163 0.0020385 0.42062 1.4435 1.4398 16.0079 144.9442 0.00038126 -84.7136 0.19694
5.301 0.98809 5.4899e-005 3.8183 0.011973 6.9286e-005 0.0011614 0.2319 0.0006593 0.23255 0.21454 0 0.032349 0.0389 0 1.2957 0.43497 0.13168 0.016377 9.3425 0.10206 0.00012934 0.78807 0.0079545 0.0088505 0.001619 0.98384 0.98937 3.5247e-006 1.4099e-005 0.15357 0.67967 0.77301 0.0015157 0.78477 0.41649 0.0020373 0.42062 1.4455 1.4417 16.008 144.9443 0.00038022 -84.7206 0.19794
5.302 0.98809 5.4899e-005 3.8183 0.011973 6.9299e-005 0.0011614 0.2319 0.0006593 0.23255 0.21455 0 0.032349 0.0389 0 1.2958 0.43502 0.1317 0.016378 9.3445 0.10207 0.00012935 0.78806 0.0079551 0.0088511 0.0016171 0.98387 0.98941 3.5204e-006 1.4082e-005 0.15358 0.68061 0.77375 0.0015148 0.78603 0.41669 0.0020361 0.42063 1.4474 1.4437 16.008 144.9443 0.00037919 -84.7276 0.19894
5.303 0.98809 5.4899e-005 3.8183 0.011973 6.9312e-005 0.0011614 0.2319 0.0006593 0.23255 0.21455 0 0.032349 0.0389 0 1.2959 0.43507 0.13172 0.01638 9.3466 0.10208 0.00012937 0.78805 0.0079557 0.0088517 0.0016153 0.98389 0.98944 3.5161e-006 1.4065e-005 0.15358 0.68155 0.77449 0.0015139 0.78727 0.41689 0.0020349 0.42063 1.4493 1.4456 16.0081 144.9443 0.00037816 -84.7345 0.19994
5.304 0.98809 5.4899e-005 3.8183 0.011973 6.9325e-005 0.0011614 0.2319 0.0006593 0.23256 0.21455 0 0.032349 0.0389 0 1.296 0.43511 0.13173 0.016381 9.3486 0.10209 0.00012938 0.78804 0.0079563 0.0088524 0.0016134 0.98392 0.98947 3.5118e-006 1.4048e-005 0.15359 0.68249 0.77522 0.0015129 0.78851 0.41708 0.0020337 0.42064 1.4512 1.4475 16.0081 144.9443 0.00037714 -84.7413 0.20094
5.305 0.98809 5.4899e-005 3.8183 0.011973 6.9338e-005 0.0011614 0.2319 0.0006593 0.23256 0.21455 0 0.032349 0.0389 0 1.2961 0.43516 0.13175 0.016383 9.3506 0.10209 0.00012939 0.78803 0.0079569 0.008853 0.0016116 0.98394 0.9895 3.5076e-006 1.4031e-005 0.15359 0.68343 0.77595 0.001512 0.78975 0.41728 0.0020326 0.42065 1.453 1.4494 16.0082 144.9443 0.00037612 -84.7481 0.20194
5.306 0.98809 5.4899e-005 3.8183 0.011973 6.935e-005 0.0011614 0.23191 0.0006593 0.23256 0.21455 0 0.032349 0.0389 0 1.2962 0.43521 0.13176 0.016384 9.3526 0.1021 0.00012941 0.78803 0.0079575 0.0088537 0.0016098 0.98397 0.98953 3.5035e-006 1.4014e-005 0.1536 0.68436 0.77667 0.0015112 0.79098 0.41748 0.0020314 0.42065 1.4549 1.4513 16.0082 144.9443 0.00037511 -84.7548 0.20294
5.307 0.98809 5.4899e-005 3.8183 0.011973 6.9363e-005 0.0011614 0.23191 0.0006593 0.23256 0.21456 0 0.032349 0.0389 0 1.2963 0.43525 0.13178 0.016386 9.3546 0.10211 0.00012942 0.78802 0.0079581 0.0088543 0.001608 0.98399 0.98955 3.4993e-006 1.3998e-005 0.1536 0.68529 0.77739 0.0015103 0.7922 0.41767 0.0020303 0.42066 1.4568 1.4532 16.0083 144.9443 0.00037411 -84.7615 0.20394
5.308 0.98809 5.4899e-005 3.8183 0.011973 6.9376e-005 0.0011614 0.23191 0.0006593 0.23256 0.21456 0 0.032348 0.0389 0 1.2964 0.4353 0.13179 0.016387 9.3566 0.10212 0.00012943 0.78801 0.0079587 0.008855 0.0016063 0.98402 0.98958 3.4952e-006 1.3981e-005 0.15361 0.68622 0.77811 0.0015094 0.79341 0.41787 0.0020291 0.42066 1.4587 1.4551 16.0083 144.9444 0.0003731 -84.7681 0.20494
5.309 0.98809 5.4899e-005 3.8183 0.011973 6.9389e-005 0.0011614 0.23191 0.0006593 0.23257 0.21456 0 0.032348 0.0389 0 1.2965 0.43535 0.13181 0.016388 9.3586 0.10213 0.00012944 0.788 0.0079592 0.0088556 0.0016045 0.98404 0.98961 3.4911e-006 1.3965e-005 0.15361 0.68714 0.77882 0.0015085 0.79462 0.41807 0.002028 0.42067 1.4606 1.457 16.0084 144.9444 0.00037211 -84.7747 0.20594
5.31 0.98809 5.4899e-005 3.8183 0.011973 6.9402e-005 0.0011614 0.23191 0.0006593 0.23257 0.21456 0 0.032348 0.0389 0 1.2965 0.43539 0.13182 0.01639 9.3607 0.10214 0.00012946 0.78799 0.0079598 0.0088563 0.0016028 0.98406 0.98963 3.4871e-006 1.3949e-005 0.15362 0.68806 0.77952 0.0015077 0.79583 0.41827 0.0020268 0.42068 1.4624 1.4588 16.0084 144.9444 0.00037111 -84.7812 0.20694
5.311 0.98809 5.4899e-005 3.8183 0.011973 6.9415e-005 0.0011614 0.23192 0.0006593 0.23257 0.21456 0 0.032348 0.0389 0 1.2966 0.43544 0.13184 0.016391 9.3627 0.10215 0.00012947 0.78798 0.0079604 0.0088569 0.0016011 0.98409 0.98966 3.4831e-006 1.3933e-005 0.15362 0.68898 0.78023 0.0015068 0.79702 0.41846 0.0020257 0.42068 1.4643 1.4607 16.0085 144.9444 0.00037013 -84.7877 0.20794
5.312 0.98809 5.4899e-005 3.8183 0.011973 6.9428e-005 0.0011614 0.23192 0.0006593 0.23257 0.21457 0 0.032348 0.0389 0 1.2967 0.43549 0.13185 0.016393 9.3647 0.10216 0.00012948 0.78797 0.007961 0.0088575 0.0015994 0.98411 0.98968 3.4792e-006 1.3917e-005 0.15363 0.68989 0.78092 0.001506 0.79821 0.41866 0.0020246 0.42069 1.4662 1.4626 16.0085 144.9444 0.00036915 -84.7942 0.20894
5.313 0.98809 5.4898e-005 3.8183 0.011973 6.9441e-005 0.0011614 0.23192 0.0006593 0.23258 0.21457 0 0.032348 0.0389 0 1.2968 0.43553 0.13187 0.016394 9.3667 0.10217 0.0001295 0.78796 0.0079616 0.0088582 0.0015977 0.98413 0.98971 3.4752e-006 1.3901e-005 0.15363 0.69081 0.78162 0.0015051 0.79939 0.41886 0.0020235 0.4207 1.468 1.4645 16.0085 144.9444 0.00036817 -84.8005 0.20994
5.314 0.98809 5.4898e-005 3.8183 0.011973 6.9454e-005 0.0011614 0.23192 0.0006593 0.23258 0.21457 0 0.032348 0.0389 0 1.2969 0.43558 0.13189 0.016396 9.3687 0.10218 0.00012951 0.78795 0.0079622 0.0088588 0.001596 0.98416 0.98973 3.4713e-006 1.3886e-005 0.15363 0.69172 0.78231 0.0015043 0.80057 0.41905 0.0020224 0.4207 1.4699 1.4663 16.0086 144.9444 0.0003672 -84.8069 0.21094
5.315 0.98809 5.4898e-005 3.8183 0.011973 6.9467e-005 0.0011614 0.23192 0.0006593 0.23258 0.21457 0 0.032348 0.0389 0 1.297 0.43562 0.1319 0.016397 9.3707 0.10219 0.00012952 0.78794 0.0079628 0.0088595 0.0015943 0.98418 0.98975 3.4675e-006 1.387e-005 0.15364 0.69262 0.78299 0.0015035 0.80174 0.41925 0.0020213 0.42071 1.4717 1.4682 16.0086 144.9445 0.00036623 -84.8131 0.21194
5.316 0.98809 5.4898e-005 3.8183 0.011973 6.948e-005 0.0011614 0.23193 0.0006593 0.23258 0.21457 0 0.032348 0.0389 0 1.2971 0.43567 0.13192 0.016399 9.3728 0.10219 0.00012953 0.78794 0.0079634 0.0088601 0.0015927 0.9842 0.98977 3.4637e-006 1.3855e-005 0.15364 0.69353 0.78367 0.0015027 0.80291 0.41945 0.0020203 0.42072 1.4736 1.4701 16.0087 144.9445 0.00036527 -84.8194 0.21294
5.317 0.98809 5.4898e-005 3.8183 0.011973 6.9493e-005 0.0011614 0.23193 0.0006593 0.23258 0.21458 0 0.032347 0.0389 0 1.2972 0.43572 0.13193 0.0164 9.3748 0.1022 0.00012955 0.78793 0.007964 0.0088608 0.001591 0.98423 0.9898 3.4599e-006 1.384e-005 0.15365 0.69443 0.78435 0.0015018 0.80407 0.41964 0.0020192 0.42072 1.4754 1.4719 16.0087 144.9445 0.00036431 -84.8256 0.21394
5.318 0.98809 5.4898e-005 3.8183 0.011973 6.9506e-005 0.0011614 0.23193 0.0006593 0.23259 0.21458 0 0.032347 0.0389 0 1.2973 0.43576 0.13195 0.016402 9.3768 0.10221 0.00012956 0.78792 0.0079646 0.0088614 0.0015894 0.98425 0.98982 3.4561e-006 1.3825e-005 0.15365 0.69533 0.78502 0.001501 0.80522 0.41984 0.0020182 0.42073 1.4772 1.4738 16.0088 144.9445 0.00036336 -84.8317 0.21494
5.319 0.98809 5.4898e-005 3.8183 0.011973 6.9519e-005 0.0011614 0.23193 0.0006593 0.23259 0.21458 0 0.032347 0.0389 0 1.2974 0.43581 0.13196 0.016403 9.3788 0.10222 0.00012957 0.78791 0.0079652 0.008862 0.0015878 0.98427 0.98984 3.4524e-006 1.381e-005 0.15366 0.69622 0.78569 0.0015002 0.80637 0.42004 0.0020171 0.42074 1.4791 1.4756 16.0088 144.9445 0.00036241 -84.8378 0.21594
5.32 0.98809 5.4898e-005 3.8183 0.011973 6.9532e-005 0.0011614 0.23194 0.0006593 0.23259 0.21458 0 0.032347 0.0389 0 1.2975 0.43586 0.13198 0.016405 9.3808 0.10223 0.00012959 0.7879 0.0079658 0.0088627 0.0015862 0.98429 0.98986 3.4487e-006 1.3795e-005 0.15366 0.69712 0.78635 0.0014994 0.80751 0.42023 0.0020161 0.42075 1.4809 1.4774 16.0089 144.9445 0.00036146 -84.8438 0.21694
5.321 0.98809 5.4898e-005 3.8183 0.011973 6.9545e-005 0.0011614 0.23194 0.0006593 0.23259 0.21458 0 0.032347 0.0389 0 1.2976 0.4359 0.13199 0.016406 9.3829 0.10224 0.0001296 0.78789 0.0079664 0.0088633 0.0015846 0.98431 0.98988 3.445e-006 1.3781e-005 0.15367 0.69801 0.78701 0.0014987 0.80864 0.42043 0.002015 0.42075 1.4827 1.4793 16.0089 144.9445 0.00036052 -84.8498 0.21794
5.322 0.98809 5.4898e-005 3.8183 0.011973 6.9558e-005 0.0011614 0.23194 0.0006593 0.23259 0.21459 0 0.032347 0.0389 0 1.2977 0.43595 0.13201 0.016408 9.3849 0.10225 0.00012961 0.78788 0.007967 0.008864 0.001583 0.98433 0.98989 3.4414e-006 1.3766e-005 0.15367 0.6989 0.78767 0.0014979 0.80977 0.42063 0.002014 0.42076 1.4845 1.4811 16.0089 144.9446 0.00035959 -84.8558 0.21894
5.323 0.98809 5.4898e-005 3.8183 0.011973 6.9571e-005 0.0011614 0.23194 0.0006593 0.2326 0.21459 0 0.032347 0.0389 0 1.2978 0.436 0.13202 0.016409 9.3869 0.10226 0.00012962 0.78787 0.0079676 0.0088646 0.0015815 0.98436 0.98991 3.4378e-006 1.3752e-005 0.15368 0.69978 0.78832 0.0014971 0.81089 0.42082 0.002013 0.42077 1.4864 1.4829 16.009 144.9446 0.00035866 -84.8617 0.21994
5.324 0.98809 5.4898e-005 3.8183 0.011973 6.9584e-005 0.0011614 0.23194 0.0006593 0.2326 0.21459 0 0.032347 0.0389 0 1.2979 0.43604 0.13204 0.016411 9.3889 0.10227 0.00012964 0.78786 0.0079682 0.0088653 0.0015799 0.98438 0.98993 3.4343e-006 1.3737e-005 0.15368 0.70066 0.78897 0.0014963 0.81201 0.42102 0.002012 0.42078 1.4882 1.4847 16.009 144.9446 0.00035774 -84.8676 0.22094
5.325 0.98809 5.4898e-005 3.8183 0.011973 6.9597e-005 0.0011614 0.23195 0.0006593 0.2326 0.21459 0 0.032347 0.0389 0 1.298 0.43609 0.13205 0.016412 9.3909 0.10228 0.00012965 0.78785 0.0079688 0.0088659 0.0015784 0.9844 0.98995 3.4307e-006 1.3723e-005 0.15369 0.70154 0.78961 0.0014956 0.81312 0.42122 0.002011 0.42078 1.49 1.4866 16.0091 144.9446 0.00035682 -84.8734 0.22194
5.326 0.98809 5.4898e-005 3.8183 0.011973 6.9609e-005 0.0011614 0.23195 0.0006593 0.2326 0.21459 0 0.032347 0.0389 0 1.2981 0.43614 0.13207 0.016413 9.393 0.10228 0.00012966 0.78785 0.0079694 0.0088666 0.0015769 0.98442 0.98997 3.4272e-006 1.3709e-005 0.15369 0.70242 0.79025 0.0014948 0.81422 0.42141 0.00201 0.42079 1.4918 1.4884 16.0091 144.9446 0.0003559 -84.8792 0.22294
5.327 0.98809 5.4897e-005 3.8183 0.011973 6.9622e-005 0.0011614 0.23195 0.0006593 0.2326 0.2146 0 0.032346 0.0389 0 1.2982 0.43618 0.13209 0.016415 9.395 0.10229 0.00012968 0.78784 0.00797 0.0088672 0.0015754 0.98444 0.98998 3.4237e-006 1.3695e-005 0.1537 0.70329 0.79089 0.0014941 0.81532 0.42161 0.002009 0.4208 1.4936 1.4902 16.0091 144.9446 0.00035499 -84.8849 0.22394
5.328 0.98809 5.4897e-005 3.8183 0.011973 6.9635e-005 0.0011614 0.23195 0.0006593 0.23261 0.2146 0 0.032346 0.0389 0 1.2983 0.43623 0.1321 0.016416 9.397 0.1023 0.00012969 0.78783 0.0079706 0.0088678 0.0015739 0.98446 0.99 3.4203e-006 1.3682e-005 0.1537 0.70416 0.79152 0.0014933 0.81641 0.42181 0.0020081 0.42081 1.4954 1.492 16.0092 144.9446 0.00035408 -84.8906 0.22494
5.329 0.98809 5.4897e-005 3.8183 0.011973 6.9648e-005 0.0011614 0.23195 0.0006593 0.23261 0.2146 0 0.032346 0.0389 0 1.2984 0.43628 0.13212 0.016418 9.399 0.10231 0.0001297 0.78782 0.0079712 0.0088685 0.0015724 0.98448 0.99002 3.4169e-006 1.3668e-005 0.15371 0.70503 0.79215 0.0014926 0.8175 0.422 0.0020071 0.42081 1.4971 1.4938 16.0092 144.9447 0.00035318 -84.8962 0.22594
5.33 0.98809 5.4897e-005 3.8183 0.011973 6.9661e-005 0.0011614 0.23196 0.0006593 0.23261 0.2146 0 0.032346 0.0389 0 1.2985 0.43632 0.13213 0.016419 9.401 0.10232 0.00012971 0.78781 0.0079718 0.0088691 0.001571 0.9845 0.99003 3.4135e-006 1.3654e-005 0.15371 0.7059 0.79277 0.0014919 0.81858 0.4222 0.0020062 0.42082 1.4989 1.4956 16.0093 144.9447 0.00035228 -84.9018 0.22694
5.331 0.98809 5.4897e-005 3.8183 0.011973 6.9674e-005 0.0011614 0.23196 0.0006593 0.23261 0.2146 0 0.032346 0.0389 0 1.2985 0.43637 0.13215 0.016421 9.4031 0.10233 0.00012973 0.7878 0.0079724 0.0088698 0.0015695 0.98452 0.99005 3.4102e-006 1.3641e-005 0.15371 0.70676 0.7934 0.0014911 0.81965 0.4224 0.0020052 0.42083 1.5007 1.4974 16.0093 144.9447 0.00035139 -84.9074 0.22794
5.332 0.98809 5.4897e-005 3.8183 0.011973 6.9687e-005 0.0011614 0.23196 0.0006593 0.23262 0.21461 0 0.032346 0.0389 0 1.2986 0.43642 0.13216 0.016422 9.4051 0.10234 0.00012974 0.78779 0.007973 0.0088704 0.0015681 0.98454 0.99007 3.4068e-006 1.3628e-005 0.15372 0.70762 0.79401 0.0014904 0.82072 0.42259 0.0020043 0.42084 1.5025 1.4992 16.0093 144.9447 0.0003505 -84.9129 0.22894
5.333 0.98809 5.4897e-005 3.8183 0.011973 6.97e-005 0.0011615 0.23196 0.0006593 0.23262 0.21461 0 0.032346 0.0389 0 1.2987 0.43646 0.13218 0.016424 9.4071 0.10235 0.00012975 0.78778 0.0079736 0.008871 0.0015666 0.98456 0.99008 3.4035e-006 1.3614e-005 0.15372 0.70848 0.79463 0.0014897 0.82178 0.42279 0.0020033 0.42085 1.5043 1.5009 16.0094 144.9447 0.00034961 -84.9183 0.22994
5.334 0.98809 5.4897e-005 3.8183 0.011973 6.9713e-005 0.0011615 0.23196 0.0006593 0.23262 0.21461 0 0.032346 0.0389 0 1.2988 0.43651 0.13219 0.016425 9.4091 0.10236 0.00012977 0.78777 0.0079742 0.0088717 0.0015652 0.98458 0.9901 3.4003e-006 1.3601e-005 0.15373 0.70934 0.79524 0.001489 0.82284 0.42298 0.0020024 0.42085 1.506 1.5027 16.0094 144.9447 0.00034873 -84.9238 0.23094
5.335 0.98809 5.4897e-005 3.8183 0.011973 6.9726e-005 0.0011615 0.23197 0.0006593 0.23262 0.21461 0 0.032346 0.0389 0 1.2989 0.43656 0.13221 0.016427 9.4112 0.10237 0.00012978 0.78776 0.0079748 0.0088723 0.0015638 0.9846 0.99011 3.397e-006 1.3588e-005 0.15373 0.71019 0.79585 0.0014883 0.82389 0.42318 0.0020015 0.42086 1.5078 1.5045 16.0095 144.9447 0.00034786 -84.9292 0.23194
5.336 0.98809 5.4897e-005 3.8183 0.011973 6.9739e-005 0.0011615 0.23197 0.0006593 0.23262 0.21461 0 0.032345 0.0389 0 1.299 0.4366 0.13222 0.016428 9.4132 0.10237 0.00012979 0.78776 0.0079754 0.008873 0.0015624 0.98461 0.99013 3.3938e-006 1.3575e-005 0.15374 0.71104 0.79645 0.0014876 0.82494 0.42338 0.0020006 0.42087 1.5095 1.5063 16.0095 144.9448 0.00034698 -84.9345 0.23294
5.337 0.98809 5.4897e-005 3.8183 0.011973 6.9752e-005 0.0011615 0.23197 0.0006593 0.23263 0.21462 0 0.032345 0.0389 0 1.2991 0.43665 0.13224 0.01643 9.4152 0.10238 0.0001298 0.78775 0.0079759 0.0088736 0.001561 0.98463 0.99014 3.3906e-006 1.3563e-005 0.15374 0.71189 0.79705 0.0014869 0.82598 0.42357 0.0019997 0.42088 1.5113 1.508 16.0095 144.9448 0.00034612 -84.9398 0.23394
5.338 0.98809 5.4897e-005 3.8183 0.011973 6.9765e-005 0.0011615 0.23197 0.0006593 0.23263 0.21462 0 0.032345 0.0389 0 1.2992 0.43669 0.13225 0.016431 9.4172 0.10239 0.00012982 0.78774 0.0079765 0.0088743 0.0015596 0.98465 0.99015 3.3875e-006 1.355e-005 0.15375 0.71273 0.79765 0.0014862 0.82701 0.42377 0.0019988 0.42089 1.513 1.5098 16.0096 144.9448 0.00034525 -84.9451 0.23494
5.339 0.98809 5.4897e-005 3.8183 0.011973 6.9778e-005 0.0011615 0.23197 0.0006593 0.23263 0.21462 0 0.032345 0.0389 0 1.2993 0.43674 0.13227 0.016433 9.4193 0.1024 0.00012983 0.78773 0.0079771 0.0088749 0.0015583 0.98467 0.99017 3.3843e-006 1.3538e-005 0.15375 0.71357 0.79824 0.0014855 0.82804 0.42397 0.0019979 0.42089 1.5148 1.5115 16.0096 144.9448 0.00034439 -84.9503 0.23594
5.34 0.98809 5.4896e-005 3.8183 0.011973 6.9791e-005 0.0011615 0.23198 0.0006593 0.23263 0.21462 0 0.032345 0.0389 0 1.2994 0.43679 0.13229 0.016434 9.4213 0.10241 0.00012984 0.78772 0.0079777 0.0088755 0.001557 0.98469 0.99018 3.3812e-006 1.3525e-005 0.15376 0.71441 0.79883 0.0014849 0.82906 0.42416 0.001997 0.4209 1.5165 1.5133 16.0096 144.9448 0.00034354 -84.9555 0.23694
5.341 0.98809 5.4896e-005 3.8183 0.011973 6.9804e-005 0.0011615 0.23198 0.0006593 0.23263 0.21462 0 0.032345 0.0389 0 1.2995 0.43683 0.1323 0.016435 9.4233 0.10242 0.00012986 0.78771 0.0079783 0.0088762 0.0015556 0.98471 0.9902 3.3781e-006 1.3513e-005 0.15376 0.71525 0.79942 0.0014842 0.83008 0.42436 0.0019961 0.42091 1.5183 1.515 16.0097 144.9448 0.00034269 -84.9607 0.23794
5.342 0.98809 5.4896e-005 3.8183 0.011973 6.9817e-005 0.0011615 0.23198 0.0006593 0.23264 0.21463 0 0.032345 0.0389 0 1.2996 0.43688 0.13232 0.016437 9.4253 0.10243 0.00012987 0.7877 0.0079789 0.0088768 0.0015543 0.98472 0.99021 3.3751e-006 1.3501e-005 0.15377 0.71608 0.8 0.0014835 0.83109 0.42455 0.0019953 0.42092 1.52 1.5168 16.0097 144.9448 0.00034184 -84.9658 0.23894
5.343 0.98809 5.4896e-005 3.8183 0.011973 6.983e-005 0.0011615 0.23198 0.0006593 0.23264 0.21463 0 0.032345 0.0389 0 1.2997 0.43693 0.13233 0.016438 9.4274 0.10244 0.00012988 0.78769 0.0079795 0.0088775 0.001553 0.98474 0.99022 3.3721e-006 1.3489e-005 0.15377 0.71692 0.80058 0.0014829 0.8321 0.42475 0.0019944 0.42093 1.5217 1.5185 16.0097 144.9449 0.000341 -84.9708 0.23994
5.344 0.98809 5.4896e-005 3.8183 0.011973 6.9843e-005 0.0011615 0.23199 0.0006593 0.23264 0.21463 0 0.032345 0.0389 0 1.2998 0.43697 0.13235 0.01644 9.4294 0.10245 0.0001299 0.78768 0.0079801 0.0088781 0.0015517 0.98476 0.99024 3.3691e-006 1.3476e-005 0.15378 0.71775 0.80115 0.0014822 0.8331 0.42495 0.0019936 0.42094 1.5234 1.5202 16.0098 144.9449 0.00034016 -84.9759 0.24094
5.345 0.98809 5.4896e-005 3.8183 0.011973 6.9856e-005 0.0011615 0.23199 0.0006593 0.23264 0.21463 0 0.032345 0.0389 0 1.2999 0.43702 0.13236 0.016441 9.4314 0.10246 0.00012991 0.78767 0.0079807 0.0088787 0.0015504 0.98478 0.99025 3.3661e-006 1.3465e-005 0.15378 0.71857 0.80173 0.0014816 0.83409 0.42514 0.0019927 0.42095 1.5252 1.522 16.0098 144.9449 0.00033933 -84.9809 0.24194
5.346 0.98809 5.4896e-005 3.8183 0.011973 6.9868e-005 0.0011615 0.23199 0.0006593 0.23264 0.21463 0 0.032344 0.0389 0 1.3 0.43707 0.13238 0.016443 9.4334 0.10246 0.00012992 0.78767 0.0079813 0.0088794 0.0015491 0.98479 0.99026 3.3631e-006 1.3453e-005 0.15379 0.7194 0.8023 0.0014809 0.83508 0.42534 0.0019919 0.42095 1.5269 1.5237 16.0099 144.9449 0.0003385 -84.9858 0.24294
5.347 0.98809 5.4896e-005 3.8183 0.011973 6.9881e-005 0.0011615 0.23199 0.0006593 0.23265 0.21464 0 0.032344 0.0389 0 1.3001 0.43711 0.13239 0.016444 9.4355 0.10247 0.00012993 0.78766 0.0079819 0.00888 0.0015478 0.98481 0.99027 3.3602e-006 1.3441e-005 0.15379 0.72022 0.80286 0.0014803 0.83607 0.42553 0.001991 0.42096 1.5286 1.5254 16.0099 144.9449 0.00033767 -84.9907 0.24394
5.348 0.98809 5.4896e-005 3.8183 0.011973 6.9894e-005 0.0011615 0.23199 0.0006593 0.23265 0.21464 0 0.032344 0.0389 0 1.3002 0.43716 0.13241 0.016446 9.4375 0.10248 0.00012995 0.78765 0.0079825 0.0088807 0.0015466 0.98483 0.99029 3.3573e-006 1.3429e-005 0.15379 0.72104 0.80343 0.0014797 0.83704 0.42573 0.0019902 0.42097 1.5303 1.5271 16.0099 144.9449 0.00033685 -84.9956 0.24494
5.349 0.98809 5.4896e-005 3.8183 0.011973 6.9907e-005 0.0011615 0.232 0.0006593 0.23265 0.21464 0 0.032344 0.0389 0 1.3003 0.43721 0.13242 0.016447 9.4395 0.10249 0.00012996 0.78764 0.0079831 0.0088813 0.0015453 0.98485 0.9903 3.3544e-006 1.3418e-005 0.1538 0.72185 0.80399 0.001479 0.83802 0.42593 0.0019894 0.42098 1.532 1.5289 16.01 144.945 0.00033603 -85.0005 0.24594
5.35 0.98809 5.4896e-005 3.8183 0.011973 6.992e-005 0.0011615 0.232 0.0006593 0.23265 0.21464 0 0.032344 0.0389 0 1.3004 0.43725 0.13244 0.016449 9.4416 0.1025 0.00012997 0.78763 0.0079837 0.008882 0.0015441 0.98486 0.99031 3.3516e-006 1.3407e-005 0.1538 0.72267 0.80454 0.0014784 0.83898 0.42612 0.0019886 0.42099 1.5337 1.5306 16.01 144.945 0.00033521 -85.0053 0.24694
5.351 0.98809 5.4896e-005 3.8183 0.011973 6.9933e-005 0.0011615 0.232 0.0006593 0.23265 0.21464 0 0.032344 0.0389 0 1.3005 0.4373 0.13245 0.01645 9.4436 0.10251 0.00012999 0.78762 0.0079843 0.0088826 0.0015429 0.98488 0.99032 3.3487e-006 1.3395e-005 0.15381 0.72348 0.8051 0.0014778 0.83995 0.42632 0.0019878 0.421 1.5354 1.5323 16.01 144.945 0.0003344 -85.01 0.24794
5.352 0.98809 5.4896e-005 3.8183 0.011973 6.9946e-005 0.0011615 0.232 0.0006593 0.23266 0.21465 0 0.032344 0.0389 0 1.3005 0.43735 0.13247 0.016452 9.4456 0.10252 0.00013 0.78761 0.0079849 0.0088832 0.0015416 0.9849 0.99034 3.3459e-006 1.3384e-005 0.15381 0.72429 0.80565 0.0014772 0.8409 0.42651 0.001987 0.42101 1.5371 1.534 16.0101 144.945 0.0003336 -85.0148 0.24894
5.353 0.98809 5.4896e-005 3.8183 0.011973 6.9959e-005 0.0011615 0.232 0.0006593 0.23266 0.21465 0 0.032344 0.0389 0 1.3006 0.43739 0.13249 0.016453 9.4477 0.10253 0.00013001 0.7876 0.0079855 0.0088839 0.0015404 0.98491 0.99035 3.3431e-006 1.3373e-005 0.15382 0.72509 0.8062 0.0014766 0.84185 0.42671 0.0019862 0.42102 1.5387 1.5357 16.0101 144.945 0.0003328 -85.0195 0.24994
5.354 0.98809 5.4895e-005 3.8183 0.011973 6.9972e-005 0.0011615 0.23201 0.0006593 0.23266 0.21465 0 0.032344 0.0389 0 1.3007 0.43744 0.1325 0.016455 9.4497 0.10254 0.00013002 0.78759 0.0079861 0.0088845 0.0015393 0.98493 0.99036 3.3404e-006 1.3362e-005 0.15382 0.7259 0.80674 0.001476 0.8428 0.4269 0.0019854 0.42103 1.5404 1.5374 16.0101 144.945 0.000332 -85.0242 0.25094
5.355 0.98809 5.4895e-005 3.8183 0.011972 6.9985e-005 0.0011615 0.23201 0.0006593 0.23266 0.21465 0 0.032344 0.0389 0 1.3008 0.43748 0.13252 0.016456 9.4517 0.10254 0.00013004 0.78759 0.0079866 0.0088852 0.0015381 0.98494 0.99037 3.3377e-006 1.3351e-005 0.15383 0.7267 0.80728 0.0014754 0.84374 0.4271 0.0019846 0.42103 1.5421 1.539 16.0102 144.945 0.0003312 -85.0288 0.25194
5.356 0.98809 5.4895e-005 3.8183 0.011972 6.9998e-005 0.0011615 0.23201 0.0006593 0.23266 0.21465 0 0.032343 0.0389 0 1.3009 0.43753 0.13253 0.016457 9.4537 0.10255 0.00013005 0.78758 0.0079872 0.0088858 0.0015369 0.98496 0.99038 3.3349e-006 1.334e-005 0.15383 0.7275 0.80782 0.0014748 0.84468 0.42729 0.0019838 0.42104 1.5438 1.5407 16.0102 144.9451 0.00033041 -85.0334 0.25294
5.357 0.98809 5.4895e-005 3.8183 0.011972 7.0011e-005 0.0011615 0.23201 0.0006593 0.23267 0.21465 0 0.032343 0.0389 0 1.301 0.43758 0.13255 0.016459 9.4558 0.10256 0.00013006 0.78757 0.0079878 0.0088864 0.0015357 0.98498 0.99039 3.3323e-006 1.3329e-005 0.15384 0.7283 0.80836 0.0014742 0.84561 0.42749 0.0019831 0.42105 1.5454 1.5424 16.0102 144.9451 0.00032962 -85.0379 0.25394
5.358 0.98809 5.4895e-005 3.8183 0.011972 7.0024e-005 0.0011615 0.23201 0.0006593 0.23267 0.21466 0 0.032343 0.0389 0 1.3011 0.43762 0.13256 0.01646 9.4578 0.10257 0.00013008 0.78756 0.0079884 0.0088871 0.0015346 0.98499 0.9904 3.3296e-006 1.3319e-005 0.15384 0.72909 0.80889 0.0014736 0.84653 0.42769 0.0019823 0.42106 1.5471 1.5441 16.0102 144.9451 0.00032884 -85.0425 0.25494
5.359 0.98809 5.4895e-005 3.8183 0.011972 7.0037e-005 0.0011615 0.23202 0.0006593 0.23267 0.21466 0 0.032343 0.0389 0 1.3012 0.43767 0.13258 0.016462 9.4598 0.10258 0.00013009 0.78755 0.007989 0.0088877 0.0015334 0.98501 0.99041 3.3269e-006 1.3308e-005 0.15385 0.72988 0.80942 0.001473 0.84745 0.42788 0.0019815 0.42107 1.5488 1.5457 16.0103 144.9451 0.00032806 -85.047 0.25594
5.36 0.98809 5.4895e-005 3.8183 0.011972 7.005e-005 0.0011615 0.23202 0.0006593 0.23267 0.21466 0 0.032343 0.0389 0 1.3013 0.43772 0.13259 0.016463 9.4619 0.10259 0.0001301 0.78754 0.0079896 0.0088884 0.0015323 0.98502 0.99043 3.3243e-006 1.3297e-005 0.15385 0.73067 0.80995 0.0014725 0.84837 0.42808 0.0019808 0.42108 1.5504 1.5474 16.0103 144.9451 0.00032728 -85.0514 0.25694
5.361 0.98809 5.4895e-005 3.8183 0.011972 7.0063e-005 0.0011615 0.23202 0.0006593 0.23267 0.21466 0 0.032343 0.0389 0 1.3014 0.43776 0.13261 0.016465 9.4639 0.1026 0.00013011 0.78753 0.0079902 0.008889 0.0015312 0.98504 0.99044 3.3217e-006 1.3287e-005 0.15386 0.73146 0.81047 0.0014719 0.84928 0.42827 0.00198 0.42109 1.5521 1.5491 16.0103 144.9451 0.00032651 -85.0558 0.25794
5.362 0.98809 5.4895e-005 3.8183 0.011972 7.0076e-005 0.0011615 0.23202 0.0006593 0.23268 0.21466 0 0.032343 0.0389 0 1.3015 0.43781 0.13262 0.016466 9.4659 0.10261 0.00013013 0.78752 0.0079908 0.0088896 0.00153 0.98505 0.99045 3.3191e-006 1.3277e-005 0.15386 0.73224 0.81099 0.0014713 0.85018 0.42847 0.0019793 0.4211 1.5537 1.5507 16.0104 144.9452 0.00032574 -85.0602 0.25894
5.363 0.98809 5.4895e-005 3.8183 0.011972 7.0089e-005 0.0011615 0.23202 0.0006593 0.23268 0.21467 0 0.032343 0.0389 0 1.3016 0.43786 0.13264 0.016468 9.468 0.10262 0.00013014 0.78751 0.0079914 0.0088903 0.0015289 0.98507 0.99046 3.3166e-006 1.3266e-005 0.15386 0.73302 0.81151 0.0014708 0.85108 0.42866 0.0019786 0.42111 1.5554 1.5524 16.0104 144.9452 0.00032498 -85.0646 0.25994
5.364 0.98809 5.4895e-005 3.8183 0.011972 7.0102e-005 0.0011615 0.23203 0.0006593 0.23268 0.21467 0 0.032343 0.0389 0 1.3017 0.4379 0.13265 0.016469 9.47 0.10263 0.00013015 0.7875 0.007992 0.0088909 0.0015278 0.98508 0.99047 3.314e-006 1.3256e-005 0.15387 0.7338 0.81202 0.0014702 0.85197 0.42886 0.0019778 0.42112 1.557 1.554 16.0104 144.9452 0.00032422 -85.0689 0.26094
5.365 0.98809 5.4895e-005 3.8183 0.011972 7.0114e-005 0.0011616 0.23203 0.0006593 0.23268 0.21467 0 0.032343 0.0389 0 1.3018 0.43795 0.13267 0.016471 9.472 0.10263 0.00013017 0.7875 0.0079926 0.0088916 0.0015267 0.9851 0.99048 3.3115e-006 1.3246e-005 0.15387 0.73458 0.81254 0.0014697 0.85286 0.42905 0.0019771 0.42113 1.5586 1.5557 16.0105 144.9452 0.00032346 -85.0732 0.26194
5.366 0.98809 5.4895e-005 3.8183 0.011972 7.0127e-005 0.0011616 0.23203 0.0006593 0.23268 0.21467 0 0.032342 0.0389 0 1.3019 0.438 0.13269 0.016472 9.4741 0.10264 0.00013018 0.78749 0.0079932 0.0088922 0.0015257 0.98511 0.99049 3.309e-006 1.3236e-005 0.15388 0.73536 0.81305 0.0014691 0.85375 0.42925 0.0019764 0.42114 1.5603 1.5573 16.0105 144.9452 0.00032271 -85.0775 0.26294
5.367 0.98809 5.4894e-005 3.8183 0.011972 7.014e-005 0.0011616 0.23203 0.0006593 0.23269 0.21467 0 0.032342 0.0389 0 1.302 0.43804 0.1327 0.016474 9.4761 0.10265 0.00013019 0.78748 0.0079938 0.0088928 0.0015246 0.98513 0.9905 3.3065e-006 1.3226e-005 0.15388 0.73613 0.81355 0.0014686 0.85462 0.42944 0.0019757 0.42115 1.5619 1.5589 16.0105 144.9452 0.00032195 -85.0817 0.26394
5.368 0.98809 5.4894e-005 3.8183 0.011972 7.0153e-005 0.0011616 0.23203 0.0006593 0.23269 0.21468 0 0.032342 0.0389 0 1.3021 0.43809 0.13272 0.016475 9.4782 0.10266 0.0001302 0.78747 0.0079944 0.0088935 0.0015235 0.98514 0.99051 3.3041e-006 1.3217e-005 0.15389 0.7369 0.81406 0.001468 0.8555 0.42964 0.001975 0.42116 1.5635 1.5606 16.0105 144.9452 0.00032121 -85.0859 0.26494
5.369 0.98809 5.4894e-005 3.8183 0.011972 7.0166e-005 0.0011616 0.23204 0.0006593 0.23269 0.21468 0 0.032342 0.0389 0 1.3022 0.43814 0.13273 0.016476 9.4802 0.10267 0.00013022 0.78746 0.0079949 0.0088941 0.0015224 0.98515 0.99052 3.3016e-006 1.3207e-005 0.15389 0.73767 0.81456 0.0014675 0.85637 0.42983 0.0019743 0.42117 1.5651 1.5622 16.0106 144.9453 0.00032046 -85.0901 0.26594
5.37 0.98809 5.4894e-005 3.8183 0.011972 7.0179e-005 0.0011616 0.23204 0.0006593 0.23269 0.21468 0 0.032342 0.0389 0 1.3023 0.43818 0.13275 0.016478 9.4822 0.10268 0.00013023 0.78745 0.0079955 0.0088947 0.0015214 0.98517 0.99053 3.2992e-006 1.3197e-005 0.1539 0.73843 0.81506 0.0014669 0.85723 0.43003 0.0019736 0.42118 1.5667 1.5638 16.0106 144.9453 0.00031972 -85.0942 0.26694
5.371 0.98809 5.4894e-005 3.8183 0.011972 7.0192e-005 0.0011616 0.23204 0.0006593 0.23269 0.21468 0 0.032342 0.0389 0 1.3024 0.43823 0.13276 0.016479 9.4843 0.10269 0.00013024 0.78744 0.0079961 0.0088954 0.0015203 0.98518 0.99054 3.2968e-006 1.3188e-005 0.1539 0.73919 0.81555 0.0014664 0.85809 0.43022 0.0019729 0.42119 1.5683 1.5654 16.0106 144.9453 0.00031899 -85.0983 0.26794
5.372 0.98809 5.4894e-005 3.8183 0.011972 7.0205e-005 0.0011616 0.23204 0.0006593 0.2327 0.21468 0 0.032342 0.0389 0 1.3025 0.43828 0.13278 0.016481 9.4863 0.1027 0.00013026 0.78743 0.0079967 0.008896 0.0015193 0.9852 0.99055 3.2945e-006 1.3178e-005 0.15391 0.73995 0.81605 0.0014659 0.85894 0.43042 0.0019722 0.4212 1.57 1.5671 16.0107 144.9453 0.00031826 -85.1024 0.26894
5.373 0.98809 5.4894e-005 3.8183 0.011972 7.0218e-005 0.0011616 0.23204 0.0006593 0.2327 0.21469 0 0.032342 0.0389 0 1.3025 0.43832 0.13279 0.016482 9.4883 0.10271 0.00013027 0.78742 0.0079973 0.0088967 0.0015183 0.98521 0.99056 3.2921e-006 1.3169e-005 0.15391 0.74071 0.81654 0.0014654 0.85979 0.43061 0.0019715 0.42121 1.5716 1.5687 16.0107 144.9453 0.00031753 -85.1064 0.26994
5.374 0.98809 5.4894e-005 3.8183 0.011972 7.0231e-005 0.0011616 0.23205 0.0006593 0.2327 0.21469 0 0.032342 0.0389 0 1.3026 0.43837 0.13281 0.016484 9.4904 0.10272 0.00013028 0.78742 0.0079979 0.0088973 0.0015172 0.98522 0.99056 3.2898e-006 1.3159e-005 0.15392 0.74147 0.81703 0.0014649 0.86064 0.43081 0.0019709 0.42122 1.5731 1.5703 16.0107 144.9453 0.0003168 -85.1105 0.27094
5.375 0.98809 5.4894e-005 3.8183 0.011972 7.0244e-005 0.0011616 0.23205 0.0006593 0.2327 0.21469 0 0.032342 0.0389 0 1.3027 0.43841 0.13282 0.016485 9.4924 0.10272 0.00013029 0.78741 0.0079985 0.0088979 0.0015162 0.98524 0.99057 3.2874e-006 1.315e-005 0.15392 0.74222 0.81751 0.0014643 0.86148 0.431 0.0019702 0.42123 1.5747 1.5719 16.0107 144.9454 0.00031608 -85.1144 0.27194
5.376 0.98809 5.4894e-005 3.8183 0.011972 7.0257e-005 0.0011616 0.23205 0.0006593 0.2327 0.21469 0 0.032341 0.0389 0 1.3028 0.43846 0.13284 0.016487 9.4945 0.10273 0.00013031 0.7874 0.0079991 0.0088986 0.0015153 0.98525 0.99058 3.2851e-006 1.3141e-005 0.15393 0.74297 0.818 0.0014638 0.86231 0.4312 0.0019695 0.42124 1.5763 1.5735 16.0108 144.9454 0.00031536 -85.1184 0.27294
5.377 0.98809 5.4894e-005 3.8183 0.011972 7.027e-005 0.0011616 0.23205 0.0006593 0.23271 0.21469 0 0.032341 0.0389 0 1.3029 0.43851 0.13285 0.016488 9.4965 0.10274 0.00013032 0.78739 0.0079997 0.0088992 0.0015143 0.98526 0.99059 3.2829e-006 1.3132e-005 0.15393 0.74372 0.81848 0.0014633 0.86314 0.43139 0.0019689 0.42125 1.5779 1.5751 16.0108 144.9454 0.00031464 -85.1223 0.27394
5.378 0.98809 5.4894e-005 3.8183 0.011972 7.0283e-005 0.0011616 0.23205 0.0006593 0.23271 0.2147 0 0.032341 0.0389 0 1.303 0.43855 0.13287 0.01649 9.4985 0.10275 0.00013033 0.78738 0.0080003 0.0088999 0.0015133 0.98528 0.9906 3.2806e-006 1.3123e-005 0.15394 0.74447 0.81895 0.0014628 0.86397 0.43159 0.0019682 0.42126 1.5795 1.5767 16.0108 144.9454 0.00031393 -85.1262 0.27494
5.379 0.98809 5.4894e-005 3.8183 0.011972 7.0296e-005 0.0011616 0.23206 0.0006593 0.23271 0.2147 0 0.032341 0.0389 0 1.3031 0.4386 0.13289 0.016491 9.5006 0.10276 0.00013034 0.78737 0.0080009 0.0089005 0.0015123 0.98529 0.99061 3.2784e-006 1.3114e-005 0.15394 0.74521 0.81943 0.0014624 0.86479 0.43178 0.0019676 0.42127 1.5811 1.5782 16.0108 144.9454 0.00031322 -85.1301 0.27594
5.38 0.98809 5.4893e-005 3.8183 0.011972 7.0309e-005 0.0011616 0.23206 0.0006593 0.23271 0.2147 0 0.032341 0.0389 0 1.3032 0.43865 0.1329 0.016493 9.5026 0.10277 0.00013036 0.78736 0.0080015 0.0089011 0.0015114 0.9853 0.99062 3.2761e-006 1.3105e-005 0.15394 0.74595 0.8199 0.0014619 0.8656 0.43198 0.0019669 0.42128 1.5826 1.5798 16.0109 144.9454 0.00031252 -85.1339 0.27694
5.381 0.98809 5.4893e-005 3.8183 0.011972 7.0322e-005 0.0011616 0.23206 0.0006593 0.23271 0.2147 0 0.032341 0.0389 0 1.3033 0.43869 0.13292 0.016494 9.5047 0.10278 0.00013037 0.78735 0.0080021 0.0089018 0.0015104 0.98532 0.99063 3.2739e-006 1.3096e-005 0.15395 0.74669 0.82037 0.0014614 0.86641 0.43217 0.0019663 0.42129 1.5842 1.5814 16.0109 144.9455 0.00031182 -85.1377 0.27794
5.382 0.98809 5.4893e-005 3.8183 0.011972 7.0335e-005 0.0011616 0.23206 0.0006593 0.23272 0.2147 0 0.032341 0.0389 0 1.3034 0.43874 0.13293 0.016495 9.5067 0.10279 0.00013038 0.78734 0.0080026 0.0089024 0.0015095 0.98533 0.99064 3.2717e-006 1.3087e-005 0.15395 0.74743 0.82084 0.0014609 0.86722 0.43236 0.0019657 0.4213 1.5858 1.583 16.0109 144.9455 0.00031112 -85.1415 0.27894
5.383 0.98809 5.4893e-005 3.8183 0.011972 7.0348e-005 0.0011616 0.23206 0.0006593 0.23272 0.2147 0 0.032341 0.0389 0 1.3035 0.43879 0.13295 0.016497 9.5087 0.1028 0.0001304 0.78733 0.0080032 0.008903 0.0015085 0.98534 0.99064 3.2696e-006 1.3078e-005 0.15396 0.74817 0.82131 0.0014604 0.86802 0.43256 0.001965 0.42131 1.5873 1.5845 16.0109 144.9455 0.00031042 -85.1453 0.27994
5.384 0.98809 5.4893e-005 3.8183 0.011972 7.036e-005 0.0011616 0.23207 0.0006593 0.23272 0.21471 0 0.032341 0.0389 0 1.3036 0.43883 0.13296 0.016498 9.5108 0.1028 0.00013041 0.78733 0.0080038 0.0089037 0.0015076 0.98535 0.99065 3.2674e-006 1.307e-005 0.15396 0.7489 0.82177 0.0014599 0.86882 0.43275 0.0019644 0.42132 1.5889 1.5861 16.011 144.9455 0.00030973 -85.149 0.28094
5.385 0.98809 5.4893e-005 3.8183 0.011972 7.0373e-005 0.0011616 0.23207 0.0006593 0.23272 0.21471 0 0.032341 0.0389 0 1.3037 0.43888 0.13298 0.0165 9.5128 0.10281 0.00013042 0.78732 0.0080044 0.0089043 0.0015066 0.98537 0.99066 3.2653e-006 1.3061e-005 0.15397 0.74963 0.82223 0.0014595 0.86961 0.43295 0.0019638 0.42133 1.5904 1.5877 16.011 144.9455 0.00030904 -85.1527 0.28194
5.386 0.98809 5.4893e-005 3.8183 0.011972 7.0386e-005 0.0011616 0.23207 0.0006593 0.23272 0.21471 0 0.03234 0.0389 0 1.3038 0.43893 0.13299 0.016501 9.5149 0.10282 0.00013043 0.78731 0.008005 0.008905 0.0015057 0.98538 0.99067 3.2631e-006 1.3053e-005 0.15397 0.75036 0.82269 0.001459 0.8704 0.43314 0.0019632 0.42134 1.592 1.5892 16.011 144.9455 0.00030835 -85.1564 0.28294
5.387 0.98809 5.4893e-005 3.8183 0.011972 7.0399e-005 0.0011616 0.23207 0.0006593 0.23273 0.21471 0 0.03234 0.0389 0 1.3039 0.43897 0.13301 0.016503 9.5169 0.10283 0.00013045 0.7873 0.0080056 0.0089056 0.0015048 0.98539 0.99068 3.261e-006 1.3044e-005 0.15398 0.75108 0.82314 0.0014585 0.87118 0.43334 0.0019626 0.42135 1.5935 1.5908 16.011 144.9456 0.00030767 -85.16 0.28394
5.388 0.98809 5.4893e-005 3.8183 0.011972 7.0412e-005 0.0011616 0.23207 0.0006593 0.23273 0.21471 0 0.03234 0.0389 0 1.304 0.43902 0.13302 0.016504 9.5189 0.10284 0.00013046 0.78729 0.0080062 0.0089062 0.0015039 0.9854 0.99069 3.259e-006 1.3036e-005 0.15398 0.75181 0.8236 0.0014581 0.87196 0.43353 0.001962 0.42136 1.5951 1.5923 16.0111 144.9456 0.00030699 -85.1636 0.28494
5.389 0.98809 5.4893e-005 3.8183 0.011972 7.0425e-005 0.0011616 0.23208 0.0006593 0.23273 0.21472 0 0.03234 0.0389 0 1.3041 0.43907 0.13304 0.016506 9.521 0.10285 0.00013047 0.78728 0.0080068 0.0089069 0.001503 0.98541 0.99069 3.2569e-006 1.3028e-005 0.15399 0.75253 0.82405 0.0014576 0.87274 0.43373 0.0019614 0.42137 1.5966 1.5939 16.0111 144.9456 0.00030632 -85.1672 0.28594
5.39 0.98809 5.4893e-005 3.8183 0.011972 7.0438e-005 0.0011616 0.23208 0.0006593 0.23273 0.21472 0 0.03234 0.0389 0 1.3042 0.43911 0.13305 0.016507 9.523 0.10286 0.00013049 0.78727 0.0080074 0.0089075 0.0015021 0.98543 0.9907 3.2548e-006 1.3019e-005 0.15399 0.75325 0.8245 0.0014571 0.87351 0.43392 0.0019608 0.42138 1.5981 1.5954 16.0111 144.9456 0.00030564 -85.1708 0.28694
5.391 0.98809 5.4893e-005 3.8183 0.011972 7.0451e-005 0.0011616 0.23208 0.0006593 0.23273 0.21472 0 0.03234 0.0389 0 1.3043 0.43916 0.13307 0.016509 9.5251 0.10287 0.0001305 0.78726 0.008008 0.0089081 0.0015012 0.98544 0.99071 3.2528e-006 1.3011e-005 0.154 0.75397 0.82494 0.0014567 0.87427 0.43411 0.0019602 0.42139 1.5997 1.597 16.0111 144.9456 0.00030497 -85.1743 0.28794
5.392 0.98809 5.4893e-005 3.8183 0.011972 7.0464e-005 0.0011616 0.23208 0.0006593 0.23274 0.21472 0 0.03234 0.0389 0 1.3044 0.43921 0.13308 0.01651 9.5271 0.10288 0.00013051 0.78725 0.0080086 0.0089088 0.0015003 0.98545 0.99072 3.2508e-006 1.3003e-005 0.154 0.75468 0.82539 0.0014562 0.87503 0.43431 0.0019596 0.4214 1.6012 1.5985 16.0111 144.9456 0.00030431 -85.1778 0.28894
5.393 0.98809 5.4893e-005 3.8183 0.011972 7.0477e-005 0.0011616 0.23208 0.0006593 0.23274 0.21472 0 0.03234 0.0389 0 1.3044 0.43925 0.1331 0.016511 9.5292 0.10289 0.00013052 0.78725 0.0080091 0.0089094 0.0014995 0.98546 0.99073 3.2488e-006 1.2995e-005 0.15401 0.75539 0.82583 0.0014558 0.87579 0.4345 0.001959 0.42141 1.6027 1.6 16.0112 144.9457 0.00030364 -85.1813 0.28994
5.394 0.98809 5.4892e-005 3.8183 0.011972 7.049e-005 0.0011616 0.23209 0.0006593 0.23274 0.21472 0 0.03234 0.0389 0 1.3045 0.4393 0.13312 0.016513 9.5312 0.10289 0.00013054 0.78724 0.0080097 0.00891 0.0014986 0.98547 0.99073 3.2468e-006 1.2987e-005 0.15401 0.7561 0.82627 0.0014554 0.87654 0.4347 0.0019585 0.42143 1.6042 1.6015 16.0112 144.9457 0.00030298 -85.1848 0.29094
5.395 0.98809 5.4892e-005 3.8183 0.011972 7.0503e-005 0.0011616 0.23209 0.0006593 0.23274 0.21473 0 0.03234 0.0389 0 1.3046 0.43934 0.13313 0.016514 9.5333 0.1029 0.00013055 0.78723 0.0080103 0.0089107 0.0014978 0.98548 0.99074 3.2448e-006 1.2979e-005 0.15401 0.75681 0.82671 0.0014549 0.87729 0.43489 0.0019579 0.42144 1.6057 1.6031 16.0112 144.9457 0.00030232 -85.1882 0.29194
5.396 0.98809 5.4892e-005 3.8183 0.011972 7.0516e-005 0.0011617 0.23209 0.0006593 0.23274 0.21473 0 0.032339 0.0389 0 1.3047 0.43939 0.13315 0.016516 9.5353 0.10291 0.00013056 0.78722 0.0080109 0.0089113 0.0014969 0.9855 0.99075 3.2429e-006 1.2972e-005 0.15402 0.75752 0.82714 0.0014545 0.87803 0.43508 0.0019573 0.42145 1.6072 1.6046 16.0112 144.9457 0.00030167 -85.1916 0.29294
5.397 0.98809 5.4892e-005 3.8183 0.011972 7.0529e-005 0.0011617 0.23209 0.0006593 0.23275 0.21473 0 0.032339 0.0389 0 1.3048 0.43944 0.13316 0.016517 9.5373 0.10292 0.00013058 0.78721 0.0080115 0.008912 0.0014961 0.98551 0.99076 3.2409e-006 1.2964e-005 0.15402 0.75822 0.82758 0.0014541 0.87877 0.43528 0.0019568 0.42146 1.6087 1.6061 16.0113 144.9457 0.00030102 -85.195 0.29394
5.398 0.98809 5.4892e-005 3.8183 0.011972 7.0542e-005 0.0011617 0.23209 0.0006593 0.23275 0.21473 0 0.032339 0.0389 0 1.3049 0.43948 0.13318 0.016519 9.5394 0.10293 0.00013059 0.7872 0.0080121 0.0089126 0.0014952 0.98552 0.99076 3.239e-006 1.2956e-005 0.15403 0.75892 0.82801 0.0014536 0.87951 0.43547 0.0019562 0.42147 1.6102 1.6076 16.0113 144.9457 0.00030037 -85.1983 0.29494
5.399 0.98809 5.4892e-005 3.8183 0.011972 7.0555e-005 0.0011617 0.2321 0.0006593 0.23275 0.21473 0 0.032339 0.0389 0 1.305 0.43953 0.13319 0.01652 9.5414 0.10294 0.0001306 0.78719 0.0080127 0.0089132 0.0014944 0.98553 0.99077 3.2371e-006 1.2948e-005 0.15403 0.75962 0.82844 0.0014532 0.88024 0.43566 0.0019556 0.42148 1.6117 1.6091 16.0113 144.9458 0.00029972 -85.2017 0.29594
5.4 0.98809 5.4892e-005 3.8183 0.011972 7.0568e-005 0.0011617 0.2321 0.0006593 0.23275 0.21474 0 0.032339 0.0389 0 1.3051 0.43958 0.13321 0.016522 9.5435 0.10295 0.00013061 0.78718 0.0080133 0.0089139 0.0014935 0.98554 0.99078 3.2352e-006 1.2941e-005 0.15404 0.76032 0.82886 0.0014528 0.88096 0.43586 0.0019551 0.42149 1.6132 1.6106 16.0113 144.9458 0.00029908 -85.205 0.29694
5.401 0.98809 5.4892e-005 3.8183 0.011972 7.0581e-005 0.0011617 0.2321 0.0006593 0.23275 0.21474 0 0.032339 0.0389 0 1.3052 0.43962 0.13322 0.016523 9.5455 0.10296 0.00013063 0.78717 0.0080139 0.0089145 0.0014927 0.98555 0.99079 3.2333e-006 1.2933e-005 0.15404 0.76102 0.82929 0.0014524 0.88168 0.43605 0.0019545 0.4215 1.6147 1.6121 16.0113 144.9458 0.00029844 -85.2083 0.29794
5.402 0.98809 5.4892e-005 3.8183 0.011972 7.0594e-005 0.0011617 0.2321 0.0006593 0.23276 0.21474 0 0.032339 0.0389 0 1.3053 0.43967 0.13324 0.016525 9.5476 0.10297 0.00013064 0.78716 0.0080145 0.0089151 0.0014919 0.98556 0.99079 3.2314e-006 1.2926e-005 0.15405 0.76171 0.82971 0.001452 0.8824 0.43625 0.001954 0.42151 1.6162 1.6136 16.0114 144.9458 0.00029781 -85.2115 0.29894
5.403 0.98809 5.4892e-005 3.8183 0.011972 7.0606e-005 0.0011617 0.2321 0.0006593 0.23276 0.21474 0 0.032339 0.0389 0 1.3054 0.43972 0.13325 0.016526 9.5496 0.10297 0.00013065 0.78716 0.008015 0.0089158 0.0014911 0.98557 0.9908 3.2296e-006 1.2919e-005 0.15405 0.7624 0.83013 0.0014515 0.88311 0.43644 0.0019535 0.42152 1.6177 1.6151 16.0114 144.9458 0.00029717 -85.2147 0.29994
5.404 0.98809 5.4892e-005 3.8183 0.011972 7.0619e-005 0.0011617 0.2321 0.0006593 0.23276 0.21474 0 0.032339 0.0389 0 1.3055 0.43976 0.13327 0.016528 9.5517 0.10298 0.00013067 0.78715 0.0080156 0.0089164 0.0014903 0.98558 0.99081 3.2278e-006 1.2911e-005 0.15406 0.76309 0.83055 0.0014511 0.88382 0.43663 0.0019529 0.42153 1.6191 1.6166 16.0114 144.9458 0.00029654 -85.218 0.30094
5.405 0.98809 5.4892e-005 3.8183 0.011972 7.0632e-005 0.0011617 0.23211 0.0006593 0.23276 0.21475 0 0.032339 0.0389 0 1.3056 0.43981 0.13328 0.016529 9.5537 0.10299 0.00013068 0.78714 0.0080162 0.008917 0.0014895 0.98559 0.99082 3.2259e-006 1.2904e-005 0.15406 0.76377 0.83096 0.0014507 0.88453 0.43683 0.0019524 0.42155 1.6206 1.618 16.0114 144.9459 0.00029592 -85.2211 0.30194
5.406 0.98809 5.4892e-005 3.8183 0.011972 7.0645e-005 0.0011617 0.23211 0.0006593 0.23276 0.21475 0 0.032338 0.0389 0 1.3057 0.43986 0.1333 0.01653 9.5558 0.103 0.00013069 0.78713 0.0080168 0.0089177 0.0014887 0.9856 0.99082 3.2241e-006 1.2897e-005 0.15407 0.76446 0.83138 0.0014503 0.88523 0.43702 0.0019519 0.42156 1.6221 1.6195 16.0114 144.9459 0.00029529 -85.2243 0.30294
5.407 0.98809 5.4891e-005 3.8183 0.011972 7.0658e-005 0.0011617 0.23211 0.0006593 0.23277 0.21475 0 0.032338 0.0389 0 1.3058 0.4399 0.13332 0.016532 9.5578 0.10301 0.0001307 0.78712 0.0080174 0.0089183 0.001488 0.98561 0.99083 3.2223e-006 1.289e-005 0.15407 0.76514 0.83179 0.0014499 0.88593 0.43721 0.0019514 0.42157 1.6235 1.621 16.0115 144.9459 0.00029467 -85.2275 0.30394
5.408 0.98809 5.4891e-005 3.8183 0.011972 7.0671e-005 0.0011617 0.23211 0.0006593 0.23277 0.21475 0 0.032338 0.0389 0 1.3059 0.43995 0.13333 0.016533 9.5599 0.10302 0.00013072 0.78711 0.008018 0.008919 0.0014872 0.98562 0.99084 3.2206e-006 1.2882e-005 0.15407 0.76582 0.8322 0.0014495 0.88662 0.43741 0.0019508 0.42158 1.625 1.6225 16.0115 144.9459 0.00029405 -85.2306 0.30494
5.409 0.98809 5.4891e-005 3.8183 0.011972 7.0684e-005 0.0011617 0.23211 0.0006593 0.23277 0.21475 0 0.032338 0.0389 0 1.306 0.44 0.13335 0.016535 9.5619 0.10303 0.00013073 0.7871 0.0080186 0.0089196 0.0014864 0.98563 0.99084 3.2188e-006 1.2875e-005 0.15408 0.7665 0.8326 0.0014492 0.88731 0.4376 0.0019503 0.42159 1.6265 1.6239 16.0115 144.9459 0.00029343 -85.2337 0.30594
5.41 0.98809 5.4891e-005 3.8183 0.011972 7.0697e-005 0.0011617 0.23212 0.0006593 0.23277 0.21475 0 0.032338 0.0389 0 1.3061 0.44004 0.13336 0.016536 9.564 0.10304 0.00013074 0.78709 0.0080192 0.0089202 0.0014857 0.98564 0.99085 3.2171e-006 1.2868e-005 0.15408 0.76718 0.83301 0.0014488 0.88799 0.43779 0.0019498 0.4216 1.6279 1.6254 16.0115 144.9459 0.00029282 -85.2367 0.30694
5.411 0.98809 5.4891e-005 3.8183 0.011972 7.071e-005 0.0011617 0.23212 0.0006593 0.23277 0.21476 0 0.032338 0.0389 0 1.3062 0.44009 0.13338 0.016538 9.566 0.10305 0.00013075 0.78708 0.0080198 0.0089209 0.0014849 0.98565 0.99086 3.2153e-006 1.2861e-005 0.15409 0.76785 0.83341 0.0014484 0.88867 0.43799 0.0019493 0.42161 1.6294 1.6268 16.0115 144.946 0.00029221 -85.2398 0.30794
5.412 0.98809 5.4891e-005 3.8183 0.011972 7.0723e-005 0.0011617 0.23212 0.0006593 0.23277 0.21476 0 0.032338 0.0389 0 1.3063 0.44013 0.13339 0.016539 9.5681 0.10305 0.00013077 0.78708 0.0080203 0.0089215 0.0014842 0.98566 0.99086 3.2136e-006 1.2855e-005 0.15409 0.76852 0.83381 0.001448 0.88935 0.43818 0.0019488 0.42162 1.6308 1.6283 16.0115 144.946 0.0002916 -85.2428 0.30894
5.413 0.98809 5.4891e-005 3.8183 0.011972 7.0736e-005 0.0011617 0.23212 0.0006593 0.23278 0.21476 0 0.032338 0.0389 0 1.3063 0.44018 0.13341 0.016541 9.5701 0.10306 0.00013078 0.78707 0.0080209 0.0089221 0.0014834 0.98567 0.99087 3.2119e-006 1.2848e-005 0.1541 0.76919 0.83421 0.0014476 0.89002 0.43837 0.0019483 0.42164 1.6322 1.6297 16.0116 144.946 0.000291 -85.2458 0.30994
5.414 0.98809 5.4891e-005 3.8183 0.011972 7.0749e-005 0.0011617 0.23212 0.0006593 0.23278 0.21476 0 0.032338 0.0389 0 1.3064 0.44023 0.13342 0.016542 9.5722 0.10307 0.00013079 0.78706 0.0080215 0.0089228 0.0014827 0.98568 0.99088 3.2102e-006 1.2841e-005 0.1541 0.76986 0.83461 0.0014472 0.89069 0.43857 0.0019478 0.42165 1.6337 1.6312 16.0116 144.946 0.0002904 -85.2488 0.31094
5.415 0.98809 5.4891e-005 3.8183 0.011972 7.0762e-005 0.0011617 0.23213 0.0006593 0.23278 0.21476 0 0.032338 0.0389 0 1.3065 0.44027 0.13344 0.016544 9.5742 0.10308 0.00013081 0.78705 0.0080221 0.0089234 0.0014819 0.98569 0.99088 3.2085e-006 1.2834e-005 0.15411 0.77052 0.83501 0.0014469 0.89135 0.43876 0.0019473 0.42166 1.6351 1.6326 16.0116 144.946 0.0002898 -85.2518 0.31194
5.416 0.98809 5.4891e-005 3.8183 0.011972 7.0775e-005 0.0011617 0.23213 0.0006593 0.23278 0.21477 0 0.032338 0.0389 0 1.3066 0.44032 0.13345 0.016545 9.5763 0.10309 0.00013082 0.78704 0.0080227 0.008924 0.0014812 0.9857 0.99089 3.2068e-006 1.2827e-005 0.15411 0.77119 0.8354 0.0014465 0.89201 0.43895 0.0019468 0.42167 1.6365 1.6341 16.0116 144.9461 0.0002892 -85.2547 0.31294
5.417 0.98809 5.4891e-005 3.8183 0.011971 7.0788e-005 0.0011617 0.23213 0.0006593 0.23278 0.21477 0 0.032337 0.0389 0 1.3067 0.44037 0.13347 0.016546 9.5783 0.1031 0.00013083 0.78703 0.0080233 0.0089247 0.0014805 0.98571 0.9909 3.2052e-006 1.2821e-005 0.15412 0.77185 0.83579 0.0014461 0.89267 0.43914 0.0019464 0.42168 1.638 1.6355 16.0116 144.9461 0.00028861 -85.2576 0.31394
5.418 0.98809 5.4891e-005 3.8183 0.011971 7.0801e-005 0.0011617 0.23213 0.0006593 0.23279 0.21477 0 0.032337 0.0389 0 1.3068 0.44041 0.13348 0.016548 9.5804 0.10311 0.00013084 0.78702 0.0080239 0.0089253 0.0014798 0.98572 0.9909 3.2036e-006 1.2814e-005 0.15412 0.77251 0.83618 0.0014457 0.89332 0.43934 0.0019459 0.42169 1.6394 1.6369 16.0116 144.9461 0.00028801 -85.2605 0.31494
5.419 0.98809 5.4891e-005 3.8183 0.011971 7.0814e-005 0.0011617 0.23213 0.0006593 0.23279 0.21477 0 0.032337 0.0389 0 1.3069 0.44046 0.1335 0.016549 9.5824 0.10312 0.00013086 0.78701 0.0080245 0.0089259 0.0014791 0.98573 0.99091 3.2019e-006 1.2808e-005 0.15413 0.77317 0.83657 0.0014454 0.89397 0.43953 0.0019454 0.4217 1.6408 1.6384 16.0117 144.9461 0.00028743 -85.2634 0.31594
5.42 0.98809 5.489e-005 3.8183 0.011971 7.0827e-005 0.0011617 0.23214 0.0006593 0.23279 0.21477 0 0.032337 0.0389 0 1.307 0.44051 0.13351 0.016551 9.5845 0.10313 0.00013087 0.787 0.008025 0.0089266 0.0014784 0.98574 0.99091 3.2003e-006 1.2801e-005 0.15413 0.77382 0.83696 0.001445 0.89462 0.43972 0.0019449 0.42172 1.6422 1.6398 16.0117 144.9461 0.00028684 -85.2662 0.31694
5.421 0.98809 5.489e-005 3.8183 0.011971 7.0839e-005 0.0011617 0.23214 0.0006593 0.23279 0.21477 0 0.032337 0.0389 0 1.3071 0.44055 0.13353 0.016552 9.5866 0.10314 0.00013088 0.787 0.0080256 0.0089272 0.0014777 0.98575 0.99092 3.1987e-006 1.2795e-005 0.15414 0.77447 0.83734 0.0014447 0.89526 0.43992 0.0019445 0.42173 1.6436 1.6412 16.0117 144.9461 0.00028626 -85.2691 0.31794
5.422 0.98809 5.489e-005 3.8183 0.011971 7.0852e-005 0.0011617 0.23214 0.0006593 0.23279 0.21478 0 0.032337 0.0389 0 1.3072 0.4406 0.13355 0.016554 9.5886 0.10314 0.0001309 0.78699 0.0080262 0.0089278 0.001477 0.98576 0.99093 3.1971e-006 1.2789e-005 0.15414 0.77513 0.83772 0.0014443 0.89589 0.44011 0.001944 0.42174 1.645 1.6426 16.0117 144.9462 0.00028568 -85.2719 0.31894
5.423 0.98809 5.489e-005 3.8183 0.011971 7.0865e-005 0.0011617 0.23214 0.0006593 0.2328 0.21478 0 0.032337 0.0389 0 1.3073 0.44065 0.13356 0.016555 9.5907 0.10315 0.00013091 0.78698 0.0080268 0.0089285 0.0014763 0.98577 0.99093 3.1955e-006 1.2782e-005 0.15414 0.77578 0.8381 0.001444 0.89653 0.4403 0.0019435 0.42175 1.6464 1.644 16.0117 144.9462 0.0002851 -85.2747 0.31994
5.424 0.98809 5.489e-005 3.8183 0.011971 7.0878e-005 0.0011617 0.23214 0.0006593 0.2328 0.21478 0 0.032337 0.0389 0 1.3074 0.44069 0.13358 0.016557 9.5927 0.10316 0.00013092 0.78697 0.0080274 0.0089291 0.0014756 0.98578 0.99094 3.194e-006 1.2776e-005 0.15415 0.77642 0.83848 0.0014436 0.89716 0.44049 0.0019431 0.42176 1.6478 1.6454 16.0117 144.9462 0.00028452 -85.2775 0.32094
5.425 0.98809 5.489e-005 3.8183 0.011971 7.0891e-005 0.0011617 0.23215 0.0006593 0.2328 0.21478 0 0.032337 0.0389 0 1.3075 0.44074 0.13359 0.016558 9.5948 0.10317 0.00013093 0.78696 0.008028 0.0089297 0.001475 0.98579 0.99094 3.1924e-006 1.277e-005 0.15415 0.77707 0.83886 0.0014433 0.89778 0.44069 0.0019426 0.42177 1.6492 1.6468 16.0118 144.9462 0.00028395 -85.2802 0.32194
5.426 0.98809 5.489e-005 3.8183 0.011971 7.0904e-005 0.0011617 0.23215 0.0006593 0.2328 0.21478 0 0.032337 0.0389 0 1.3076 0.44079 0.13361 0.01656 9.5968 0.10318 0.00013095 0.78695 0.0080286 0.0089304 0.0014743 0.9858 0.99095 3.1909e-006 1.2764e-005 0.15416 0.77771 0.83923 0.0014429 0.89841 0.44088 0.0019422 0.42179 1.6506 1.6482 16.0118 144.9462 0.00028338 -85.2829 0.32294
5.427 0.98809 5.489e-005 3.8183 0.011971 7.0917e-005 0.0011617 0.23215 0.0006593 0.2328 0.21479 0 0.032336 0.0389 0 1.3077 0.44083 0.13362 0.016561 9.5989 0.10319 0.00013096 0.78694 0.0080292 0.008931 0.0014736 0.9858 0.99096 3.1893e-006 1.2757e-005 0.15416 0.77835 0.83961 0.0014426 0.89902 0.44107 0.0019417 0.4218 1.652 1.6496 16.0118 144.9462 0.00028281 -85.2856 0.32394
5.428 0.98809 5.489e-005 3.8183 0.011971 7.093e-005 0.0011618 0.23215 0.0006593 0.23281 0.21479 0 0.032336 0.0389 0 1.3078 0.44088 0.13364 0.016562 9.6009 0.1032 0.00013097 0.78693 0.0080298 0.0089316 0.001473 0.98581 0.99096 3.1878e-006 1.2751e-005 0.15417 0.77899 0.83998 0.0014423 0.89964 0.44126 0.0019413 0.42181 1.6534 1.651 16.0118 144.9463 0.00028225 -85.2883 0.32494
5.429 0.98809 5.489e-005 3.8183 0.011971 7.0943e-005 0.0011618 0.23215 0.0006593 0.23281 0.21479 0 0.032336 0.0389 0 1.3079 0.44092 0.13365 0.016564 9.603 0.10321 0.00013099 0.78692 0.0080303 0.0089323 0.0014723 0.98582 0.99097 3.1863e-006 1.2745e-005 0.15417 0.77963 0.84035 0.0014419 0.90025 0.44146 0.0019408 0.42182 1.6548 1.6524 16.0118 144.9463 0.00028169 -85.291 0.32594
5.43 0.98809 5.489e-005 3.8183 0.011971 7.0956e-005 0.0011618 0.23215 0.0006593 0.23281 0.21479 0 0.032336 0.0389 0 1.308 0.44097 0.13367 0.016565 9.6051 0.10322 0.000131 0.78692 0.0080309 0.0089329 0.0014717 0.98583 0.99097 3.1848e-006 1.2739e-005 0.15418 0.78026 0.84071 0.0014416 0.90086 0.44165 0.0019404 0.42183 1.6561 1.6538 16.0118 144.9463 0.00028113 -85.2937 0.32694
5.431 0.98809 5.489e-005 3.8183 0.011971 7.0969e-005 0.0011618 0.23216 0.0006593 0.23281 0.21479 0 0.032336 0.0389 0 1.3081 0.44102 0.13368 0.016567 9.6071 0.10322 0.00013101 0.78691 0.0080315 0.0089335 0.001471 0.98584 0.99098 3.1833e-006 1.2733e-005 0.15418 0.7809 0.84108 0.0014412 0.90146 0.44184 0.00194 0.42184 1.6575 1.6552 16.0118 144.9463 0.00028057 -85.2963 0.32794
5.432 0.98809 5.489e-005 3.8183 0.011971 7.0982e-005 0.0011618 0.23216 0.0006593 0.23281 0.21479 0 0.032336 0.0389 0 1.3082 0.44106 0.1337 0.016568 9.6092 0.10323 0.00013102 0.7869 0.0080321 0.0089342 0.0014704 0.98585 0.99099 3.1819e-006 1.2728e-005 0.15419 0.78153 0.84144 0.0014409 0.90206 0.44203 0.0019395 0.42186 1.6589 1.6565 16.0119 144.9463 0.00028002 -85.2989 0.32894
5.433 0.98809 5.4889e-005 3.8183 0.011971 7.0995e-005 0.0011618 0.23216 0.0006593 0.23282 0.2148 0 0.032336 0.0389 0 1.3082 0.44111 0.13371 0.01657 9.6112 0.10324 0.00013104 0.78689 0.0080327 0.0089348 0.0014697 0.98586 0.99099 3.1804e-006 1.2722e-005 0.15419 0.78216 0.84181 0.0014406 0.90266 0.44223 0.0019391 0.42187 1.6603 1.6579 16.0119 144.9464 0.00027946 -85.3015 0.32994
5.434 0.98809 5.4889e-005 3.8183 0.011971 7.1008e-005 0.0011618 0.23216 0.0006593 0.23282 0.2148 0 0.032336 0.0389 0 1.3083 0.44116 0.13373 0.016571 9.6133 0.10325 0.00013105 0.78688 0.0080333 0.0089354 0.0014691 0.98586 0.991 3.1789e-006 1.2716e-005 0.1542 0.78279 0.84217 0.0014403 0.90325 0.44242 0.0019387 0.42188 1.6616 1.6593 16.0119 144.9464 0.00027891 -85.3041 0.33094
5.435 0.98809 5.4889e-005 3.8183 0.011971 7.1021e-005 0.0011618 0.23216 0.0006593 0.23282 0.2148 0 0.032336 0.0389 0 1.3084 0.4412 0.13374 0.016573 9.6154 0.10326 0.00013106 0.78687 0.0080339 0.0089361 0.0014685 0.98587 0.991 3.1775e-006 1.271e-005 0.1542 0.78341 0.84253 0.0014399 0.90384 0.44261 0.0019383 0.42189 1.663 1.6607 16.0119 144.9464 0.00027837 -85.3066 0.33194
5.436 0.98809 5.4889e-005 3.8183 0.011971 7.1034e-005 0.0011618 0.23217 0.0006593 0.23282 0.2148 0 0.032336 0.0389 0 1.3085 0.44125 0.13376 0.016574 9.6174 0.10327 0.00013107 0.78686 0.0080344 0.0089367 0.0014678 0.98588 0.99101 3.1761e-006 1.2704e-005 0.1542 0.78404 0.84288 0.0014396 0.90443 0.4428 0.0019378 0.4219 1.6643 1.662 16.0119 144.9464 0.00027782 -85.3092 0.33294
5.437 0.98809 5.4889e-005 3.8183 0.011971 7.1047e-005 0.0011618 0.23217 0.0006593 0.23282 0.2148 0 0.032336 0.0389 0 1.3086 0.4413 0.13378 0.016575 9.6195 0.10328 0.00013109 0.78685 0.008035 0.0089373 0.0014672 0.98589 0.99101 3.1747e-006 1.2699e-005 0.15421 0.78466 0.84324 0.0014393 0.90501 0.44299 0.0019374 0.42192 1.6657 1.6634 16.0119 144.9464 0.00027728 -85.3117 0.33394
5.438 0.98809 5.4889e-005 3.8183 0.011971 7.106e-005 0.0011618 0.23217 0.0006593 0.23282 0.21481 0 0.032335 0.0389 0 1.3087 0.44134 0.13379 0.016577 9.6215 0.10329 0.0001311 0.78684 0.0080356 0.008938 0.0014666 0.9859 0.99102 3.1733e-006 1.2693e-005 0.15421 0.78528 0.84359 0.001439 0.90559 0.44319 0.001937 0.42193 1.667 1.6647 16.0119 144.9464 0.00027674 -85.3142 0.33494
5.439 0.98809 5.4889e-005 3.8183 0.011971 7.1072e-005 0.0011618 0.23217 0.0006593 0.23283 0.21481 0 0.032335 0.0389 0 1.3088 0.44139 0.13381 0.016578 9.6236 0.1033 0.00013111 0.78684 0.0080362 0.0089386 0.001466 0.9859 0.99102 3.1719e-006 1.2688e-005 0.15422 0.78589 0.84394 0.0014387 0.90616 0.44338 0.0019366 0.42194 1.6684 1.6661 16.0119 144.9465 0.0002762 -85.3167 0.33594
5.44 0.98809 5.4889e-005 3.8183 0.011971 7.1085e-005 0.0011618 0.23217 0.0006593 0.23283 0.21481 0 0.032335 0.0389 0 1.3089 0.44144 0.13382 0.01658 9.6257 0.1033 0.00013113 0.78683 0.0080368 0.0089392 0.0014654 0.98591 0.99103 3.1705e-006 1.2682e-005 0.15422 0.78651 0.84429 0.0014384 0.90674 0.44357 0.0019362 0.42195 1.6697 1.6674 16.012 144.9465 0.00027567 -85.3191 0.33694
5.441 0.98809 5.4889e-005 3.8183 0.011971 7.1098e-005 0.0011618 0.23218 0.0006593 0.23283 0.21481 0 0.032335 0.0389 0 1.309 0.44148 0.13384 0.016581 9.6277 0.10331 0.00013114 0.78682 0.0080374 0.0089399 0.0014648 0.98592 0.99103 3.1691e-006 1.2677e-005 0.15423 0.78712 0.84464 0.0014381 0.9073 0.44376 0.0019358 0.42196 1.671 1.6688 16.012 144.9465 0.00027514 -85.3216 0.33794
5.442 0.98809 5.4889e-005 3.8183 0.011971 7.1111e-005 0.0011618 0.23218 0.0006593 0.23283 0.21481 0 0.032335 0.0389 0 1.3091 0.44153 0.13385 0.016583 9.6298 0.10332 0.00013115 0.78681 0.008038 0.0089405 0.0014642 0.98593 0.99104 3.1678e-006 1.2671e-005 0.15423 0.78774 0.84499 0.0014378 0.90787 0.44395 0.0019354 0.42198 1.6724 1.6701 16.012 144.9465 0.00027461 -85.324 0.33894
5.443 0.98809 5.4889e-005 3.8183 0.011971 7.1124e-005 0.0011618 0.23218 0.0006593 0.23283 0.21481 0 0.032335 0.0389 0 1.3092 0.44158 0.13387 0.016584 9.6318 0.10333 0.00013116 0.7868 0.0080386 0.0089411 0.0014636 0.98594 0.99104 3.1664e-006 1.2666e-005 0.15424 0.78835 0.84534 0.0014375 0.90843 0.44414 0.001935 0.42199 1.6737 1.6714 16.012 144.9465 0.00027408 -85.3264 0.33994
5.444 0.98809 5.4889e-005 3.8183 0.011971 7.1137e-005 0.0011618 0.23218 0.0006593 0.23284 0.21482 0 0.032335 0.0389 0 1.3093 0.44162 0.13388 0.016586 9.6339 0.10334 0.00013118 0.78679 0.0080391 0.0089418 0.0014631 0.98594 0.99105 3.1651e-006 1.266e-005 0.15424 0.78896 0.84568 0.0014372 0.90899 0.44434 0.0019346 0.422 1.675 1.6728 16.012 144.9465 0.00027355 -85.3288 0.34094
5.445 0.98809 5.4889e-005 3.8183 0.011971 7.115e-005 0.0011618 0.23218 0.0006593 0.23284 0.21482 0 0.032335 0.0389 0 1.3094 0.44167 0.1339 0.016587 9.636 0.10335 0.00013119 0.78678 0.0080397 0.0089424 0.0014625 0.98595 0.99105 3.1637e-006 1.2655e-005 0.15425 0.78956 0.84602 0.0014369 0.90954 0.44453 0.0019342 0.42201 1.6763 1.6741 16.012 144.9466 0.00027303 -85.3312 0.34194
5.446 0.98809 5.4889e-005 3.8183 0.011971 7.1163e-005 0.0011618 0.23218 0.0006593 0.23284 0.21482 0 0.032335 0.0389 0 1.3095 0.44171 0.13391 0.016589 9.638 0.10336 0.0001312 0.78677 0.0080403 0.008943 0.0014619 0.98596 0.99106 3.1624e-006 1.265e-005 0.15425 0.79017 0.84636 0.0014366 0.9101 0.44472 0.0019338 0.42202 1.6777 1.6754 16.012 144.9466 0.00027251 -85.3336 0.34294
5.447 0.98809 5.4888e-005 3.8183 0.011971 7.1176e-005 0.0011618 0.23219 0.0006593 0.23284 0.21482 0 0.032335 0.0389 0 1.3096 0.44176 0.13393 0.01659 9.6401 0.10337 0.00013121 0.78676 0.0080409 0.0089437 0.0014613 0.98597 0.99106 3.1611e-006 1.2644e-005 0.15426 0.79077 0.8467 0.0014363 0.91064 0.44491 0.0019334 0.42204 1.679 1.6768 16.012 144.9466 0.00027199 -85.3359 0.34394
5.448 0.98809 5.4888e-005 3.8183 0.011971 7.1189e-005 0.0011618 0.23219 0.0006593 0.23284 0.21482 0 0.032335 0.0389 0 1.3097 0.44181 0.13394 0.016591 9.6422 0.10338 0.00013123 0.78676 0.0080415 0.0089443 0.0014608 0.98597 0.99107 3.1598e-006 1.2639e-005 0.15426 0.79137 0.84704 0.001436 0.91119 0.4451 0.0019331 0.42205 1.6803 1.6781 16.012 144.9466 0.00027147 -85.3382 0.34494
5.449 0.98809 5.4888e-005 3.8183 0.011971 7.1202e-005 0.0011618 0.23219 0.0006593 0.23285 0.21482 0 0.032334 0.0389 0 1.3098 0.44185 0.13396 0.016593 9.6442 0.10338 0.00013124 0.78675 0.0080421 0.0089449 0.0014602 0.98598 0.99107 3.1585e-006 1.2634e-005 0.15426 0.79197 0.84738 0.0014357 0.91173 0.44529 0.0019327 0.42206 1.6816 1.6794 16.0121 144.9466 0.00027096 -85.3405 0.34594
5.45 0.98809 5.4888e-005 3.8183 0.011971 7.1215e-005 0.0011618 0.23219 0.0006593 0.23285 0.21483 0 0.032334 0.0389 0 1.3099 0.4419 0.13397 0.016594 9.6463 0.10339 0.00013125 0.78674 0.0080427 0.0089455 0.0014597 0.98599 0.99108 3.1572e-006 1.2629e-005 0.15427 0.79257 0.84771 0.0014354 0.91227 0.44548 0.0019323 0.42207 1.6829 1.6807 16.0121 144.9467 0.00027045 -85.3428 0.34694
5.451 0.98809 5.4888e-005 3.8183 0.011971 7.1228e-005 0.0011618 0.23219 0.0006593 0.23285 0.21483 0 0.032334 0.0389 0 1.31 0.44195 0.13399 0.016596 9.6484 0.1034 0.00013127 0.78673 0.0080432 0.0089462 0.0014591 0.986 0.99108 3.156e-006 1.2624e-005 0.15427 0.79316 0.84804 0.0014351 0.9128 0.44568 0.0019319 0.42209 1.6842 1.682 16.0121 144.9467 0.00026994 -85.3451 0.34794
5.452 0.98809 5.4888e-005 3.8183 0.011971 7.1241e-005 0.0011618 0.2322 0.0006593 0.23285 0.21483 0 0.032334 0.0389 0 1.3101 0.44199 0.13401 0.016597 9.6504 0.10341 0.00013128 0.78672 0.0080438 0.0089468 0.0014585 0.986 0.99109 3.1547e-006 1.2619e-005 0.15428 0.79375 0.84837 0.0014348 0.91333 0.44587 0.0019316 0.4221 1.6855 1.6833 16.0121 144.9467 0.00026943 -85.3474 0.34894
5.453 0.98809 5.4888e-005 3.8183 0.011971 7.1254e-005 0.0011618 0.2322 0.0006593 0.23285 0.21483 0 0.032334 0.0389 0 1.3101 0.44204 0.13402 0.016599 9.6525 0.10342 0.00013129 0.78671 0.0080444 0.0089474 0.001458 0.98601 0.99109 3.1534e-006 1.2614e-005 0.15428 0.79435 0.8487 0.0014345 0.91386 0.44606 0.0019312 0.42211 1.6868 1.6846 16.0121 144.9467 0.00026893 -85.3496 0.34994
5.454 0.98809 5.4888e-005 3.8183 0.011971 7.1267e-005 0.0011618 0.2322 0.0006593 0.23285 0.21483 0 0.032334 0.0389 0 1.3102 0.44209 0.13404 0.0166 9.6546 0.10343 0.0001313 0.7867 0.008045 0.0089481 0.0014574 0.98602 0.9911 3.1522e-006 1.2609e-005 0.15429 0.79494 0.84903 0.0014343 0.91439 0.44625 0.0019308 0.42212 1.6881 1.6859 16.0121 144.9467 0.00026843 -85.3518 0.35094
5.455 0.98809 5.4888e-005 3.8183 0.011971 7.128e-005 0.0011618 0.2322 0.0006593 0.23286 0.21484 0 0.032334 0.0389 0 1.3103 0.44213 0.13405 0.016602 9.6566 0.10344 0.00013132 0.78669 0.0080456 0.0089487 0.0014569 0.98602 0.9911 3.151e-006 1.2604e-005 0.15429 0.79552 0.84936 0.001434 0.91491 0.44644 0.0019305 0.42214 1.6894 1.6872 16.0121 144.9467 0.00026793 -85.354 0.35194
5.456 0.98809 5.4888e-005 3.8183 0.011971 7.1293e-005 0.0011618 0.2322 0.0006593 0.23286 0.21484 0 0.032334 0.0389 0 1.3104 0.44218 0.13407 0.016603 9.6587 0.10345 0.00013133 0.78668 0.0080462 0.0089493 0.0014564 0.98603 0.99111 3.1497e-006 1.2599e-005 0.1543 0.79611 0.84968 0.0014337 0.91543 0.44663 0.0019301 0.42215 1.6906 1.6885 16.0121 144.9468 0.00026743 -85.3562 0.35294
5.457 0.98809 5.4888e-005 3.8183 0.011971 7.1305e-005 0.0011618 0.23221 0.0006593 0.23286 0.21484 0 0.032334 0.0389 0 1.3105 0.44223 0.13408 0.016604 9.6608 0.10346 0.00013134 0.78668 0.0080467 0.00895 0.0014558 0.98604 0.99111 3.1485e-006 1.2594e-005 0.1543 0.79669 0.85001 0.0014334 0.91595 0.44682 0.0019298 0.42216 1.6919 1.6898 16.0121 144.9468 0.00026693 -85.3584 0.35394
5.458 0.98809 5.4888e-005 3.8183 0.011971 7.1318e-005 0.0011618 0.23221 0.0006593 0.23286 0.21484 0 0.032334 0.0389 0 1.3106 0.44227 0.1341 0.016606 9.6628 0.10346 0.00013136 0.78667 0.0080473 0.0089506 0.0014553 0.98605 0.99112 3.1473e-006 1.2589e-005 0.15431 0.79728 0.85033 0.0014331 0.91646 0.44701 0.0019294 0.42217 1.6932 1.6911 16.0121 144.9468 0.00026644 -85.3606 0.35494
5.459 0.98809 5.4888e-005 3.8183 0.011971 7.1331e-005 0.0011619 0.23221 0.0006593 0.23286 0.21484 0 0.032333 0.0389 0 1.3107 0.44232 0.13411 0.016607 9.6649 0.10347 0.00013137 0.78666 0.0080479 0.0089512 0.0014548 0.98605 0.99112 3.1461e-006 1.2585e-005 0.15431 0.79786 0.85065 0.0014329 0.91697 0.4472 0.001929 0.42219 1.6945 1.6923 16.0121 144.9468 0.00026595 -85.3627 0.35594
5.46 0.98809 5.4887e-005 3.8183 0.011971 7.1344e-005 0.0011619 0.23221 0.0006593 0.23287 0.21484 0 0.032333 0.0389 0 1.3108 0.44236 0.13413 0.016609 9.667 0.10348 0.00013138 0.78665 0.0080485 0.0089519 0.0014543 0.98606 0.99113 3.1449e-006 1.258e-005 0.15432 0.79844 0.85097 0.0014326 0.91747 0.44739 0.0019287 0.4222 1.6957 1.6936 16.0122 144.9468 0.00026546 -85.3649 0.35694
5.461 0.98809 5.4887e-005 3.8183 0.011971 7.1357e-005 0.0011619 0.23221 0.0006593 0.23287 0.21485 0 0.032333 0.0389 0 1.3109 0.44241 0.13414 0.01661 9.669 0.10349 0.00013139 0.78664 0.0080491 0.0089525 0.0014538 0.98607 0.99113 3.1438e-006 1.2575e-005 0.15432 0.79901 0.85129 0.0014323 0.91798 0.44759 0.0019283 0.42221 1.697 1.6949 16.0122 144.9469 0.00026497 -85.367 0.35794
5.462 0.98809 5.4887e-005 3.8183 0.011971 7.137e-005 0.0011619 0.23221 0.0006593 0.23287 0.21485 0 0.032333 0.0389 0 1.311 0.44246 0.13416 0.016612 9.6711 0.1035 0.00013141 0.78663 0.0080497 0.0089531 0.0014532 0.98607 0.99113 3.1426e-006 1.257e-005 0.15432 0.79959 0.8516 0.0014321 0.91848 0.44778 0.001928 0.42222 1.6983 1.6961 16.0122 144.9469 0.00026449 -85.3691 0.35894
5.463 0.98809 5.4887e-005 3.8183 0.011971 7.1383e-005 0.0011619 0.23222 0.0006593 0.23287 0.21485 0 0.032333 0.0389 0 1.3111 0.4425 0.13417 0.016613 9.6732 0.10351 0.00013142 0.78662 0.0080503 0.0089537 0.0014527 0.98608 0.99114 3.1414e-006 1.2566e-005 0.15433 0.80016 0.85192 0.0014318 0.91898 0.44797 0.0019277 0.42223 1.6995 1.6974 16.0122 144.9469 0.000264 -85.3712 0.35994
5.464 0.98809 5.4887e-005 3.8183 0.011971 7.1396e-005 0.0011619 0.23222 0.0006593 0.23287 0.21485 0 0.032333 0.0389 0 1.3112 0.44255 0.13419 0.016615 9.6752 0.10352 0.00013143 0.78661 0.0080508 0.0089544 0.0014523 0.98609 0.99114 3.1403e-006 1.2561e-005 0.15433 0.80073 0.85223 0.0014316 0.91947 0.44816 0.0019273 0.42225 1.7008 1.6987 16.0122 144.9469 0.00026352 -85.3732 0.36094
5.465 0.98809 5.4887e-005 3.8183 0.011971 7.1409e-005 0.0011619 0.23222 0.0006593 0.23287 0.21485 0 0.032333 0.0389 0 1.3113 0.4426 0.1342 0.016616 9.6773 0.10353 0.00013144 0.78661 0.0080514 0.008955 0.0014518 0.98609 0.99115 3.1391e-006 1.2557e-005 0.15434 0.8013 0.85254 0.0014313 0.91996 0.44835 0.001927 0.42226 1.702 1.6999 16.0122 144.9469 0.00026304 -85.3753 0.36194
5.466 0.98809 5.4887e-005 3.8183 0.011971 7.1422e-005 0.0011619 0.23222 0.0006593 0.23288 0.21485 0 0.032333 0.0389 0 1.3114 0.44264 0.13422 0.016618 9.6794 0.10354 0.00013146 0.7866 0.008052 0.0089556 0.0014513 0.9861 0.99115 3.138e-006 1.2552e-005 0.15434 0.80187 0.85285 0.0014311 0.92045 0.44854 0.0019267 0.42227 1.7033 1.7012 16.0122 144.9469 0.00026257 -85.3773 0.36294
5.467 0.98809 5.4887e-005 3.8183 0.011971 7.1435e-005 0.0011619 0.23222 0.0006593 0.23288 0.21486 0 0.032333 0.0389 0 1.3115 0.44269 0.13423 0.016619 9.6814 0.10354 0.00013147 0.78659 0.0080526 0.0089563 0.0014508 0.98611 0.99116 3.1369e-006 1.2548e-005 0.15435 0.80244 0.85316 0.0014308 0.92093 0.44873 0.0019263 0.42229 1.7045 1.7024 16.0122 144.947 0.00026209 -85.3794 0.36394
5.468 0.98809 5.4887e-005 3.8183 0.011971 7.1448e-005 0.0011619 0.23223 0.0006593 0.23288 0.21486 0 0.032333 0.0389 0 1.3116 0.44274 0.13425 0.01662 9.6835 0.10355 0.00013148 0.78658 0.0080532 0.0089569 0.0014503 0.98611 0.99116 3.1358e-006 1.2543e-005 0.15435 0.803 0.85347 0.0014306 0.92142 0.44892 0.001926 0.4223 1.7058 1.7037 16.0122 144.947 0.00026162 -85.3814 0.36494
5.469 0.98809 5.4887e-005 3.8183 0.011971 7.1461e-005 0.0011619 0.23223 0.0006593 0.23288 0.21486 0 0.032333 0.0389 0 1.3117 0.44278 0.13427 0.016622 9.6856 0.10356 0.0001315 0.78657 0.0080538 0.0089575 0.0014498 0.98612 0.99116 3.1347e-006 1.2539e-005 0.15436 0.80356 0.85378 0.0014303 0.9219 0.44911 0.0019257 0.42231 1.707 1.7049 16.0122 144.947 0.00026115 -85.3834 0.36594
5.47 0.98809 5.4887e-005 3.8183 0.011971 7.1474e-005 0.0011619 0.23223 0.0006593 0.23288 0.21486 0 0.032332 0.0389 0 1.3118 0.44283 0.13428 0.016623 9.6877 0.10357 0.00013151 0.78656 0.0080543 0.0089581 0.0014493 0.98612 0.99117 3.1336e-006 1.2534e-005 0.15436 0.80413 0.85408 0.00143 0.92237 0.4493 0.0019253 0.42232 1.7082 1.7062 16.0122 144.947 0.00026068 -85.3853 0.36694
5.471 0.98809 5.4887e-005 3.8183 0.011971 7.1487e-005 0.0011619 0.23223 0.0006593 0.23289 0.21486 0 0.032332 0.0389 0 1.3119 0.44288 0.1343 0.016625 9.6897 0.10358 0.00013152 0.78655 0.0080549 0.0089588 0.0014488 0.98613 0.99117 3.1325e-006 1.253e-005 0.15437 0.80468 0.85438 0.0014298 0.92285 0.44949 0.001925 0.42234 1.7095 1.7074 16.0122 144.947 0.00026022 -85.3873 0.36794
5.472 0.98809 5.4887e-005 3.8183 0.011971 7.15e-005 0.0011619 0.23223 0.0006593 0.23289 0.21486 0 0.032332 0.0389 0 1.3119 0.44292 0.13431 0.016626 9.6918 0.10359 0.00013153 0.78654 0.0080555 0.0089594 0.0014483 0.98614 0.99118 3.1314e-006 1.2526e-005 0.15437 0.80524 0.85469 0.0014295 0.92332 0.44968 0.0019247 0.42235 1.7107 1.7086 16.0122 144.9471 0.00025975 -85.3893 0.36894
5.473 0.98809 5.4886e-005 3.8183 0.011971 7.1513e-005 0.0011619 0.23223 0.0006593 0.23289 0.21487 0 0.032332 0.0389 0 1.312 0.44297 0.13433 0.016628 9.6939 0.1036 0.00013155 0.78653 0.0080561 0.00896 0.0014479 0.98614 0.99118 3.1303e-006 1.2521e-005 0.15438 0.8058 0.85499 0.0014293 0.92378 0.44987 0.0019244 0.42236 1.7119 1.7099 16.0122 144.9471 0.00025929 -85.3912 0.36994
5.474 0.98809 5.4886e-005 3.8183 0.011971 7.1526e-005 0.0011619 0.23224 0.0006593 0.23289 0.21487 0 0.032332 0.0389 0 1.3121 0.44302 0.13434 0.016629 9.6959 0.10361 0.00013156 0.78653 0.0080567 0.0089607 0.0014474 0.98615 0.99119 3.1292e-006 1.2517e-005 0.15438 0.80635 0.85529 0.0014291 0.92425 0.45006 0.0019241 0.42237 1.7131 1.7111 16.0123 144.9471 0.00025883 -85.3931 0.37094
5.475 0.98809 5.4886e-005 3.8183 0.011971 7.1538e-005 0.0011619 0.23224 0.0006593 0.23289 0.21487 0 0.032332 0.0389 0 1.3122 0.44306 0.13436 0.016631 9.698 0.10361 0.00013157 0.78652 0.0080573 0.0089613 0.001447 0.98615 0.99119 3.1282e-006 1.2513e-005 0.15438 0.8069 0.85558 0.0014288 0.92471 0.45025 0.0019238 0.42239 1.7143 1.7123 16.0123 144.9471 0.00025837 -85.395 0.37194
5.476 0.98809 5.4886e-005 3.8183 0.011971 7.1551e-005 0.0011619 0.23224 0.0006593 0.23289 0.21487 0 0.032332 0.0389 0 1.3123 0.44311 0.13437 0.016632 9.7001 0.10362 0.00013158 0.78651 0.0080578 0.0089619 0.0014465 0.98616 0.99119 3.1271e-006 1.2509e-005 0.15439 0.80746 0.85588 0.0014286 0.92517 0.45044 0.0019234 0.4224 1.7156 1.7135 16.0123 144.9471 0.00025792 -85.3969 0.37294
5.477 0.98809 5.4886e-005 3.8183 0.011971 7.1564e-005 0.0011619 0.23224 0.0006593 0.2329 0.21487 0 0.032332 0.0389 0 1.3124 0.44315 0.13439 0.016633 9.7022 0.10363 0.0001316 0.7865 0.0080584 0.0089626 0.001446 0.98617 0.9912 3.1261e-006 1.2504e-005 0.15439 0.808 0.85618 0.0014283 0.92563 0.45063 0.0019231 0.42241 1.7168 1.7148 16.0123 144.9471 0.00025746 -85.3988 0.37394
5.478 0.98809 5.4886e-005 3.8183 0.011971 7.1577e-005 0.0011619 0.23224 0.0006593 0.2329 0.21488 0 0.032332 0.0389 0 1.3125 0.4432 0.1344 0.016635 9.7042 0.10364 0.00013161 0.78649 0.008059 0.0089632 0.0014456 0.98617 0.9912 3.1251e-006 1.25e-005 0.1544 0.80855 0.85647 0.0014281 0.92608 0.45082 0.0019228 0.42242 1.718 1.716 16.0123 144.9472 0.00025701 -85.4007 0.37494
5.479 0.98809 5.4886e-005 3.8183 0.01197 7.159e-005 0.0011619 0.23225 0.0006593 0.2329 0.21488 0 0.032332 0.0389 0 1.3126 0.44325 0.13442 0.016636 9.7063 0.10365 0.00013162 0.78648 0.0080596 0.0089638 0.0014452 0.98618 0.9912 3.124e-006 1.2496e-005 0.1544 0.8091 0.85676 0.0014279 0.92653 0.45101 0.0019225 0.42244 1.7192 1.7172 16.0123 144.9472 0.00025656 -85.4026 0.37594
5.48 0.98809 5.4886e-005 3.8183 0.01197 7.1603e-005 0.0011619 0.23225 0.0006593 0.2329 0.21488 0 0.032332 0.0389 0 1.3127 0.44329 0.13443 0.016638 9.7084 0.10366 0.00013164 0.78647 0.0080602 0.0089644 0.0014447 0.98618 0.99121 3.123e-006 1.2492e-005 0.15441 0.80964 0.85705 0.0014277 0.92698 0.4512 0.0019222 0.42245 1.7204 1.7184 16.0123 144.9472 0.00025611 -85.4044 0.37694
5.481 0.98809 5.4886e-005 3.8183 0.01197 7.1616e-005 0.0011619 0.23225 0.0006593 0.2329 0.21488 0 0.032331 0.0389 0 1.3128 0.44334 0.13445 0.016639 9.7105 0.10367 0.00013165 0.78646 0.0080608 0.0089651 0.0014443 0.98619 0.99121 3.122e-006 1.2488e-005 0.15441 0.81018 0.85734 0.0014275 0.92742 0.45139 0.0019219 0.42246 1.7216 1.7196 16.0123 144.9472 0.00025567 -85.4062 0.37794
5.482 0.98809 5.4886e-005 3.8183 0.01197 7.1629e-005 0.0011619 0.23225 0.0006593 0.23291 0.21488 0 0.032331 0.0389 0 1.3129 0.44339 0.13446 0.016641 9.7125 0.10368 0.00013166 0.78645 0.0080613 0.0089657 0.0014439 0.9862 0.99122 3.121e-006 1.2484e-005 0.15442 0.81072 0.85763 0.0014272 0.92787 0.45158 0.0019216 0.42248 1.7228 1.7208 16.0123 144.9472 0.00025522 -85.4081 0.37894
5.483 0.98809 5.4886e-005 3.8183 0.01197 7.1642e-005 0.0011619 0.23225 0.0006593 0.23291 0.21488 0 0.032331 0.0389 0 1.313 0.44343 0.13448 0.016642 9.7146 0.10369 0.00013167 0.78645 0.0080619 0.0089663 0.0014434 0.9862 0.99122 3.12e-006 1.248e-005 0.15442 0.81126 0.85792 0.001427 0.92831 0.45177 0.0019213 0.42249 1.724 1.722 16.0123 144.9473 0.00025478 -85.4099 0.37994
5.484 0.98809 5.4886e-005 3.8183 0.01197 7.1655e-005 0.0011619 0.23225 0.0006593 0.23291 0.21489 0 0.032331 0.0389 0 1.3131 0.44348 0.1345 0.016644 9.7167 0.10369 0.00013169 0.78644 0.0080625 0.008967 0.001443 0.98621 0.99122 3.119e-006 1.2476e-005 0.15443 0.8118 0.85821 0.0014268 0.92874 0.45196 0.001921 0.4225 1.7252 1.7232 16.0123 144.9473 0.00025434 -85.4117 0.38094
5.485 0.98809 5.4886e-005 3.8183 0.01197 7.1668e-005 0.0011619 0.23226 0.0006593 0.23291 0.21489 0 0.032331 0.0389 0 1.3132 0.44353 0.13451 0.016645 9.7188 0.1037 0.0001317 0.78643 0.0080631 0.0089676 0.0014426 0.98621 0.99123 3.118e-006 1.2472e-005 0.15443 0.81234 0.85849 0.0014266 0.92918 0.45215 0.0019207 0.42251 1.7263 1.7244 16.0123 144.9473 0.0002539 -85.4134 0.38194
5.486 0.98809 5.4886e-005 3.8183 0.01197 7.1681e-005 0.0011619 0.23226 0.0006593 0.23291 0.21489 0 0.032331 0.0389 0 1.3133 0.44357 0.13453 0.016646 9.7209 0.10371 0.00013171 0.78642 0.0080637 0.0089682 0.0014421 0.98622 0.99123 3.117e-006 1.2468e-005 0.15444 0.81287 0.85878 0.0014263 0.92961 0.45234 0.0019205 0.42253 1.7275 1.7256 16.0123 144.9473 0.00025346 -85.4152 0.38294
5.487 0.98809 5.4885e-005 3.8183 0.01197 7.1694e-005 0.0011619 0.23226 0.0006593 0.23291 0.21489 0 0.032331 0.0389 0 1.3134 0.44362 0.13454 0.016648 9.7229 0.10372 0.00013172 0.78641 0.0080643 0.0089688 0.0014417 0.98622 0.99123 3.1161e-006 1.2464e-005 0.15444 0.8134 0.85906 0.0014261 0.93004 0.45253 0.0019202 0.42254 1.7287 1.7268 16.0123 144.9473 0.00025303 -85.417 0.38394
5.488 0.98809 5.4885e-005 3.8183 0.01197 7.1707e-005 0.0011619 0.23226 0.0006593 0.23292 0.21489 0 0.032331 0.0389 0 1.3135 0.44367 0.13456 0.016649 9.725 0.10373 0.00013174 0.7864 0.0080648 0.0089695 0.0014413 0.98623 0.99124 3.1151e-006 1.246e-005 0.15444 0.81393 0.85934 0.0014259 0.93047 0.45272 0.0019199 0.42255 1.7299 1.7279 16.0123 144.9474 0.0002526 -85.4187 0.38494
5.489 0.98809 5.4885e-005 3.8183 0.01197 7.172e-005 0.0011619 0.23226 0.0006593 0.23292 0.21489 0 0.032331 0.0389 0 1.3136 0.44371 0.13457 0.016651 9.7271 0.10374 0.00013175 0.78639 0.0080654 0.0089701 0.0014409 0.98624 0.99124 3.1142e-006 1.2457e-005 0.15445 0.81446 0.85962 0.0014257 0.93089 0.4529 0.0019196 0.42257 1.731 1.7291 16.0123 144.9474 0.00025217 -85.4204 0.38594
5.49 0.98809 5.4885e-005 3.8183 0.01197 7.1733e-005 0.001162 0.23227 0.0006593 0.23292 0.2149 0 0.032331 0.0389 0 1.3137 0.44376 0.13459 0.016652 9.7292 0.10375 0.00013176 0.78638 0.008066 0.0089707 0.0014404 0.98624 0.99125 3.1132e-006 1.2453e-005 0.15445 0.81499 0.8599 0.0014254 0.93131 0.45309 0.0019193 0.42258 1.7322 1.7303 16.0123 144.9474 0.00025174 -85.4221 0.38694
5.491 0.98809 5.4885e-005 3.8183 0.01197 7.1746e-005 0.001162 0.23227 0.0006593 0.23292 0.2149 0 0.032331 0.0389 0 1.3137 0.4438 0.1346 0.016654 9.7312 0.10376 0.00013178 0.78638 0.0080666 0.0089713 0.00144 0.98625 0.99125 3.1123e-006 1.2449e-005 0.15446 0.81551 0.86018 0.0014252 0.93173 0.45328 0.001919 0.42259 1.7334 1.7315 16.0123 144.9474 0.00025131 -85.4238 0.38794
5.492 0.98809 5.4885e-005 3.8183 0.01197 7.1758e-005 0.001162 0.23227 0.0006593 0.23292 0.2149 0 0.032331 0.0389 0 1.3138 0.44385 0.13462 0.016655 9.7333 0.10377 0.00013179 0.78637 0.0080672 0.008972 0.0014396 0.98625 0.99125 3.1113e-006 1.2445e-005 0.15446 0.81604 0.86045 0.001425 0.93214 0.45347 0.0019188 0.4226 1.7345 1.7326 16.0123 144.9474 0.00025088 -85.4255 0.38894
5.493 0.98809 5.4885e-005 3.8183 0.01197 7.1771e-005 0.001162 0.23227 0.0006593 0.23293 0.2149 0 0.03233 0.0389 0 1.3139 0.4439 0.13463 0.016657 9.7354 0.10377 0.0001318 0.78636 0.0080677 0.0089726 0.0014392 0.98626 0.99126 3.1104e-006 1.2442e-005 0.15447 0.81656 0.86073 0.0014248 0.93256 0.45366 0.0019185 0.42262 1.7357 1.7338 16.0123 144.9474 0.00025046 -85.4272 0.38994
5.494 0.98809 5.4885e-005 3.8183 0.01197 7.1784e-005 0.001162 0.23227 0.0006593 0.23293 0.2149 0 0.03233 0.0389 0 1.314 0.44394 0.13465 0.016658 9.7375 0.10378 0.00013181 0.78635 0.0080683 0.0089732 0.0014388 0.98626 0.99126 3.1095e-006 1.2438e-005 0.15447 0.81708 0.861 0.0014246 0.93297 0.45385 0.0019182 0.42263 1.7369 1.735 16.0123 144.9475 0.00025004 -85.4289 0.39094
5.495 0.98809 5.4885e-005 3.8183 0.01197 7.1797e-005 0.001162 0.23227 0.0006593 0.23293 0.2149 0 0.03233 0.0389 0 1.3141 0.44399 0.13466 0.016659 9.7396 0.10379 0.00013183 0.78634 0.0080689 0.0089739 0.0014384 0.98627 0.99126 3.1086e-006 1.2434e-005 0.15448 0.8176 0.86127 0.0014244 0.93338 0.45404 0.001918 0.42264 1.738 1.7361 16.0123 144.9475 0.00024962 -85.4305 0.39194
5.496 0.98809 5.4885e-005 3.8183 0.01197 7.181e-005 0.001162 0.23228 0.0006593 0.23293 0.21491 0 0.03233 0.0389 0 1.3142 0.44404 0.13468 0.016661 9.7416 0.1038 0.00013184 0.78633 0.0080695 0.0089745 0.0014381 0.98627 0.99127 3.1077e-006 1.2431e-005 0.15448 0.81812 0.86154 0.0014242 0.93378 0.45423 0.0019177 0.42266 1.7392 1.7373 16.0123 144.9475 0.0002492 -85.4322 0.39294
5.497 0.98809 5.4885e-005 3.8183 0.01197 7.1823e-005 0.001162 0.23228 0.0006593 0.23293 0.21491 0 0.03233 0.0389 0 1.3143 0.44408 0.13469 0.016662 9.7437 0.10381 0.00013185 0.78632 0.0080701 0.0089751 0.0014377 0.98628 0.99127 3.1068e-006 1.2427e-005 0.15449 0.81863 0.86181 0.001424 0.93419 0.45442 0.0019174 0.42267 1.7403 1.7384 16.0123 144.9475 0.00024879 -85.4338 0.39394
5.498 0.98809 5.4885e-005 3.8183 0.01197 7.1836e-005 0.001162 0.23228 0.0006593 0.23293 0.21491 0 0.03233 0.0389 0 1.3144 0.44413 0.13471 0.016664 9.7458 0.10382 0.00013186 0.78631 0.0080707 0.0089757 0.0014373 0.98628 0.99127 3.1059e-006 1.2424e-005 0.15449 0.81915 0.86208 0.0014238 0.93459 0.45461 0.0019172 0.42268 1.7414 1.7396 16.0123 144.9475 0.00024837 -85.4354 0.39494
5.499 0.98809 5.4885e-005 3.8183 0.01197 7.1849e-005 0.001162 0.23228 0.0006593 0.23294 0.21491 0 0.03233 0.0389 0 1.3145 0.44418 0.13472 0.016665 9.7479 0.10383 0.00013188 0.7863 0.0080712 0.0089764 0.0014369 0.98629 0.99128 3.105e-006 1.242e-005 0.15449 0.81966 0.86235 0.0014236 0.93499 0.45479 0.0019169 0.4227 1.7426 1.7407 16.0123 144.9476 0.00024796 -85.4371 0.39594
5.5 0.98809 5.4884e-005 3.8183 0.01197 7.1862e-005 0.001162 0.23228 0.0006593 0.23294 0.21491 0 0.03233 0.0389 0 1.3146 0.44422 0.13474 0.016667 9.75 0.10384 0.00013189 0.7863 0.0080718 0.008977 0.0014365 0.98629 0.99128 3.1041e-006 1.2417e-005 0.1545 0.82017 0.86262 0.0014234 0.93538 0.45498 0.0019166 0.42271 1.7437 1.7419 16.0123 144.9476 0.00024755 -85.4387 0.39694
5.501 0.98809 5.4884e-005 3.8183 0.01197 7.1875e-005 0.001162 0.23228 0.0006593 0.23294 0.21491 0 0.03233 0.0389 0 1.3147 0.44427 0.13476 0.016668 9.7521 0.10384 0.0001319 0.78629 0.0080724 0.0089776 0.0014361 0.9863 0.99128 3.1033e-006 1.2413e-005 0.1545 0.82068 0.86288 0.0014232 0.93577 0.45517 0.0019164 0.42272 1.7449 1.743 16.0123 144.9476 0.00024714 -85.4402 0.39794
5.502 0.98809 5.4884e-005 3.8183 0.01197 7.1888e-005 0.001162 0.23229 0.0006593 0.23294 0.21492 0 0.03233 0.0389 0 1.3148 0.44432 0.13477 0.01667 9.7541 0.10385 0.00013192 0.78628 0.008073 0.0089782 0.0014357 0.9863 0.99129 3.1024e-006 1.241e-005 0.15451 0.82119 0.86315 0.001423 0.93617 0.45536 0.0019161 0.42273 1.746 1.7441 16.0123 144.9476 0.00024673 -85.4418 0.39894
5.503 0.98809 5.4884e-005 3.8183 0.01197 7.1901e-005 0.001162 0.23229 0.0006593 0.23294 0.21492 0 0.03233 0.0389 0 1.3149 0.44436 0.13479 0.016671 9.7562 0.10386 0.00013193 0.78627 0.0080736 0.0089789 0.0014354 0.98631 0.99129 3.1015e-006 1.2406e-005 0.15451 0.82169 0.86341 0.0014228 0.93655 0.45555 0.0019159 0.42275 1.7471 1.7453 16.0123 144.9476 0.00024633 -85.4434 0.39994
5.504 0.98809 5.4884e-005 3.8183 0.01197 7.1914e-005 0.001162 0.23229 0.0006593 0.23294 0.21492 0 0.032329 0.0389 0 1.315 0.44441 0.1348 0.016672 9.7583 0.10387 0.00013194 0.78626 0.0080741 0.0089795 0.001435 0.98631 0.99129 3.1007e-006 1.2403e-005 0.15452 0.8222 0.86367 0.0014226 0.93694 0.45574 0.0019156 0.42276 1.7482 1.7464 16.0124 144.9477 0.00024592 -85.4449 0.40094
5.505 0.98809 5.4884e-005 3.8183 0.01197 7.1927e-005 0.001162 0.23229 0.0006593 0.23295 0.21492 0 0.032329 0.0389 0 1.3151 0.44446 0.13482 0.016674 9.7604 0.10388 0.00013195 0.78625 0.0080747 0.0089801 0.0014346 0.98632 0.9913 3.0998e-006 1.2399e-005 0.15452 0.8227 0.86393 0.0014224 0.93732 0.45592 0.0019154 0.42277 1.7494 1.7475 16.0124 144.9477 0.00024552 -85.4465 0.40194
5.506 0.98809 5.4884e-005 3.8183 0.01197 7.194e-005 0.001162 0.23229 0.0006593 0.23295 0.21492 0 0.032329 0.0389 0 1.3152 0.4445 0.13483 0.016675 9.7625 0.10389 0.00013197 0.78624 0.0080753 0.0089807 0.0014342 0.98632 0.9913 3.099e-006 1.2396e-005 0.15453 0.8232 0.86419 0.0014222 0.93771 0.45611 0.0019151 0.42279 1.7505 1.7487 16.0124 144.9477 0.00024512 -85.448 0.40294
5.507 0.98809 5.4884e-005 3.8183 0.01197 7.1953e-005 0.001162 0.2323 0.0006593 0.23295 0.21492 0 0.032329 0.0389 0 1.3153 0.44455 0.13485 0.016677 9.7646 0.1039 0.00013198 0.78623 0.0080759 0.0089814 0.0014339 0.98633 0.9913 3.0982e-006 1.2393e-005 0.15453 0.8237 0.86445 0.001422 0.93808 0.4563 0.0019149 0.4228 1.7516 1.7498 16.0124 144.9477 0.00024472 -85.4495 0.40394
5.508 0.98809 5.4884e-005 3.8183 0.01197 7.1966e-005 0.001162 0.2323 0.0006593 0.23295 0.21493 0 0.032329 0.0389 0 1.3154 0.44459 0.13486 0.016678 9.7666 0.10391 0.00013199 0.78623 0.0080765 0.008982 0.0014335 0.98633 0.99131 3.0973e-006 1.2389e-005 0.15454 0.8242 0.86471 0.0014218 0.93846 0.45649 0.0019146 0.42281 1.7527 1.7509 16.0124 144.9477 0.00024432 -85.451 0.40494
5.509 0.98809 5.4884e-005 3.8183 0.01197 7.1978e-005 0.001162 0.2323 0.0006593 0.23295 0.21493 0 0.032329 0.0389 0 1.3155 0.44464 0.13488 0.01668 9.7687 0.10392 0.000132 0.78622 0.008077 0.0089826 0.0014332 0.98634 0.99131 3.0965e-006 1.2386e-005 0.15454 0.8247 0.86497 0.0014217 0.93884 0.45668 0.0019144 0.42283 1.7538 1.752 16.0124 144.9477 0.00024393 -85.4525 0.40594
5.51 0.98809 5.4884e-005 3.8183 0.01197 7.1991e-005 0.001162 0.2323 0.0006593 0.23296 0.21493 0 0.032329 0.0389 0 1.3155 0.44469 0.13489 0.016681 9.7708 0.10392 0.00013202 0.78621 0.0080776 0.0089832 0.0014328 0.98634 0.99131 3.0957e-006 1.2383e-005 0.15455 0.8252 0.86522 0.0014215 0.93921 0.45687 0.0019141 0.42284 1.7549 1.7531 16.0124 144.9478 0.00024353 -85.454 0.40694
5.511 0.98809 5.4884e-005 3.8183 0.01197 7.2004e-005 0.001162 0.2323 0.0006593 0.23296 0.21493 0 0.032329 0.0389 0 1.3156 0.44473 0.13491 0.016683 9.7729 0.10393 0.00013203 0.7862 0.0080782 0.0089839 0.0014325 0.98634 0.99131 3.0949e-006 1.238e-005 0.15455 0.82569 0.86548 0.0014213 0.93958 0.45705 0.0019139 0.42285 1.756 1.7542 16.0124 144.9478 0.00024314 -85.4555 0.40794
5.512 0.98809 5.4884e-005 3.8183 0.01197 7.2017e-005 0.001162 0.2323 0.0006593 0.23296 0.21493 0 0.032329 0.0389 0 1.3157 0.44478 0.13492 0.016684 9.775 0.10394 0.00013204 0.78619 0.0080788 0.0089845 0.0014321 0.98635 0.99132 3.0941e-006 1.2376e-005 0.15455 0.82618 0.86573 0.0014211 0.93994 0.45724 0.0019137 0.42287 1.7571 1.7553 16.0124 144.9478 0.00024275 -85.457 0.40894
5.513 0.98809 5.4883e-005 3.8183 0.01197 7.203e-005 0.001162 0.23231 0.0006593 0.23296 0.21493 0 0.032329 0.0389 0 1.3158 0.44483 0.13494 0.016685 9.7771 0.10395 0.00013205 0.78618 0.0080794 0.0089851 0.0014318 0.98635 0.99132 3.0933e-006 1.2373e-005 0.15456 0.82667 0.86598 0.0014209 0.94031 0.45743 0.0019134 0.42288 1.7582 1.7564 16.0124 144.9478 0.00024236 -85.4584 0.40994
5.514 0.98809 5.4883e-005 3.8183 0.01197 7.2043e-005 0.001162 0.23231 0.0006593 0.23296 0.21494 0 0.032329 0.0389 0 1.3159 0.44487 0.13495 0.016687 9.7792 0.10396 0.00013207 0.78617 0.0080799 0.0089857 0.0014314 0.98636 0.99132 3.0925e-006 1.237e-005 0.15456 0.82716 0.86623 0.0014208 0.94067 0.45762 0.0019132 0.42289 1.7593 1.7575 16.0124 144.9478 0.00024198 -85.4599 0.41094
5.515 0.98809 5.4883e-005 3.8183 0.01197 7.2056e-005 0.001162 0.23231 0.0006593 0.23296 0.21494 0 0.032328 0.0389 0 1.316 0.44492 0.13497 0.016688 9.7812 0.10397 0.00013208 0.78616 0.0080805 0.0089864 0.0014311 0.98636 0.99133 3.0917e-006 1.2367e-005 0.15457 0.82765 0.86648 0.0014206 0.94103 0.45781 0.0019129 0.42291 1.7604 1.7586 16.0124 144.9479 0.00024159 -85.4613 0.41194
5.516 0.98809 5.4883e-005 3.8183 0.01197 7.2069e-005 0.001162 0.23231 0.0006593 0.23297 0.21494 0 0.032328 0.0389 0 1.3161 0.44497 0.13498 0.01669 9.7833 0.10398 0.00013209 0.78615 0.0080811 0.008987 0.0014307 0.98637 0.99133 3.0909e-006 1.2364e-005 0.15457 0.82814 0.86673 0.0014204 0.94139 0.45799 0.0019127 0.42292 1.7615 1.7597 16.0124 144.9479 0.00024121 -85.4627 0.41294
5.517 0.98809 5.4883e-005 3.8183 0.01197 7.2082e-005 0.001162 0.23231 0.0006593 0.23297 0.21494 0 0.032328 0.0389 0 1.3162 0.44501 0.135 0.016691 9.7854 0.10399 0.00013211 0.78615 0.0080817 0.0089876 0.0014304 0.98637 0.99133 3.0902e-006 1.2361e-005 0.15458 0.82862 0.86698 0.0014202 0.94175 0.45818 0.0019125 0.42293 1.7626 1.7608 16.0123 144.9479 0.00024082 -85.4642 0.41394
5.518 0.98809 5.4883e-005 3.8183 0.01197 7.2095e-005 0.001162 0.23231 0.0006593 0.23297 0.21494 0 0.032328 0.0389 0 1.3163 0.44506 0.13501 0.016693 9.7875 0.10399 0.00013212 0.78614 0.0080823 0.0089882 0.0014301 0.98638 0.99133 3.0894e-006 1.2358e-005 0.15458 0.8291 0.86722 0.0014201 0.9421 0.45837 0.0019123 0.42295 1.7637 1.7619 16.0123 144.9479 0.00024044 -85.4656 0.41494
5.519 0.98809 5.4883e-005 3.8183 0.01197 7.2108e-005 0.001162 0.23232 0.0006593 0.23297 0.21494 0 0.032328 0.0389 0 1.3164 0.44511 0.13503 0.016694 9.7896 0.104 0.00013213 0.78613 0.0080828 0.0089889 0.0014297 0.98638 0.99134 3.0886e-006 1.2354e-005 0.15459 0.82959 0.86747 0.0014199 0.94245 0.45856 0.001912 0.42296 1.7647 1.763 16.0123 144.9479 0.00024006 -85.467 0.41594
5.52 0.98809 5.4883e-005 3.8183 0.01197 7.2121e-005 0.0011621 0.23232 0.0006593 0.23297 0.21495 0 0.032328 0.0389 0 1.3165 0.44515 0.13505 0.016695 9.7917 0.10401 0.00013214 0.78612 0.0080834 0.0089895 0.0014294 0.98638 0.99134 3.0879e-006 1.2351e-005 0.15459 0.83007 0.86771 0.0014197 0.9428 0.45874 0.0019118 0.42297 1.7658 1.7641 16.0123 144.948 0.00023969 -85.4683 0.41694
5.521 0.98809 5.4883e-005 3.8183 0.01197 7.2134e-005 0.0011621 0.23232 0.0006593 0.23297 0.21495 0 0.032328 0.0389 0 1.3166 0.4452 0.13506 0.016697 9.7938 0.10402 0.00013216 0.78611 0.008084 0.0089901 0.0014291 0.98639 0.99134 3.0871e-006 1.2348e-005 0.1546 0.83054 0.86796 0.0014195 0.94315 0.45893 0.0019116 0.42299 1.7669 1.7652 16.0123 144.948 0.00023931 -85.4697 0.41794
5.522 0.98809 5.4883e-005 3.8183 0.01197 7.2147e-005 0.0011621 0.23232 0.0006593 0.23298 0.21495 0 0.032328 0.0389 0 1.3167 0.44524 0.13508 0.016698 9.7959 0.10403 0.00013217 0.7861 0.0080846 0.0089907 0.0014287 0.98639 0.99135 3.0864e-006 1.2345e-005 0.1546 0.83102 0.8682 0.0014194 0.94349 0.45912 0.0019114 0.423 1.768 1.7662 16.0123 144.948 0.00023894 -85.4711 0.41894
5.523 0.98809 5.4883e-005 3.8183 0.01197 7.216e-005 0.0011621 0.23232 0.0006593 0.23298 0.21495 0 0.032328 0.0389 0 1.3168 0.44529 0.13509 0.0167 9.798 0.10404 0.00013218 0.78609 0.0080852 0.0089914 0.0014284 0.9864 0.99135 3.0856e-006 1.2342e-005 0.1546 0.8315 0.86844 0.0014192 0.94384 0.45931 0.0019111 0.42301 1.769 1.7673 16.0123 144.948 0.00023857 -85.4724 0.41994
5.524 0.98809 5.4883e-005 3.8183 0.01197 7.2173e-005 0.0011621 0.23233 0.0006593 0.23298 0.21495 0 0.032328 0.0389 0 1.3169 0.44534 0.13511 0.016701 9.8 0.10405 0.00013219 0.78608 0.0080857 0.008992 0.0014281 0.9864 0.99135 3.0849e-006 1.234e-005 0.15461 0.83197 0.86868 0.001419 0.94418 0.45949 0.0019109 0.42303 1.7701 1.7684 16.0123 144.948 0.00023819 -85.4738 0.42094
5.525 0.98809 5.4883e-005 3.8183 0.01197 7.2186e-005 0.0011621 0.23233 0.0006593 0.23298 0.21495 0 0.032328 0.0389 0 1.317 0.44538 0.13512 0.016703 9.8021 0.10406 0.00013221 0.78608 0.0080863 0.0089926 0.0014278 0.98641 0.99135 3.0842e-006 1.2337e-005 0.15461 0.83244 0.86892 0.0014189 0.94452 0.45968 0.0019107 0.42304 1.7712 1.7694 16.0123 144.9481 0.00023782 -85.4751 0.42194
5.526 0.98809 5.4882e-005 3.8183 0.01197 7.2198e-005 0.0011621 0.23233 0.0006593 0.23298 0.21496 0 0.032328 0.0389 0 1.3171 0.44543 0.13514 0.016704 9.8042 0.10407 0.00013222 0.78607 0.0080869 0.0089932 0.0014275 0.98641 0.99136 3.0834e-006 1.2334e-005 0.15462 0.83292 0.86916 0.0014187 0.94485 0.45987 0.0019105 0.42305 1.7722 1.7705 16.0123 144.9481 0.00023746 -85.4765 0.42294
5.527 0.98809 5.4882e-005 3.8183 0.01197 7.2211e-005 0.0011621 0.23233 0.0006593 0.23298 0.21496 0 0.032327 0.0389 0 1.3172 0.44548 0.13515 0.016706 9.8063 0.10407 0.00013223 0.78606 0.0080875 0.0089939 0.0014271 0.98641 0.99136 3.0827e-006 1.2331e-005 0.15462 0.83339 0.8694 0.0014185 0.94519 0.46005 0.0019103 0.42307 1.7733 1.7716 16.0123 144.9481 0.00023709 -85.4778 0.42394
5.528 0.98809 5.4882e-005 3.8183 0.01197 7.2224e-005 0.0011621 0.23233 0.0006593 0.23299 0.21496 0 0.032327 0.0389 0 1.3173 0.44552 0.13517 0.016707 9.8084 0.10408 0.00013224 0.78605 0.0080881 0.0089945 0.0014268 0.98642 0.99136 3.082e-006 1.2328e-005 0.15463 0.83385 0.86963 0.0014184 0.94552 0.46024 0.0019101 0.42308 1.7743 1.7726 16.0123 144.9481 0.00023673 -85.4791 0.42494
5.529 0.98809 5.4882e-005 3.8183 0.01197 7.2237e-005 0.0011621 0.23233 0.0006593 0.23299 0.21496 0 0.032327 0.0389 0 1.3173 0.44557 0.13518 0.016708 9.8105 0.10409 0.00013226 0.78604 0.0080886 0.0089951 0.0014265 0.98642 0.99136 3.0813e-006 1.2325e-005 0.15463 0.83432 0.86987 0.0014182 0.94585 0.46043 0.0019098 0.42309 1.7754 1.7737 16.0123 144.9481 0.00023636 -85.4804 0.42594
5.53 0.98809 5.4882e-005 3.8183 0.01197 7.225e-005 0.0011621 0.23234 0.0006593 0.23299 0.21496 0 0.032327 0.0389 0 1.3174 0.44562 0.1352 0.01671 9.8126 0.1041 0.00013227 0.78603 0.0080892 0.0089957 0.0014262 0.98643 0.99137 3.0806e-006 1.2322e-005 0.15464 0.83479 0.8701 0.0014181 0.94618 0.46062 0.0019096 0.42311 1.7764 1.7747 16.0123 144.9481 0.000236 -85.4817 0.42694
5.531 0.98809 5.4882e-005 3.8183 0.01197 7.2263e-005 0.0011621 0.23234 0.0006593 0.23299 0.21496 0 0.032327 0.0389 0 1.3175 0.44566 0.13521 0.016711 9.8147 0.10411 0.00013228 0.78602 0.0080898 0.0089964 0.0014259 0.98643 0.99137 3.0799e-006 1.232e-005 0.15464 0.83525 0.87033 0.0014179 0.9465 0.4608 0.0019094 0.42312 1.7775 1.7758 16.0123 144.9482 0.00023564 -85.483 0.42794
5.532 0.98809 5.4882e-005 3.8183 0.01197 7.2276e-005 0.0011621 0.23234 0.0006593 0.23299 0.21497 0 0.032327 0.0389 0 1.3176 0.44571 0.13523 0.016713 9.8168 0.10412 0.0001323 0.78601 0.0080904 0.008997 0.0014256 0.98643 0.99137 3.0792e-006 1.2317e-005 0.15465 0.83571 0.87057 0.0014178 0.94683 0.46099 0.0019092 0.42313 1.7785 1.7768 16.0123 144.9482 0.00023528 -85.4842 0.42894
5.533 0.98809 5.4882e-005 3.8183 0.01197 7.2289e-005 0.0011621 0.23234 0.0006593 0.233 0.21497 0 0.032327 0.0389 0 1.3177 0.44576 0.13524 0.016714 9.8189 0.10413 0.00013231 0.78601 0.0080909 0.0089976 0.0014253 0.98644 0.99138 3.0785e-006 1.2314e-005 0.15465 0.83617 0.8708 0.0014176 0.94715 0.46118 0.001909 0.42315 1.7795 1.7779 16.0123 144.9482 0.00023492 -85.4855 0.42994
5.534 0.98809 5.4882e-005 3.8183 0.01197 7.2302e-005 0.0011621 0.23234 0.0006593 0.233 0.21497 0 0.032327 0.0389 0 1.3178 0.4458 0.13526 0.016716 9.821 0.10414 0.00013232 0.786 0.0080915 0.0089982 0.001425 0.98644 0.99138 3.0778e-006 1.2311e-005 0.15465 0.83663 0.87103 0.0014174 0.94747 0.46136 0.0019088 0.42316 1.7806 1.7789 16.0123 144.9482 0.00023457 -85.4867 0.43094
5.535 0.98809 5.4882e-005 3.8183 0.01197 7.2315e-005 0.0011621 0.23234 0.0006593 0.233 0.21497 0 0.032327 0.0389 0 1.3179 0.44585 0.13527 0.016717 9.8231 0.10414 0.00013233 0.78599 0.0080921 0.0089989 0.0014247 0.98645 0.99138 3.0771e-006 1.2309e-005 0.15466 0.83709 0.87126 0.0014173 0.94779 0.46155 0.0019086 0.42317 1.7816 1.78 16.0123 144.9482 0.00023421 -85.488 0.43194
5.536 0.98809 5.4882e-005 3.8183 0.01197 7.2328e-005 0.0011621 0.23235 0.0006593 0.233 0.21497 0 0.032327 0.0389 0 1.318 0.44589 0.13529 0.016718 9.8252 0.10415 0.00013235 0.78598 0.0080927 0.0089995 0.0014244 0.98645 0.99138 3.0765e-006 1.2306e-005 0.15466 0.83755 0.87149 0.0014171 0.9481 0.46174 0.0019084 0.42319 1.7826 1.781 16.0123 144.9483 0.00023386 -85.4892 0.43294
5.537 0.98809 5.4882e-005 3.8183 0.01197 7.2341e-005 0.0011621 0.23235 0.0006593 0.233 0.21497 0 0.032327 0.0389 0 1.3181 0.44594 0.13531 0.01672 9.8273 0.10416 0.00013236 0.78597 0.0080933 0.0090001 0.0014241 0.98645 0.99139 3.0758e-006 1.2303e-005 0.15467 0.83801 0.87171 0.001417 0.94842 0.46192 0.0019082 0.4232 1.7837 1.782 16.0123 144.9483 0.00023351 -85.4905 0.43394
5.538 0.98809 5.4882e-005 3.8183 0.01197 7.2354e-005 0.0011621 0.23235 0.0006593 0.233 0.21498 0 0.032326 0.0389 0 1.3182 0.44599 0.13532 0.016721 9.8294 0.10417 0.00013237 0.78596 0.0080938 0.0090007 0.0014238 0.98646 0.99139 3.0751e-006 1.2301e-005 0.15467 0.83846 0.87194 0.0014168 0.94873 0.46211 0.001908 0.42321 1.7847 1.7831 16.0123 144.9483 0.00023316 -85.4917 0.43494
5.539 0.98809 5.4882e-005 3.8183 0.01197 7.2367e-005 0.0011621 0.23235 0.0006593 0.23301 0.21498 0 0.032326 0.0389 0 1.3183 0.44603 0.13534 0.016723 9.8315 0.10418 0.00013238 0.78595 0.0080944 0.0090014 0.0014236 0.98646 0.99139 3.0745e-006 1.2298e-005 0.15468 0.83891 0.87217 0.0014167 0.94904 0.4623 0.0019078 0.42323 1.7857 1.7841 16.0123 144.9483 0.00023281 -85.4929 0.43594
5.54 0.98809 5.4881e-005 3.8183 0.01197 7.238e-005 0.0011621 0.23235 0.0006593 0.23301 0.21498 0 0.032326 0.0389 0 1.3184 0.44608 0.13535 0.016724 9.8335 0.10419 0.0001324 0.78594 0.008095 0.009002 0.0014233 0.98646 0.99139 3.0738e-006 1.2295e-005 0.15468 0.83936 0.87239 0.0014165 0.94935 0.46248 0.0019076 0.42324 1.7867 1.7851 16.0123 144.9483 0.00023246 -85.4941 0.43694
5.541 0.98809 5.4881e-005 3.8183 0.011969 7.2393e-005 0.0011621 0.23235 0.0006593 0.23301 0.21498 0 0.032326 0.0389 0 1.3185 0.44613 0.13537 0.016726 9.8356 0.1042 0.00013241 0.78593 0.0080956 0.0090026 0.001423 0.98647 0.9914 3.0732e-006 1.2293e-005 0.15469 0.83981 0.87261 0.0014164 0.94966 0.46267 0.0019074 0.42325 1.7878 1.7861 16.0123 144.9484 0.00023212 -85.4953 0.43794
5.542 0.98809 5.4881e-005 3.8183 0.011969 7.2406e-005 0.0011621 0.23236 0.0006593 0.23301 0.21498 0 0.032326 0.0389 0 1.3186 0.44617 0.13538 0.016727 9.8377 0.10421 0.00013242 0.78593 0.0080961 0.0090032 0.0014227 0.98647 0.9914 3.0725e-006 1.229e-005 0.15469 0.84026 0.87284 0.0014162 0.94996 0.46285 0.0019072 0.42327 1.7888 1.7871 16.0123 144.9484 0.00023178 -85.4965 0.43894
5.543 0.98809 5.4881e-005 3.8183 0.011969 7.2418e-005 0.0011621 0.23236 0.0006593 0.23301 0.21498 0 0.032326 0.0389 0 1.3187 0.44622 0.1354 0.016729 9.8398 0.10422 0.00013243 0.78592 0.0080967 0.0090038 0.0014224 0.98648 0.9914 3.0719e-006 1.2288e-005 0.1547 0.84071 0.87306 0.0014161 0.95026 0.46304 0.001907 0.42328 1.7898 1.7882 16.0123 144.9484 0.00023143 -85.4977 0.43994
5.544 0.98809 5.4881e-005 3.8183 0.011969 7.2431e-005 0.0011621 0.23236 0.0006593 0.23301 0.21499 0 0.032326 0.0389 0 1.3188 0.44627 0.13541 0.01673 9.8419 0.10422 0.00013245 0.78591 0.0080973 0.0090045 0.0014221 0.98648 0.9914 3.0713e-006 1.2285e-005 0.1547 0.84115 0.87328 0.0014159 0.95056 0.46323 0.0019069 0.42329 1.7908 1.7892 16.0123 144.9484 0.00023109 -85.4988 0.44094
5.545 0.98809 5.4881e-005 3.8183 0.011969 7.2444e-005 0.0011621 0.23236 0.0006593 0.23302 0.21499 0 0.032326 0.0389 0 1.3189 0.44631 0.13543 0.016731 9.844 0.10423 0.00013246 0.7859 0.0080979 0.0090051 0.0014219 0.98648 0.9914 3.0706e-006 1.2282e-005 0.1547 0.8416 0.8735 0.0014158 0.95086 0.46341 0.0019067 0.42331 1.7918 1.7902 16.0123 144.9484 0.00023075 -85.5 0.44194
5.546 0.98809 5.4881e-005 3.8183 0.011969 7.2457e-005 0.0011621 0.23236 0.0006593 0.23302 0.21499 0 0.032326 0.0389 0 1.319 0.44636 0.13544 0.016733 9.8461 0.10424 0.00013247 0.78589 0.0080985 0.0090057 0.0014216 0.98649 0.99141 3.07e-006 1.228e-005 0.15471 0.84204 0.87372 0.0014156 0.95116 0.4636 0.0019065 0.42332 1.7928 1.7912 16.0123 144.9485 0.00023041 -85.5011 0.44294
5.547 0.98809 5.4881e-005 3.8183 0.011969 7.247e-005 0.0011621 0.23236 0.0006593 0.23302 0.21499 0 0.032326 0.0389 0 1.319 0.44641 0.13546 0.016734 9.8482 0.10425 0.00013249 0.78588 0.008099 0.0090063 0.0014213 0.98649 0.99141 3.0694e-006 1.2277e-005 0.15471 0.84248 0.87394 0.0014155 0.95145 0.46379 0.0019063 0.42333 1.7938 1.7922 16.0123 144.9485 0.00023008 -85.5023 0.44394
5.548 0.98809 5.4881e-005 3.8183 0.011969 7.2483e-005 0.0011621 0.23237 0.0006593 0.23302 0.21499 0 0.032326 0.0389 0 1.3191 0.44645 0.13547 0.016736 9.8503 0.10426 0.0001325 0.78587 0.0080996 0.009007 0.0014211 0.98649 0.99141 3.0688e-006 1.2275e-005 0.15472 0.84292 0.87415 0.0014154 0.95175 0.46397 0.0019061 0.42335 1.7948 1.7932 16.0123 144.9485 0.00022974 -85.5034 0.44494
5.549 0.98809 5.4881e-005 3.8183 0.011969 7.2496e-005 0.0011621 0.23237 0.0006593 0.23302 0.21499 0 0.032326 0.0389 0 1.3192 0.4465 0.13549 0.016737 9.8524 0.10427 0.00013251 0.78586 0.0081002 0.0090076 0.0014208 0.9865 0.99141 3.0681e-006 1.2273e-005 0.15472 0.84336 0.87437 0.0014152 0.95204 0.46416 0.0019059 0.42336 1.7958 1.7942 16.0122 144.9485 0.00022941 -85.5046 0.44594
5.55 0.98809 5.4881e-005 3.8183 0.011969 7.2509e-005 0.0011621 0.23237 0.0006593 0.23302 0.215 0 0.032325 0.0389 0 1.3193 0.44654 0.1355 0.016739 9.8545 0.10428 0.00013252 0.78586 0.0081008 0.0090082 0.0014205 0.9865 0.99142 3.0675e-006 1.227e-005 0.15473 0.8438 0.87458 0.0014151 0.95233 0.46434 0.0019057 0.42337 1.7968 1.7952 16.0122 144.9485 0.00022907 -85.5057 0.44694
5.551 0.98809 5.4881e-005 3.8183 0.011969 7.2522e-005 0.0011622 0.23237 0.0006593 0.23303 0.215 0 0.032325 0.0389 0 1.3194 0.44659 0.13552 0.01674 9.8566 0.10429 0.00013254 0.78585 0.0081013 0.0090088 0.0014203 0.9865 0.99142 3.0669e-006 1.2268e-005 0.15473 0.84424 0.8748 0.0014149 0.95261 0.46453 0.0019056 0.42339 1.7978 1.7962 16.0122 144.9486 0.00022874 -85.5068 0.44794
5.552 0.98809 5.4881e-005 3.8183 0.011969 7.2535e-005 0.0011622 0.23237 0.0006593 0.23303 0.215 0 0.032325 0.0389 0 1.3195 0.44664 0.13553 0.016741 9.8587 0.10429 0.00013255 0.78584 0.0081019 0.0090094 0.00142 0.98651 0.99142 3.0663e-006 1.2265e-005 0.15474 0.84467 0.87501 0.0014148 0.9529 0.46471 0.0019054 0.4234 1.7988 1.7972 16.0122 144.9486 0.00022841 -85.5079 0.44894
5.553 0.98809 5.488e-005 3.8183 0.011969 7.2548e-005 0.0011622 0.23237 0.0006593 0.23303 0.215 0 0.032325 0.0389 0 1.3196 0.44668 0.13555 0.016743 9.8608 0.1043 0.00013256 0.78583 0.0081025 0.0090101 0.0014197 0.98651 0.99142 3.0657e-006 1.2263e-005 0.15474 0.8451 0.87522 0.0014147 0.95318 0.4649 0.0019052 0.42341 1.7997 1.7982 16.0122 144.9486 0.00022808 -85.509 0.44994
5.554 0.98809 5.488e-005 3.8183 0.011969 7.2561e-005 0.0011622 0.23238 0.0006593 0.23303 0.215 0 0.032325 0.0389 0 1.3197 0.44673 0.13556 0.016744 9.8629 0.10431 0.00013257 0.78582 0.0081031 0.0090107 0.0014195 0.98651 0.99143 3.0651e-006 1.2261e-005 0.15475 0.84554 0.87544 0.0014145 0.95347 0.46509 0.001905 0.42343 1.8007 1.7992 16.0122 144.9486 0.00022776 -85.5101 0.45094
5.555 0.98809 5.488e-005 3.8183 0.011969 7.2574e-005 0.0011622 0.23238 0.0006593 0.23303 0.215 0 0.032325 0.0389 0 1.3198 0.44678 0.13558 0.016746 9.865 0.10432 0.00013259 0.78581 0.0081036 0.0090113 0.0014192 0.98652 0.99143 3.0645e-006 1.2258e-005 0.15475 0.84597 0.87565 0.0014144 0.95375 0.46527 0.0019049 0.42344 1.8017 1.8001 16.0122 144.9486 0.00022743 -85.5112 0.45194
5.556 0.98809 5.488e-005 3.8183 0.011969 7.2587e-005 0.0011622 0.23238 0.0006593 0.23303 0.215 0 0.032325 0.0389 0 1.3199 0.44682 0.1356 0.016747 9.8671 0.10433 0.0001326 0.7858 0.0081042 0.0090119 0.001419 0.98652 0.99143 3.064e-006 1.2256e-005 0.15475 0.8464 0.87586 0.0014143 0.95403 0.46546 0.0019047 0.42346 1.8027 1.8011 16.0122 144.9486 0.0002271 -85.5122 0.45294
5.557 0.98809 5.488e-005 3.8183 0.011969 7.26e-005 0.0011622 0.23238 0.0006593 0.23304 0.21501 0 0.032325 0.0389 0 1.32 0.44687 0.13561 0.016749 9.8692 0.10434 0.00013261 0.78579 0.0081048 0.0090125 0.0014187 0.98652 0.99143 3.0634e-006 1.2254e-005 0.15476 0.84682 0.87607 0.0014141 0.9543 0.46564 0.0019045 0.42347 1.8037 1.8021 16.0122 144.9487 0.00022678 -85.5133 0.45394
5.558 0.98809 5.488e-005 3.8183 0.011969 7.2613e-005 0.0011622 0.23238 0.0006593 0.23304 0.21501 0 0.032325 0.0389 0 1.3201 0.44692 0.13563 0.01675 9.8713 0.10435 0.00013262 0.78579 0.0081054 0.0090132 0.0014185 0.98653 0.99143 3.0628e-006 1.2251e-005 0.15476 0.84725 0.87627 0.001414 0.95458 0.46583 0.0019043 0.42348 1.8046 1.8031 16.0122 144.9487 0.00022646 -85.5144 0.45494
5.559 0.98809 5.488e-005 3.8183 0.011969 7.2626e-005 0.0011622 0.23238 0.0006593 0.23304 0.21501 0 0.032325 0.0389 0 1.3202 0.44696 0.13564 0.016752 9.8734 0.10436 0.00013264 0.78578 0.008106 0.0090138 0.0014182 0.98653 0.99144 3.0623e-006 1.2249e-005 0.15477 0.84768 0.87648 0.0014138 0.95485 0.46601 0.0019042 0.4235 1.8056 1.8041 16.0122 144.9487 0.00022614 -85.5154 0.45594
5.56 0.98809 5.488e-005 3.8183 0.011969 7.2638e-005 0.0011622 0.23239 0.0006593 0.23304 0.21501 0 0.032325 0.0389 0 1.3203 0.44701 0.13566 0.016753 9.8755 0.10436 0.00013265 0.78577 0.0081065 0.0090144 0.001418 0.98653 0.99144 3.0617e-006 1.2247e-005 0.15477 0.8481 0.87669 0.0014137 0.95512 0.4662 0.001904 0.42351 1.8066 1.805 16.0122 144.9487 0.00022582 -85.5165 0.45694
5.561 0.98809 5.488e-005 3.8183 0.011969 7.2651e-005 0.0011622 0.23239 0.0006593 0.23304 0.21501 0 0.032325 0.0389 0 1.3204 0.44705 0.13567 0.016754 9.8777 0.10437 0.00013266 0.78576 0.0081071 0.009015 0.0014177 0.98654 0.99144 3.0611e-006 1.2244e-005 0.15478 0.84852 0.87689 0.0014135 0.95539 0.46638 0.0019038 0.42352 1.8075 1.806 16.0122 144.9487 0.0002255 -85.5175 0.45794
5.562 0.98809 5.488e-005 3.8183 0.011969 7.2664e-005 0.0011622 0.23239 0.0006593 0.23304 0.21501 0 0.032324 0.0389 0 1.3205 0.4471 0.13569 0.016756 9.8798 0.10438 0.00013267 0.78575 0.0081077 0.0090157 0.0014175 0.98654 0.99144 3.0606e-006 1.2242e-005 0.15478 0.84894 0.8771 0.0014134 0.95566 0.46657 0.0019037 0.42354 1.8085 1.807 16.0122 144.9488 0.00022518 -85.5185 0.45894
5.563 0.98809 5.488e-005 3.8183 0.011969 7.2677e-005 0.0011622 0.23239 0.0006593 0.23305 0.21502 0 0.032324 0.0389 0 1.3206 0.44715 0.1357 0.016757 9.8819 0.10439 0.00013269 0.78574 0.0081083 0.0090163 0.0014172 0.98654 0.99144 3.06e-006 1.224e-005 0.15479 0.84936 0.8773 0.0014134 0.95593 0.46675 0.0019035 0.42355 1.8094 1.8079 16.0122 144.9488 0.00022487 -85.5196 0.45994
5.564 0.98809 5.488e-005 3.8183 0.011969 7.269e-005 0.0011622 0.23239 0.0006593 0.23305 0.21502 0 0.032324 0.0389 0 1.3207 0.44719 0.13572 0.016759 9.884 0.1044 0.0001327 0.78573 0.0081088 0.0090169 0.001417 0.98655 0.99145 3.0594e-006 1.2238e-005 0.15479 0.84978 0.87751 0.0014133 0.95619 0.46694 0.0019033 0.42356 1.8104 1.8089 16.0122 144.9488 0.00022455 -85.5206 0.46094
5.565 0.98809 5.488e-005 3.8183 0.011969 7.2703e-005 0.0011622 0.23239 0.0006593 0.23305 0.21502 0 0.032324 0.0389 0 1.3208 0.44724 0.13573 0.01676 9.8861 0.10441 0.00013271 0.78572 0.0081094 0.0090175 0.0014168 0.98655 0.99145 3.0589e-006 1.2236e-005 0.1548 0.8502 0.87771 0.0014132 0.95646 0.46712 0.0019032 0.42358 1.8113 1.8098 16.0122 144.9488 0.00022424 -85.5216 0.46194
5.566 0.98809 5.4879e-005 3.8183 0.011969 7.2716e-005 0.0011622 0.2324 0.0006593 0.23305 0.21502 0 0.032324 0.0389 0 1.3208 0.44729 0.13575 0.016762 9.8882 0.10442 0.00013273 0.78572 0.00811 0.0090181 0.0014165 0.98655 0.99145 3.0583e-006 1.2233e-005 0.1548 0.85062 0.87791 0.0014131 0.95672 0.46731 0.001903 0.42359 1.8123 1.8108 16.0121 144.9488 0.00022393 -85.5226 0.46294
5.567 0.98809 5.4879e-005 3.8183 0.011969 7.2729e-005 0.0011622 0.2324 0.0006593 0.23305 0.21502 0 0.032324 0.0389 0 1.3209 0.44733 0.13576 0.016763 9.8903 0.10443 0.00013274 0.78571 0.0081106 0.0090188 0.0014163 0.98656 0.99145 3.0578e-006 1.2231e-005 0.1548 0.85103 0.87811 0.0014129 0.95698 0.46749 0.0019029 0.4236 1.8132 1.8118 16.0121 144.9489 0.00022362 -85.5236 0.46394
5.568 0.98809 5.4879e-005 3.8183 0.011969 7.2742e-005 0.0011622 0.2324 0.0006593 0.23305 0.21502 0 0.032324 0.0389 0 1.321 0.44738 0.13578 0.016764 9.8924 0.10443 0.00013275 0.7857 0.0081111 0.0090194 0.001416 0.98656 0.99145 3.0573e-006 1.2229e-005 0.15481 0.85144 0.87831 0.0014127 0.95723 0.46768 0.0019027 0.42362 1.8142 1.8127 16.0121 144.9489 0.00022331 -85.5246 0.46494
5.569 0.98809 5.4879e-005 3.8183 0.011969 7.2755e-005 0.0011622 0.2324 0.0006593 0.23306 0.21503 0 0.032324 0.0389 0 1.3211 0.44743 0.13579 0.016766 9.8945 0.10444 0.00013276 0.78569 0.0081117 0.00902 0.0014158 0.98656 0.99146 3.0568e-006 1.2227e-005 0.15481 0.85186 0.87851 0.0014125 0.95749 0.46786 0.0019025 0.42363 1.8151 1.8136 16.0121 144.9489 0.000223 -85.5255 0.46594
5.57 0.98809 5.4879e-005 3.8183 0.011969 7.2768e-005 0.0011622 0.2324 0.0006593 0.23306 0.21503 0 0.032324 0.0389 0 1.3212 0.44747 0.13581 0.016767 9.8966 0.10445 0.00013278 0.78568 0.0081123 0.0090206 0.0014155 0.98656 0.99146 3.0563e-006 1.2225e-005 0.15482 0.85227 0.87871 0.0014123 0.95775 0.46805 0.0019024 0.42365 1.8161 1.8146 16.0121 144.9489 0.0002227 -85.5265 0.46694
5.571 0.98809 5.4879e-005 3.8183 0.011969 7.2781e-005 0.0011622 0.2324 0.0006593 0.23306 0.21503 0 0.032324 0.0389 0 1.3213 0.44752 0.13582 0.016769 9.8987 0.10446 0.00013279 0.78567 0.0081129 0.0090212 0.0014153 0.98657 0.99146 3.0558e-006 1.2223e-005 0.15482 0.85268 0.8789 0.0014121 0.958 0.46823 0.0019022 0.42366 1.817 1.8155 16.0121 144.9489 0.00022239 -85.5275 0.46794
5.572 0.98809 5.4879e-005 3.8183 0.011969 7.2794e-005 0.0011622 0.23241 0.0006593 0.23306 0.21503 0 0.032324 0.0389 0 1.3214 0.44757 0.13584 0.01677 9.9008 0.10447 0.0001328 0.78566 0.0081134 0.0090219 0.0014151 0.98657 0.99146 3.0552e-006 1.2221e-005 0.15483 0.85309 0.8791 0.001412 0.95825 0.46842 0.0019021 0.42367 1.8179 1.8165 16.0121 144.949 0.00022209 -85.5284 0.46894
5.573 0.98809 5.4879e-005 3.8183 0.011969 7.2807e-005 0.0011622 0.23241 0.0006593 0.23306 0.21503 0 0.032324 0.0389 0 1.3215 0.44761 0.13585 0.016772 9.9029 0.10448 0.00013281 0.78565 0.008114 0.0090225 0.0014149 0.98657 0.99146 3.0547e-006 1.2219e-005 0.15483 0.85349 0.8793 0.0014119 0.9585 0.4686 0.0019019 0.42369 1.8189 1.8174 16.0121 144.949 0.00022178 -85.5294 0.46994
5.574 0.98809 5.4879e-005 3.8183 0.011969 7.282e-005 0.0011622 0.23241 0.0006593 0.23306 0.21503 0 0.032323 0.0389 0 1.3216 0.44766 0.13587 0.016773 9.905 0.10449 0.00013283 0.78565 0.0081146 0.0090231 0.0014146 0.98658 0.99147 3.0542e-006 1.2217e-005 0.15484 0.8539 0.87949 0.0014118 0.95875 0.46879 0.0019018 0.4237 1.8198 1.8183 16.0121 144.949 0.00022148 -85.5303 0.47094
5.575 0.98809 5.4879e-005 3.8183 0.011969 7.2833e-005 0.0011622 0.23241 0.0006593 0.23307 0.21503 0 0.032323 0.0389 0 1.3217 0.4477 0.13588 0.016774 9.9071 0.1045 0.00013284 0.78564 0.0081152 0.0090237 0.0014144 0.98658 0.99147 3.0537e-006 1.2215e-005 0.15484 0.8543 0.87969 0.0014117 0.959 0.46897 0.0019016 0.42371 1.8207 1.8193 16.0121 144.949 0.00022118 -85.5313 0.47194
5.576 0.98809 5.4879e-005 3.8183 0.011969 7.2845e-005 0.0011622 0.23241 0.0006593 0.23307 0.21504 0 0.032323 0.0389 0 1.3218 0.44775 0.1359 0.016776 9.9092 0.1045 0.00013285 0.78563 0.0081157 0.0090243 0.0014142 0.98658 0.99147 3.0532e-006 1.2213e-005 0.15485 0.85471 0.87988 0.0014116 0.95924 0.46915 0.0019015 0.42373 1.8217 1.8202 16.0121 144.949 0.00022088 -85.5322 0.47294
5.577 0.98809 5.4879e-005 3.8183 0.011969 7.2858e-005 0.0011622 0.23241 0.0006593 0.23307 0.21504 0 0.032323 0.0389 0 1.3219 0.4478 0.13592 0.016777 9.9114 0.10451 0.00013286 0.78562 0.0081163 0.009025 0.001414 0.98658 0.99147 3.0527e-006 1.2211e-005 0.15485 0.85511 0.88007 0.0014115 0.95949 0.46934 0.0019013 0.42374 1.8226 1.8211 16.0121 144.9491 0.00022058 -85.5331 0.47394
5.578 0.98809 5.4879e-005 3.8183 0.011969 7.2871e-005 0.0011622 0.23242 0.0006593 0.23307 0.21504 0 0.032323 0.0389 0 1.322 0.44784 0.13593 0.016779 9.9135 0.10452 0.00013288 0.78561 0.0081169 0.0090256 0.0014138 0.98659 0.99147 3.0522e-006 1.2209e-005 0.15485 0.85551 0.88026 0.0014115 0.95973 0.46952 0.0019012 0.42375 1.8235 1.8221 16.012 144.9491 0.00022029 -85.5341 0.47494
5.579 0.98809 5.4878e-005 3.8183 0.011969 7.2884e-005 0.0011622 0.23242 0.0006593 0.23307 0.21504 0 0.032323 0.0389 0 1.3221 0.44789 0.13595 0.01678 9.9156 0.10453 0.00013289 0.7856 0.0081175 0.0090262 0.0014136 0.98659 0.99148 3.0517e-006 1.2207e-005 0.15486 0.85591 0.88045 0.0014114 0.95997 0.46971 0.001901 0.42377 1.8244 1.823 16.012 144.9491 0.00021999 -85.535 0.47594
5.58 0.98809 5.4878e-005 3.8183 0.011969 7.2897e-005 0.0011622 0.23242 0.0006593 0.23307 0.21504 0 0.032323 0.0389 0 1.3222 0.44794 0.13596 0.016782 9.9177 0.10454 0.0001329 0.78559 0.008118 0.0090268 0.0014134 0.98659 0.99148 3.0512e-006 1.2205e-005 0.15486 0.85631 0.88065 0.0014114 0.96021 0.46989 0.0019009 0.42378 1.8253 1.8239 16.012 144.9491 0.0002197 -85.5359 0.47694
5.581 0.98809 5.4878e-005 3.8183 0.011969 7.291e-005 0.0011623 0.23242 0.0006593 0.23308 0.21504 0 0.032323 0.0389 0 1.3223 0.44798 0.13598 0.016783 9.9198 0.10455 0.00013291 0.78558 0.0081186 0.0090274 0.0014132 0.9866 0.99148 3.0507e-006 1.2203e-005 0.15487 0.8567 0.88083 0.0014113 0.96045 0.47007 0.0019007 0.4238 1.8263 1.8248 16.012 144.9491 0.0002194 -85.5368 0.47794
5.582 0.98809 5.4878e-005 3.8183 0.011969 7.2923e-005 0.0011623 0.23242 0.0006593 0.23308 0.21505 0 0.032323 0.0389 0 1.3224 0.44803 0.13599 0.016784 9.9219 0.10456 0.00013293 0.78558 0.0081192 0.009028 0.001413 0.9866 0.99148 3.0502e-006 1.2201e-005 0.15487 0.8571 0.88102 0.0014112 0.96068 0.47026 0.0019006 0.42381 1.8272 1.8257 16.012 144.9492 0.00021911 -85.5377 0.47894
5.583 0.98809 5.4878e-005 3.8183 0.011969 7.2936e-005 0.0011623 0.23242 0.0006593 0.23308 0.21505 0 0.032323 0.0389 0 1.3225 0.44808 0.13601 0.016786 9.924 0.10457 0.00013294 0.78557 0.0081198 0.0090287 0.0014128 0.9866 0.99148 3.0497e-006 1.2199e-005 0.15488 0.85749 0.88121 0.0014111 0.96092 0.47044 0.0019004 0.42382 1.8281 1.8267 16.012 144.9492 0.00021882 -85.5386 0.47994
5.584 0.98809 5.4878e-005 3.8183 0.011969 7.2949e-005 0.0011623 0.23243 0.0006593 0.23308 0.21505 0 0.032323 0.0389 0 1.3225 0.44812 0.13602 0.016787 9.9261 0.10457 0.00013295 0.78556 0.0081203 0.0090293 0.0014126 0.9866 0.99148 3.0492e-006 1.2197e-005 0.15488 0.85789 0.8814 0.001411 0.96115 0.47063 0.0019003 0.42384 1.829 1.8276 16.012 144.9492 0.00021853 -85.5395 0.48094
5.585 0.98809 5.4878e-005 3.8183 0.011969 7.2962e-005 0.0011623 0.23243 0.0006593 0.23308 0.21505 0 0.032323 0.0389 0 1.3226 0.44817 0.13604 0.016789 9.9282 0.10458 0.00013297 0.78555 0.0081209 0.0090299 0.0014123 0.98661 0.99149 3.0488e-006 1.2195e-005 0.15489 0.85828 0.88158 0.0014109 0.96138 0.47081 0.0019001 0.42385 1.8299 1.8285 16.012 144.9492 0.00021824 -85.5403 0.48194
5.586 0.98809 5.4878e-005 3.8183 0.011969 7.2975e-005 0.0011623 0.23243 0.0006593 0.23308 0.21505 0 0.032322 0.0389 0 1.3227 0.44822 0.13605 0.01679 9.9304 0.10459 0.00013298 0.78554 0.0081215 0.0090305 0.0014121 0.98661 0.99149 3.0483e-006 1.2193e-005 0.15489 0.85867 0.88177 0.0014107 0.96161 0.47099 0.0019 0.42386 1.8308 1.8294 16.012 144.9492 0.00021796 -85.5412 0.48294
5.587 0.98809 5.4878e-005 3.8183 0.011969 7.2988e-005 0.0011623 0.23243 0.0006593 0.23309 0.21505 0 0.032322 0.0389 0 1.3228 0.44826 0.13607 0.016792 9.9325 0.1046 0.00013299 0.78553 0.0081221 0.0090311 0.0014119 0.98661 0.99149 3.0478e-006 1.2191e-005 0.15489 0.85906 0.88196 0.0014106 0.96184 0.47118 0.0018999 0.42388 1.8317 1.8303 16.012 144.9493 0.00021767 -85.5421 0.48394
5.588 0.98809 5.4878e-005 3.8183 0.011969 7.3001e-005 0.0011623 0.23243 0.0006593 0.23309 0.21506 0 0.032322 0.0389 0 1.3229 0.44831 0.13608 0.016793 9.9346 0.10461 0.000133 0.78552 0.0081226 0.0090318 0.0014117 0.98661 0.99149 3.0474e-006 1.2189e-005 0.1549 0.85945 0.88214 0.0014105 0.96207 0.47136 0.0018997 0.42389 1.8326 1.8312 16.012 144.9493 0.00021738 -85.5429 0.48494
5.589 0.98809 5.4878e-005 3.8183 0.011969 7.3014e-005 0.0011623 0.23243 0.0006593 0.23309 0.21506 0 0.032322 0.0389 0 1.323 0.44835 0.1361 0.016794 9.9367 0.10462 0.00013302 0.78551 0.0081232 0.0090324 0.0014115 0.98662 0.99149 3.0469e-006 1.2188e-005 0.1549 0.85984 0.88232 0.0014103 0.9623 0.47154 0.0018996 0.4239 1.8335 1.8321 16.0119 144.9493 0.0002171 -85.5438 0.48594
5.59 0.98809 5.4878e-005 3.8183 0.011969 7.3027e-005 0.0011623 0.23244 0.0006593 0.23309 0.21506 0 0.032322 0.0389 0 1.3231 0.4484 0.13611 0.016796 9.9388 0.10463 0.00013303 0.78551 0.0081238 0.009033 0.0014113 0.98662 0.99149 3.0465e-006 1.2186e-005 0.15491 0.86022 0.88251 0.0014102 0.96252 0.47173 0.0018995 0.42392 1.8344 1.833 16.0119 144.9493 0.00021682 -85.5446 0.48694
5.591 0.98809 5.4878e-005 3.8183 0.011969 7.304e-005 0.0011623 0.23244 0.0006593 0.23309 0.21506 0 0.032322 0.0389 0 1.3232 0.44845 0.13613 0.016797 9.9409 0.10464 0.00013304 0.7855 0.0081243 0.0090336 0.0014111 0.98662 0.9915 3.046e-006 1.2184e-005 0.15491 0.86061 0.88269 0.0014101 0.96274 0.47191 0.0018993 0.42393 1.8353 1.8339 16.0119 144.9493 0.00021654 -85.5455 0.48794
5.592 0.98809 5.4878e-005 3.8183 0.011969 7.3052e-005 0.0011623 0.23244 0.0006593 0.23309 0.21506 0 0.032322 0.0389 0 1.3233 0.44849 0.13614 0.016799 9.943 0.10464 0.00013305 0.78549 0.0081249 0.0090342 0.0014109 0.98663 0.9915 3.0456e-006 1.2182e-005 0.15492 0.86099 0.88287 0.0014099 0.96297 0.47209 0.0018992 0.42395 1.8361 1.8348 16.0119 144.9494 0.00021626 -85.5463 0.48894
5.593 0.98809 5.4877e-005 3.8183 0.011969 7.3065e-005 0.0011623 0.23244 0.0006593 0.2331 0.21506 0 0.032322 0.0389 0 1.3234 0.44854 0.13616 0.0168 9.9452 0.10465 0.00013307 0.78548 0.0081255 0.0090348 0.0014107 0.98663 0.9915 3.0451e-006 1.218e-005 0.15492 0.86137 0.88305 0.0014098 0.96319 0.47228 0.001899 0.42396 1.837 1.8356 16.0119 144.9494 0.00021598 -85.5471 0.48994
5.594 0.98809 5.4877e-005 3.8183 0.011969 7.3078e-005 0.0011623 0.23244 0.0006593 0.2331 0.21506 0 0.032322 0.0389 0 1.3235 0.44859 0.13617 0.016802 9.9473 0.10466 0.00013308 0.78547 0.0081261 0.0090355 0.0014105 0.98663 0.9915 3.0447e-006 1.2179e-005 0.15493 0.86176 0.88323 0.0014098 0.9634 0.47246 0.0018989 0.42397 1.8379 1.8365 16.0119 144.9494 0.0002157 -85.548 0.49094
5.595 0.98809 5.4877e-005 3.8183 0.011969 7.3091e-005 0.0011623 0.23244 0.0006593 0.2331 0.21507 0 0.032322 0.0389 0 1.3236 0.44863 0.13619 0.016803 9.9494 0.10467 0.00013309 0.78546 0.0081266 0.0090361 0.0014103 0.98663 0.9915 3.0442e-006 1.2177e-005 0.15493 0.86214 0.88341 0.0014097 0.96362 0.47264 0.0018988 0.42399 1.8388 1.8374 16.0119 144.9494 0.00021542 -85.5488 0.49194
5.596 0.98809 5.4877e-005 3.8183 0.011969 7.3104e-005 0.0011623 0.23245 0.0006593 0.2331 0.21507 0 0.032322 0.0389 0 1.3237 0.44868 0.1362 0.016804 9.9515 0.10468 0.0001331 0.78545 0.0081272 0.0090367 0.0014102 0.98664 0.9915 3.0438e-006 1.2175e-005 0.15494 0.86251 0.88359 0.0014096 0.96384 0.47283 0.0018987 0.424 1.8397 1.8383 16.0119 144.9494 0.00021514 -85.5496 0.49294
5.597 0.98809 5.4877e-005 3.8183 0.011969 7.3117e-005 0.0011623 0.23245 0.0006593 0.2331 0.21507 0 0.032322 0.0389 0 1.3238 0.44873 0.13622 0.016806 9.9536 0.10469 0.00013312 0.78544 0.0081278 0.0090373 0.00141 0.98664 0.99151 3.0434e-006 1.2173e-005 0.15494 0.86289 0.88376 0.0014095 0.96405 0.47301 0.0018985 0.42401 1.8405 1.8392 16.0119 144.9494 0.00021487 -85.5504 0.49394
5.598 0.98809 5.4877e-005 3.8183 0.011969 7.313e-005 0.0011623 0.23245 0.0006593 0.2331 0.21507 0 0.032322 0.0389 0 1.3239 0.44877 0.13624 0.016807 9.9557 0.1047 0.00013313 0.78544 0.0081284 0.0090379 0.0014098 0.98664 0.99151 3.0429e-006 1.2172e-005 0.15494 0.86327 0.88394 0.0014095 0.96427 0.47319 0.0018984 0.42403 1.8414 1.8401 16.0119 144.9495 0.0002146 -85.5512 0.49494
5.599 0.98809 5.4877e-005 3.8183 0.011969 7.3143e-005 0.0011623 0.23245 0.0006593 0.23311 0.21507 0 0.032321 0.0389 0 1.324 0.44882 0.13625 0.016809 9.9578 0.10471 0.00013314 0.78543 0.0081289 0.0090386 0.0014096 0.98664 0.99151 3.0425e-006 1.217e-005 0.15495 0.86364 0.88412 0.0014094 0.96448 0.47338 0.0018983 0.42404 1.8423 1.8409 16.0118 144.9495 0.00021432 -85.552 0.49594
5.6 0.98809 5.4877e-005 3.8183 0.011969 7.3156e-005 0.0011623 0.23245 0.0006593 0.23311 0.21507 0 0.032321 0.0389 0 1.3241 0.44886 0.13627 0.01681 9.96 0.10471 0.00013315 0.78542 0.0081295 0.0090392 0.0014094 0.98664 0.99151 3.0421e-006 1.2168e-005 0.15495 0.86402 0.88429 0.0014093 0.96469 0.47356 0.0018981 0.42406 1.8431 1.8418 16.0118 144.9495 0.00021405 -85.5528 0.49694
5.601 0.98809 5.4877e-005 3.8183 0.011969 7.3169e-005 0.0011623 0.23245 0.0006593 0.23311 0.21508 0 0.032321 0.0389 0 1.3242 0.44891 0.13628 0.016812 9.9621 0.10472 0.00013317 0.78541 0.0081301 0.0090398 0.0014092 0.98665 0.99151 3.0416e-006 1.2167e-005 0.15496 0.86439 0.88447 0.0014092 0.9649 0.47374 0.001898 0.42407 1.844 1.8427 16.0118 144.9495 0.00021378 -85.5536 0.49794
5.602 0.98809 5.4877e-005 3.8183 0.011968 7.3182e-005 0.0011623 0.23246 0.0006593 0.23311 0.21508 0 0.032321 0.0389 0 1.3242 0.44896 0.1363 0.016813 9.9642 0.10473 0.00013318 0.7854 0.0081306 0.0090404 0.001409 0.98665 0.99151 3.0412e-006 1.2165e-005 0.15496 0.86476 0.88464 0.0014092 0.96511 0.47393 0.0018979 0.42408 1.8449 1.8435 16.0118 144.9495 0.00021351 -85.5543 0.49894
5.603 0.98809 5.4877e-005 3.8183 0.011968 7.3195e-005 0.0011623 0.23246 0.0006593 0.23311 0.21508 0 0.032321 0.0389 0 1.3243 0.449 0.13631 0.016814 9.9663 0.10474 0.00013319 0.78539 0.0081312 0.009041 0.0014089 0.98665 0.99152 3.0408e-006 1.2163e-005 0.15497 0.86513 0.88481 0.0014091 0.96531 0.47411 0.0018978 0.4241 1.8457 1.8444 16.0118 144.9496 0.00021324 -85.5551 0.49994
5.604 0.98809 5.4877e-005 3.8183 0.011968 7.3208e-005 0.0011623 0.23246 0.0006593 0.23311 0.21508 0 0.032321 0.0389 0 1.3244 0.44905 0.13633 0.016816 9.9684 0.10475 0.0001332 0.78538 0.0081318 0.0090416 0.0014087 0.98665 0.99152 3.0404e-006 1.2162e-005 0.15497 0.8655 0.88499 0.0014089 0.96552 0.47429 0.0018976 0.42411 1.8466 1.8453 16.0118 144.9496 0.00021298 -85.5559 0.50094
5.605 0.98809 5.4877e-005 3.8183 0.011968 7.3221e-005 0.0011623 0.23246 0.0006593 0.23311 0.21508 0 0.032321 0.0389 0 1.3245 0.4491 0.13634 0.016817 9.9706 0.10476 0.00013322 0.78537 0.0081324 0.0090423 0.0014085 0.98666 0.99152 3.04e-006 1.216e-005 0.15498 0.86587 0.88516 0.0014088 0.96572 0.47447 0.0018975 0.42412 1.8475 1.8461 16.0118 144.9496 0.00021271 -85.5566 0.50194
5.606 0.98809 5.4876e-005 3.8183 0.011968 7.3234e-005 0.0011623 0.23246 0.0006593 0.23312 0.21508 0 0.032321 0.0389 0 1.3246 0.44914 0.13636 0.016819 9.9727 0.10477 0.00013323 0.78537 0.0081329 0.0090429 0.0014083 0.98666 0.99152 3.0396e-006 1.2158e-005 0.15498 0.86624 0.88533 0.0014087 0.96592 0.47466 0.0018974 0.42414 1.8483 1.847 16.0118 144.9496 0.00021244 -85.5574 0.50294
5.607 0.98809 5.4876e-005 3.8183 0.011968 7.3247e-005 0.0011623 0.23246 0.0006593 0.23312 0.21508 0 0.032321 0.0389 0 1.3247 0.44919 0.13637 0.01682 9.9748 0.10478 0.00013324 0.78536 0.0081335 0.0090435 0.0014081 0.98666 0.99152 3.0392e-006 1.2157e-005 0.15499 0.86661 0.8855 0.0014086 0.96613 0.47484 0.0018973 0.42415 1.8492 1.8478 16.0118 144.9496 0.00021218 -85.5582 0.50394
5.608 0.98809 5.4876e-005 3.8183 0.011968 7.3259e-005 0.0011623 0.23247 0.0006593 0.23312 0.21509 0 0.032321 0.0389 0 1.3248 0.44924 0.13639 0.016822 9.9769 0.10478 0.00013325 0.78535 0.0081341 0.0090441 0.001408 0.98666 0.99152 3.0388e-006 1.2155e-005 0.15499 0.86697 0.88567 0.0014085 0.96633 0.47502 0.0018971 0.42417 1.85 1.8487 16.0117 144.9497 0.00021192 -85.5589 0.50494
5.609 0.98809 5.4876e-005 3.8183 0.011968 7.3272e-005 0.0011623 0.23247 0.0006593 0.23312 0.21509 0 0.032321 0.0389 0 1.3249 0.44928 0.1364 0.016823 9.979 0.10479 0.00013327 0.78534 0.0081347 0.0090447 0.0014078 0.98667 0.99152 3.0384e-006 1.2153e-005 0.15499 0.86733 0.88584 0.0014084 0.96653 0.4752 0.001897 0.42418 1.8509 1.8495 16.0117 144.9497 0.00021165 -85.5596 0.50594
5.61 0.98809 5.4876e-005 3.8183 0.011968 7.3285e-005 0.0011623 0.23247 0.0006593 0.23312 0.21509 0 0.032321 0.0389 0 1.325 0.44933 0.13642 0.016824 9.9812 0.1048 0.00013328 0.78533 0.0081352 0.0090453 0.0014076 0.98667 0.99153 3.038e-006 1.2152e-005 0.155 0.8677 0.88601 0.0014083 0.96672 0.47539 0.0018969 0.42419 1.8517 1.8504 16.0117 144.9497 0.00021139 -85.5604 0.50694
5.611 0.98809 5.4876e-005 3.8183 0.011968 7.3298e-005 0.0011624 0.23247 0.0006593 0.23312 0.21509 0 0.03232 0.0389 0 1.3251 0.44938 0.13643 0.016826 9.9833 0.10481 0.00013329 0.78532 0.0081358 0.009046 0.0014074 0.98667 0.99153 3.0376e-006 1.215e-005 0.155 0.86806 0.88618 0.0014082 0.96692 0.47557 0.0018968 0.42421 1.8525 1.8512 16.0117 144.9497 0.00021113 -85.5611 0.50794
5.612 0.98809 5.4876e-005 3.8183 0.011968 7.3311e-005 0.0011624 0.23247 0.0006593 0.23313 0.21509 0 0.03232 0.0389 0 1.3252 0.44942 0.13645 0.016827 9.9854 0.10482 0.0001333 0.78531 0.0081364 0.0090466 0.0014073 0.98667 0.99153 3.0372e-006 1.2149e-005 0.15501 0.86842 0.88634 0.0014081 0.96711 0.47575 0.0018967 0.42422 1.8534 1.8521 16.0117 144.9497 0.00021087 -85.5618 0.50894
5.613 0.98809 5.4876e-005 3.8183 0.011968 7.3324e-005 0.0011624 0.23247 0.0006593 0.23313 0.21509 0 0.03232 0.0389 0 1.3253 0.44947 0.13646 0.016829 9.9875 0.10483 0.00013332 0.78531 0.0081369 0.0090472 0.0014071 0.98667 0.99153 3.0368e-006 1.2147e-005 0.15501 0.86878 0.88651 0.001408 0.96731 0.47593 0.0018966 0.42423 1.8542 1.8529 16.0117 144.9498 0.00021062 -85.5626 0.50994
5.614 0.98809 5.4876e-005 3.8183 0.011968 7.3337e-005 0.0011624 0.23247 0.0006593 0.23313 0.21509 0 0.03232 0.0389 0 1.3254 0.44951 0.13648 0.01683 9.9896 0.10484 0.00013333 0.7853 0.0081375 0.0090478 0.0014069 0.98668 0.99153 3.0364e-006 1.2146e-005 0.15502 0.86914 0.88668 0.0014079 0.9675 0.47611 0.0018964 0.42425 1.8551 1.8538 16.0117 144.9498 0.00021036 -85.5633 0.51094
5.615 0.98809 5.4876e-005 3.8183 0.011968 7.335e-005 0.0011624 0.23248 0.0006593 0.23313 0.2151 0 0.03232 0.0389 0 1.3255 0.44956 0.13649 0.016832 9.9918 0.10485 0.00013334 0.78529 0.0081381 0.0090484 0.0014068 0.98668 0.99153 3.036e-006 1.2144e-005 0.15502 0.86949 0.88684 0.0014078 0.96769 0.4763 0.0018963 0.42426 1.8559 1.8546 16.0117 144.9498 0.0002101 -85.564 0.51194
5.616 0.98809 5.4876e-005 3.8183 0.011968 7.3363e-005 0.0011624 0.23248 0.0006593 0.23313 0.2151 0 0.03232 0.0389 0 1.3256 0.44961 0.13651 0.016833 9.9939 0.10485 0.00013336 0.78528 0.0081387 0.009049 0.0014066 0.98668 0.99153 3.0357e-006 1.2143e-005 0.15503 0.86985 0.88701 0.0014078 0.96788 0.47648 0.0018962 0.42428 1.8567 1.8554 16.0116 144.9498 0.00020985 -85.5647 0.51294
5.617 0.98809 5.4876e-005 3.8183 0.011968 7.3376e-005 0.0011624 0.23248 0.0006593 0.23313 0.2151 0 0.03232 0.0389 0 1.3257 0.44965 0.13652 0.016834 9.996 0.10486 0.00013337 0.78527 0.0081392 0.0090496 0.0014064 0.98668 0.99154 3.0353e-006 1.2141e-005 0.15503 0.87021 0.88717 0.0014077 0.96807 0.47666 0.0018961 0.42429 1.8576 1.8563 16.0116 144.9498 0.00020959 -85.5654 0.51394
5.618 0.98809 5.4876e-005 3.8183 0.011968 7.3389e-005 0.0011624 0.23248 0.0006593 0.23314 0.2151 0 0.03232 0.0389 0 1.3258 0.4497 0.13654 0.016836 9.9981 0.10487 0.00013338 0.78526 0.0081398 0.0090503 0.0014063 0.98669 0.99154 3.0349e-006 1.214e-005 0.15503 0.87056 0.88733 0.0014076 0.96826 0.47684 0.001896 0.4243 1.8584 1.8571 16.0116 144.9499 0.00020934 -85.5661 0.51494
5.619 0.98809 5.4875e-005 3.8183 0.011968 7.3402e-005 0.0011624 0.23248 0.0006593 0.23314 0.2151 0 0.03232 0.0389 0 1.3259 0.44975 0.13655 0.016837 10.0003 0.10488 0.00013339 0.78525 0.0081404 0.0090509 0.0014061 0.98669 0.99154 3.0345e-006 1.2138e-005 0.15504 0.87091 0.8875 0.0014075 0.96845 0.47702 0.0018959 0.42432 1.8592 1.8579 16.0116 144.9499 0.00020909 -85.5668 0.51594
5.62 0.98809 5.4875e-005 3.8183 0.011968 7.3415e-005 0.0011624 0.23248 0.0006593 0.23314 0.2151 0 0.03232 0.0389 0 1.3259 0.44979 0.13657 0.016839 10.0024 0.10489 0.00013341 0.78524 0.0081409 0.0090515 0.001406 0.98669 0.99154 3.0342e-006 1.2137e-005 0.15504 0.87126 0.88766 0.0014075 0.96863 0.47721 0.0018958 0.42433 1.86 1.8588 16.0116 144.9499 0.00020884 -85.5675 0.51694
5.621 0.98809 5.4875e-005 3.8183 0.011968 7.3428e-005 0.0011624 0.23249 0.0006593 0.23314 0.21511 0 0.03232 0.0389 0 1.326 0.44984 0.13659 0.01684 10.0045 0.1049 0.00013342 0.78524 0.0081415 0.0090521 0.0014058 0.98669 0.99154 3.0338e-006 1.2135e-005 0.15505 0.87161 0.88782 0.0014074 0.96882 0.47739 0.0018957 0.42434 1.8609 1.8596 16.0116 144.9499 0.00020859 -85.5682 0.51794
5.622 0.98809 5.4875e-005 3.8183 0.011968 7.3441e-005 0.0011624 0.23249 0.0006593 0.23314 0.21511 0 0.03232 0.0389 0 1.3261 0.44989 0.1366 0.016842 10.0066 0.10491 0.00013343 0.78523 0.0081421 0.0090527 0.0014056 0.98669 0.99154 3.0334e-006 1.2134e-005 0.15505 0.87196 0.88798 0.0014073 0.969 0.47757 0.0018955 0.42436 1.8617 1.8604 16.0116 144.9499 0.00020834 -85.5688 0.51894
5.623 0.98809 5.4875e-005 3.8183 0.011968 7.3454e-005 0.0011624 0.23249 0.0006593 0.23314 0.21511 0 0.03232 0.0389 0 1.3262 0.44993 0.13662 0.016843 10.0088 0.10492 0.00013344 0.78522 0.0081426 0.0090533 0.0014055 0.9867 0.99154 3.0331e-006 1.2132e-005 0.15506 0.87231 0.88814 0.0014072 0.96918 0.47775 0.0018954 0.42437 1.8625 1.8612 16.0116 144.95 0.00020809 -85.5695 0.51994
5.624 0.98809 5.4875e-005 3.8183 0.011968 7.3466e-005 0.0011624 0.23249 0.0006593 0.23315 0.21511 0 0.032319 0.0389 0 1.3263 0.44998 0.13663 0.016844 10.0109 0.10492 0.00013346 0.78521 0.0081432 0.009054 0.0014053 0.9867 0.99154 3.0327e-006 1.2131e-005 0.15506 0.87266 0.8883 0.0014071 0.96936 0.47793 0.0018953 0.42439 1.8633 1.8621 16.0115 144.95 0.00020784 -85.5702 0.52094
5.625 0.98809 5.4875e-005 3.8183 0.011968 7.3479e-005 0.0011624 0.23249 0.0006593 0.23315 0.21511 0 0.032319 0.0389 0 1.3264 0.45002 0.13665 0.016846 10.013 0.10493 0.00013347 0.7852 0.0081438 0.0090546 0.0014052 0.9867 0.99155 3.0324e-006 1.2129e-005 0.15507 0.87301 0.88846 0.001407 0.96954 0.47811 0.0018952 0.4244 1.8641 1.8629 16.0115 144.95 0.0002076 -85.5708 0.52194
5.626 0.98809 5.4875e-005 3.8183 0.011968 7.3492e-005 0.0011624 0.23249 0.0006593 0.23315 0.21511 0 0.032319 0.0389 0 1.3265 0.45007 0.13666 0.016847 10.0151 0.10494 0.00013348 0.78519 0.0081444 0.0090552 0.001405 0.9867 0.99155 3.032e-006 1.2128e-005 0.15507 0.87335 0.88862 0.001407 0.96972 0.47829 0.0018951 0.42441 1.8649 1.8637 16.0115 144.95 0.00020735 -85.5715 0.52294
5.627 0.98809 5.4875e-005 3.8183 0.011968 7.3505e-005 0.0011624 0.2325 0.0006593 0.23315 0.21511 0 0.032319 0.0389 0 1.3266 0.45012 0.13668 0.016849 10.0173 0.10495 0.00013349 0.78518 0.0081449 0.0090558 0.0014049 0.9867 0.99155 3.0317e-006 1.2127e-005 0.15508 0.87369 0.88878 0.0014069 0.9699 0.47848 0.001895 0.42443 1.8658 1.8645 16.0115 144.95 0.00020711 -85.5722 0.52394
5.628 0.98809 5.4875e-005 3.8183 0.011968 7.3518e-005 0.0011624 0.2325 0.0006593 0.23315 0.21512 0 0.032319 0.0389 0 1.3267 0.45016 0.13669 0.01685 10.0194 0.10496 0.00013351 0.78517 0.0081455 0.0090564 0.0014047 0.98671 0.99155 3.0313e-006 1.2125e-005 0.15508 0.87404 0.88893 0.0014068 0.97007 0.47866 0.0018949 0.42444 1.8666 1.8653 16.0115 144.9501 0.00020687 -85.5728 0.52494
5.629 0.98809 5.4875e-005 3.8183 0.011968 7.3531e-005 0.0011624 0.2325 0.0006593 0.23315 0.21512 0 0.032319 0.0389 0 1.3268 0.45021 0.13671 0.016852 10.0215 0.10497 0.00013352 0.78517 0.0081461 0.009057 0.0014045 0.98671 0.99155 3.031e-006 1.2124e-005 0.15508 0.87438 0.88909 0.0014067 0.97025 0.47884 0.0018948 0.42445 1.8674 1.8661 16.0115 144.9501 0.00020662 -85.5735 0.52594
5.63 0.98809 5.4875e-005 3.8183 0.011968 7.3544e-005 0.0011624 0.2325 0.0006593 0.23315 0.21512 0 0.032319 0.0389 0 1.3269 0.45026 0.13672 0.016853 10.0236 0.10498 0.00013353 0.78516 0.0081466 0.0090576 0.0014044 0.98671 0.99155 3.0306e-006 1.2122e-005 0.15509 0.87472 0.88924 0.0014066 0.97042 0.47902 0.0018947 0.42447 1.8682 1.8669 16.0115 144.9501 0.00020638 -85.5741 0.52694
5.631 0.98809 5.4875e-005 3.8183 0.011968 7.3557e-005 0.0011624 0.2325 0.0006593 0.23316 0.21512 0 0.032319 0.0389 0 1.327 0.4503 0.13674 0.016854 10.0258 0.10499 0.00013354 0.78515 0.0081472 0.0090583 0.0014042 0.98671 0.99155 3.0303e-006 1.2121e-005 0.15509 0.87506 0.8894 0.0014065 0.97059 0.4792 0.0018946 0.42448 1.869 1.8677 16.0115 144.9501 0.00020614 -85.5747 0.52794
5.632 0.98809 5.4874e-005 3.8183 0.011968 7.357e-005 0.0011624 0.2325 0.0006593 0.23316 0.21512 0 0.032319 0.0389 0 1.3271 0.45035 0.13675 0.016856 10.0279 0.10499 0.00013356 0.78514 0.0081478 0.0090589 0.0014041 0.98671 0.99156 3.0299e-006 1.212e-005 0.1551 0.8754 0.88955 0.0014065 0.97077 0.47938 0.0018945 0.4245 1.8698 1.8685 16.0114 144.9501 0.0002059 -85.5754 0.52894
5.633 0.98809 5.4874e-005 3.8183 0.011968 7.3583e-005 0.0011624 0.2325 0.0006593 0.23316 0.21512 0 0.032319 0.0389 0 1.3272 0.4504 0.13677 0.016857 10.03 0.105 0.00013357 0.78513 0.0081483 0.0090595 0.001404 0.98672 0.99156 3.0296e-006 1.2118e-005 0.1551 0.87574 0.88971 0.0014064 0.97094 0.47956 0.0018944 0.42451 1.8706 1.8693 16.0114 144.9502 0.00020566 -85.576 0.52994
5.634 0.98809 5.4874e-005 3.8183 0.011968 7.3596e-005 0.0011624 0.23251 0.0006593 0.23316 0.21512 0 0.032319 0.0389 0 1.3273 0.45044 0.13678 0.016859 10.0322 0.10501 0.00013358 0.78512 0.0081489 0.0090601 0.0014038 0.98672 0.99156 3.0293e-006 1.2117e-005 0.15511 0.87607 0.88986 0.0014063 0.97111 0.47974 0.0018943 0.42452 1.8714 1.8701 16.0114 144.9502 0.00020543 -85.5766 0.53094
5.635 0.98809 5.4874e-005 3.8183 0.011968 7.3609e-005 0.0011624 0.23251 0.0006593 0.23316 0.21513 0 0.032319 0.0389 0 1.3274 0.45049 0.1368 0.01686 10.0343 0.10502 0.00013359 0.78511 0.0081495 0.0090607 0.0014037 0.98672 0.99156 3.0289e-006 1.2116e-005 0.15511 0.87641 0.89001 0.0014063 0.97127 0.47992 0.0018942 0.42454 1.8721 1.8709 16.0114 144.9502 0.00020519 -85.5772 0.53194
5.636 0.98809 5.4874e-005 3.8183 0.011968 7.3622e-005 0.0011624 0.23251 0.0006593 0.23316 0.21513 0 0.032318 0.0389 0 1.3275 0.45053 0.13681 0.016862 10.0364 0.10503 0.00013361 0.7851 0.0081501 0.0090613 0.0014035 0.98672 0.99156 3.0286e-006 1.2114e-005 0.15512 0.87674 0.89017 0.0014062 0.97144 0.4801 0.0018941 0.42455 1.8729 1.8717 16.0114 144.9502 0.00020495 -85.5779 0.53294
5.637 0.98809 5.4874e-005 3.8183 0.011968 7.3635e-005 0.0011624 0.23251 0.0006593 0.23317 0.21513 0 0.032318 0.0389 0 1.3275 0.45058 0.13683 0.016863 10.0386 0.10504 0.00013362 0.7851 0.0081506 0.0090619 0.0014034 0.98672 0.99156 3.0283e-006 1.2113e-005 0.15512 0.87708 0.89032 0.0014061 0.97161 0.48029 0.001894 0.42456 1.8737 1.8725 16.0114 144.9502 0.00020472 -85.5785 0.53394
5.638 0.98809 5.4874e-005 3.8183 0.011968 7.3648e-005 0.0011624 0.23251 0.0006593 0.23317 0.21513 0 0.032318 0.0389 0 1.3276 0.45063 0.13684 0.016864 10.0407 0.10505 0.00013363 0.78509 0.0081512 0.0090626 0.0014032 0.98672 0.99156 3.0279e-006 1.2112e-005 0.15512 0.87741 0.89047 0.001406 0.97177 0.48047 0.0018939 0.42458 1.8745 1.8733 16.0114 144.9503 0.00020449 -85.5791 0.53494
5.639 0.98809 5.4874e-005 3.8183 0.011968 7.366e-005 0.0011624 0.23251 0.0006593 0.23317 0.21513 0 0.032318 0.0389 0 1.3277 0.45067 0.13686 0.016866 10.0428 0.10505 0.00013364 0.78508 0.0081518 0.0090632 0.0014031 0.98673 0.99156 3.0276e-006 1.211e-005 0.15513 0.87774 0.89062 0.001406 0.97194 0.48065 0.0018938 0.42459 1.8753 1.8741 16.0113 144.9503 0.00020425 -85.5797 0.53594
5.64 0.98809 5.4874e-005 3.8183 0.011968 7.3673e-005 0.0011624 0.23252 0.0006593 0.23317 0.21513 0 0.032318 0.0389 0 1.3278 0.45072 0.13687 0.016867 10.0449 0.10506 0.00013366 0.78507 0.0081523 0.0090638 0.001403 0.98673 0.99156 3.0273e-006 1.2109e-005 0.15513 0.87807 0.89077 0.0014059 0.9721 0.48083 0.0018937 0.42461 1.8761 1.8749 16.0113 144.9503 0.00020402 -85.5803 0.53694
5.641 0.98809 5.4874e-005 3.8183 0.011968 7.3686e-005 0.0011624 0.23252 0.0006593 0.23317 0.21514 0 0.032318 0.0389 0 1.3279 0.45077 0.13689 0.016869 10.0471 0.10507 0.00013367 0.78506 0.0081529 0.0090644 0.0014028 0.98673 0.99157 3.027e-006 1.2108e-005 0.15514 0.8784 0.89092 0.0014058 0.97226 0.48101 0.0018936 0.42462 1.8769 1.8757 16.0113 144.9503 0.00020379 -85.5809 0.53794
5.642 0.98809 5.4874e-005 3.8183 0.011968 7.3699e-005 0.0011625 0.23252 0.0006593 0.23317 0.21514 0 0.032318 0.0389 0 1.328 0.45081 0.1369 0.01687 10.0492 0.10508 0.00013368 0.78505 0.0081535 0.009065 0.0014027 0.98673 0.99157 3.0267e-006 1.2107e-005 0.15514 0.87873 0.89107 0.0014057 0.97242 0.48119 0.0018935 0.42463 1.8776 1.8764 16.0113 144.9503 0.00020356 -85.5815 0.53894
5.643 0.98809 5.4874e-005 3.8183 0.011968 7.3712e-005 0.0011625 0.23252 0.0006593 0.23317 0.21514 0 0.032318 0.0389 0 1.3281 0.45086 0.13692 0.016871 10.0513 0.10509 0.00013369 0.78504 0.008154 0.0090656 0.0014025 0.98673 0.99157 3.0264e-006 1.2105e-005 0.15515 0.87906 0.89122 0.0014057 0.97258 0.48137 0.0018934 0.42465 1.8784 1.8772 16.0113 144.9504 0.00020333 -85.582 0.53994
5.644 0.98809 5.4874e-005 3.8183 0.011968 7.3725e-005 0.0011625 0.23252 0.0006593 0.23318 0.21514 0 0.032318 0.0389 0 1.3282 0.45091 0.13694 0.016873 10.0535 0.1051 0.00013371 0.78504 0.0081546 0.0090662 0.0014024 0.98674 0.99157 3.026e-006 1.2104e-005 0.15515 0.87938 0.89136 0.0014056 0.97274 0.48155 0.0018933 0.42466 1.8792 1.878 16.0113 144.9504 0.0002031 -85.5826 0.54094
5.645 0.98809 5.4873e-005 3.8183 0.011968 7.3738e-005 0.0011625 0.23252 0.0006593 0.23318 0.21514 0 0.032318 0.0389 0 1.3283 0.45095 0.13695 0.016874 10.0556 0.10511 0.00013372 0.78503 0.0081552 0.0090668 0.0014023 0.98674 0.99157 3.0257e-006 1.2103e-005 0.15516 0.87971 0.89151 0.0014055 0.9729 0.48173 0.0018932 0.42467 1.88 1.8788 16.0112 144.9504 0.00020287 -85.5832 0.54194
5.646 0.98809 5.4873e-005 3.8183 0.011968 7.3751e-005 0.0011625 0.23252 0.0006593 0.23318 0.21514 0 0.032318 0.0389 0 1.3284 0.451 0.13697 0.016876 10.0577 0.10512 0.00013373 0.78502 0.0081557 0.0090675 0.0014021 0.98674 0.99157 3.0254e-006 1.2102e-005 0.15516 0.88003 0.89166 0.0014054 0.97306 0.48191 0.0018931 0.42469 1.8807 1.8796 16.0112 144.9504 0.00020265 -85.5838 0.54294
5.647 0.98809 5.4873e-005 3.8183 0.011968 7.3764e-005 0.0011625 0.23253 0.0006593 0.23318 0.21514 0 0.032318 0.0389 0 1.3285 0.45105 0.13698 0.016877 10.0599 0.10512 0.00013374 0.78501 0.0081563 0.0090681 0.001402 0.98674 0.99157 3.0251e-006 1.21e-005 0.15516 0.88035 0.8918 0.0014054 0.97321 0.48209 0.0018931 0.4247 1.8815 1.8803 16.0112 144.9504 0.00020242 -85.5843 0.54394
5.648 0.98809 5.4873e-005 3.8183 0.011968 7.3777e-005 0.0011625 0.23253 0.0006593 0.23318 0.21515 0 0.032318 0.0389 0 1.3286 0.45109 0.137 0.016879 10.062 0.10513 0.00013376 0.785 0.0081569 0.0090687 0.0014019 0.98674 0.99157 3.0248e-006 1.2099e-005 0.15517 0.88068 0.89195 0.0014053 0.97337 0.48227 0.001893 0.42472 1.8823 1.8811 16.0112 144.9505 0.0002022 -85.5849 0.54494
5.649 0.98809 5.4873e-005 3.8183 0.011968 7.379e-005 0.0011625 0.23253 0.0006593 0.23318 0.21515 0 0.032317 0.0389 0 1.3287 0.45114 0.13701 0.01688 10.0641 0.10514 0.00013377 0.78499 0.0081575 0.0090693 0.0014017 0.98674 0.99158 3.0245e-006 1.2098e-005 0.15517 0.881 0.89209 0.0014052 0.97352 0.48245 0.0018929 0.42473 1.883 1.8819 16.0112 144.9505 0.00020197 -85.5855 0.54594
5.65 0.98809 5.4873e-005 3.8183 0.011968 7.3803e-005 0.0011625 0.23253 0.0006593 0.23319 0.21515 0 0.032317 0.0389 0 1.3288 0.45118 0.13703 0.016881 10.0663 0.10515 0.00013378 0.78498 0.008158 0.0090699 0.0014016 0.98675 0.99158 3.0242e-006 1.2097e-005 0.15518 0.88132 0.89224 0.0014052 0.97368 0.48263 0.0018928 0.42474 1.8838 1.8826 16.0112 144.9505 0.00020175 -85.586 0.54694
5.651 0.98809 5.4873e-005 3.8183 0.011968 7.3816e-005 0.0011625 0.23253 0.0006593 0.23319 0.21515 0 0.032317 0.0389 0 1.3289 0.45123 0.13704 0.016883 10.0684 0.10516 0.00013379 0.78497 0.0081586 0.0090705 0.0014015 0.98675 0.99158 3.0239e-006 1.2096e-005 0.15518 0.88164 0.89238 0.0014051 0.97383 0.48281 0.0018927 0.42476 1.8846 1.8834 16.0112 144.9505 0.00020153 -85.5866 0.54794
5.652 0.98809 5.4873e-005 3.8183 0.011968 7.3829e-005 0.0011625 0.23253 0.0006593 0.23319 0.21515 0 0.032317 0.0389 0 1.329 0.45128 0.13706 0.016884 10.0705 0.10517 0.00013381 0.78497 0.0081592 0.0090711 0.0014013 0.98675 0.99158 3.0236e-006 1.2094e-005 0.15519 0.88196 0.89252 0.001405 0.97398 0.48299 0.0018926 0.42477 1.8853 1.8842 16.0111 144.9505 0.0002013 -85.5871 0.54894
5.653 0.98809 5.4873e-005 3.8183 0.011968 7.3842e-005 0.0011625 0.23254 0.0006593 0.23319 0.21515 0 0.032317 0.0389 0 1.3291 0.45132 0.13707 0.016886 10.0727 0.10518 0.00013382 0.78496 0.0081597 0.0090717 0.0014012 0.98675 0.99158 3.0233e-006 1.2093e-005 0.15519 0.88227 0.89267 0.001405 0.97413 0.48317 0.0018925 0.42479 1.8861 1.8849 16.0111 144.9506 0.00020108 -85.5877 0.54994
5.654 0.98809 5.4873e-005 3.8183 0.011968 7.3854e-005 0.0011625 0.23254 0.0006593 0.23319 0.21515 0 0.032317 0.0389 0 1.3292 0.45137 0.13709 0.016887 10.0748 0.10519 0.00013383 0.78495 0.0081603 0.0090724 0.0014011 0.98675 0.99158 3.023e-006 1.2092e-005 0.1552 0.88259 0.89281 0.0014049 0.97428 0.48335 0.0018924 0.4248 1.8868 1.8857 16.0111 144.9506 0.00020086 -85.5882 0.55094
5.655 0.98809 5.4873e-005 3.8183 0.011968 7.3867e-005 0.0011625 0.23254 0.0006593 0.23319 0.21516 0 0.032317 0.0389 0 1.3292 0.45142 0.1371 0.016889 10.077 0.10519 0.00013384 0.78494 0.0081609 0.009073 0.001401 0.98675 0.99158 3.0228e-006 1.2091e-005 0.1552 0.8829 0.89295 0.0014048 0.97443 0.48353 0.0018923 0.42481 1.8876 1.8864 16.0111 144.9506 0.00020065 -85.5888 0.55194
5.656 0.98809 5.4873e-005 3.8183 0.011968 7.388e-005 0.0011625 0.23254 0.0006593 0.23319 0.21516 0 0.032317 0.0389 0 1.3293 0.45146 0.13712 0.01689 10.0791 0.1052 0.00013386 0.78493 0.0081614 0.0090736 0.0014008 0.98676 0.99158 3.0225e-006 1.209e-005 0.1552 0.88322 0.89309 0.0014047 0.97457 0.48371 0.0018923 0.42483 1.8883 1.8872 16.0111 144.9506 0.00020043 -85.5893 0.55294
5.657 0.98809 5.4873e-005 3.8183 0.011968 7.3893e-005 0.0011625 0.23254 0.0006593 0.2332 0.21516 0 0.032317 0.0389 0 1.3294 0.45151 0.13713 0.016891 10.0812 0.10521 0.00013387 0.78492 0.008162 0.0090742 0.0014007 0.98676 0.99158 3.0222e-006 1.2089e-005 0.15521 0.88353 0.89323 0.0014047 0.97472 0.48389 0.0018922 0.42484 1.8891 1.8879 16.0111 144.9506 0.00020021 -85.5898 0.55394
5.658 0.98809 5.4873e-005 3.8183 0.011968 7.3906e-005 0.0011625 0.23254 0.0006593 0.2332 0.21516 0 0.032317 0.0389 0 1.3295 0.45156 0.13715 0.016893 10.0834 0.10522 0.00013388 0.78491 0.0081626 0.0090748 0.0014006 0.98676 0.99158 3.0219e-006 1.2088e-005 0.15521 0.88384 0.89337 0.0014046 0.97486 0.48407 0.0018921 0.42485 1.8898 1.8887 16.011 144.9507 0.00019999 -85.5904 0.55494
5.659 0.98809 5.4872e-005 3.8183 0.011968 7.3919e-005 0.0011625 0.23254 0.0006593 0.2332 0.21516 0 0.032317 0.0389 0 1.3296 0.4516 0.13716 0.016894 10.0855 0.10523 0.00013389 0.78491 0.0081631 0.0090754 0.0014005 0.98676 0.99159 3.0216e-006 1.2086e-005 0.15522 0.88416 0.89351 0.0014045 0.97501 0.48425 0.001892 0.42487 1.8906 1.8894 16.011 144.9507 0.00019978 -85.5909 0.55594
5.66 0.98809 5.4872e-005 3.8183 0.011968 7.3932e-005 0.0011625 0.23255 0.0006593 0.2332 0.21516 0 0.032317 0.0389 0 1.3297 0.45165 0.13718 0.016896 10.0876 0.10524 0.00013391 0.7849 0.0081637 0.009076 0.0014003 0.98676 0.99159 3.0213e-006 1.2085e-005 0.15522 0.88447 0.89365 0.0014045 0.97515 0.48443 0.0018919 0.42488 1.8913 1.8902 16.011 144.9507 0.00019956 -85.5914 0.55694
5.661 0.98809 5.4872e-005 3.8183 0.011968 7.3945e-005 0.0011625 0.23255 0.0006593 0.2332 0.21516 0 0.032317 0.0389 0 1.3298 0.45169 0.13719 0.016897 10.0898 0.10525 0.00013392 0.78489 0.0081643 0.0090766 0.0014002 0.98676 0.99159 3.0211e-006 1.2084e-005 0.15523 0.88478 0.89378 0.0014044 0.97529 0.4846 0.0018918 0.4249 1.8921 1.8909 16.011 144.9507 0.00019935 -85.5919 0.55794
5.662 0.98809 5.4872e-005 3.8183 0.011968 7.3958e-005 0.0011625 0.23255 0.0006593 0.2332 0.21517 0 0.032316 0.0389 0 1.3299 0.45174 0.13721 0.016898 10.0919 0.10525 0.00013393 0.78488 0.0081648 0.0090773 0.0014001 0.98677 0.99159 3.0208e-006 1.2083e-005 0.15523 0.88508 0.89392 0.0014044 0.97544 0.48478 0.0018918 0.42491 1.8928 1.8917 16.011 144.9507 0.00019914 -85.5924 0.55894
5.663 0.98809 5.4872e-005 3.8183 0.011968 7.3971e-005 0.0011625 0.23255 0.0006593 0.23321 0.21517 0 0.032316 0.0389 0 1.33 0.45179 0.13722 0.0169 10.0941 0.10526 0.00013394 0.78487 0.0081654 0.0090779 0.0014 0.98677 0.99159 3.0205e-006 1.2082e-005 0.15524 0.88539 0.89406 0.0014043 0.97558 0.48496 0.0018917 0.42492 1.8935 1.8924 16.011 144.9508 0.00019892 -85.593 0.55994
5.664 0.98809 5.4872e-005 3.8183 0.011967 7.3984e-005 0.0011625 0.23255 0.0006593 0.23321 0.21517 0 0.032316 0.0389 0 1.3301 0.45183 0.13724 0.016901 10.0962 0.10527 0.00013396 0.78486 0.008166 0.0090785 0.0013999 0.98677 0.99159 3.0202e-006 1.2081e-005 0.15524 0.8857 0.8942 0.0014042 0.97572 0.48514 0.0018916 0.42494 1.8943 1.8932 16.0109 144.9508 0.00019871 -85.5935 0.56094
5.665 0.98809 5.4872e-005 3.8183 0.011967 7.3997e-005 0.0011625 0.23255 0.0006593 0.23321 0.21517 0 0.032316 0.0389 0 1.3302 0.45188 0.13725 0.016903 10.0983 0.10528 0.00013397 0.78485 0.0081665 0.0090791 0.0013997 0.98677 0.99159 3.02e-006 1.208e-005 0.15525 0.886 0.89433 0.0014042 0.97586 0.48532 0.0018915 0.42495 1.895 1.8939 16.0109 144.9508 0.0001985 -85.594 0.56194
5.666 0.98809 5.4872e-005 3.8183 0.011967 7.401e-005 0.0011625 0.23256 0.0006593 0.23321 0.21517 0 0.032316 0.0389 0 1.3303 0.45193 0.13727 0.016904 10.1005 0.10529 0.00013398 0.78484 0.0081671 0.0090797 0.0013996 0.98677 0.99159 3.0197e-006 1.2079e-005 0.15525 0.88631 0.89447 0.0014041 0.97599 0.4855 0.0018914 0.42496 1.8957 1.8946 16.0109 144.9508 0.00019829 -85.5945 0.56294
5.667 0.98809 5.4872e-005 3.8183 0.011967 7.4023e-005 0.0011625 0.23256 0.0006593 0.23321 0.21517 0 0.032316 0.0389 0 1.3304 0.45197 0.13728 0.016906 10.1026 0.1053 0.00013399 0.78484 0.0081677 0.0090803 0.0013995 0.98677 0.99159 3.0194e-006 1.2078e-005 0.15525 0.88661 0.8946 0.0014041 0.97613 0.48568 0.0018913 0.42498 1.8965 1.8954 16.0109 144.9508 0.00019808 -85.595 0.56394
5.668 0.98809 5.4872e-005 3.8183 0.011967 7.4036e-005 0.0011625 0.23256 0.0006593 0.23321 0.21517 0 0.032316 0.0389 0 1.3305 0.45202 0.1373 0.016907 10.1048 0.10531 0.00013401 0.78483 0.0081682 0.0090809 0.0013994 0.98677 0.99159 3.0192e-006 1.2077e-005 0.15526 0.88691 0.89474 0.001404 0.97627 0.48586 0.0018913 0.42499 1.8972 1.8961 16.0109 144.9509 0.00019787 -85.5955 0.56494
5.669 0.98809 5.4872e-005 3.8183 0.011967 7.4049e-005 0.0011625 0.23256 0.0006593 0.23321 0.21518 0 0.032316 0.0389 0 1.3306 0.45207 0.13731 0.016908 10.1069 0.10532 0.00013402 0.78482 0.0081688 0.0090815 0.0013993 0.98678 0.9916 3.0189e-006 1.2076e-005 0.15526 0.88722 0.89487 0.0014039 0.9764 0.48604 0.0018912 0.42501 1.8979 1.8968 16.0109 144.9509 0.00019767 -85.5959 0.56594
5.67 0.98809 5.4872e-005 3.8183 0.011967 7.4061e-005 0.0011625 0.23256 0.0006593 0.23322 0.21518 0 0.032316 0.0389 0 1.3307 0.45211 0.13733 0.01691 10.109 0.10532 0.00013403 0.78481 0.0081694 0.0090821 0.0013992 0.98678 0.9916 3.0187e-006 1.2075e-005 0.15527 0.88752 0.895 0.0014039 0.97654 0.48622 0.0018911 0.42502 1.8986 1.8975 16.0108 144.9509 0.00019746 -85.5964 0.56694
5.671 0.98809 5.4872e-005 3.8183 0.011967 7.4074e-005 0.0011626 0.23256 0.0006593 0.23322 0.21518 0 0.032316 0.0389 0 1.3308 0.45216 0.13735 0.016911 10.1112 0.10533 0.00013404 0.7848 0.0081699 0.0090827 0.0013991 0.98678 0.9916 3.0184e-006 1.2074e-005 0.15527 0.88782 0.89514 0.0014038 0.97667 0.48639 0.001891 0.42503 1.8994 1.8983 16.0108 144.9509 0.00019725 -85.5969 0.56794
5.672 0.98809 5.4871e-005 3.8183 0.011967 7.4087e-005 0.0011626 0.23256 0.0006593 0.23322 0.21518 0 0.032316 0.0389 0 1.3308 0.4522 0.13736 0.016913 10.1133 0.10534 0.00013406 0.78479 0.0081705 0.0090834 0.0013989 0.98678 0.9916 3.0181e-006 1.2073e-005 0.15528 0.88812 0.89527 0.0014038 0.9768 0.48657 0.001891 0.42505 1.9001 1.899 16.0108 144.9509 0.00019705 -85.5974 0.56894
5.673 0.98809 5.4871e-005 3.8183 0.011967 7.41e-005 0.0011626 0.23257 0.0006593 0.23322 0.21518 0 0.032316 0.0389 0 1.3309 0.45225 0.13738 0.016914 10.1155 0.10535 0.00013407 0.78478 0.0081711 0.009084 0.0013988 0.98678 0.9916 3.0179e-006 1.2071e-005 0.15528 0.88841 0.8954 0.0014037 0.97693 0.48675 0.0018909 0.42506 1.9008 1.8997 16.0108 144.951 0.00019684 -85.5979 0.56994
5.674 0.98809 5.4871e-005 3.8183 0.011967 7.4113e-005 0.0011626 0.23257 0.0006593 0.23322 0.21518 0 0.032316 0.0389 0 1.331 0.4523 0.13739 0.016915 10.1176 0.10536 0.00013408 0.78478 0.0081716 0.0090846 0.0013987 0.98678 0.9916 3.0176e-006 1.207e-005 0.15529 0.88871 0.89553 0.0014036 0.97707 0.48693 0.0018908 0.42507 1.9015 1.9004 16.0108 144.951 0.00019664 -85.5983 0.57094
5.675 0.98809 5.4871e-005 3.8183 0.011967 7.4126e-005 0.0011626 0.23257 0.0006593 0.23322 0.21518 0 0.032316 0.0389 0 1.3311 0.45234 0.13741 0.016917 10.1198 0.10537 0.00013409 0.78477 0.0081722 0.0090852 0.0013986 0.98678 0.9916 3.0174e-006 1.2069e-005 0.15529 0.88901 0.89566 0.0014036 0.9772 0.48711 0.0018907 0.42509 1.9022 1.9012 16.0108 144.951 0.00019644 -85.5988 0.57194
5.676 0.98809 5.4871e-005 3.8183 0.011967 7.4139e-005 0.0011626 0.23257 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3312 0.45239 0.13742 0.016918 10.1219 0.10538 0.00013411 0.78476 0.0081728 0.0090858 0.0013985 0.98679 0.9916 3.0171e-006 1.2068e-005 0.15529 0.8893 0.89579 0.0014035 0.97733 0.48729 0.0018907 0.4251 1.903 1.9019 16.0107 144.951 0.00019624 -85.5993 0.57294
5.677 0.98809 5.4871e-005 3.8183 0.011967 7.4152e-005 0.0011626 0.23257 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3313 0.45244 0.13744 0.01692 10.124 0.10538 0.00013412 0.78475 0.0081733 0.0090864 0.0013984 0.98679 0.9916 3.0169e-006 1.2067e-005 0.1553 0.8896 0.89592 0.0014035 0.97745 0.48747 0.0018906 0.42512 1.9037 1.9026 16.0107 144.951 0.00019603 -85.5997 0.57394
5.678 0.98809 5.4871e-005 3.8183 0.011967 7.4165e-005 0.0011626 0.23257 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3314 0.45248 0.13745 0.016921 10.1262 0.10539 0.00013413 0.78474 0.0081739 0.009087 0.0013983 0.98679 0.9916 3.0166e-006 1.2066e-005 0.1553 0.88989 0.89605 0.0014034 0.97758 0.48764 0.0018905 0.42513 1.9044 1.9033 16.0107 144.9511 0.00019583 -85.6002 0.57494
5.679 0.98809 5.4871e-005 3.8183 0.011967 7.4178e-005 0.0011626 0.23257 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3315 0.45253 0.13747 0.016923 10.1283 0.1054 0.00013414 0.78473 0.0081745 0.0090876 0.0013982 0.98679 0.9916 3.0164e-006 1.2066e-005 0.15531 0.89018 0.89618 0.0014034 0.97771 0.48782 0.0018904 0.42514 1.9051 1.904 16.0107 144.9511 0.00019563 -85.6007 0.57594
5.68 0.98809 5.4871e-005 3.8183 0.011967 7.4191e-005 0.0011626 0.23258 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3316 0.45258 0.13748 0.016924 10.1305 0.10541 0.00013416 0.78472 0.008175 0.0090882 0.0013981 0.98679 0.99161 3.0162e-006 1.2065e-005 0.15531 0.89047 0.89631 0.0014033 0.97783 0.488 0.0018904 0.42516 1.9058 1.9047 16.0107 144.9511 0.00019543 -85.6011 0.57694
5.681 0.98809 5.4871e-005 3.8183 0.011967 7.4204e-005 0.0011626 0.23258 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3317 0.45262 0.1375 0.016925 10.1326 0.10542 0.00013417 0.78471 0.0081756 0.0090888 0.001398 0.98679 0.99161 3.0159e-006 1.2064e-005 0.15532 0.89076 0.89644 0.0014033 0.97796 0.48818 0.0018903 0.42517 1.9065 1.9054 16.0107 144.9511 0.00019524 -85.6016 0.57794
5.682 0.98809 5.4871e-005 3.8183 0.011967 7.4217e-005 0.0011626 0.23258 0.0006593 0.23323 0.21519 0 0.032315 0.0389 0 1.3318 0.45267 0.13751 0.016927 10.1348 0.10543 0.00013418 0.78471 0.0081762 0.0090895 0.0013979 0.98679 0.99161 3.0157e-006 1.2063e-005 0.15532 0.89105 0.89657 0.0014032 0.97808 0.48836 0.0018902 0.42518 1.9072 1.9061 16.0106 144.9511 0.00019504 -85.602 0.57894
5.683 0.98809 5.4871e-005 3.8183 0.011967 7.423e-005 0.0011626 0.23258 0.0006593 0.23324 0.2152 0 0.032315 0.0389 0 1.3319 0.45271 0.13753 0.016928 10.1369 0.10544 0.00013419 0.7847 0.0081767 0.0090901 0.0013978 0.9868 0.99161 3.0154e-006 1.2062e-005 0.15533 0.89134 0.89669 0.0014032 0.97821 0.48853 0.0018901 0.4252 1.9079 1.9069 16.0106 144.9512 0.00019484 -85.6025 0.57994
5.684 0.98809 5.4871e-005 3.8183 0.011967 7.4243e-005 0.0011626 0.23258 0.0006593 0.23324 0.2152 0 0.032315 0.0389 0 1.332 0.45276 0.13754 0.01693 10.1391 0.10545 0.00013421 0.78469 0.0081773 0.0090907 0.0013977 0.9868 0.99161 3.0152e-006 1.2061e-005 0.15533 0.89163 0.89682 0.0014031 0.97833 0.48871 0.0018901 0.42521 1.9086 1.9076 16.0106 144.9512 0.00019465 -85.6029 0.58094
5.685 0.98809 5.487e-005 3.8183 0.011967 7.4255e-005 0.0011626 0.23258 0.0006593 0.23324 0.2152 0 0.032315 0.0389 0 1.3321 0.45281 0.13756 0.016931 10.1412 0.10545 0.00013422 0.78468 0.0081779 0.0090913 0.0013976 0.9868 0.99161 3.015e-006 1.206e-005 0.15533 0.89192 0.89695 0.001403 0.97845 0.48889 0.00189 0.42523 1.9093 1.9083 16.0106 144.9512 0.00019445 -85.6033 0.58194
5.686 0.98809 5.487e-005 3.8183 0.011967 7.4268e-005 0.0011626 0.23259 0.0006593 0.23324 0.2152 0 0.032315 0.0389 0 1.3322 0.45285 0.13757 0.016932 10.1434 0.10546 0.00013423 0.78467 0.0081784 0.0090919 0.0013975 0.9868 0.99161 3.0147e-006 1.2059e-005 0.15534 0.8922 0.89707 0.001403 0.97857 0.48907 0.0018899 0.42524 1.91 1.909 16.0106 144.9512 0.00019426 -85.6038 0.58294
5.687 0.98809 5.487e-005 3.8183 0.011967 7.4281e-005 0.0011626 0.23259 0.0006593 0.23324 0.2152 0 0.032315 0.0389 0 1.3323 0.4529 0.13759 0.016934 10.1455 0.10547 0.00013424 0.78466 0.008179 0.0090925 0.0013974 0.9868 0.99161 3.0145e-006 1.2058e-005 0.15534 0.89249 0.8972 0.0014029 0.97869 0.48925 0.0018899 0.42525 1.9107 1.9097 16.0105 144.9512 0.00019406 -85.6042 0.58394
5.688 0.98809 5.487e-005 3.8183 0.011967 7.4294e-005 0.0011626 0.23259 0.0006593 0.23324 0.2152 0 0.032315 0.0389 0 1.3324 0.45295 0.1376 0.016935 10.1477 0.10548 0.00013426 0.78465 0.0081796 0.0090931 0.0013973 0.9868 0.99161 3.0143e-006 1.2057e-005 0.15535 0.89277 0.89732 0.0014029 0.97881 0.48942 0.0018898 0.42527 1.9114 1.9103 16.0105 144.9513 0.00019387 -85.6046 0.58494
5.689 0.98809 5.487e-005 3.8183 0.011967 7.4307e-005 0.0011626 0.23259 0.0006593 0.23324 0.2152 0 0.032314 0.0389 0 1.3324 0.45299 0.13762 0.016937 10.1498 0.10549 0.00013427 0.78465 0.0081801 0.0090937 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.15535 0.89306 0.89744 0.0014028 0.97893 0.4896 0.0018897 0.42528 1.9121 1.911 16.0105 144.9513 0.00019368 -85.6051 0.58594
5.69 0.98809 5.487e-005 3.8183 0.011967 7.432e-005 0.0011626 0.23259 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.3325 0.45304 0.13763 0.016938 10.152 0.1055 0.00013428 0.78464 0.0081807 0.0090943 0.0013971 0.9868 0.99161 3.0138e-006 1.2055e-005 0.15536 0.89334 0.89757 0.0014028 0.97905 0.48978 0.0018897 0.42529 1.9128 1.9117 16.0105 144.9513 0.00019348 -85.6055 0.58694
5.691 0.98809 5.487e-005 3.8183 0.011967 7.4333e-005 0.0011626 0.23259 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.3326 0.45309 0.13765 0.01694 10.1541 0.10551 0.00013429 0.78463 0.0081812 0.0090949 0.001397 0.98681 0.99162 3.0136e-006 1.2054e-005 0.15536 0.89362 0.89769 0.0014027 0.97917 0.48996 0.0018896 0.42531 1.9135 1.9124 16.0105 144.9513 0.00019329 -85.6059 0.58794
5.692 0.98809 5.487e-005 3.8183 0.011967 7.4346e-005 0.0011626 0.23259 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.3327 0.45313 0.13766 0.016941 10.1563 0.10551 0.00013431 0.78462 0.0081818 0.0090955 0.0013969 0.98681 0.99162 3.0134e-006 1.2053e-005 0.15537 0.8939 0.89781 0.0014027 0.97929 0.49013 0.0018895 0.42532 1.9141 1.9131 16.0105 144.9513 0.0001931 -85.6063 0.58894
5.693 0.98809 5.487e-005 3.8183 0.011967 7.4359e-005 0.0011626 0.2326 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.3328 0.45318 0.13768 0.016942 10.1584 0.10552 0.00013432 0.78461 0.0081824 0.0090962 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.15537 0.89418 0.89794 0.0014026 0.9794 0.49031 0.0018895 0.42534 1.9148 1.9138 16.0104 144.9514 0.00019291 -85.6068 0.58994
5.694 0.98809 5.487e-005 3.8183 0.011967 7.4372e-005 0.0011626 0.2326 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.3329 0.45322 0.13769 0.016944 10.1606 0.10553 0.00013433 0.7846 0.0081829 0.0090968 0.0013967 0.98681 0.99162 3.0129e-006 1.2052e-005 0.15537 0.89446 0.89806 0.0014026 0.97952 0.49049 0.0018894 0.42535 1.9155 1.9145 16.0104 144.9514 0.00019273 -85.6072 0.59094
5.695 0.98809 5.487e-005 3.8183 0.011967 7.4385e-005 0.0011626 0.2326 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.333 0.45327 0.13771 0.016945 10.1627 0.10554 0.00013434 0.78459 0.0081835 0.0090974 0.0013966 0.98681 0.99162 3.0127e-006 1.2051e-005 0.15538 0.89474 0.89818 0.0014025 0.97963 0.49067 0.0018893 0.42536 1.9162 1.9152 16.0104 144.9514 0.00019254 -85.6076 0.59194
5.696 0.98809 5.487e-005 3.8183 0.011967 7.4398e-005 0.0011626 0.2326 0.0006593 0.23325 0.21521 0 0.032314 0.0389 0 1.3331 0.45332 0.13772 0.016947 10.1649 0.10555 0.00013436 0.78459 0.0081841 0.009098 0.0013965 0.98681 0.99162 3.0125e-006 1.205e-005 0.15538 0.89502 0.8983 0.0014025 0.97975 0.49084 0.0018893 0.42538 1.9169 1.9159 16.0104 144.9514 0.00019235 -85.608 0.59294
5.697 0.98809 5.487e-005 3.8183 0.011967 7.4411e-005 0.0011626 0.2326 0.0006593 0.23326 0.21522 0 0.032314 0.0389 0 1.3332 0.45336 0.13774 0.016948 10.167 0.10556 0.00013437 0.78458 0.0081846 0.0090986 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.15539 0.89529 0.89842 0.0014024 0.97986 0.49102 0.0018892 0.42539 1.9176 1.9165 16.0104 144.9514 0.00019216 -85.6084 0.59394
5.698 0.98809 5.4869e-005 3.8183 0.011967 7.4424e-005 0.0011626 0.2326 0.0006593 0.23326 0.21522 0 0.032314 0.0389 0 1.3333 0.45341 0.13776 0.016949 10.1692 0.10557 0.00013438 0.78457 0.0081852 0.0090992 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.15539 0.89557 0.89854 0.0014024 0.97997 0.4912 0.0018891 0.4254 1.9182 1.9172 16.0103 144.9515 0.00019198 -85.6088 0.59494
5.699 0.98809 5.4869e-005 3.8183 0.011967 7.4437e-005 0.0011626 0.2326 0.0006593 0.23326 0.21522 0 0.032314 0.0389 0 1.3334 0.45346 0.13777 0.016951 10.1713 0.10558 0.00013439 0.78456 0.0081858 0.0090998 0.0013962 0.98682 0.99162 3.0119e-006 1.2047e-005 0.1554 0.89584 0.89866 0.0014023 0.98008 0.49137 0.0018891 0.42542 1.9189 1.9179 16.0103 144.9515 0.00019179 -85.6092 0.59594
5.7 0.98809 5.4869e-005 3.8183 0.011967 7.4449e-005 0.0011626 0.23261 0.0006593 0.23326 0.21522 0 0.032314 0.0389 0 1.3335 0.4535 0.13779 0.016952 10.1735 0.10558 0.00013441 0.78455 0.0081863 0.0091004 0.0013961 0.98682 0.99162 3.0116e-006 1.2046e-005 0.1554 0.89612 0.89878 0.0014023 0.98019 0.49155 0.001889 0.42543 1.9196 1.9186 16.0103 144.9515 0.00019161 -85.6096 0.59694
5.701 0.98809 5.4869e-005 3.8183 0.011967 7.4462e-005 0.0011627 0.23261 0.0006593 0.23326 0.21522 0 0.032314 0.0389 0 1.3336 0.45355 0.1378 0.016954 10.1756 0.10559 0.00013442 0.78454 0.0081869 0.009101 0.001396 0.98682 0.99162 3.0114e-006 1.2046e-005 0.15541 0.89639 0.8989 0.0014022 0.9803 0.49173 0.0018889 0.42545 1.9203 1.9192 16.0103 144.9515 0.00019142 -85.61 0.59794
5.702 0.98809 5.4869e-005 3.8183 0.011967 7.4475e-005 0.0011627 0.23261 0.0006593 0.23326 0.21522 0 0.032314 0.0389 0 1.3337 0.4536 0.13782 0.016955 10.1778 0.1056 0.00013443 0.78453 0.0081875 0.0091016 0.0013959 0.98682 0.99162 3.0112e-006 1.2045e-005 0.15541 0.89666 0.89902 0.0014022 0.98041 0.4919 0.0018889 0.42546 1.9209 1.9199 16.0103 144.9515 0.00019124 -85.6104 0.59894
5.703 0.98809 5.4869e-005 3.8183 0.011967 7.4488e-005 0.0011627 0.23261 0.0006593 0.23326 0.21522 0 0.032313 0.0389 0 1.3338 0.45364 0.13783 0.016957 10.1799 0.10561 0.00013444 0.78452 0.008188 0.0091022 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.15541 0.89693 0.89913 0.0014021 0.98052 0.49208 0.0018888 0.42547 1.9216 1.9206 16.0102 144.9516 0.00019106 -85.6108 0.59994
5.704 0.98809 5.4869e-005 3.8183 0.011967 7.4501e-005 0.0011627 0.23261 0.0006593 0.23327 0.21523 0 0.032313 0.0389 0 1.3339 0.45369 0.13785 0.016958 10.1821 0.10562 0.00013446 0.78452 0.0081886 0.0091028 0.0013957 0.98682 0.99163 3.0108e-006 1.2043e-005 0.15542 0.8972 0.89925 0.0014021 0.98063 0.49226 0.0018888 0.42549 1.9223 1.9213 16.0102 144.9516 0.00019088 -85.6111 0.60094
5.705 0.98809 5.4869e-005 3.8183 0.011967 7.4514e-005 0.0011627 0.23261 0.0006593 0.23327 0.21523 0 0.032313 0.0389 0 1.334 0.45373 0.13786 0.016959 10.1842 0.10563 0.00013447 0.78451 0.0081891 0.0091035 0.0013957 0.98682 0.99163 3.0106e-006 1.2042e-005 0.15542 0.89747 0.89937 0.001402 0.98074 0.49243 0.0018887 0.4255 1.9229 1.9219 16.0102 144.9516 0.00019069 -85.6115 0.60194
5.706 0.98809 5.4869e-005 3.8183 0.011967 7.4527e-005 0.0011627 0.23261 0.0006593 0.23327 0.21523 0 0.032313 0.0389 0 1.334 0.45378 0.13788 0.016961 10.1864 0.10564 0.00013448 0.7845 0.0081897 0.0091041 0.0013956 0.98682 0.99163 3.0104e-006 1.2042e-005 0.15543 0.89774 0.89948 0.001402 0.98084 0.49261 0.0018886 0.42551 1.9236 1.9226 16.0102 144.9516 0.00019051 -85.6119 0.60294
5.707 0.98809 5.4869e-005 3.8183 0.011967 7.454e-005 0.0011627 0.23262 0.0006593 0.23327 0.21523 0 0.032313 0.0389 0 1.3341 0.45383 0.13789 0.016962 10.1885 0.10564 0.00013449 0.78449 0.0081903 0.0091047 0.0013955 0.98683 0.99163 3.0102e-006 1.2041e-005 0.15543 0.89801 0.8996 0.0014019 0.98095 0.49279 0.0018886 0.42553 1.9242 1.9233 16.0102 144.9516 0.00019033 -85.6123 0.60394
5.708 0.98809 5.4869e-005 3.8183 0.011967 7.4553e-005 0.0011627 0.23262 0.0006593 0.23327 0.21523 0 0.032313 0.0389 0 1.3342 0.45387 0.13791 0.016964 10.1907 0.10565 0.00013451 0.78448 0.0081908 0.0091053 0.0013954 0.98683 0.99163 3.01e-006 1.204e-005 0.15544 0.89828 0.89972 0.0014019 0.98105 0.49296 0.0018885 0.42554 1.9249 1.9239 16.0101 144.9517 0.00019016 -85.6126 0.60494
5.709 0.98809 5.4869e-005 3.8183 0.011967 7.4566e-005 0.0011627 0.23262 0.0006593 0.23327 0.21523 0 0.032313 0.0389 0 1.3343 0.45392 0.13792 0.016965 10.1928 0.10566 0.00013452 0.78447 0.0081914 0.0091059 0.0013953 0.98683 0.99163 3.0098e-006 1.2039e-005 0.15544 0.89854 0.89983 0.0014019 0.98116 0.49314 0.0018884 0.42556 1.9256 1.9246 16.0101 144.9517 0.00018998 -85.613 0.60594
5.71 0.98809 5.4869e-005 3.8183 0.011967 7.4579e-005 0.0011627 0.23262 0.0006593 0.23328 0.21523 0 0.032313 0.0389 0 1.3344 0.45397 0.13794 0.016966 10.195 0.10567 0.00013453 0.78446 0.008192 0.0091065 0.0013952 0.98683 0.99163 3.0096e-006 1.2038e-005 0.15545 0.89881 0.89995 0.0014018 0.98126 0.49332 0.0018884 0.42557 1.9262 1.9252 16.0101 144.9517 0.0001898 -85.6134 0.60694
5.711 0.98809 5.4868e-005 3.8183 0.011967 7.4592e-005 0.0011627 0.23262 0.0006593 0.23328 0.21523 0 0.032313 0.0389 0 1.3345 0.45401 0.13795 0.016968 10.1972 0.10568 0.00013454 0.78446 0.0081925 0.0091071 0.0013951 0.98683 0.99163 3.0094e-006 1.2038e-005 0.15545 0.89908 0.90006 0.0014018 0.98137 0.49349 0.0018883 0.42558 1.9269 1.9259 16.0101 144.9517 0.00018962 -85.6138 0.60794
5.712 0.98809 5.4868e-005 3.8183 0.011967 7.4605e-005 0.0011627 0.23262 0.0006593 0.23328 0.21524 0 0.032313 0.0389 0 1.3346 0.45406 0.13797 0.016969 10.1993 0.10569 0.00013456 0.78445 0.0081931 0.0091077 0.001395 0.98683 0.99163 3.0092e-006 1.2037e-005 0.15545 0.89934 0.90017 0.0014017 0.98147 0.49367 0.0018883 0.4256 1.9275 1.9266 16.0101 144.9517 0.00018945 -85.6141 0.60894
5.713 0.98809 5.4868e-005 3.8183 0.011967 7.4618e-005 0.0011627 0.23262 0.0006593 0.23328 0.21524 0 0.032313 0.0389 0 1.3347 0.45411 0.13798 0.016971 10.2015 0.1057 0.00013457 0.78444 0.0081937 0.0091083 0.001395 0.98683 0.99163 3.009e-006 1.2036e-005 0.15546 0.8996 0.90029 0.0014017 0.98157 0.49385 0.0018882 0.42561 1.9282 1.9272 16.01 144.9518 0.00018927 -85.6145 0.60994
5.714 0.98809 5.4868e-005 3.8183 0.011967 7.463e-005 0.0011627 0.23263 0.0006593 0.23328 0.21524 0 0.032313 0.0389 0 1.3348 0.45415 0.138 0.016972 10.2036 0.1057 0.00013458 0.78443 0.0081942 0.0091089 0.0013949 0.98683 0.99163 3.0088e-006 1.2035e-005 0.15546 0.89986 0.9004 0.0014016 0.98167 0.49402 0.0018882 0.42562 1.9288 1.9279 16.01 144.9518 0.00018909 -85.6148 0.61094
5.715 0.98809 5.4868e-005 3.8183 0.011967 7.4643e-005 0.0011627 0.23263 0.0006593 0.23328 0.21524 0 0.032313 0.0389 0 1.3349 0.4542 0.13801 0.016973 10.2058 0.10571 0.00013459 0.78442 0.0081948 0.0091095 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.15547 0.90013 0.90051 0.0014016 0.98177 0.4942 0.0018881 0.42564 1.9295 1.9285 16.01 144.9518 0.00018892 -85.6152 0.61194
5.716 0.98809 5.4868e-005 3.8183 0.011967 7.4656e-005 0.0011627 0.23263 0.0006593 0.23328 0.21524 0 0.032313 0.0389 0 1.335 0.45424 0.13803 0.016975 10.2079 0.10572 0.00013461 0.78441 0.0081953 0.0091101 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.15547 0.90039 0.90062 0.0014015 0.98187 0.49437 0.001888 0.42565 1.9301 1.9292 16.01 144.9518 0.00018875 -85.6156 0.61294
5.717 0.98809 5.4868e-005 3.8183 0.011967 7.4669e-005 0.0011627 0.23263 0.0006593 0.23329 0.21524 0 0.032312 0.0389 0 1.3351 0.45429 0.13804 0.016976 10.2101 0.10573 0.00013462 0.7844 0.0081959 0.0091107 0.0013946 0.98684 0.99163 3.0083e-006 1.2033e-005 0.15548 0.90065 0.90074 0.0014015 0.98197 0.49455 0.001888 0.42566 1.9308 1.9298 16.01 144.9518 0.00018857 -85.6159 0.61394
5.718 0.98809 5.4868e-005 3.8183 0.011967 7.4682e-005 0.0011627 0.23263 0.0006593 0.23329 0.21524 0 0.032312 0.0389 0 1.3352 0.45434 0.13806 0.016978 10.2123 0.10574 0.00013463 0.7844 0.0081965 0.0091113 0.0013946 0.98684 0.99164 3.0081e-006 1.2032e-005 0.15548 0.9009 0.90085 0.0014015 0.98207 0.49473 0.0018879 0.42568 1.9314 1.9305 16.0099 144.9519 0.0001884 -85.6163 0.61494
5.719 0.98809 5.4868e-005 3.8183 0.011967 7.4695e-005 0.0011627 0.23263 0.0006593 0.23329 0.21525 0 0.032312 0.0389 0 1.3353 0.45438 0.13807 0.016979 10.2144 0.10575 0.00013464 0.78439 0.008197 0.0091119 0.0013945 0.98684 0.99164 3.0079e-006 1.2032e-005 0.15548 0.90116 0.90096 0.0014014 0.98217 0.4949 0.0018879 0.42569 1.9321 1.9311 16.0099 144.9519 0.00018823 -85.6166 0.61594
5.72 0.98809 5.4868e-005 3.8183 0.011967 7.4708e-005 0.0011627 0.23263 0.0006593 0.23329 0.21525 0 0.032312 0.0389 0 1.3354 0.45443 0.13809 0.016981 10.2166 0.10576 0.00013466 0.78438 0.0081976 0.0091125 0.0013944 0.98684 0.99164 3.0077e-006 1.2031e-005 0.15549 0.90142 0.90107 0.0014014 0.98226 0.49508 0.0018878 0.42571 1.9327 1.9317 16.0099 144.9519 0.00018806 -85.6169 0.61694
5.721 0.98809 5.4868e-005 3.8183 0.011967 7.4721e-005 0.0011627 0.23264 0.0006593 0.23329 0.21525 0 0.032312 0.0389 0 1.3355 0.45448 0.1381 0.016982 10.2187 0.10576 0.00013467 0.78437 0.0081982 0.0091132 0.0013943 0.98684 0.99164 3.0075e-006 1.203e-005 0.15549 0.90168 0.90118 0.0014013 0.98236 0.49525 0.0018878 0.42572 1.9333 1.9324 16.0099 144.9519 0.00018789 -85.6173 0.61794
5.722 0.98809 5.4868e-005 3.8183 0.011967 7.4734e-005 0.0011627 0.23264 0.0006593 0.23329 0.21525 0 0.032312 0.0389 0 1.3356 0.45452 0.13812 0.016983 10.2209 0.10577 0.00013468 0.78436 0.0081987 0.0091138 0.0013942 0.98684 0.99164 3.0074e-006 1.2029e-005 0.1555 0.90193 0.90129 0.0014013 0.98246 0.49543 0.0018877 0.42573 1.934 1.933 16.0099 144.9519 0.00018772 -85.6176 0.61894
5.723 0.98809 5.4868e-005 3.8183 0.011967 7.4747e-005 0.0011627 0.23264 0.0006593 0.23329 0.21525 0 0.032312 0.0389 0 1.3356 0.45457 0.13813 0.016985 10.2231 0.10578 0.00013469 0.78435 0.0081993 0.0091144 0.0013942 0.98684 0.99164 3.0072e-006 1.2029e-005 0.1555 0.90219 0.9014 0.0014012 0.98255 0.4956 0.0018877 0.42575 1.9346 1.9337 16.0098 144.952 0.00018755 -85.618 0.61994
5.724 0.98809 5.4868e-005 3.8183 0.011967 7.476e-005 0.0011627 0.23264 0.0006593 0.2333 0.21525 0 0.032312 0.0389 0 1.3357 0.45462 0.13815 0.016986 10.2252 0.10579 0.00013471 0.78434 0.0081998 0.009115 0.0013941 0.98684 0.99164 3.007e-006 1.2028e-005 0.15551 0.90244 0.90151 0.0014012 0.98265 0.49578 0.0018876 0.42576 1.9353 1.9343 16.0098 144.952 0.00018738 -85.6183 0.62094
5.725 0.98809 5.4867e-005 3.8183 0.011966 7.4773e-005 0.0011627 0.23264 0.0006593 0.2333 0.21525 0 0.032312 0.0389 0 1.3358 0.45466 0.13816 0.016988 10.2274 0.1058 0.00013472 0.78434 0.0082004 0.0091156 0.001394 0.98684 0.99164 3.0068e-006 1.2027e-005 0.15551 0.90269 0.90161 0.0014012 0.98274 0.49596 0.0018875 0.42577 1.9359 1.9349 16.0098 144.952 0.00018721 -85.6186 0.62194
5.726 0.98809 5.4867e-005 3.8183 0.011966 7.4786e-005 0.0011627 0.23264 0.0006593 0.2333 0.21526 0 0.032312 0.0389 0 1.3359 0.45471 0.13818 0.016989 10.2295 0.10581 0.00013473 0.78433 0.008201 0.0091162 0.0013939 0.98685 0.99164 3.0067e-006 1.2027e-005 0.15552 0.90295 0.90172 0.0014011 0.98284 0.49613 0.0018875 0.42579 1.9365 1.9356 16.0098 144.952 0.00018704 -85.619 0.62294
5.727 0.98809 5.4867e-005 3.8183 0.011966 7.4799e-005 0.0011627 0.23264 0.0006593 0.2333 0.21526 0 0.032312 0.0389 0 1.336 0.45475 0.13819 0.01699 10.2317 0.10582 0.00013474 0.78432 0.0082015 0.0091168 0.0013938 0.98685 0.99164 3.0065e-006 1.2026e-005 0.15552 0.9032 0.90183 0.0014011 0.98293 0.49631 0.0018874 0.4258 1.9371 1.9362 16.0098 144.9521 0.00018687 -85.6193 0.62394
5.728 0.98809 5.4867e-005 3.8183 0.011966 7.4812e-005 0.0011627 0.23265 0.0006593 0.2333 0.21526 0 0.032312 0.0389 0 1.3361 0.4548 0.13821 0.016992 10.2339 0.10583 0.00013476 0.78431 0.0082021 0.0091174 0.0013938 0.98685 0.99164 3.0063e-006 1.2025e-005 0.15552 0.90345 0.90194 0.001401 0.98302 0.49648 0.0018874 0.42581 1.9378 1.9368 16.0097 144.9521 0.00018671 -85.6196 0.62494
5.729 0.98809 5.4867e-005 3.8183 0.011966 7.4824e-005 0.0011627 0.23265 0.0006593 0.2333 0.21526 0 0.032312 0.0389 0 1.3362 0.45485 0.13822 0.016993 10.236 0.10583 0.00013477 0.7843 0.0082026 0.009118 0.0013937 0.98685 0.99164 3.0061e-006 1.2024e-005 0.15553 0.9037 0.90204 0.001401 0.98311 0.49666 0.0018873 0.42583 1.9384 1.9375 16.0097 144.9521 0.00018654 -85.62 0.62594
5.73 0.98809 5.4867e-005 3.8183 0.011966 7.4837e-005 0.0011627 0.23265 0.0006593 0.2333 0.21526 0 0.032312 0.0389 0 1.3363 0.45489 0.13824 0.016995 10.2382 0.10584 0.00013478 0.78429 0.0082032 0.0091186 0.0013936 0.98685 0.99164 3.0059e-006 1.2024e-005 0.15553 0.90395 0.90215 0.001401 0.9832 0.49683 0.0018873 0.42584 1.939 1.9381 16.0097 144.9521 0.00018638 -85.6203 0.62694
5.731 0.98809 5.4867e-005 3.8183 0.011966 7.485e-005 0.0011628 0.23265 0.0006593 0.23331 0.21526 0 0.032311 0.0389 0 1.3364 0.45494 0.13826 0.016996 10.2404 0.10585 0.00013479 0.78428 0.0082038 0.0091192 0.0013935 0.98685 0.99164 3.0058e-006 1.2023e-005 0.15554 0.9042 0.90226 0.0014009 0.98329 0.49701 0.0018872 0.42586 1.9397 1.9387 16.0097 144.9521 0.00018621 -85.6206 0.62794
5.732 0.98809 5.4867e-005 3.8183 0.011966 7.4863e-005 0.0011628 0.23265 0.0006593 0.23331 0.21526 0 0.032311 0.0389 0 1.3365 0.45499 0.13827 0.016997 10.2425 0.10586 0.00013481 0.78428 0.0082043 0.0091198 0.0013935 0.98685 0.99164 3.0056e-006 1.2022e-005 0.15554 0.90445 0.90236 0.0014009 0.98339 0.49718 0.0018872 0.42587 1.9403 1.9394 16.0096 144.9522 0.00018605 -85.6209 0.62894
5.733 0.98809 5.4867e-005 3.8183 0.011966 7.4876e-005 0.0011628 0.23265 0.0006593 0.23331 0.21526 0 0.032311 0.0389 0 1.3366 0.45503 0.13829 0.016999 10.2447 0.10587 0.00013482 0.78427 0.0082049 0.0091204 0.0013934 0.98685 0.99164 3.0054e-006 1.2022e-005 0.15555 0.90469 0.90247 0.0014008 0.98347 0.49736 0.0018871 0.42588 1.9409 1.94 16.0096 144.9522 0.00018589 -85.6212 0.62994
5.734 0.98809 5.4867e-005 3.8183 0.011966 7.4889e-005 0.0011628 0.23265 0.0006593 0.23331 0.21527 0 0.032311 0.0389 0 1.3367 0.45508 0.1383 0.017 10.2468 0.10588 0.00013483 0.78426 0.0082055 0.009121 0.0013933 0.98685 0.99165 3.0053e-006 1.2021e-005 0.15555 0.90494 0.90257 0.0014008 0.98356 0.49753 0.0018871 0.4259 1.9415 1.9406 16.0096 144.9522 0.00018572 -85.6215 0.63094
5.735 0.98809 5.4867e-005 3.8183 0.011966 7.4902e-005 0.0011628 0.23266 0.0006593 0.23331 0.21527 0 0.032311 0.0389 0 1.3368 0.45512 0.13832 0.017002 10.249 0.10589 0.00013484 0.78425 0.008206 0.0091216 0.0013933 0.98685 0.99165 3.0051e-006 1.202e-005 0.15556 0.90518 0.90268 0.0014008 0.98365 0.49771 0.001887 0.42591 1.9421 1.9412 16.0096 144.9522 0.00018556 -85.6219 0.63194
5.736 0.98809 5.4867e-005 3.8183 0.011966 7.4915e-005 0.0011628 0.23266 0.0006593 0.23331 0.21527 0 0.032311 0.0389 0 1.3369 0.45517 0.13833 0.017003 10.2512 0.10589 0.00013486 0.78424 0.0082066 0.0091222 0.0013932 0.98685 0.99165 3.005e-006 1.202e-005 0.15556 0.90543 0.90278 0.0014007 0.98374 0.49788 0.001887 0.42592 1.9428 1.9418 16.0096 144.9522 0.0001854 -85.6222 0.63294
5.737 0.98809 5.4867e-005 3.8183 0.011966 7.4928e-005 0.0011628 0.23266 0.0006593 0.23331 0.21527 0 0.032311 0.0389 0 1.337 0.45522 0.13835 0.017004 10.2533 0.1059 0.00013487 0.78423 0.0082071 0.0091228 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.15556 0.90567 0.90289 0.0014007 0.98383 0.49806 0.0018869 0.42594 1.9434 1.9425 16.0095 144.9523 0.00018524 -85.6225 0.63394
5.738 0.98809 5.4866e-005 3.8183 0.011966 7.4941e-005 0.0011628 0.23266 0.0006593 0.23332 0.21527 0 0.032311 0.0389 0 1.3371 0.45526 0.13836 0.017006 10.2555 0.10591 0.00013488 0.78422 0.0082077 0.0091234 0.001393 0.98686 0.99165 3.0046e-006 1.2018e-005 0.15557 0.90592 0.90299 0.0014006 0.98391 0.49823 0.0018869 0.42595 1.944 1.9431 16.0095 144.9523 0.00018508 -85.6228 0.63494
5.739 0.98809 5.4866e-005 3.8183 0.011966 7.4954e-005 0.0011628 0.23266 0.0006593 0.23332 0.21527 0 0.032311 0.0389 0 1.3371 0.45531 0.13838 0.017007 10.2577 0.10592 0.00013489 0.78421 0.0082083 0.009124 0.001393 0.98686 0.99165 3.0045e-006 1.2018e-005 0.15557 0.90616 0.90309 0.0014006 0.984 0.49841 0.0018868 0.42596 1.9446 1.9437 16.0095 144.9523 0.00018492 -85.6231 0.63594
5.74 0.98809 5.4866e-005 3.8183 0.011966 7.4967e-005 0.0011628 0.23266 0.0006593 0.23332 0.21527 0 0.032311 0.0389 0 1.3372 0.45536 0.13839 0.017009 10.2598 0.10593 0.00013491 0.78421 0.0082088 0.0091246 0.0013929 0.98686 0.99165 3.0043e-006 1.2017e-005 0.15558 0.9064 0.90319 0.0014006 0.98408 0.49858 0.0018868 0.42598 1.9452 1.9443 16.0095 144.9523 0.00018476 -85.6234 0.63694
5.741 0.98809 5.4866e-005 3.8183 0.011966 7.498e-005 0.0011628 0.23266 0.0006593 0.23332 0.21528 0 0.032311 0.0389 0 1.3373 0.4554 0.13841 0.01701 10.262 0.10594 0.00013492 0.7842 0.0082094 0.0091253 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.15558 0.90664 0.9033 0.0014005 0.98417 0.49876 0.0018867 0.42599 1.9458 1.9449 16.0095 144.9523 0.0001846 -85.6237 0.63794
5.742 0.98809 5.4866e-005 3.8183 0.011966 7.4993e-005 0.0011628 0.23267 0.0006593 0.23332 0.21528 0 0.032311 0.0389 0 1.3374 0.45545 0.13842 0.017012 10.2642 0.10595 0.00013493 0.78419 0.0082099 0.0091259 0.0013928 0.98686 0.99165 3.004e-006 1.2016e-005 0.15559 0.90688 0.9034 0.0014005 0.98425 0.49893 0.0018867 0.42601 1.9464 1.9455 16.0094 144.9524 0.00018444 -85.624 0.63894
5.743 0.9881 5.4866e-005 3.8183 0.011966 7.5005e-005 0.0011628 0.23267 0.0006593 0.23332 0.21528 0 0.032311 0.0389 0 1.3375 0.4555 0.13844 0.017013 10.2663 0.10595 0.00013494 0.78418 0.0082105 0.0091265 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.15559 0.90712 0.9035 0.0014005 0.98434 0.4991 0.0018866 0.42602 1.947 1.9461 16.0094 144.9524 0.00018429 -85.6243 0.63994
5.744 0.9881 5.4866e-005 3.8183 0.011966 7.5018e-005 0.0011628 0.23267 0.0006593 0.23332 0.21528 0 0.032311 0.0389 0 1.3376 0.45554 0.13845 0.017014 10.2685 0.10596 0.00013496 0.78417 0.0082111 0.0091271 0.0013926 0.98686 0.99165 3.0037e-006 1.2015e-005 0.1556 0.90736 0.9036 0.0014004 0.98442 0.49928 0.0018866 0.42603 1.9476 1.9467 16.0094 144.9524 0.00018413 -85.6246 0.64094
5.745 0.9881 5.4866e-005 3.8183 0.011966 7.5031e-005 0.0011628 0.23267 0.0006593 0.23333 0.21528 0 0.03231 0.0389 0 1.3377 0.45559 0.13847 0.017016 10.2707 0.10597 0.00013497 0.78416 0.0082116 0.0091277 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.1556 0.9076 0.9037 0.0014004 0.9845 0.49945 0.0018866 0.42605 1.9482 1.9474 16.0094 144.9524 0.00018397 -85.6248 0.64194
5.746 0.9881 5.4866e-005 3.8183 0.011966 7.5044e-005 0.0011628 0.23267 0.0006593 0.23333 0.21528 0 0.03231 0.0389 0 1.3378 0.45563 0.13848 0.017017 10.2728 0.10598 0.00013498 0.78415 0.0082122 0.0091283 0.0013925 0.98686 0.99165 3.0034e-006 1.2014e-005 0.1556 0.90784 0.9038 0.0014004 0.98459 0.49963 0.0018865 0.42606 1.9488 1.948 16.0093 144.9524 0.00018382 -85.6251 0.64294
5.747 0.9881 5.4866e-005 3.8183 0.011966 7.5057e-005 0.0011628 0.23267 0.0006593 0.23333 0.21528 0 0.03231 0.0389 0 1.3379 0.45568 0.1385 0.017019 10.275 0.10599 0.00013499 0.78415 0.0082127 0.0091289 0.0013924 0.98686 0.99165 3.0033e-006 1.2013e-005 0.15561 0.90807 0.9039 0.0014003 0.98467 0.4998 0.0018865 0.42607 1.9495 1.9486 16.0093 144.9525 0.00018366 -85.6254 0.64394
5.748 0.9881 5.4866e-005 3.8183 0.011966 7.507e-005 0.0011628 0.23267 0.0006593 0.23333 0.21528 0 0.03231 0.0389 0 1.338 0.45573 0.13851 0.01702 10.2772 0.106 0.000135 0.78414 0.0082133 0.0091295 0.0013924 0.98687 0.99165 3.0031e-006 1.2012e-005 0.15561 0.90831 0.904 0.0014003 0.98475 0.49998 0.0018864 0.42609 1.9501 1.9492 16.0093 144.9525 0.00018351 -85.6257 0.64494
5.749 0.9881 5.4866e-005 3.8183 0.011966 7.5083e-005 0.0011628 0.23268 0.0006593 0.23333 0.21529 0 0.03231 0.0389 0 1.3381 0.45577 0.13853 0.017021 10.2794 0.10601 0.00013502 0.78413 0.0082139 0.0091301 0.0013923 0.98687 0.99165 3.0029e-006 1.2012e-005 0.15562 0.90854 0.9041 0.0014002 0.98483 0.50015 0.0018864 0.4261 1.9506 1.9498 16.0093 144.9525 0.00018335 -85.626 0.64594
5.75 0.9881 5.4866e-005 3.8183 0.011966 7.5096e-005 0.0011628 0.23268 0.0006593 0.23333 0.21529 0 0.03231 0.0389 0 1.3382 0.45582 0.13854 0.017023 10.2815 0.10601 0.00013503 0.78412 0.0082144 0.0091307 0.0013922 0.98687 0.99165 3.0028e-006 1.2011e-005 0.15562 0.90878 0.9042 0.0014002 0.98491 0.50032 0.0018863 0.42611 1.9512 1.9504 16.0093 144.9525 0.0001832 -85.6263 0.64694
5.751 0.9881 5.4865e-005 3.8183 0.011966 7.5109e-005 0.0011628 0.23268 0.0006593 0.23333 0.21529 0 0.03231 0.0389 0 1.3383 0.45587 0.13856 0.017024 10.2837 0.10602 0.00013504 0.78411 0.008215 0.0091313 0.0013922 0.98687 0.99166 3.0026e-006 1.201e-005 0.15563 0.90901 0.9043 0.0014002 0.98499 0.5005 0.0018863 0.42613 1.9518 1.951 16.0092 144.9525 0.00018305 -85.6265 0.64794
5.752 0.9881 5.4865e-005 3.8183 0.011966 7.5122e-005 0.0011628 0.23268 0.0006593 0.23333 0.21529 0 0.03231 0.0389 0 1.3384 0.45591 0.13857 0.017026 10.2859 0.10603 0.00013505 0.7841 0.0082155 0.0091319 0.0013921 0.98687 0.99166 3.0025e-006 1.201e-005 0.15563 0.90924 0.9044 0.0014001 0.98507 0.50067 0.0018862 0.42614 1.9524 1.9516 16.0092 144.9526 0.00018289 -85.6268 0.64894
5.753 0.9881 5.4865e-005 3.8183 0.011966 7.5135e-005 0.0011628 0.23268 0.0006593 0.23334 0.21529 0 0.03231 0.0389 0 1.3385 0.45596 0.13859 0.017027 10.288 0.10604 0.00013507 0.78409 0.0082161 0.0091325 0.001392 0.98687 0.99166 3.0023e-006 1.2009e-005 0.15563 0.90948 0.90449 0.0014001 0.98515 0.50084 0.0018862 0.42616 1.953 1.9522 16.0092 144.9526 0.00018274 -85.6271 0.64994
5.754 0.9881 5.4865e-005 3.8183 0.011966 7.5148e-005 0.0011628 0.23268 0.0006593 0.23334 0.21529 0 0.03231 0.0389 0 1.3386 0.45601 0.1386 0.017028 10.2902 0.10605 0.00013508 0.78409 0.0082167 0.0091331 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.15564 0.90971 0.90459 0.0014001 0.98523 0.50102 0.0018861 0.42617 1.9536 1.9527 16.0092 144.9526 0.00018259 -85.6274 0.65094
5.755 0.9881 5.4865e-005 3.8183 0.011966 7.5161e-005 0.0011628 0.23268 0.0006593 0.23334 0.21529 0 0.03231 0.0389 0 1.3387 0.45605 0.13862 0.01703 10.2924 0.10606 0.00013509 0.78408 0.0082172 0.0091337 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.15564 0.90994 0.90469 0.0014 0.9853 0.50119 0.0018861 0.42618 1.9542 1.9533 16.0091 144.9526 0.00018244 -85.6276 0.65194
5.756 0.9881 5.4865e-005 3.8183 0.011966 7.5174e-005 0.0011628 0.23269 0.0006593 0.23334 0.2153 0 0.03231 0.0389 0 1.3387 0.4561 0.13863 0.017031 10.2946 0.10607 0.0001351 0.78407 0.0082178 0.0091343 0.0013918 0.98687 0.99166 3.0019e-006 1.2008e-005 0.15565 0.91017 0.90478 0.0014 0.98538 0.50137 0.0018861 0.4262 1.9548 1.9539 16.0091 144.9526 0.00018229 -85.6279 0.65294
5.757 0.9881 5.4865e-005 3.8183 0.011966 7.5187e-005 0.0011628 0.23269 0.0006593 0.23334 0.2153 0 0.03231 0.0389 0 1.3388 0.45614 0.13865 0.017033 10.2967 0.10607 0.00013512 0.78406 0.0082183 0.0091349 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.15565 0.9104 0.90488 0.0014 0.98546 0.50154 0.001886 0.42621 1.9554 1.9545 16.0091 144.9527 0.00018214 -85.6282 0.65394
5.758 0.9881 5.4865e-005 3.8183 0.011966 7.5199e-005 0.0011628 0.23269 0.0006593 0.23334 0.2153 0 0.03231 0.0389 0 1.3389 0.45619 0.13866 0.017034 10.2989 0.10608 0.00013513 0.78405 0.0082189 0.0091355 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.15566 0.91063 0.90498 0.0014 0.98553 0.50171 0.001886 0.42622 1.956 1.9551 16.0091 144.9527 0.00018199 -85.6284 0.65494
5.759 0.9881 5.4865e-005 3.8183 0.011966 7.5212e-005 0.0011628 0.23269 0.0006593 0.23334 0.2153 0 0.032309 0.0389 0 1.339 0.45624 0.13868 0.017035 10.3011 0.10609 0.00013514 0.78404 0.0082195 0.0091361 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.15566 0.91085 0.90507 0.0013999 0.98561 0.50189 0.0018859 0.42624 1.9566 1.9557 16.009 144.9527 0.00018184 -85.6287 0.65594
5.76 0.9881 5.4865e-005 3.8183 0.011966 7.5225e-005 0.0011629 0.23269 0.0006593 0.23335 0.2153 0 0.032309 0.0389 0 1.3391 0.45628 0.13869 0.017037 10.3032 0.1061 0.00013515 0.78403 0.00822 0.0091367 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.15567 0.91108 0.90517 0.0013999 0.98568 0.50206 0.0018859 0.42625 1.9571 1.9563 16.009 144.9527 0.0001817 -85.629 0.65694
5.761 0.9881 5.4865e-005 3.8183 0.011966 7.5238e-005 0.0011629 0.23269 0.0006593 0.23335 0.2153 0 0.032309 0.0389 0 1.3392 0.45633 0.13871 0.017038 10.3054 0.10611 0.00013517 0.78403 0.0082206 0.0091373 0.0013915 0.98688 0.99166 3.0012e-006 1.2005e-005 0.15567 0.91131 0.90526 0.0013999 0.98576 0.50223 0.0018858 0.42626 1.9577 1.9569 16.009 144.9527 0.00018155 -85.6292 0.65794
5.762 0.9881 5.4865e-005 3.8183 0.011966 7.5251e-005 0.0011629 0.23269 0.0006593 0.23335 0.2153 0 0.032309 0.0389 0 1.3393 0.45638 0.13872 0.01704 10.3076 0.10612 0.00013518 0.78402 0.0082211 0.0091379 0.0013915 0.98688 0.99166 3.001e-006 1.2004e-005 0.15567 0.91153 0.90536 0.0013998 0.98583 0.50241 0.0018858 0.42628 1.9583 1.9575 16.009 144.9528 0.0001814 -85.6295 0.65894
5.763 0.9881 5.4865e-005 3.8183 0.011966 7.5264e-005 0.0011629 0.2327 0.0006593 0.23335 0.2153 0 0.032309 0.0389 0 1.3394 0.45642 0.13874 0.017041 10.3098 0.10613 0.00013519 0.78401 0.0082217 0.0091385 0.0013914 0.98688 0.99166 3.0009e-006 1.2004e-005 0.15568 0.91176 0.90545 0.0013998 0.98591 0.50258 0.0018858 0.42629 1.9589 1.958 16.009 144.9528 0.00018125 -85.6297 0.65994
5.764 0.9881 5.4864e-005 3.8183 0.011966 7.5277e-005 0.0011629 0.2327 0.0006593 0.23335 0.21531 0 0.032309 0.0389 0 1.3395 0.45647 0.13875 0.017042 10.3119 0.10613 0.0001352 0.784 0.0082222 0.0091391 0.0013914 0.98688 0.99166 3.0008e-006 1.2003e-005 0.15568 0.91198 0.90555 0.0013998 0.98598 0.50275 0.0018857 0.4263 1.9595 1.9586 16.0089 144.9528 0.00018111 -85.63 0.66094
5.765 0.9881 5.4864e-005 3.8183 0.011966 7.529e-005 0.0011629 0.2327 0.0006593 0.23335 0.21531 0 0.032309 0.0389 0 1.3396 0.45651 0.13877 0.017044 10.3141 0.10614 0.00013522 0.78399 0.0082228 0.0091397 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.15569 0.91221 0.90564 0.0013997 0.98605 0.50293 0.0018857 0.42632 1.96 1.9592 16.0089 144.9528 0.00018096 -85.6303 0.66194
5.766 0.9881 5.4864e-005 3.8183 0.011966 7.5303e-005 0.0011629 0.2327 0.0006593 0.23335 0.21531 0 0.032309 0.0389 0 1.3397 0.45656 0.13878 0.017045 10.3163 0.10615 0.00013523 0.78398 0.0082234 0.0091403 0.0013912 0.98688 0.99166 3.0005e-006 1.2002e-005 0.15569 0.91243 0.90573 0.0013997 0.98612 0.5031 0.0018856 0.42633 1.9606 1.9598 16.0089 144.9528 0.00018082 -85.6305 0.66294
5.767 0.9881 5.4864e-005 3.8183 0.011966 7.5316e-005 0.0011629 0.2327 0.0006593 0.23336 0.21531 0 0.032309 0.0389 0 1.3398 0.45661 0.1388 0.017047 10.3185 0.10616 0.00013524 0.78397 0.0082239 0.0091409 0.0013912 0.98688 0.99166 3.0004e-006 1.2001e-005 0.1557 0.91265 0.90583 0.0013997 0.9862 0.50327 0.0018856 0.42635 1.9612 1.9603 16.0089 144.9529 0.00018067 -85.6308 0.66394
5.768 0.9881 5.4864e-005 3.8183 0.011966 7.5329e-005 0.0011629 0.2327 0.0006593 0.23336 0.21531 0 0.032309 0.0389 0 1.3399 0.45665 0.13882 0.017048 10.3206 0.10617 0.00013525 0.78397 0.0082245 0.0091415 0.0013911 0.98688 0.99166 3.0003e-006 1.2001e-005 0.1557 0.91287 0.90592 0.0013996 0.98627 0.50345 0.0018856 0.42636 1.9618 1.9609 16.0088 144.9529 0.00018053 -85.631 0.66494
5.769 0.9881 5.4864e-005 3.8183 0.011966 7.5342e-005 0.0011629 0.2327 0.0006593 0.23336 0.21531 0 0.032309 0.0389 0 1.34 0.4567 0.13883 0.017049 10.3228 0.10618 0.00013527 0.78396 0.008225 0.0091421 0.0013911 0.98688 0.99166 3.0001e-006 1.2e-005 0.15571 0.91309 0.90601 0.0013996 0.98634 0.50362 0.0018855 0.42637 1.9623 1.9615 16.0088 144.9529 0.00018039 -85.6313 0.66594
5.77 0.9881 5.4864e-005 3.8183 0.011966 7.5355e-005 0.0011629 0.2327 0.0006593 0.23336 0.21531 0 0.032309 0.0389 0 1.3401 0.45675 0.13885 0.017051 10.325 0.10619 0.00013528 0.78395 0.0082256 0.0091427 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.15571 0.91331 0.9061 0.0013996 0.98641 0.50379 0.0018855 0.42639 1.9629 1.9621 16.0088 144.9529 0.00018025 -85.6315 0.66694
5.771 0.9881 5.4864e-005 3.8183 0.011966 7.5368e-005 0.0011629 0.23271 0.0006593 0.23336 0.21531 0 0.032309 0.0389 0 1.3402 0.45679 0.13886 0.017052 10.3272 0.10619 0.00013529 0.78394 0.0082262 0.0091433 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.15571 0.91353 0.90619 0.0013996 0.98648 0.50396 0.0018854 0.4264 1.9635 1.9626 16.0088 144.9529 0.0001801 -85.6317 0.66794
5.772 0.9881 5.4864e-005 3.8183 0.011966 7.538e-005 0.0011629 0.23271 0.0006593 0.23336 0.21532 0 0.032309 0.0389 0 1.3402 0.45684 0.13888 0.017054 10.3293 0.1062 0.0001353 0.78393 0.0082267 0.0091439 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.15572 0.91375 0.90628 0.0013995 0.98655 0.50414 0.0018854 0.42641 1.964 1.9632 16.0087 144.953 0.00017996 -85.632 0.66894
5.773 0.9881 5.4864e-005 3.8183 0.011966 7.5393e-005 0.0011629 0.23271 0.0006593 0.23336 0.21532 0 0.032309 0.0389 0 1.3403 0.45689 0.13889 0.017055 10.3315 0.10621 0.00013532 0.78392 0.0082273 0.0091445 0.0013908 0.98688 0.99167 2.9996e-006 1.1998e-005 0.15572 0.91397 0.90638 0.0013995 0.98662 0.50431 0.0018854 0.42643 1.9646 1.9638 16.0087 144.953 0.00017982 -85.6322 0.66994
5.774 0.9881 5.4864e-005 3.8183 0.011966 7.5406e-005 0.0011629 0.23271 0.0006593 0.23337 0.21532 0 0.032308 0.0389 0 1.3404 0.45693 0.13891 0.017057 10.3337 0.10622 0.00013533 0.78391 0.0082278 0.0091451 0.0013908 0.98689 0.99167 2.9994e-006 1.1998e-005 0.15573 0.91419 0.90647 0.0013995 0.98669 0.50448 0.0018853 0.42644 1.9652 1.9643 16.0087 144.953 0.00017968 -85.6325 0.67094
5.775 0.9881 5.4864e-005 3.8183 0.011966 7.5419e-005 0.0011629 0.23271 0.0006593 0.23337 0.21532 0 0.032308 0.0389 0 1.3405 0.45698 0.13892 0.017058 10.3359 0.10623 0.00013534 0.78391 0.0082284 0.0091457 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.15573 0.9144 0.90656 0.0013994 0.98675 0.50465 0.0018853 0.42645 1.9657 1.9649 16.0087 144.953 0.00017954 -85.6327 0.67194
5.776 0.9881 5.4864e-005 3.8183 0.011966 7.5432e-005 0.0011629 0.23271 0.0006593 0.23337 0.21532 0 0.032308 0.0389 0 1.3406 0.45702 0.13894 0.017059 10.3381 0.10624 0.00013535 0.7839 0.0082289 0.0091463 0.0013907 0.98689 0.99167 2.9992e-006 1.1997e-005 0.15574 0.91462 0.90665 0.0013994 0.98682 0.50483 0.0018853 0.42647 1.9663 1.9655 16.0087 144.953 0.0001794 -85.6329 0.67294
5.777 0.9881 5.4863e-005 3.8183 0.011966 7.5445e-005 0.0011629 0.23271 0.0006593 0.23337 0.21532 0 0.032308 0.0389 0 1.3407 0.45707 0.13895 0.017061 10.3402 0.10625 0.00013536 0.78389 0.0082295 0.0091469 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.15574 0.91483 0.90674 0.0013994 0.98689 0.505 0.0018852 0.42648 1.9669 1.966 16.0086 144.9531 0.00017926 -85.6332 0.67394
5.778 0.9881 5.4863e-005 3.8183 0.011966 7.5458e-005 0.0011629 0.23272 0.0006593 0.23337 0.21532 0 0.032308 0.0389 0 1.3408 0.45712 0.13897 0.017062 10.3424 0.10625 0.00013538 0.78388 0.0082301 0.0091475 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.15574 0.91505 0.90683 0.0013994 0.98696 0.50517 0.0018852 0.42649 1.9674 1.9666 16.0086 144.9531 0.00017912 -85.6334 0.67494
5.779 0.9881 5.4863e-005 3.8183 0.011966 7.5471e-005 0.0011629 0.23272 0.0006593 0.23337 0.21533 0 0.032308 0.0389 0 1.3409 0.45716 0.13898 0.017064 10.3446 0.10626 0.00013539 0.78387 0.0082306 0.0091481 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.15575 0.91526 0.90691 0.0013993 0.98702 0.50534 0.0018851 0.42651 1.968 1.9672 16.0086 144.9531 0.00017898 -85.6336 0.67594
5.78 0.9881 5.4863e-005 3.8183 0.011966 7.5484e-005 0.0011629 0.23272 0.0006593 0.23337 0.21533 0 0.032308 0.0389 0 1.341 0.45721 0.139 0.017065 10.3468 0.10627 0.0001354 0.78386 0.0082312 0.0091487 0.0013905 0.98689 0.99167 2.9987e-006 1.1995e-005 0.15575 0.91548 0.907 0.0013993 0.98709 0.50552 0.0018851 0.42652 1.9685 1.9677 16.0086 144.9531 0.00017885 -85.6339 0.67694
5.781 0.9881 5.4863e-005 3.8183 0.011966 7.5497e-005 0.0011629 0.23272 0.0006593 0.23337 0.21533 0 0.032308 0.0389 0 1.3411 0.45726 0.13901 0.017066 10.349 0.10628 0.00013541 0.78385 0.0082317 0.0091493 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.15576 0.91569 0.90709 0.0013993 0.98715 0.50569 0.0018851 0.42653 1.9691 1.9683 16.0085 144.9531 0.00017871 -85.6341 0.67794
5.782 0.9881 5.4863e-005 3.8183 0.011966 7.551e-005 0.0011629 0.23272 0.0006593 0.23338 0.21533 0 0.032308 0.0389 0 1.3412 0.4573 0.13903 0.017068 10.3511 0.10629 0.00013543 0.78385 0.0082323 0.0091499 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.15576 0.9159 0.90718 0.0013992 0.98722 0.50586 0.001885 0.42655 1.9696 1.9688 16.0085 144.9532 0.00017857 -85.6343 0.67894
5.783 0.9881 5.4863e-005 3.8183 0.011966 7.5523e-005 0.0011629 0.23272 0.0006593 0.23338 0.21533 0 0.032308 0.0389 0 1.3413 0.45735 0.13904 0.017069 10.3533 0.1063 0.00013544 0.78384 0.0082328 0.0091505 0.0013903 0.98689 0.99167 2.9984e-006 1.1993e-005 0.15577 0.91611 0.90727 0.0013992 0.98728 0.50603 0.001885 0.42656 1.9702 1.9694 16.0085 144.9532 0.00017844 -85.6345 0.67994
5.784 0.9881 5.4863e-005 3.8183 0.011966 7.5536e-005 0.0011629 0.23272 0.0006593 0.23338 0.21533 0 0.032308 0.0389 0 1.3414 0.45739 0.13906 0.017071 10.3555 0.10631 0.00013545 0.78383 0.0082334 0.0091511 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.15577 0.91632 0.90735 0.0013992 0.98735 0.5062 0.001885 0.42657 1.9708 1.9699 16.0085 144.9532 0.0001783 -85.6347 0.68094
5.785 0.9881 5.4863e-005 3.8183 0.011966 7.5549e-005 0.0011629 0.23273 0.0006593 0.23338 0.21533 0 0.032308 0.0389 0 1.3415 0.45744 0.13907 0.017072 10.3577 0.10631 0.00013546 0.78382 0.008234 0.0091517 0.0013902 0.98689 0.99167 2.9982e-006 1.1993e-005 0.15578 0.91653 0.90744 0.0013992 0.98741 0.50638 0.0018849 0.42659 1.9713 1.9705 16.0084 144.9532 0.00017817 -85.635 0.68194
5.786 0.9881 5.4863e-005 3.8183 0.011965 7.5561e-005 0.0011629 0.23273 0.0006593 0.23338 0.21533 0 0.032308 0.0389 0 1.3416 0.45749 0.13909 0.017073 10.3599 0.10632 0.00013548 0.78381 0.0082345 0.0091523 0.0013902 0.98689 0.99167 2.998e-006 1.1992e-005 0.15578 0.91674 0.90753 0.0013991 0.98748 0.50655 0.0018849 0.4266 1.9719 1.9711 16.0084 144.9532 0.00017803 -85.6352 0.68294
5.787 0.9881 5.4863e-005 3.8183 0.011965 7.5574e-005 0.0011629 0.23273 0.0006593 0.23338 0.21534 0 0.032308 0.0389 0 1.3417 0.45753 0.1391 0.017075 10.3621 0.10633 0.00013549 0.7838 0.0082351 0.0091529 0.0013901 0.98689 0.99167 2.9979e-006 1.1992e-005 0.15578 0.91695 0.90761 0.0013991 0.98754 0.50672 0.0018849 0.42661 1.9724 1.9716 16.0084 144.9533 0.0001779 -85.6354 0.68394
5.788 0.9881 5.4863e-005 3.8183 0.011965 7.5587e-005 0.0011629 0.23273 0.0006593 0.23338 0.21534 0 0.032308 0.0389 0 1.3417 0.45758 0.13912 0.017076 10.3642 0.10634 0.0001355 0.7838 0.0082356 0.0091535 0.0013901 0.9869 0.99167 2.9978e-006 1.1991e-005 0.15579 0.91716 0.9077 0.0013991 0.9876 0.50689 0.0018848 0.42663 1.973 1.9722 16.0084 144.9533 0.00017776 -85.6356 0.68494
5.789 0.9881 5.4863e-005 3.8183 0.011965 7.56e-005 0.001163 0.23273 0.0006593 0.23339 0.21534 0 0.032307 0.0389 0 1.3418 0.45763 0.13913 0.017078 10.3664 0.10635 0.00013551 0.78379 0.0082362 0.0091541 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.15579 0.91737 0.90779 0.001399 0.98766 0.50706 0.0018848 0.42664 1.9735 1.9727 16.0083 144.9533 0.00017763 -85.6358 0.68594
5.79 0.9881 5.4862e-005 3.8183 0.011965 7.5613e-005 0.001163 0.23273 0.0006593 0.23339 0.21534 0 0.032307 0.0389 0 1.3419 0.45767 0.13915 0.017079 10.3686 0.10636 0.00013553 0.78378 0.0082367 0.0091547 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.1558 0.91757 0.90787 0.001399 0.98772 0.50723 0.0018848 0.42666 1.974 1.9732 16.0083 144.9533 0.0001775 -85.6361 0.68694
5.791 0.9881 5.4862e-005 3.8183 0.011965 7.5626e-005 0.001163 0.23273 0.0006593 0.23339 0.21534 0 0.032307 0.0389 0 1.342 0.45772 0.13916 0.01708 10.3708 0.10637 0.00013554 0.78377 0.0082373 0.0091553 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.1558 0.91778 0.90796 0.001399 0.98779 0.50741 0.0018847 0.42667 1.9746 1.9738 16.0083 144.9534 0.00017736 -85.6363 0.68794
5.792 0.9881 5.4862e-005 3.8183 0.011965 7.5639e-005 0.001163 0.23273 0.0006593 0.23339 0.21534 0 0.032307 0.0389 0 1.3421 0.45777 0.13918 0.017082 10.373 0.10637 0.00013555 0.78376 0.0082379 0.0091559 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.15581 0.91798 0.90804 0.001399 0.98785 0.50758 0.0018847 0.42668 1.9751 1.9743 16.0083 144.9534 0.00017723 -85.6365 0.68894
5.793 0.9881 5.4862e-005 3.8183 0.011965 7.5652e-005 0.001163 0.23274 0.0006593 0.23339 0.21534 0 0.032307 0.0389 0 1.3422 0.45781 0.13919 0.017083 10.3752 0.10638 0.00013556 0.78375 0.0082384 0.0091565 0.0013898 0.9869 0.99167 2.9972e-006 1.1989e-005 0.15581 0.91819 0.90813 0.0013989 0.98791 0.50775 0.0018847 0.4267 1.9757 1.9749 16.0082 144.9534 0.0001771 -85.6367 0.68994
5.794 0.9881 5.4862e-005 3.8183 0.011965 7.5665e-005 0.001163 0.23274 0.0006593 0.23339 0.21534 0 0.032307 0.0389 0 1.3423 0.45786 0.13921 0.017085 10.3773 0.10639 0.00013558 0.78374 0.008239 0.0091571 0.0013898 0.9869 0.99168 2.9971e-006 1.1988e-005 0.15581 0.91839 0.90821 0.0013989 0.98797 0.50792 0.0018846 0.42671 1.9762 1.9754 16.0082 144.9534 0.00017697 -85.6369 0.69094
5.795 0.9881 5.4862e-005 3.8183 0.011965 7.5678e-005 0.001163 0.23274 0.0006593 0.23339 0.21535 0 0.032307 0.0389 0 1.3424 0.4579 0.13922 0.017086 10.3795 0.1064 0.00013559 0.78374 0.0082395 0.0091577 0.0013897 0.9869 0.99168 2.9971e-006 1.1988e-005 0.15582 0.9186 0.90829 0.0013989 0.98803 0.50809 0.0018846 0.42672 1.9768 1.976 16.0082 144.9534 0.00017684 -85.6371 0.69194
5.796 0.9881 5.4862e-005 3.8183 0.011965 7.5691e-005 0.001163 0.23274 0.0006593 0.23339 0.21535 0 0.032307 0.0389 0 1.3425 0.45795 0.13924 0.017087 10.3817 0.10641 0.0001356 0.78373 0.0082401 0.0091583 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.15582 0.9188 0.90838 0.0013989 0.98809 0.50826 0.0018846 0.42674 1.9773 1.9765 16.0082 144.9535 0.00017671 -85.6373 0.69294
5.797 0.9881 5.4862e-005 3.8183 0.011965 7.5704e-005 0.001163 0.23274 0.0006593 0.2334 0.21535 0 0.032307 0.0389 0 1.3426 0.458 0.13925 0.017089 10.3839 0.10642 0.00013561 0.78372 0.0082406 0.0091589 0.0013896 0.9869 0.99168 2.9969e-006 1.1987e-005 0.15583 0.919 0.90846 0.0013988 0.98815 0.50843 0.0018845 0.42675 1.9778 1.977 16.0081 144.9535 0.00017658 -85.6375 0.69394
5.798 0.9881 5.4862e-005 3.8183 0.011965 7.5717e-005 0.001163 0.23274 0.0006593 0.2334 0.21535 0 0.032307 0.0389 0 1.3427 0.45804 0.13927 0.01709 10.3861 0.10643 0.00013562 0.78371 0.0082412 0.0091595 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.15583 0.9192 0.90854 0.0013988 0.98821 0.50861 0.0018845 0.42676 1.9784 1.9776 16.0081 144.9535 0.00017645 -85.6377 0.69494
5.799 0.9881 5.4862e-005 3.8183 0.011965 7.573e-005 0.001163 0.23274 0.0006593 0.2334 0.21535 0 0.032307 0.0389 0 1.3428 0.45809 0.13928 0.017092 10.3883 0.10643 0.00013564 0.7837 0.0082417 0.0091601 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.15584 0.91941 0.90863 0.0013988 0.98826 0.50878 0.0018845 0.42678 1.9789 1.9781 16.0081 144.9535 0.00017632 -85.6379 0.69594
5.8 0.9881 5.4862e-005 3.8183 0.011965 7.5742e-005 0.001163 0.23275 0.0006593 0.2334 0.21535 0 0.032307 0.0389 0 1.3429 0.45814 0.1393 0.017093 10.3905 0.10644 0.00013565 0.78369 0.0082423 0.0091607 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.15584 0.91961 0.90871 0.0013988 0.98832 0.50895 0.0018844 0.42679 1.9794 1.9787 16.0081 144.9535 0.00017619 -85.6381 0.69694
5.801 0.9881 5.4862e-005 3.8183 0.011965 7.5755e-005 0.001163 0.23275 0.0006593 0.2334 0.21535 0 0.032307 0.0389 0 1.343 0.45818 0.13931 0.017094 10.3926 0.10645 0.00013566 0.78368 0.0082429 0.0091613 0.0013894 0.9869 0.99168 2.9964e-006 1.1986e-005 0.15585 0.91981 0.90879 0.0013987 0.98838 0.50912 0.0018844 0.4268 1.98 1.9792 16.008 144.9536 0.00017607 -85.6383 0.69794
5.802 0.9881 5.4862e-005 3.8183 0.011965 7.5768e-005 0.001163 0.23275 0.0006593 0.2334 0.21535 0 0.032307 0.0389 0 1.3431 0.45823 0.13933 0.017096 10.3948 0.10646 0.00013567 0.78368 0.0082434 0.0091619 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.15585 0.92 0.90887 0.0013987 0.98844 0.50929 0.0018844 0.42682 1.9805 1.9797 16.008 144.9536 0.00017594 -85.6385 0.69894
5.803 0.9881 5.4861e-005 3.8183 0.011965 7.5781e-005 0.001163 0.23275 0.0006593 0.2334 0.21536 0 0.032307 0.0389 0 1.3432 0.45827 0.13934 0.017097 10.397 0.10647 0.00013569 0.78367 0.008244 0.0091625 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.15585 0.9202 0.90896 0.0013987 0.98849 0.50946 0.0018843 0.42683 1.981 1.9802 16.008 144.9536 0.00017581 -85.6387 0.69994
5.804 0.9881 5.4861e-005 3.8183 0.011965 7.5794e-005 0.001163 0.23275 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3432 0.45832 0.13936 0.017099 10.3992 0.10648 0.0001357 0.78366 0.0082445 0.0091631 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.15586 0.9204 0.90904 0.0013987 0.98855 0.50963 0.0018843 0.42684 1.9815 1.9808 16.008 144.9536 0.00017569 -85.6389 0.70094
5.805 0.9881 5.4861e-005 3.8183 0.011965 7.5807e-005 0.001163 0.23275 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3433 0.45837 0.13937 0.0171 10.4014 0.10649 0.00013571 0.78365 0.0082451 0.0091637 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.15586 0.9206 0.90912 0.0013987 0.98861 0.5098 0.0018843 0.42686 1.9821 1.9813 16.0079 144.9536 0.00017556 -85.6391 0.70194
5.806 0.9881 5.4861e-005 3.8183 0.011965 7.582e-005 0.001163 0.23275 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3434 0.45841 0.13939 0.017101 10.4036 0.10649 0.00013572 0.78364 0.0082456 0.0091643 0.0013892 0.98691 0.99168 2.9959e-006 1.1983e-005 0.15587 0.92079 0.9092 0.0013986 0.98866 0.50997 0.0018842 0.42687 1.9826 1.9818 16.0079 144.9537 0.00017543 -85.6393 0.70294
5.807 0.9881 5.4861e-005 3.8183 0.011965 7.5833e-005 0.001163 0.23275 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3435 0.45846 0.1394 0.017103 10.4058 0.1065 0.00013574 0.78363 0.0082462 0.0091649 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.15587 0.92099 0.90928 0.0013986 0.98872 0.51014 0.0018842 0.42688 1.9831 1.9824 16.0079 144.9537 0.00017531 -85.6395 0.70394
5.808 0.9881 5.4861e-005 3.8183 0.011965 7.5846e-005 0.001163 0.23276 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3436 0.45851 0.13942 0.017104 10.408 0.10651 0.00013575 0.78362 0.0082467 0.0091655 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.15588 0.92119 0.90936 0.0013986 0.98877 0.51031 0.0018842 0.4269 1.9837 1.9829 16.0079 144.9537 0.00017519 -85.6396 0.70494
5.809 0.9881 5.4861e-005 3.8183 0.011965 7.5859e-005 0.001163 0.23276 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3437 0.45855 0.13943 0.017106 10.4102 0.10652 0.00013576 0.78362 0.0082473 0.0091661 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.15588 0.92138 0.90944 0.0013986 0.98883 0.51048 0.0018842 0.42691 1.9842 1.9834 16.0078 144.9537 0.00017506 -85.6398 0.70594
5.81 0.9881 5.4861e-005 3.8183 0.011965 7.5872e-005 0.001163 0.23276 0.0006593 0.23341 0.21536 0 0.032306 0.0389 0 1.3438 0.4586 0.13945 0.017107 10.4124 0.10653 0.00013577 0.78361 0.0082479 0.0091667 0.001389 0.98691 0.99168 2.9955e-006 1.1982e-005 0.15588 0.92158 0.90952 0.0013985 0.98888 0.51066 0.0018841 0.42692 1.9847 1.9839 16.0078 144.9537 0.00017494 -85.64 0.70694
5.811 0.9881 5.4861e-005 3.8183 0.011965 7.5885e-005 0.001163 0.23276 0.0006593 0.23341 0.21537 0 0.032306 0.0389 0 1.3439 0.45865 0.13946 0.017108 10.4145 0.10654 0.00013579 0.7836 0.0082484 0.0091673 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.15589 0.92177 0.9096 0.0013985 0.98893 0.51083 0.0018841 0.42694 1.9852 1.9845 16.0078 144.9538 0.00017481 -85.6402 0.70794
5.812 0.9881 5.4861e-005 3.8183 0.011965 7.5898e-005 0.001163 0.23276 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.344 0.45869 0.13948 0.01711 10.4167 0.10655 0.0001358 0.78359 0.008249 0.0091679 0.0013889 0.98691 0.99168 2.9953e-006 1.1981e-005 0.15589 0.92196 0.90968 0.0013985 0.98899 0.511 0.0018841 0.42695 1.9857 1.985 16.0078 144.9538 0.00017469 -85.6404 0.70894
5.813 0.9881 5.4861e-005 3.8183 0.011965 7.5911e-005 0.001163 0.23276 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.3441 0.45874 0.13949 0.017111 10.4189 0.10655 0.00013581 0.78358 0.0082495 0.0091685 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.1559 0.92215 0.90976 0.0013985 0.98904 0.51117 0.001884 0.42696 1.9863 1.9855 16.0077 144.9538 0.00017457 -85.6406 0.70994
5.814 0.9881 5.4861e-005 3.8183 0.011965 7.5923e-005 0.001163 0.23276 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.3442 0.45878 0.13951 0.017113 10.4211 0.10656 0.00013582 0.78357 0.0082501 0.0091691 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.1559 0.92235 0.90983 0.0013984 0.98909 0.51134 0.001884 0.42698 1.9868 1.986 16.0077 144.9538 0.00017445 -85.6407 0.71094
5.815 0.9881 5.4861e-005 3.8183 0.011965 7.5936e-005 0.001163 0.23277 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.3443 0.45883 0.13952 0.017114 10.4233 0.10657 0.00013583 0.78356 0.0082506 0.0091697 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.15591 0.92254 0.90991 0.0013984 0.98915 0.51151 0.001884 0.42699 1.9873 1.9865 16.0077 144.9538 0.00017433 -85.6409 0.71194
5.816 0.9881 5.4861e-005 3.8183 0.011965 7.5949e-005 0.001163 0.23277 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.3444 0.45888 0.13954 0.017115 10.4255 0.10658 0.00013585 0.78356 0.0082512 0.0091703 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.15591 0.92273 0.90999 0.0013984 0.9892 0.51168 0.0018839 0.427 1.9878 1.9871 16.0077 144.9539 0.0001742 -85.6411 0.71294
5.817 0.9881 5.486e-005 3.8183 0.011965 7.5962e-005 0.001163 0.23277 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.3445 0.45892 0.13956 0.017117 10.4277 0.10659 0.00013586 0.78355 0.0082517 0.0091709 0.0013888 0.98691 0.99168 2.9948e-006 1.1979e-005 0.15591 0.92292 0.91007 0.0013984 0.98925 0.51185 0.0018839 0.42702 1.9883 1.9876 16.0076 144.9539 0.00017408 -85.6413 0.71394
5.818 0.9881 5.486e-005 3.8183 0.011965 7.5975e-005 0.0011631 0.23277 0.0006593 0.23342 0.21537 0 0.032306 0.0389 0 1.3446 0.45897 0.13957 0.017118 10.4299 0.1066 0.00013587 0.78354 0.0082523 0.0091715 0.0013887 0.98691 0.99168 2.9948e-006 1.1979e-005 0.15592 0.92311 0.91014 0.0013984 0.9893 0.51202 0.0018839 0.42703 1.9888 1.9881 16.0076 144.9539 0.00017396 -85.6415 0.71494
5.819 0.9881 5.486e-005 3.8183 0.011965 7.5988e-005 0.0011631 0.23277 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3447 0.45902 0.13959 0.01712 10.4321 0.10661 0.00013588 0.78353 0.0082528 0.0091721 0.0013887 0.98691 0.99168 2.9947e-006 1.1978e-005 0.15592 0.9233 0.91022 0.0013983 0.98935 0.51219 0.0018839 0.42704 1.9893 1.9886 16.0076 144.9539 0.00017384 -85.6416 0.71594
5.82 0.9881 5.486e-005 3.8183 0.011965 7.6001e-005 0.0011631 0.23277 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3447 0.45906 0.1396 0.017121 10.4343 0.10661 0.0001359 0.78352 0.0082534 0.0091727 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.15593 0.92348 0.9103 0.0013983 0.9894 0.51236 0.0018838 0.42706 1.9898 1.9891 16.0076 144.9539 0.00017372 -85.6418 0.71694
5.821 0.9881 5.486e-005 3.8183 0.011965 7.6014e-005 0.0011631 0.23277 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3448 0.45911 0.13962 0.017122 10.4365 0.10662 0.00013591 0.78351 0.0082539 0.0091733 0.0013886 0.98691 0.99169 2.9945e-006 1.1978e-005 0.15593 0.92367 0.91037 0.0013983 0.98945 0.51253 0.0018838 0.42707 1.9904 1.9896 16.0075 144.954 0.00017361 -85.642 0.71794
5.822 0.9881 5.486e-005 3.8183 0.011965 7.6027e-005 0.0011631 0.23277 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3449 0.45915 0.13963 0.017124 10.4387 0.10663 0.00013592 0.78351 0.0082545 0.0091739 0.0013885 0.98691 0.99169 2.9944e-006 1.1977e-005 0.15594 0.92386 0.91045 0.0013983 0.9895 0.5127 0.0018838 0.42708 1.9909 1.9901 16.0075 144.954 0.00017349 -85.6421 0.71894
5.823 0.9881 5.486e-005 3.8183 0.011965 7.604e-005 0.0011631 0.23278 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.345 0.4592 0.13965 0.017125 10.4409 0.10664 0.00013593 0.7835 0.0082551 0.0091745 0.0013885 0.98692 0.99169 2.9943e-006 1.1977e-005 0.15594 0.92405 0.91053 0.0013983 0.98955 0.51287 0.0018838 0.4271 1.9914 1.9906 16.0075 144.954 0.00017337 -85.6423 0.71994
5.824 0.9881 5.486e-005 3.8183 0.011965 7.6053e-005 0.0011631 0.23278 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3451 0.45925 0.13966 0.017126 10.4431 0.10665 0.00013595 0.78349 0.0082556 0.0091751 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.15595 0.92423 0.9106 0.0013982 0.9896 0.51304 0.0018837 0.42711 1.9919 1.9911 16.0074 144.954 0.00017325 -85.6425 0.72094
5.825 0.9881 5.486e-005 3.8183 0.011965 7.6066e-005 0.0011631 0.23278 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3452 0.45929 0.13968 0.017128 10.4453 0.10666 0.00013596 0.78348 0.0082562 0.0091756 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.15595 0.92442 0.91068 0.0013982 0.98965 0.51321 0.0018837 0.42712 1.9924 1.9917 16.0074 144.954 0.00017313 -85.6426 0.72194
5.826 0.9881 5.486e-005 3.8183 0.011965 7.6079e-005 0.0011631 0.23278 0.0006593 0.23343 0.21538 0 0.032305 0.0389 0 1.3453 0.45934 0.13969 0.017129 10.4474 0.10666 0.00013597 0.78347 0.0082567 0.0091762 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.15595 0.9246 0.91075 0.0013982 0.9897 0.51337 0.0018837 0.42714 1.9929 1.9922 16.0074 144.9541 0.00017302 -85.6428 0.72294
5.827 0.9881 5.486e-005 3.8183 0.011965 7.6091e-005 0.0011631 0.23278 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.3454 0.45939 0.13971 0.017131 10.4496 0.10667 0.00013598 0.78346 0.0082573 0.0091768 0.0013884 0.98692 0.99169 2.9939e-006 1.1976e-005 0.15596 0.92479 0.91083 0.0013982 0.98975 0.51354 0.0018836 0.42715 1.9934 1.9927 16.0074 144.9541 0.0001729 -85.643 0.72394
5.828 0.9881 5.486e-005 3.8183 0.011965 7.6104e-005 0.0011631 0.23278 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.3455 0.45943 0.13972 0.017132 10.4518 0.10668 0.000136 0.78345 0.0082578 0.0091774 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.15596 0.92497 0.9109 0.0013982 0.9898 0.51371 0.0018836 0.42716 1.9939 1.9932 16.0073 144.9541 0.00017278 -85.6431 0.72494
5.829 0.9881 5.486e-005 3.8183 0.011965 7.6117e-005 0.0011631 0.23278 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.3456 0.45948 0.13974 0.017133 10.454 0.10669 0.00013601 0.78345 0.0082584 0.009178 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.15597 0.92515 0.91098 0.0013981 0.98985 0.51388 0.0018836 0.42718 1.9944 1.9937 16.0073 144.9541 0.00017267 -85.6433 0.72594
5.83 0.9881 5.4859e-005 3.8183 0.011965 7.613e-005 0.0011631 0.23278 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.3457 0.45953 0.13975 0.017135 10.4562 0.1067 0.00013602 0.78344 0.0082589 0.0091786 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.15597 0.92533 0.91105 0.0013981 0.98989 0.51405 0.0018836 0.42719 1.9949 1.9942 16.0073 144.9541 0.00017255 -85.6435 0.72694
5.831 0.9881 5.4859e-005 3.8183 0.011965 7.6143e-005 0.0011631 0.23279 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.3458 0.45957 0.13977 0.017136 10.4584 0.10671 0.00013603 0.78343 0.0082595 0.0091792 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.15598 0.92552 0.91112 0.0013981 0.98994 0.51422 0.0018835 0.4272 1.9954 1.9947 16.0073 144.9542 0.00017244 -85.6436 0.72794
5.832 0.9881 5.4859e-005 3.8183 0.011965 7.6156e-005 0.0011631 0.23279 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.3459 0.45962 0.13978 0.017138 10.4606 0.10672 0.00013604 0.78342 0.00826 0.0091798 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.15598 0.9257 0.9112 0.0013981 0.98999 0.51439 0.0018835 0.42722 1.9959 1.9952 16.0072 144.9542 0.00017232 -85.6438 0.72894
5.833 0.9881 5.4859e-005 3.8183 0.011965 7.6169e-005 0.0011631 0.23279 0.0006593 0.23344 0.21539 0 0.032305 0.0389 0 1.346 0.45966 0.1398 0.017139 10.4628 0.10672 0.00013606 0.78341 0.0082606 0.0091804 0.0013881 0.98692 0.99169 2.9934e-006 1.1973e-005 0.15598 0.92588 0.91127 0.0013981 0.99004 0.51456 0.0018835 0.42723 1.9964 1.9957 16.0072 144.9542 0.00017221 -85.6439 0.72994
5.834 0.9881 5.4859e-005 3.8183 0.011965 7.6182e-005 0.0011631 0.23279 0.0006593 0.23344 0.21539 0 0.032304 0.0389 0 1.3461 0.45971 0.13981 0.01714 10.465 0.10673 0.00013607 0.7834 0.0082611 0.009181 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.15599 0.92606 0.91134 0.001398 0.99008 0.51473 0.0018835 0.42724 1.9969 1.9962 16.0072 144.9542 0.0001721 -85.6441 0.73094
5.835 0.9881 5.4859e-005 3.8183 0.011965 7.6195e-005 0.0011631 0.23279 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3462 0.45976 0.13983 0.017142 10.4672 0.10674 0.00013608 0.78339 0.0082617 0.0091816 0.0013881 0.98692 0.99169 2.9932e-006 1.1973e-005 0.15599 0.92624 0.91142 0.001398 0.99013 0.5149 0.0018834 0.42726 1.9974 1.9967 16.0072 144.9542 0.00017198 -85.6443 0.73194
5.836 0.9881 5.4859e-005 3.8183 0.011965 7.6208e-005 0.0011631 0.23279 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3462 0.4598 0.13984 0.017143 10.4694 0.10675 0.00013609 0.78339 0.0082622 0.0091822 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.156 0.92642 0.91149 0.001398 0.99017 0.51507 0.0018834 0.42727 1.9979 1.9972 16.0071 144.9543 0.00017187 -85.6444 0.73294
5.837 0.9881 5.4859e-005 3.8183 0.011965 7.6221e-005 0.0011631 0.23279 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3463 0.45985 0.13986 0.017145 10.4716 0.10676 0.00013611 0.78338 0.0082628 0.0091828 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.156 0.9266 0.91156 0.001398 0.99022 0.51524 0.0018834 0.42728 1.9984 1.9976 16.0071 144.9543 0.00017176 -85.6446 0.73394
5.838 0.9881 5.4859e-005 3.8183 0.011965 7.6234e-005 0.0011631 0.23279 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3464 0.4599 0.13987 0.017146 10.4738 0.10677 0.00013612 0.78337 0.0082633 0.0091834 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.15601 0.92677 0.91163 0.001398 0.99027 0.5154 0.0018834 0.4273 1.9988 1.9981 16.0071 144.9543 0.00017165 -85.6447 0.73494
5.839 0.9881 5.4859e-005 3.8183 0.011965 7.6247e-005 0.0011631 0.2328 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3465 0.45994 0.13989 0.017147 10.476 0.10678 0.00013613 0.78336 0.0082639 0.009184 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.15601 0.92695 0.91171 0.0013979 0.99031 0.51557 0.0018833 0.42731 1.9993 1.9986 16.0071 144.9543 0.00017153 -85.6449 0.73594
5.84 0.9881 5.4859e-005 3.8183 0.011965 7.626e-005 0.0011631 0.2328 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3466 0.45999 0.1399 0.017149 10.4782 0.10678 0.00013614 0.78335 0.0082645 0.0091846 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.15601 0.92713 0.91178 0.0013979 0.99035 0.51574 0.0018833 0.42732 1.9998 1.9991 16.007 144.9544 0.00017142 -85.645 0.73694
5.841 0.9881 5.4859e-005 3.8183 0.011965 7.6272e-005 0.0011631 0.2328 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3467 0.46003 0.13992 0.01715 10.4804 0.10679 0.00013616 0.78334 0.008265 0.0091852 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.15602 0.9273 0.91185 0.0013979 0.9904 0.51591 0.0018833 0.42734 2.0003 1.9996 16.007 144.9544 0.00017131 -85.6452 0.73794
5.842 0.9881 5.4859e-005 3.8183 0.011965 7.6285e-005 0.0011631 0.2328 0.0006593 0.23345 0.2154 0 0.032304 0.0389 0 1.3468 0.46008 0.13993 0.017152 10.4826 0.1068 0.00013617 0.78333 0.0082656 0.0091858 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.15602 0.92748 0.91192 0.0013979 0.99044 0.51608 0.0018833 0.42735 2.0008 2.0001 16.007 144.9544 0.0001712 -85.6453 0.73894
5.843 0.9881 5.4858e-005 3.8183 0.011965 7.6298e-005 0.0011631 0.2328 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.3469 0.46013 0.13995 0.017153 10.4848 0.10681 0.00013618 0.78333 0.0082661 0.0091864 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.15603 0.92766 0.91199 0.0013979 0.99049 0.51625 0.0018832 0.42736 2.0013 2.0006 16.0069 144.9544 0.00017109 -85.6455 0.73994
5.844 0.9881 5.4858e-005 3.8183 0.011965 7.6311e-005 0.0011631 0.2328 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.347 0.46017 0.13996 0.017154 10.487 0.10682 0.00013619 0.78332 0.0082667 0.009187 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.15603 0.92783 0.91206 0.0013979 0.99053 0.51642 0.0018832 0.42737 2.0018 2.0011 16.0069 144.9544 0.00017098 -85.6456 0.74094
5.845 0.9881 5.4858e-005 3.8183 0.011965 7.6324e-005 0.0011631 0.2328 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.3471 0.46022 0.13998 0.017156 10.4892 0.10683 0.0001362 0.78331 0.0082672 0.0091876 0.0013877 0.98693 0.99169 2.9925e-006 1.197e-005 0.15604 0.928 0.91213 0.0013978 0.99057 0.51658 0.0018832 0.42739 2.0023 2.0016 16.0069 144.9545 0.00017087 -85.6458 0.74194
5.846 0.9881 5.4858e-005 3.8183 0.011965 7.6337e-005 0.0011631 0.23281 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.3472 0.46027 0.13999 0.017157 10.4914 0.10684 0.00013622 0.7833 0.0082678 0.0091881 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.15604 0.92818 0.9122 0.0013978 0.99062 0.51675 0.0018832 0.4274 2.0027 2.002 16.0069 144.9545 0.00017076 -85.6459 0.74294
5.847 0.9881 5.4858e-005 3.8183 0.011964 7.635e-005 0.0011632 0.23281 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.3473 0.46031 0.14001 0.017159 10.4937 0.10684 0.00013623 0.78329 0.0082683 0.0091887 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.15605 0.92835 0.91227 0.0013978 0.99066 0.51692 0.0018832 0.42741 2.0032 2.0025 16.0068 144.9545 0.00017066 -85.646 0.74394
5.848 0.9881 5.4858e-005 3.8183 0.011964 7.6363e-005 0.0011632 0.23281 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.3474 0.46036 0.14002 0.01716 10.4959 0.10685 0.00013624 0.78328 0.0082689 0.0091893 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.15605 0.92852 0.91234 0.0013978 0.9907 0.51709 0.0018831 0.42743 2.0037 2.003 16.0068 144.9545 0.00017055 -85.6462 0.74494
5.849 0.9881 5.4858e-005 3.8183 0.011964 7.6376e-005 0.0011632 0.23281 0.0006593 0.23346 0.21541 0 0.032304 0.0389 0 1.3475 0.4604 0.14004 0.017161 10.4981 0.10686 0.00013625 0.78328 0.0082694 0.0091899 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.15605 0.9287 0.91241 0.0013978 0.99074 0.51726 0.0018831 0.42744 2.0042 2.0035 16.0068 144.9545 0.00017044 -85.6463 0.74594
5.85 0.9881 5.4858e-005 3.8183 0.011964 7.6389e-005 0.0011632 0.23281 0.0006593 0.23346 0.21541 0 0.032303 0.0389 0 1.3476 0.46045 0.14005 0.017163 10.5003 0.10687 0.00013627 0.78327 0.00827 0.0091905 0.0013875 0.98693 0.99169 2.9921e-006 1.1968e-005 0.15606 0.92887 0.91248 0.0013977 0.99079 0.51743 0.0018831 0.42745 2.0047 2.004 16.0068 144.9546 0.00017033 -85.6465 0.74694
5.851 0.9881 5.4858e-005 3.8183 0.011964 7.6402e-005 0.0011632 0.23281 0.0006593 0.23347 0.21541 0 0.032303 0.0389 0 1.3477 0.4605 0.14007 0.017164 10.5025 0.10688 0.00013628 0.78326 0.0082705 0.0091911 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.15606 0.92904 0.91255 0.0013977 0.99083 0.51759 0.0018831 0.42747 2.0051 2.0044 16.0067 144.9546 0.00017022 -85.6466 0.74794
5.852 0.9881 5.4858e-005 3.8183 0.011964 7.6415e-005 0.0011632 0.23281 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.3477 0.46054 0.14008 0.017166 10.5047 0.10689 0.00013629 0.78325 0.0082711 0.0091917 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.15607 0.92921 0.91262 0.0013977 0.99087 0.51776 0.001883 0.42748 2.0056 2.0049 16.0067 144.9546 0.00017012 -85.6467 0.74894
5.853 0.9881 5.4858e-005 3.8183 0.011964 7.6428e-005 0.0011632 0.23281 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.3478 0.46059 0.1401 0.017167 10.5069 0.10689 0.0001363 0.78324 0.0082716 0.0091923 0.0013874 0.98693 0.99169 2.9919e-006 1.1967e-005 0.15607 0.92938 0.91268 0.0013977 0.99091 0.51793 0.001883 0.42749 2.0061 2.0054 16.0067 144.9546 0.00017001 -85.6469 0.74994
5.854 0.9881 5.4858e-005 3.8183 0.011964 7.644e-005 0.0011632 0.23282 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.3479 0.46064 0.14011 0.017168 10.5091 0.1069 0.00013632 0.78323 0.0082722 0.0091929 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.15608 0.92955 0.91275 0.0013977 0.99095 0.5181 0.001883 0.42751 2.0066 2.0059 16.0066 144.9546 0.00016991 -85.647 0.75094
5.855 0.9881 5.4858e-005 3.8183 0.011964 7.6453e-005 0.0011632 0.23282 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.348 0.46068 0.14013 0.01717 10.5113 0.10691 0.00013633 0.78322 0.0082727 0.0091935 0.0013874 0.98693 0.9917 2.9917e-006 1.1967e-005 0.15608 0.92972 0.91282 0.0013977 0.99099 0.51827 0.001883 0.42752 2.007 2.0064 16.0066 144.9547 0.0001698 -85.6472 0.75194
5.856 0.9881 5.4857e-005 3.8183 0.011964 7.6466e-005 0.0011632 0.23282 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.3481 0.46073 0.14014 0.017171 10.5135 0.10692 0.00013634 0.78322 0.0082733 0.0091941 0.0013874 0.98693 0.9917 2.9917e-006 1.1966e-005 0.15608 0.92988 0.91289 0.0013976 0.99103 0.51843 0.001883 0.42753 2.0075 2.0068 16.0066 144.9547 0.0001697 -85.6473 0.75294
5.857 0.9881 5.4857e-005 3.8183 0.011964 7.6479e-005 0.0011632 0.23282 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.3482 0.46077 0.14016 0.017172 10.5157 0.10693 0.00013635 0.78321 0.0082738 0.0091947 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.15609 0.93005 0.91296 0.0013976 0.99107 0.5186 0.0018829 0.42755 2.008 2.0073 16.0066 144.9547 0.00016959 -85.6474 0.75394
5.858 0.9881 5.4857e-005 3.8183 0.011964 7.6492e-005 0.0011632 0.23282 0.0006593 0.23347 0.21542 0 0.032303 0.0389 0 1.3483 0.46082 0.14017 0.017174 10.5179 0.10694 0.00013636 0.7832 0.0082744 0.0091953 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.15609 0.93022 0.91302 0.0013976 0.99111 0.51877 0.0018829 0.42756 2.0085 2.0078 16.0065 144.9547 0.00016949 -85.6476 0.75494
5.859 0.9881 5.4857e-005 3.8183 0.011964 7.6505e-005 0.0011632 0.23282 0.0006593 0.23348 0.21542 0 0.032303 0.0389 0 1.3484 0.46087 0.14019 0.017175 10.5201 0.10695 0.00013638 0.78319 0.0082749 0.0091959 0.0013873 0.98693 0.9917 2.9914e-006 1.1966e-005 0.1561 0.93039 0.91309 0.0013976 0.99115 0.51894 0.0018829 0.42757 2.0089 2.0082 16.0065 144.9547 0.00016938 -85.6477 0.75594
5.86 0.9881 5.4857e-005 3.8183 0.011964 7.6518e-005 0.0011632 0.23282 0.0006593 0.23348 0.21543 0 0.032303 0.0389 0 1.3485 0.46091 0.1402 0.017177 10.5223 0.10695 0.00013639 0.78318 0.0082755 0.0091965 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.1561 0.93055 0.91316 0.0013976 0.99119 0.5191 0.0018829 0.42759 2.0094 2.0087 16.0065 144.9548 0.00016928 -85.6478 0.75694
5.861 0.9881 5.4857e-005 3.8183 0.011964 7.6531e-005 0.0011632 0.23282 0.0006593 0.23348 0.21543 0 0.032303 0.0389 0 1.3486 0.46096 0.14022 0.017178 10.5245 0.10696 0.0001364 0.78317 0.008276 0.009197 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.15611 0.93072 0.91322 0.0013976 0.99123 0.51927 0.0018829 0.4276 2.0099 2.0092 16.0064 144.9548 0.00016917 -85.6479 0.75794
5.862 0.9881 5.4857e-005 3.8183 0.011964 7.6544e-005 0.0011632 0.23283 0.0006593 0.23348 0.21543 0 0.032303 0.0389 0 1.3487 0.46101 0.14023 0.017179 10.5268 0.10697 0.00013641 0.78317 0.0082766 0.0091976 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.15611 0.93088 0.91329 0.0013976 0.99127 0.51944 0.0018828 0.42761 2.0103 2.0097 16.0064 144.9548 0.00016907 -85.6481 0.75894
5.863 0.9881 5.4857e-005 3.8183 0.011964 7.6557e-005 0.0011632 0.23283 0.0006593 0.23348 0.21543 0 0.032303 0.0389 0 1.3488 0.46105 0.14025 0.017181 10.529 0.10698 0.00013643 0.78316 0.0082771 0.0091982 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.15611 0.93105 0.91336 0.0013975 0.99131 0.51961 0.0018828 0.42763 2.0108 2.0101 16.0064 144.9548 0.00016897 -85.6482 0.75994
5.864 0.9881 5.4857e-005 3.8183 0.011964 7.657e-005 0.0011632 0.23283 0.0006593 0.23348 0.21543 0 0.032303 0.0389 0 1.3489 0.4611 0.14026 0.017182 10.5312 0.10699 0.00013644 0.78315 0.0082777 0.0091988 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.15612 0.93121 0.91342 0.0013975 0.99134 0.51977 0.0018828 0.42764 2.0113 2.0106 16.0064 144.9548 0.00016887 -85.6483 0.76094
5.865 0.9881 5.4857e-005 3.8183 0.011964 7.6583e-005 0.0011632 0.23283 0.0006593 0.23348 0.21543 0 0.032303 0.0389 0 1.349 0.46115 0.14028 0.017184 10.5334 0.107 0.00013645 0.78314 0.0082782 0.0091994 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.15612 0.93137 0.91349 0.0013975 0.99138 0.51994 0.0018828 0.42765 2.0117 2.0111 16.0063 144.9549 0.00016876 -85.6485 0.76194
5.866 0.9881 5.4857e-005 3.8183 0.011964 7.6596e-005 0.0011632 0.23283 0.0006593 0.23348 0.21543 0 0.032302 0.0389 0 1.3491 0.46119 0.14029 0.017185 10.5356 0.10701 0.00013646 0.78313 0.0082788 0.0092 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.15613 0.93154 0.91355 0.0013975 0.99142 0.52011 0.0018828 0.42766 2.0122 2.0115 16.0063 144.9549 0.00016866 -85.6486 0.76294
5.867 0.9881 5.4857e-005 3.8183 0.011964 7.6609e-005 0.0011632 0.23283 0.0006593 0.23349 0.21543 0 0.032302 0.0389 0 1.3491 0.46124 0.14031 0.017186 10.5378 0.10701 0.00013648 0.78312 0.0082793 0.0092006 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.15613 0.9317 0.91362 0.0013975 0.99146 0.52028 0.0018827 0.42768 2.0126 2.012 16.0063 144.9549 0.00016856 -85.6487 0.76394
5.868 0.9881 5.4857e-005 3.8183 0.011964 7.6621e-005 0.0011632 0.23283 0.0006593 0.23349 0.21543 0 0.032302 0.0389 0 1.3492 0.46128 0.14032 0.017188 10.54 0.10702 0.00013649 0.78311 0.0082799 0.0092012 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.15614 0.93186 0.91368 0.0013975 0.99149 0.52044 0.0018827 0.42769 2.0131 2.0124 16.0063 144.9549 0.00016846 -85.6488 0.76494
5.869 0.9881 5.4856e-005 3.8183 0.011964 7.6634e-005 0.0011632 0.23283 0.0006593 0.23349 0.21544 0 0.032302 0.0389 0 1.3493 0.46133 0.14034 0.017189 10.5422 0.10703 0.0001365 0.78311 0.0082804 0.0092018 0.001387 0.98693 0.9917 2.9907e-006 1.1963e-005 0.15614 0.93202 0.91375 0.0013974 0.99153 0.52061 0.0018827 0.4277 2.0136 2.0129 16.0062 144.9549 0.00016836 -85.649 0.76594
5.87 0.9881 5.4856e-005 3.8183 0.011964 7.6647e-005 0.0011632 0.23284 0.0006593 0.23349 0.21544 0 0.032302 0.0389 0 1.3494 0.46138 0.14035 0.017191 10.5444 0.10704 0.00013651 0.7831 0.008281 0.0092024 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.15614 0.93218 0.91381 0.0013974 0.99157 0.52078 0.0018827 0.42772 2.014 2.0134 16.0062 144.955 0.00016826 -85.6491 0.76694
5.871 0.9881 5.4856e-005 3.8183 0.011964 7.666e-005 0.0011632 0.23284 0.0006593 0.23349 0.21544 0 0.032302 0.0389 0 1.3495 0.46142 0.14037 0.017192 10.5466 0.10705 0.00013652 0.78309 0.0082815 0.009203 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.15615 0.93234 0.91387 0.0013974 0.9916 0.52094 0.0018827 0.42773 2.0145 2.0138 16.0062 144.955 0.00016816 -85.6492 0.76794
5.872 0.9881 5.4856e-005 3.8183 0.011964 7.6673e-005 0.0011632 0.23284 0.0006593 0.23349 0.21544 0 0.032302 0.0389 0 1.3496 0.46147 0.14038 0.017193 10.5489 0.10706 0.00013654 0.78308 0.0082821 0.0092036 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.15615 0.9325 0.91394 0.0013974 0.99164 0.52111 0.0018826 0.42774 2.0149 2.0143 16.0061 144.955 0.00016806 -85.6493 0.76894
5.873 0.9881 5.4856e-005 3.8183 0.011964 7.6686e-005 0.0011632 0.23284 0.0006593 0.23349 0.21544 0 0.032302 0.0389 0 1.3497 0.46152 0.1404 0.017195 10.5511 0.10706 0.00013655 0.78307 0.0082826 0.0092042 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.15616 0.93266 0.914 0.0013974 0.99168 0.52128 0.0018826 0.42776 2.0154 2.0147 16.0061 144.955 0.00016796 -85.6494 0.76994
5.874 0.9881 5.4856e-005 3.8183 0.011964 7.6699e-005 0.0011632 0.23284 0.0006593 0.23349 0.21544 0 0.032302 0.0389 0 1.3498 0.46156 0.14041 0.017196 10.5533 0.10707 0.00013656 0.78306 0.0082832 0.0092047 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.15616 0.93282 0.91407 0.0013974 0.99171 0.52144 0.0018826 0.42777 2.0159 2.0152 16.0061 144.955 0.00016786 -85.6496 0.77094
5.875 0.9881 5.4856e-005 3.8183 0.011964 7.6712e-005 0.0011632 0.23284 0.0006593 0.2335 0.21544 0 0.032302 0.0389 0 1.3499 0.46161 0.14043 0.017197 10.5555 0.10708 0.00013657 0.78306 0.0082837 0.0092053 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.15617 0.93298 0.91413 0.0013974 0.99175 0.52161 0.0018826 0.42778 2.0163 2.0157 16.0061 144.9551 0.00016776 -85.6497 0.77194
5.876 0.9881 5.4856e-005 3.8183 0.011964 7.6725e-005 0.0011633 0.23284 0.0006593 0.2335 0.21544 0 0.032302 0.0389 0 1.35 0.46165 0.14044 0.017199 10.5577 0.10709 0.00013659 0.78305 0.0082843 0.0092059 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.15617 0.93314 0.91419 0.0013973 0.99178 0.52178 0.0018826 0.4278 2.0168 2.0161 16.006 144.9551 0.00016767 -85.6498 0.77294
5.877 0.9881 5.4856e-005 3.8183 0.011964 7.6738e-005 0.0011633 0.23284 0.0006593 0.2335 0.21545 0 0.032302 0.0389 0 1.3501 0.4617 0.14046 0.0172 10.5599 0.1071 0.0001366 0.78304 0.0082848 0.0092065 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.15617 0.9333 0.91425 0.0013973 0.99182 0.52194 0.0018825 0.42781 2.0172 2.0166 16.006 144.9551 0.00016757 -85.6499 0.77394
5.878 0.9881 5.4856e-005 3.8183 0.011964 7.6751e-005 0.0011633 0.23284 0.0006593 0.2335 0.21545 0 0.032302 0.0389 0 1.3502 0.46175 0.14047 0.017202 10.5621 0.10711 0.00013661 0.78303 0.0082854 0.0092071 0.0013867 0.98694 0.9917 2.9903e-006 1.1961e-005 0.15618 0.93345 0.91432 0.0013973 0.99185 0.52211 0.0018825 0.42782 2.0177 2.017 16.006 144.9551 0.00016747 -85.65 0.77494
5.879 0.9881 5.4856e-005 3.8183 0.011964 7.6764e-005 0.0011633 0.23285 0.0006593 0.2335 0.21545 0 0.032302 0.0389 0 1.3503 0.46179 0.14049 0.017203 10.5644 0.10712 0.00013662 0.78302 0.0082859 0.0092077 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.15618 0.93361 0.91438 0.0013973 0.99189 0.52228 0.0018825 0.42783 2.0181 2.0175 16.0059 144.9551 0.00016737 -85.6501 0.77594
5.88 0.9881 5.4856e-005 3.8183 0.011964 7.6777e-005 0.0011633 0.23285 0.0006593 0.2335 0.21545 0 0.032302 0.0389 0 1.3504 0.46184 0.1405 0.017204 10.5666 0.10712 0.00013664 0.78301 0.0082865 0.0092083 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.15619 0.93377 0.91444 0.0013973 0.99192 0.52244 0.0018825 0.42785 2.0186 2.0179 16.0059 144.9552 0.00016728 -85.6502 0.77694
5.881 0.9881 5.4856e-005 3.8183 0.011964 7.6789e-005 0.0011633 0.23285 0.0006593 0.2335 0.21545 0 0.032302 0.0389 0 1.3505 0.46189 0.14052 0.017206 10.5688 0.10713 0.00013665 0.783 0.008287 0.0092089 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.15619 0.93392 0.9145 0.0013973 0.99196 0.52261 0.0018825 0.42786 2.019 2.0184 16.0059 144.9552 0.00016718 -85.6504 0.77794
5.882 0.9881 5.4855e-005 3.8183 0.011964 7.6802e-005 0.0011633 0.23285 0.0006593 0.2335 0.21545 0 0.032301 0.0389 0 1.3506 0.46193 0.14053 0.017207 10.571 0.10714 0.00013666 0.783 0.0082876 0.0092095 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.1562 0.93408 0.91457 0.0013973 0.99199 0.52278 0.0018824 0.42787 2.0195 2.0188 16.0059 144.9552 0.00016708 -85.6505 0.77894
5.883 0.9881 5.4855e-005 3.8183 0.011964 7.6815e-005 0.0011633 0.23285 0.0006593 0.23351 0.21545 0 0.032301 0.0389 0 1.3506 0.46198 0.14055 0.017209 10.5732 0.10715 0.00013667 0.78299 0.0082881 0.0092101 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.1562 0.93423 0.91463 0.0013972 0.99202 0.52294 0.0018824 0.42789 2.0199 2.0193 16.0058 144.9552 0.00016699 -85.6506 0.77994
5.884 0.9881 5.4855e-005 3.8183 0.011964 7.6828e-005 0.0011633 0.23285 0.0006593 0.23351 0.21545 0 0.032301 0.0389 0 1.3507 0.46202 0.14056 0.01721 10.5754 0.10716 0.00013668 0.78298 0.0082887 0.0092107 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.1562 0.93439 0.91469 0.0013972 0.99206 0.52311 0.0018824 0.4279 2.0204 2.0197 16.0058 144.9553 0.00016689 -85.6507 0.78094
5.885 0.9881 5.4855e-005 3.8183 0.011964 7.6841e-005 0.0011633 0.23285 0.0006593 0.23351 0.21545 0 0.032301 0.0389 0 1.3508 0.46207 0.14058 0.017211 10.5777 0.10717 0.0001367 0.78297 0.0082892 0.0092112 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.15621 0.93454 0.91475 0.0013972 0.99209 0.52327 0.0018824 0.42791 2.0208 2.0202 16.0058 144.9553 0.0001668 -85.6508 0.78194
5.886 0.9881 5.4855e-005 3.8183 0.011964 7.6854e-005 0.0011633 0.23285 0.0006593 0.23351 0.21546 0 0.032301 0.0389 0 1.3509 0.46212 0.14059 0.017213 10.5799 0.10717 0.00013671 0.78296 0.0082898 0.0092118 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.15621 0.93469 0.91481 0.0013972 0.99212 0.52344 0.0018824 0.42793 2.0213 2.0206 16.0057 144.9553 0.0001667 -85.6509 0.78294
5.887 0.9881 5.4855e-005 3.8183 0.011964 7.6867e-005 0.0011633 0.23286 0.0006593 0.23351 0.21546 0 0.032301 0.0389 0 1.351 0.46216 0.14061 0.017214 10.5821 0.10718 0.00013672 0.78295 0.0082903 0.0092124 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.15622 0.93485 0.91487 0.0013972 0.99216 0.52361 0.0018824 0.42794 2.0217 2.0211 16.0057 144.9553 0.00016661 -85.651 0.78394
5.888 0.9881 5.4855e-005 3.8183 0.011964 7.688e-005 0.0011633 0.23286 0.0006593 0.23351 0.21546 0 0.032301 0.0389 0 1.3511 0.46221 0.14062 0.017216 10.5843 0.10719 0.00013673 0.78295 0.0082909 0.009213 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.15622 0.935 0.91493 0.0013972 0.99219 0.52377 0.0018823 0.42795 2.0221 2.0215 16.0057 144.9553 0.00016651 -85.6511 0.78494
5.889 0.9881 5.4855e-005 3.8183 0.011964 7.6893e-005 0.0011633 0.23286 0.0006593 0.23351 0.21546 0 0.032301 0.0389 0 1.3512 0.46226 0.14064 0.017217 10.5865 0.1072 0.00013675 0.78294 0.0082914 0.0092136 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.15623 0.93515 0.91499 0.0013972 0.99222 0.52394 0.0018823 0.42796 2.0226 2.0219 16.0057 144.9554 0.00016642 -85.6512 0.78594
5.89 0.9881 5.4855e-005 3.8183 0.011964 7.6906e-005 0.0011633 0.23286 0.0006593 0.23351 0.21546 0 0.032301 0.0389 0 1.3513 0.4623 0.14065 0.017218 10.5887 0.10721 0.00013676 0.78293 0.008292 0.0092142 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.15623 0.9353 0.91505 0.0013972 0.99225 0.5241 0.0018823 0.42798 2.023 2.0224 16.0056 144.9554 0.00016633 -85.6513 0.78694
5.891 0.9881 5.4855e-005 3.8183 0.011964 7.6919e-005 0.0011633 0.23286 0.0006593 0.23352 0.21546 0 0.032301 0.0389 0 1.3514 0.46235 0.14067 0.01722 10.591 0.10722 0.00013677 0.78292 0.0082925 0.0092148 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.15623 0.93545 0.91511 0.0013971 0.99229 0.52427 0.0018823 0.42799 2.0235 2.0228 16.0056 144.9554 0.00016623 -85.6514 0.78794
5.892 0.9881 5.4855e-005 3.8183 0.011964 7.6932e-005 0.0011633 0.23286 0.0006593 0.23352 0.21546 0 0.032301 0.0389 0 1.3515 0.46239 0.14068 0.017221 10.5932 0.10723 0.00013678 0.78291 0.008293 0.0092154 0.0013864 0.98694 0.9917 2.9893e-006 1.1957e-005 0.15624 0.9356 0.91517 0.0013971 0.99232 0.52444 0.0018823 0.428 2.0239 2.0233 16.0056 144.9554 0.00016614 -85.6515 0.78894
5.893 0.9881 5.4855e-005 3.8183 0.011964 7.6945e-005 0.0011633 0.23286 0.0006593 0.23352 0.21546 0 0.032301 0.0389 0 1.3516 0.46244 0.1407 0.017222 10.5954 0.10723 0.00013679 0.7829 0.0082936 0.009216 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.15624 0.93575 0.91523 0.0013971 0.99235 0.5246 0.0018823 0.42802 2.0243 2.0237 16.0055 144.9554 0.00016605 -85.6517 0.78994
5.894 0.9881 5.4855e-005 3.8183 0.011964 7.6957e-005 0.0011633 0.23286 0.0006593 0.23352 0.21547 0 0.032301 0.0389 0 1.3517 0.46249 0.14072 0.017224 10.5976 0.10724 0.00013681 0.78289 0.0082941 0.0092166 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.15625 0.9359 0.91529 0.0013971 0.99238 0.52477 0.0018822 0.42803 2.0248 2.0242 16.0055 144.9555 0.00016596 -85.6518 0.79094
5.895 0.9881 5.4854e-005 3.8183 0.011964 7.697e-005 0.0011633 0.23287 0.0006593 0.23352 0.21547 0 0.032301 0.0389 0 1.3518 0.46253 0.14073 0.017225 10.5998 0.10725 0.00013682 0.78289 0.0082947 0.0092171 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.15625 0.93605 0.91535 0.0013971 0.99241 0.52493 0.0018822 0.42804 2.0252 2.0246 16.0055 144.9555 0.00016586 -85.6519 0.79194
5.896 0.9881 5.4854e-005 3.8183 0.011964 7.6983e-005 0.0011633 0.23287 0.0006593 0.23352 0.21547 0 0.032301 0.0389 0 1.3519 0.46258 0.14075 0.017227 10.6021 0.10726 0.00013683 0.78288 0.0082952 0.0092177 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.15626 0.9362 0.91541 0.0013971 0.99244 0.5251 0.0018822 0.42806 2.0257 2.025 16.0055 144.9555 0.00016577 -85.652 0.79294
5.897 0.9881 5.4854e-005 3.8183 0.011964 7.6996e-005 0.0011633 0.23287 0.0006593 0.23352 0.21547 0 0.032301 0.0389 0 1.352 0.46263 0.14076 0.017228 10.6043 0.10727 0.00013684 0.78287 0.0082958 0.0092183 0.0013862 0.98694 0.9917 2.9891e-006 1.1956e-005 0.15626 0.93635 0.91547 0.0013971 0.99247 0.52526 0.0018822 0.42807 2.0261 2.0255 16.0054 144.9555 0.00016568 -85.6521 0.79394
5.898 0.9881 5.4854e-005 3.8183 0.011964 7.7009e-005 0.0011633 0.23287 0.0006593 0.23352 0.21547 0 0.032301 0.0389 0 1.352 0.46267 0.14078 0.017229 10.6065 0.10728 0.00013686 0.78286 0.0082963 0.0092189 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.15627 0.93649 0.91552 0.0013971 0.9925 0.52543 0.0018822 0.42808 2.0265 2.0259 16.0054 144.9555 0.00016559 -85.6522 0.79494
5.899 0.9881 5.4854e-005 3.8183 0.011964 7.7022e-005 0.0011633 0.23287 0.0006593 0.23353 0.21547 0 0.0323 0.0389 0 1.3521 0.46272 0.14079 0.017231 10.6087 0.10728 0.00013687 0.78285 0.0082969 0.0092195 0.0013862 0.98694 0.9917 2.9889e-006 1.1956e-005 0.15627 0.93664 0.91558 0.001397 0.99253 0.52559 0.0018822 0.42809 2.027 2.0263 16.0054 144.9556 0.0001655 -85.6523 0.79594
5.9 0.9881 5.4854e-005 3.8183 0.011964 7.7035e-005 0.0011633 0.23287 0.0006593 0.23353 0.21547 0 0.0323 0.0389 0 1.3522 0.46276 0.14081 0.017232 10.6109 0.10729 0.00013688 0.78284 0.0082974 0.0092201 0.0013862 0.98695 0.99171 2.9888e-006 1.1955e-005 0.15627 0.93679 0.91564 0.001397 0.99256 0.52576 0.0018821 0.42811 2.0274 2.0268 16.0053 144.9556 0.00016541 -85.6524 0.79694
5.901 0.9881 5.4854e-005 3.8183 0.011964 7.7048e-005 0.0011633 0.23287 0.0006593 0.23353 0.21547 0 0.0323 0.0389 0 1.3523 0.46281 0.14082 0.017234 10.6132 0.1073 0.00013689 0.78284 0.008298 0.0092207 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.15628 0.93693 0.9157 0.001397 0.99259 0.52592 0.0018821 0.42812 2.0278 2.0272 16.0053 144.9556 0.00016532 -85.6525 0.79794
5.902 0.9881 5.4854e-005 3.8183 0.011964 7.7061e-005 0.0011633 0.23287 0.0006593 0.23353 0.21547 0 0.0323 0.0389 0 1.3524 0.46286 0.14084 0.017235 10.6154 0.10731 0.0001369 0.78283 0.0082985 0.0092213 0.0013861 0.98695 0.99171 2.9886e-006 1.1955e-005 0.15628 0.93708 0.91576 0.001397 0.99262 0.52609 0.0018821 0.42813 2.0283 2.0276 16.0053 144.9556 0.00016523 -85.6526 0.79894
5.903 0.9881 5.4854e-005 3.8183 0.011964 7.7074e-005 0.0011633 0.23288 0.0006593 0.23353 0.21548 0 0.0323 0.0389 0 1.3525 0.4629 0.14085 0.017236 10.6176 0.10732 0.00013692 0.78282 0.0082991 0.0092219 0.0013861 0.98695 0.99171 2.9886e-006 1.1955e-005 0.15629 0.93722 0.91581 0.001397 0.99265 0.52625 0.0018821 0.42815 2.0287 2.0281 16.0053 144.9556 0.00016514 -85.6526 0.79994
5.904 0.9881 5.4854e-005 3.8183 0.011964 7.7087e-005 0.0011634 0.23288 0.0006593 0.23353 0.21548 0 0.0323 0.0389 0 1.3526 0.46295 0.14087 0.017238 10.6198 0.10733 0.00013693 0.78281 0.0082996 0.0092224 0.0013861 0.98695 0.99171 2.9886e-006 1.1955e-005 0.15629 0.93737 0.91587 0.001397 0.99268 0.52642 0.0018821 0.42816 2.0291 2.0285 16.0052 144.9557 0.00016505 -85.6527 0.80094
5.905 0.9881 5.4854e-005 3.8183 0.011964 7.71e-005 0.0011634 0.23288 0.0006593 0.23353 0.21548 0 0.0323 0.0389 0 1.3527 0.463 0.14088 0.017239 10.6221 0.10734 0.00013694 0.7828 0.0083002 0.009223 0.0013861 0.98695 0.99171 2.9886e-006 1.1954e-005 0.1563 0.93751 0.91593 0.001397 0.99271 0.52658 0.0018821 0.42817 2.0295 2.0289 16.0052 144.9557 0.00016496 -85.6528 0.80194
5.906 0.9881 5.4854e-005 3.8183 0.011964 7.7113e-005 0.0011634 0.23288 0.0006593 0.23353 0.21548 0 0.0323 0.0389 0 1.3528 0.46304 0.1409 0.01724 10.6243 0.10734 0.00013695 0.78279 0.0083007 0.0092236 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.1563 0.93766 0.91598 0.001397 0.99274 0.52675 0.0018821 0.42818 2.03 2.0294 16.0052 144.9557 0.00016487 -85.6529 0.80294
5.907 0.9881 5.4854e-005 3.8183 0.011964 7.7125e-005 0.0011634 0.23288 0.0006593 0.23353 0.21548 0 0.0323 0.0389 0 1.3529 0.46309 0.14091 0.017242 10.6265 0.10735 0.00013697 0.78278 0.0083013 0.0092242 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.1563 0.9378 0.91604 0.0013969 0.99277 0.52691 0.001882 0.4282 2.0304 2.0298 16.0051 144.9557 0.00016478 -85.653 0.80394
5.908 0.9881 5.4853e-005 3.8183 0.011963 7.7138e-005 0.0011634 0.23288 0.0006593 0.23354 0.21548 0 0.0323 0.0389 0 1.353 0.46313 0.14093 0.017243 10.6287 0.10736 0.00013698 0.78278 0.0083018 0.0092248 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.15631 0.93794 0.9161 0.0013969 0.9928 0.52708 0.001882 0.42821 2.0308 2.0302 16.0051 144.9557 0.0001647 -85.6531 0.80494
5.909 0.9881 5.4853e-005 3.8183 0.011963 7.7151e-005 0.0011634 0.23288 0.0006593 0.23354 0.21548 0 0.0323 0.0389 0 1.3531 0.46318 0.14094 0.017245 10.631 0.10737 0.00013699 0.78277 0.0083023 0.0092254 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.15631 0.93809 0.91615 0.0013969 0.99283 0.52724 0.001882 0.42822 2.0312 2.0306 16.0051 144.9558 0.00016461 -85.6532 0.80594
5.91 0.9881 5.4853e-005 3.8183 0.011963 7.7164e-005 0.0011634 0.23288 0.0006593 0.23354 0.21548 0 0.0323 0.0389 0 1.3532 0.46323 0.14096 0.017246 10.6332 0.10738 0.000137 0.78276 0.0083029 0.009226 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15632 0.93823 0.91621 0.0013969 0.99286 0.52741 0.001882 0.42824 2.0317 2.0311 16.005 144.9558 0.00016452 -85.6533 0.80694
5.911 0.9881 5.4853e-005 3.8183 0.011963 7.7177e-005 0.0011634 0.23288 0.0006593 0.23354 0.21548 0 0.0323 0.0389 0 1.3533 0.46327 0.14097 0.017247 10.6354 0.10739 0.00013702 0.78275 0.0083034 0.0092266 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15632 0.93837 0.91627 0.0013969 0.99288 0.52757 0.001882 0.42825 2.0321 2.0315 16.005 144.9558 0.00016443 -85.6534 0.80794
5.912 0.9881 5.4853e-005 3.8183 0.011963 7.719e-005 0.0011634 0.23289 0.0006593 0.23354 0.21549 0 0.0323 0.0389 0 1.3534 0.46332 0.14099 0.017249 10.6376 0.10739 0.00013703 0.78274 0.008304 0.0092272 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15633 0.93851 0.91632 0.0013969 0.99291 0.52774 0.001882 0.42826 2.0325 2.0319 16.005 144.9558 0.00016435 -85.6535 0.80894
5.913 0.9881 5.4853e-005 3.8183 0.011963 7.7203e-005 0.0011634 0.23289 0.0006593 0.23354 0.21549 0 0.0323 0.0389 0 1.3534 0.46337 0.141 0.01725 10.6399 0.1074 0.00013704 0.78273 0.0083045 0.0092277 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15633 0.93865 0.91638 0.0013969 0.99294 0.5279 0.001882 0.42827 2.0329 2.0323 16.005 144.9558 0.00016426 -85.6536 0.80994
5.914 0.9881 5.4853e-005 3.8183 0.011963 7.7216e-005 0.0011634 0.23289 0.0006593 0.23354 0.21549 0 0.0323 0.0389 0 1.3535 0.46341 0.14102 0.017252 10.6421 0.10741 0.00013705 0.78273 0.0083051 0.0092283 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15633 0.93879 0.91643 0.0013969 0.99297 0.52807 0.0018819 0.42829 2.0334 2.0328 16.0049 144.9559 0.00016417 -85.6537 0.81094
5.915 0.9881 5.4853e-005 3.8183 0.011963 7.7229e-005 0.0011634 0.23289 0.0006593 0.23354 0.21549 0 0.0323 0.0389 0 1.3536 0.46346 0.14103 0.017253 10.6443 0.10742 0.00013706 0.78272 0.0083056 0.0092289 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.15634 0.93893 0.91649 0.0013969 0.99299 0.52823 0.0018819 0.4283 2.0338 2.0332 16.0049 144.9559 0.00016409 -85.6537 0.81194
5.916 0.9881 5.4853e-005 3.8183 0.011963 7.7242e-005 0.0011634 0.23289 0.0006593 0.23355 0.21549 0 0.032299 0.0389 0 1.3537 0.4635 0.14105 0.017254 10.6465 0.10743 0.00013708 0.78271 0.0083062 0.0092295 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.15634 0.93907 0.91654 0.0013968 0.99302 0.52839 0.0018819 0.42831 2.0342 2.0336 16.0049 144.9559 0.000164 -85.6538 0.81294
5.917 0.9881 5.4853e-005 3.8183 0.011963 7.7255e-005 0.0011634 0.23289 0.0006593 0.23355 0.21549 0 0.032299 0.0389 0 1.3538 0.46355 0.14106 0.017256 10.6488 0.10744 0.00013709 0.7827 0.0083067 0.0092301 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.15635 0.93921 0.9166 0.0013968 0.99305 0.52856 0.0018819 0.42833 2.0346 2.034 16.0048 144.9559 0.00016392 -85.6539 0.81394
5.918 0.9881 5.4853e-005 3.8183 0.011963 7.7268e-005 0.0011634 0.23289 0.0006593 0.23355 0.21549 0 0.032299 0.0389 0 1.3539 0.4636 0.14108 0.017257 10.651 0.10744 0.0001371 0.78269 0.0083073 0.0092307 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.15635 0.93935 0.91665 0.0013968 0.99308 0.52872 0.0018819 0.42834 2.035 2.0344 16.0048 144.9559 0.00016383 -85.654 0.81494
5.919 0.9881 5.4853e-005 3.8183 0.011963 7.7281e-005 0.0011634 0.23289 0.0006593 0.23355 0.21549 0 0.032299 0.0389 0 1.354 0.46364 0.14109 0.017258 10.6532 0.10745 0.00013711 0.78268 0.0083078 0.0092313 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.15636 0.93949 0.91671 0.0013968 0.9931 0.52889 0.0018819 0.42835 2.0354 2.0349 16.0048 144.956 0.00016375 -85.6541 0.81594
5.92 0.9881 5.4853e-005 3.8183 0.011963 7.7293e-005 0.0011634 0.2329 0.0006593 0.23355 0.21549 0 0.032299 0.0389 0 1.3541 0.46369 0.14111 0.01726 10.6555 0.10746 0.00013713 0.78268 0.0083083 0.0092319 0.0013857 0.98695 0.99171 2.9878e-006 1.1952e-005 0.15636 0.93962 0.91676 0.0013968 0.99313 0.52905 0.0018819 0.42836 2.0359 2.0353 16.0048 144.956 0.00016366 -85.6542 0.81694
5.921 0.9881 5.4852e-005 3.8183 0.011963 7.7306e-005 0.0011634 0.2329 0.0006593 0.23355 0.2155 0 0.032299 0.0389 0 1.3542 0.46374 0.14112 0.017261 10.6577 0.10747 0.00013714 0.78267 0.0083089 0.0092324 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.15636 0.93976 0.91681 0.0013968 0.99315 0.52922 0.0018818 0.42838 2.0363 2.0357 16.0047 144.956 0.00016358 -85.6543 0.81794
5.922 0.9881 5.4852e-005 3.8183 0.011963 7.7319e-005 0.0011634 0.2329 0.0006593 0.23355 0.2155 0 0.032299 0.0389 0 1.3543 0.46378 0.14114 0.017263 10.6599 0.10748 0.00013715 0.78266 0.0083094 0.009233 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.15637 0.9399 0.91687 0.0013968 0.99318 0.52938 0.0018818 0.42839 2.0367 2.0361 16.0047 144.956 0.0001635 -85.6543 0.81894
5.923 0.9881 5.4852e-005 3.8183 0.011963 7.7332e-005 0.0011634 0.2329 0.0006593 0.23355 0.2155 0 0.032299 0.0389 0 1.3544 0.46383 0.14115 0.017264 10.6622 0.10749 0.00013716 0.78265 0.00831 0.0092336 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.15637 0.94003 0.91692 0.0013968 0.99321 0.52954 0.0018818 0.4284 2.0371 2.0365 16.0047 144.9561 0.00016341 -85.6544 0.81994
5.924 0.9881 5.4852e-005 3.8183 0.011963 7.7345e-005 0.0011634 0.2329 0.0006593 0.23355 0.2155 0 0.032299 0.0389 0 1.3545 0.46387 0.14117 0.017265 10.6644 0.1075 0.00013717 0.78264 0.0083105 0.0092342 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.15638 0.94017 0.91697 0.0013968 0.99323 0.52971 0.0018818 0.42842 2.0375 2.0369 16.0046 144.9561 0.00016333 -85.6545 0.82094
5.925 0.9881 5.4852e-005 3.8183 0.011963 7.7358e-005 0.0011634 0.2329 0.0006593 0.23356 0.2155 0 0.032299 0.0389 0 1.3546 0.46392 0.14118 0.017267 10.6666 0.1075 0.00013719 0.78263 0.0083111 0.0092348 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.15638 0.94031 0.91703 0.0013968 0.99326 0.52987 0.0018818 0.42843 2.0379 2.0373 16.0046 144.9561 0.00016325 -85.6546 0.82194
5.926 0.9881 5.4852e-005 3.8183 0.011963 7.7371e-005 0.0011634 0.2329 0.0006593 0.23356 0.2155 0 0.032299 0.0389 0 1.3547 0.46397 0.1412 0.017268 10.6688 0.10751 0.0001372 0.78262 0.0083116 0.0092354 0.0013856 0.98695 0.99171 2.9876e-006 1.1951e-005 0.15638 0.94044 0.91708 0.0013967 0.99328 0.53004 0.0018818 0.42844 2.0383 2.0378 16.0046 144.9561 0.00016316 -85.6547 0.82294
5.927 0.9881 5.4852e-005 3.8183 0.011963 7.7384e-005 0.0011634 0.2329 0.0006593 0.23356 0.2155 0 0.032299 0.0389 0 1.3548 0.46401 0.14121 0.01727 10.6711 0.10752 0.00013721 0.78262 0.0083122 0.009236 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.15639 0.94058 0.91713 0.0013967 0.99331 0.5302 0.0018818 0.42845 2.0388 2.0382 16.0045 144.9561 0.00016308 -85.6548 0.82394
5.928 0.9881 5.4852e-005 3.8183 0.011963 7.7397e-005 0.0011634 0.2329 0.0006593 0.23356 0.2155 0 0.032299 0.0389 0 1.3548 0.46406 0.14123 0.017271 10.6733 0.10753 0.00013722 0.78261 0.0083127 0.0092365 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.15639 0.94071 0.91719 0.0013967 0.99333 0.53036 0.0018818 0.42847 2.0392 2.0386 16.0045 144.9562 0.000163 -85.6548 0.82494
5.929 0.9881 5.4852e-005 3.8183 0.011963 7.741e-005 0.0011634 0.23291 0.0006593 0.23356 0.2155 0 0.032299 0.0389 0 1.3549 0.46411 0.14124 0.017272 10.6755 0.10754 0.00013724 0.7826 0.0083133 0.0092371 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.1564 0.94084 0.91724 0.0013967 0.99336 0.53053 0.0018817 0.42848 2.0396 2.039 16.0045 144.9562 0.00016292 -85.6549 0.82594
5.93 0.9881 5.4852e-005 3.8183 0.011963 7.7423e-005 0.0011634 0.23291 0.0006593 0.23356 0.21551 0 0.032299 0.0389 0 1.355 0.46415 0.14126 0.017274 10.6778 0.10755 0.00013725 0.78259 0.0083138 0.0092377 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.1564 0.94098 0.91729 0.0013967 0.99338 0.53069 0.0018817 0.42849 2.04 2.0394 16.0045 144.9562 0.00016284 -85.655 0.82694
5.931 0.9881 5.4852e-005 3.8183 0.011963 7.7436e-005 0.0011634 0.23291 0.0006593 0.23356 0.21551 0 0.032299 0.0389 0 1.3551 0.4642 0.14127 0.017275 10.68 0.10755 0.00013726 0.78258 0.0083143 0.0092383 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.15641 0.94111 0.91734 0.0013967 0.99341 0.53085 0.0018817 0.42851 2.0404 2.0398 16.0044 144.9562 0.00016275 -85.6551 0.82794
5.932 0.9881 5.4852e-005 3.8183 0.011963 7.7449e-005 0.0011634 0.23291 0.0006593 0.23356 0.21551 0 0.032299 0.0389 0 1.3552 0.46424 0.14129 0.017276 10.6822 0.10756 0.00013727 0.78257 0.0083149 0.0092389 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.15641 0.94124 0.91739 0.0013967 0.99343 0.53102 0.0018817 0.42852 2.0408 2.0402 16.0044 144.9562 0.00016267 -85.6552 0.82894
5.933 0.9881 5.4852e-005 3.8183 0.011963 7.7461e-005 0.0011635 0.23291 0.0006593 0.23357 0.21551 0 0.032298 0.0389 0 1.3553 0.46429 0.1413 0.017278 10.6845 0.10757 0.00013728 0.78257 0.0083154 0.0092395 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.15641 0.94137 0.91745 0.0013967 0.99346 0.53118 0.0018817 0.42853 2.0412 2.0406 16.0044 144.9563 0.00016259 -85.6552 0.82994
5.934 0.9881 5.4851e-005 3.8183 0.011963 7.7474e-005 0.0011635 0.23291 0.0006593 0.23357 0.21551 0 0.032298 0.0389 0 1.3554 0.46434 0.14132 0.017279 10.6867 0.10758 0.0001373 0.78256 0.008316 0.0092401 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.15642 0.94151 0.9175 0.0013967 0.99348 0.53134 0.0018817 0.42854 2.0416 2.041 16.0043 144.9563 0.00016251 -85.6553 0.83094
5.935 0.9881 5.4851e-005 3.8183 0.011963 7.7487e-005 0.0011635 0.23291 0.0006593 0.23357 0.21551 0 0.032298 0.0389 0 1.3555 0.46438 0.14133 0.017281 10.6889 0.10759 0.00013731 0.78255 0.0083165 0.0092406 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.15642 0.94164 0.91755 0.0013967 0.99351 0.53151 0.0018817 0.42856 2.042 2.0414 16.0043 144.9563 0.00016243 -85.6554 0.83194
5.936 0.9881 5.4851e-005 3.8183 0.011963 7.75e-005 0.0011635 0.23291 0.0006593 0.23357 0.21551 0 0.032298 0.0389 0 1.3556 0.46443 0.14135 0.017282 10.6912 0.1076 0.00013732 0.78254 0.0083171 0.0092412 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.15643 0.94177 0.9176 0.0013966 0.99353 0.53167 0.0018817 0.42857 2.0424 2.0418 16.0043 144.9563 0.00016235 -85.6555 0.83294
5.937 0.9881 5.4851e-005 3.8183 0.011963 7.7513e-005 0.0011635 0.23292 0.0006593 0.23357 0.21551 0 0.032298 0.0389 0 1.3557 0.46448 0.14136 0.017283 10.6934 0.1076 0.00013733 0.78253 0.0083176 0.0092418 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.15643 0.9419 0.91765 0.0013966 0.99355 0.53183 0.0018816 0.42858 2.0428 2.0422 16.0042 144.9563 0.00016227 -85.6555 0.83394
5.938 0.9881 5.4851e-005 3.8183 0.011963 7.7526e-005 0.0011635 0.23292 0.0006593 0.23357 0.21551 0 0.032298 0.0389 0 1.3558 0.46452 0.14138 0.017285 10.6956 0.10761 0.00013735 0.78252 0.0083182 0.0092424 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.15644 0.94203 0.9177 0.0013966 0.99358 0.532 0.0018816 0.4286 2.0432 2.0427 16.0042 144.9564 0.00016219 -85.6556 0.83494
5.939 0.9881 5.4851e-005 3.8183 0.011963 7.7539e-005 0.0011635 0.23292 0.0006593 0.23357 0.21552 0 0.032298 0.0389 0 1.3559 0.46457 0.14139 0.017286 10.6979 0.10762 0.00013736 0.78252 0.0083187 0.009243 0.0013854 0.98695 0.99171 2.9871e-006 1.1949e-005 0.15644 0.94216 0.91775 0.0013966 0.9936 0.53216 0.0018816 0.42861 2.0436 2.0431 16.0042 144.9564 0.00016211 -85.6557 0.83594
5.94 0.9881 5.4851e-005 3.8183 0.011963 7.7552e-005 0.0011635 0.23292 0.0006593 0.23357 0.21552 0 0.032298 0.0389 0 1.356 0.46461 0.14141 0.017287 10.7001 0.10763 0.00013737 0.78251 0.0083192 0.0092436 0.0013854 0.98696 0.99171 2.987e-006 1.1948e-005 0.15644 0.94229 0.9178 0.0013966 0.99362 0.53232 0.0018816 0.42862 2.044 2.0435 16.0041 144.9564 0.00016203 -85.6558 0.83694
5.941 0.9881 5.4851e-005 3.8183 0.011963 7.7565e-005 0.0011635 0.23292 0.0006593 0.23357 0.21552 0 0.032298 0.0389 0 1.3561 0.46466 0.14142 0.017289 10.7024 0.10764 0.00013738 0.7825 0.0083198 0.0092442 0.0013854 0.98696 0.99171 2.987e-006 1.1948e-005 0.15645 0.94242 0.91785 0.0013966 0.99365 0.53248 0.0018816 0.42863 2.0444 2.0439 16.0041 144.9564 0.00016196 -85.6558 0.83794
5.942 0.9881 5.4851e-005 3.8183 0.011963 7.7578e-005 0.0011635 0.23292 0.0006593 0.23358 0.21552 0 0.032298 0.0389 0 1.3562 0.46471 0.14144 0.01729 10.7046 0.10765 0.00013739 0.78249 0.0083203 0.0092447 0.0013854 0.98696 0.99171 2.987e-006 1.1948e-005 0.15645 0.94255 0.9179 0.0013966 0.99367 0.53265 0.0018816 0.42865 2.0448 2.0443 16.0041 144.9564 0.00016188 -85.6559 0.83894
5.943 0.9881 5.4851e-005 3.8183 0.011963 7.7591e-005 0.0011635 0.23292 0.0006593 0.23358 0.21552 0 0.032298 0.0389 0 1.3562 0.46475 0.14145 0.017292 10.7068 0.10766 0.00013741 0.78248 0.0083209 0.0092453 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.15646 0.94267 0.91795 0.0013966 0.99369 0.53281 0.0018816 0.42866 2.0452 2.0447 16.0041 144.9565 0.0001618 -85.656 0.83994
5.944 0.9881 5.4851e-005 3.8183 0.011963 7.7604e-005 0.0011635 0.23292 0.0006593 0.23358 0.21552 0 0.032298 0.0389 0 1.3563 0.4648 0.14147 0.017293 10.7091 0.10766 0.00013742 0.78247 0.0083214 0.0092459 0.0013853 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15646 0.9428 0.918 0.0013966 0.99372 0.53297 0.0018816 0.42867 2.0456 2.0451 16.004 144.9565 0.00016172 -85.656 0.84094
5.945 0.9881 5.4851e-005 3.8183 0.011963 7.7617e-005 0.0011635 0.23292 0.0006593 0.23358 0.21552 0 0.032298 0.0389 0 1.3564 0.46485 0.14148 0.017294 10.7113 0.10767 0.00013743 0.78247 0.008322 0.0092465 0.0013853 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15647 0.94293 0.91805 0.0013966 0.99374 0.53314 0.0018815 0.42868 2.046 2.0455 16.004 144.9565 0.00016164 -85.6561 0.84194
5.946 0.9881 5.4851e-005 3.8183 0.011963 7.7629e-005 0.0011635 0.23293 0.0006593 0.23358 0.21552 0 0.032298 0.0389 0 1.3565 0.46489 0.1415 0.017296 10.7135 0.10768 0.00013744 0.78246 0.0083225 0.0092471 0.0013853 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15647 0.94306 0.9181 0.0013966 0.99376 0.5333 0.0018815 0.4287 2.0464 2.0459 16.004 144.9565 0.00016157 -85.6562 0.84294
5.947 0.9881 5.485e-005 3.8183 0.011963 7.7642e-005 0.0011635 0.23293 0.0006593 0.23358 0.21552 0 0.032298 0.0389 0 1.3566 0.46494 0.14151 0.017297 10.7158 0.10769 0.00013746 0.78245 0.008323 0.0092477 0.0013853 0.98696 0.99171 2.9871e-006 1.1948e-005 0.15647 0.94318 0.91815 0.0013966 0.99378 0.53346 0.0018815 0.42871 2.0468 2.0462 16.0039 144.9565 0.00016149 -85.6563 0.84394
5.948 0.9881 5.485e-005 3.8183 0.011963 7.7655e-005 0.0011635 0.23293 0.0006593 0.23358 0.21553 0 0.032298 0.0389 0 1.3567 0.46498 0.14153 0.017299 10.718 0.1077 0.00013747 0.78244 0.0083236 0.0092483 0.0013853 0.98696 0.99171 2.987e-006 1.1947e-005 0.15648 0.94331 0.9182 0.0013965 0.9938 0.53362 0.0018815 0.42872 2.0472 2.0466 16.0039 144.9566 0.00016141 -85.6563 0.84494
5.949 0.9881 5.485e-005 3.8183 0.011963 7.7668e-005 0.0011635 0.23293 0.0006593 0.23358 0.21553 0 0.032298 0.0389 0 1.3568 0.46503 0.14154 0.0173 10.7203 0.10771 0.00013748 0.78243 0.0083241 0.0092488 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.15648 0.94343 0.91825 0.0013965 0.99383 0.53379 0.0018815 0.42873 2.0476 2.047 16.0039 144.9566 0.00016134 -85.6564 0.84594
5.95 0.9881 5.485e-005 3.8183 0.011963 7.7681e-005 0.0011635 0.23293 0.0006593 0.23358 0.21553 0 0.032297 0.0389 0 1.3569 0.46508 0.14156 0.017301 10.7225 0.10771 0.00013749 0.78242 0.0083247 0.0092494 0.0013852 0.98696 0.99171 2.9869e-006 1.1947e-005 0.15649 0.94356 0.9183 0.0013965 0.99385 0.53395 0.0018815 0.42875 2.048 2.0474 16.0038 144.9566 0.00016126 -85.6565 0.84694
5.951 0.9881 5.485e-005 3.8183 0.011963 7.7694e-005 0.0011635 0.23293 0.0006593 0.23359 0.21553 0 0.032297 0.0389 0 1.357 0.46512 0.14157 0.017303 10.7247 0.10772 0.0001375 0.78241 0.0083252 0.00925 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.15649 0.94368 0.91835 0.0013965 0.99387 0.53411 0.0018815 0.42876 2.0484 2.0478 16.0038 144.9566 0.00016118 -85.6565 0.84794
5.952 0.9881 5.485e-005 3.8183 0.011963 7.7707e-005 0.0011635 0.23293 0.0006593 0.23359 0.21553 0 0.032297 0.0389 0 1.3571 0.46517 0.14159 0.017304 10.727 0.10773 0.00013752 0.78241 0.0083258 0.0092506 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.1565 0.94381 0.9184 0.0013965 0.99389 0.53427 0.0018815 0.42877 2.0488 2.0482 16.0038 144.9566 0.00016111 -85.6566 0.84894
5.953 0.9881 5.485e-005 3.8183 0.011963 7.772e-005 0.0011635 0.23293 0.0006593 0.23359 0.21553 0 0.032297 0.0389 0 1.3572 0.46522 0.1416 0.017305 10.7292 0.10774 0.00013753 0.7824 0.0083263 0.0092512 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.1565 0.94393 0.91845 0.0013965 0.99391 0.53444 0.0018815 0.42879 2.0492 2.0486 16.0038 144.9567 0.00016103 -85.6567 0.84994
5.954 0.9881 5.485e-005 3.8183 0.011963 7.7733e-005 0.0011635 0.23293 0.0006593 0.23359 0.21553 0 0.032297 0.0389 0 1.3573 0.46526 0.14162 0.017307 10.7315 0.10775 0.00013754 0.78239 0.0083268 0.0092518 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.1565 0.94406 0.91849 0.0013965 0.99393 0.5346 0.0018814 0.4288 2.0496 2.049 16.0037 144.9567 0.00016096 -85.6567 0.85094
5.955 0.9881 5.485e-005 3.8183 0.011963 7.7746e-005 0.0011635 0.23294 0.0006593 0.23359 0.21553 0 0.032297 0.0389 0 1.3574 0.46531 0.14163 0.017308 10.7337 0.10776 0.00013755 0.78238 0.0083274 0.0092523 0.0013852 0.98696 0.99171 2.9867e-006 1.1946e-005 0.15651 0.94418 0.91854 0.0013965 0.99395 0.53476 0.0018814 0.42881 2.0499 2.0494 16.0037 144.9567 0.00016088 -85.6568 0.85194
5.956 0.9881 5.485e-005 3.8183 0.011963 7.7759e-005 0.0011635 0.23294 0.0006593 0.23359 0.21553 0 0.032297 0.0389 0 1.3575 0.46535 0.14165 0.01731 10.7359 0.10776 0.00013757 0.78237 0.0083279 0.0092529 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.15651 0.9443 0.91859 0.0013965 0.99398 0.53492 0.0018814 0.42882 2.0503 2.0498 16.0037 144.9567 0.00016081 -85.6569 0.85294
5.957 0.9881 5.485e-005 3.8183 0.011963 7.7772e-005 0.0011635 0.23294 0.0006593 0.23359 0.21554 0 0.032297 0.0389 0 1.3576 0.4654 0.14166 0.017311 10.7382 0.10777 0.00013758 0.78236 0.0083285 0.0092535 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.15652 0.94443 0.91864 0.0013965 0.994 0.53508 0.0018814 0.42884 2.0507 2.0502 16.0036 144.9568 0.00016073 -85.6569 0.85394
5.958 0.9881 5.485e-005 3.8183 0.011963 7.7784e-005 0.0011635 0.23294 0.0006593 0.23359 0.21554 0 0.032297 0.0389 0 1.3576 0.46545 0.14168 0.017312 10.7404 0.10778 0.00013759 0.78236 0.008329 0.0092541 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.15652 0.94455 0.91869 0.0013965 0.99402 0.53525 0.0018814 0.42885 2.0511 2.0506 16.0036 144.9568 0.00016066 -85.657 0.85494
5.959 0.9881 5.485e-005 3.8183 0.011963 7.7797e-005 0.0011635 0.23294 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3577 0.46549 0.14169 0.017314 10.7427 0.10779 0.0001376 0.78235 0.0083296 0.0092547 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.15653 0.94467 0.91873 0.0013965 0.99404 0.53541 0.0018814 0.42886 2.0515 2.051 16.0036 144.9568 0.00016059 -85.6571 0.85594
5.96 0.9881 5.485e-005 3.8183 0.011963 7.781e-005 0.0011635 0.23294 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3578 0.46554 0.14171 0.017315 10.7449 0.1078 0.00013761 0.78234 0.0083301 0.0092553 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.15653 0.94479 0.91878 0.0013964 0.99406 0.53557 0.0018814 0.42887 2.0519 2.0513 16.0035 144.9568 0.00016051 -85.6571 0.85694
5.961 0.9881 5.4849e-005 3.8183 0.011963 7.7823e-005 0.0011636 0.23294 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3579 0.46559 0.14172 0.017316 10.7472 0.10781 0.00013763 0.78233 0.0083306 0.0092558 0.0013851 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15653 0.94491 0.91883 0.0013964 0.99408 0.53573 0.0018814 0.42889 2.0523 2.0517 16.0035 144.9568 0.00016044 -85.6572 0.85794
5.962 0.9881 5.4849e-005 3.8183 0.011963 7.7836e-005 0.0011636 0.23294 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.358 0.46563 0.14174 0.017318 10.7494 0.10782 0.00013764 0.78232 0.0083312 0.0092564 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15654 0.94503 0.91887 0.0013964 0.9941 0.53589 0.0018814 0.4289 2.0527 2.0521 16.0035 144.9569 0.00016036 -85.6572 0.85894
5.963 0.9881 5.4849e-005 3.8183 0.011963 7.7849e-005 0.0011636 0.23294 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3581 0.46568 0.14175 0.017319 10.7516 0.10782 0.00013765 0.78231 0.0083317 0.009257 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15654 0.94515 0.91892 0.0013964 0.99412 0.53605 0.0018814 0.42891 2.053 2.0525 16.0034 144.9569 0.00016029 -85.6573 0.85994
5.964 0.9881 5.4849e-005 3.8183 0.011963 7.7862e-005 0.0011636 0.23295 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3582 0.46572 0.14177 0.017321 10.7539 0.10783 0.00013766 0.78231 0.0083323 0.0092576 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.15655 0.94527 0.91897 0.0013964 0.99414 0.53622 0.0018813 0.42892 2.0534 2.0529 16.0034 144.9569 0.00016022 -85.6574 0.86094
5.965 0.9881 5.4849e-005 3.8183 0.011963 7.7875e-005 0.0011636 0.23295 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3583 0.46577 0.14178 0.017322 10.7561 0.10784 0.00013767 0.7823 0.0083328 0.0092582 0.001385 0.98696 0.99171 2.9864e-006 1.1945e-005 0.15655 0.94539 0.91901 0.0013964 0.99416 0.53638 0.0018813 0.42894 2.0538 2.0533 16.0034 144.9569 0.00016015 -85.6574 0.86194
5.966 0.9881 5.4849e-005 3.8183 0.011963 7.7888e-005 0.0011636 0.23295 0.0006593 0.2336 0.21554 0 0.032297 0.0389 0 1.3584 0.46582 0.1418 0.017323 10.7584 0.10785 0.00013769 0.78229 0.0083333 0.0092588 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.15656 0.94551 0.91906 0.0013964 0.99418 0.53654 0.0018813 0.42895 2.0542 2.0536 16.0033 144.9569 0.00016007 -85.6575 0.86294
5.967 0.9881 5.4849e-005 3.8183 0.011963 7.7901e-005 0.0011636 0.23295 0.0006593 0.2336 0.21555 0 0.032297 0.0389 0 1.3585 0.46586 0.14181 0.017325 10.7606 0.10786 0.0001377 0.78228 0.0083339 0.0092593 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.15656 0.94563 0.91911 0.0013964 0.9942 0.5367 0.0018813 0.42896 2.0546 2.054 16.0033 144.957 0.00016 -85.6575 0.86394
5.968 0.9881 5.4849e-005 3.8183 0.011963 7.7914e-005 0.0011636 0.23295 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.3586 0.46591 0.14183 0.017326 10.7629 0.10787 0.00013771 0.78227 0.0083344 0.0092599 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.15656 0.94575 0.91915 0.0013964 0.99422 0.53686 0.0018813 0.42897 2.055 2.0544 16.0033 144.957 0.00015993 -85.6576 0.86494
5.969 0.9881 5.4849e-005 3.8183 0.011962 7.7927e-005 0.0011636 0.23295 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.3587 0.46596 0.14184 0.017327 10.7651 0.10787 0.00013772 0.78226 0.008335 0.0092605 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.15657 0.94587 0.9192 0.0013964 0.99424 0.53702 0.0018813 0.42899 2.0553 2.0548 16.0033 144.957 0.00015986 -85.6577 0.86594
5.97 0.9881 5.4849e-005 3.8183 0.011962 7.794e-005 0.0011636 0.23295 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.3588 0.466 0.14186 0.017329 10.7674 0.10788 0.00013774 0.78226 0.0083355 0.0092611 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.15657 0.94599 0.91924 0.0013964 0.99426 0.53718 0.0018813 0.429 2.0557 2.0552 16.0032 144.957 0.00015979 -85.6577 0.86694
5.971 0.9881 5.4849e-005 3.8183 0.011962 7.7952e-005 0.0011636 0.23295 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.3589 0.46605 0.14187 0.01733 10.7696 0.10789 0.00013775 0.78225 0.0083361 0.0092617 0.0013849 0.98696 0.99172 2.9858e-006 1.1944e-005 0.15658 0.9461 0.91929 0.0013964 0.99427 0.53735 0.0018813 0.42901 2.0561 2.0556 16.0032 144.957 0.00015972 -85.6578 0.86794
5.972 0.9881 5.4849e-005 3.8183 0.011962 7.7965e-005 0.0011636 0.23295 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.359 0.46609 0.14189 0.017332 10.7719 0.1079 0.00013776 0.78224 0.0083366 0.0092623 0.0013849 0.98696 0.99172 2.9858e-006 1.1944e-005 0.15658 0.94622 0.91933 0.0013964 0.99429 0.53751 0.0018813 0.42903 2.0565 2.0559 16.0032 144.9571 0.00015965 -85.6578 0.86894
5.973 0.9881 5.4849e-005 3.8183 0.011962 7.7978e-005 0.0011636 0.23296 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.359 0.46614 0.1419 0.017333 10.7741 0.10791 0.00013777 0.78223 0.0083371 0.0092628 0.0013849 0.98696 0.99172 2.9858e-006 1.1944e-005 0.15659 0.94634 0.91938 0.0013964 0.99431 0.53767 0.0018813 0.42904 2.0568 2.0563 16.0031 144.9571 0.00015958 -85.6579 0.86994
5.974 0.9881 5.4848e-005 3.8183 0.011962 7.7991e-005 0.0011636 0.23296 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.3591 0.46619 0.14192 0.017334 10.7764 0.10792 0.00013778 0.78222 0.0083377 0.0092634 0.0013849 0.98696 0.99172 2.9858e-006 1.1944e-005 0.15659 0.94645 0.91942 0.0013963 0.99433 0.53783 0.0018813 0.42905 2.0572 2.0567 16.0031 144.9571 0.0001595 -85.658 0.87094
5.975 0.9881 5.4848e-005 3.8183 0.011962 7.8004e-005 0.0011636 0.23296 0.0006593 0.23361 0.21555 0 0.032296 0.0389 0 1.3592 0.46623 0.14193 0.017336 10.7786 0.10792 0.0001378 0.78221 0.0083382 0.009264 0.0013849 0.98696 0.99172 2.9858e-006 1.1944e-005 0.15659 0.94657 0.91947 0.0013963 0.99435 0.53799 0.0018812 0.42906 2.0576 2.0571 16.0031 144.9571 0.00015943 -85.658 0.87194
5.976 0.9881 5.4848e-005 3.8183 0.011962 7.8017e-005 0.0011636 0.23296 0.0006593 0.23361 0.21556 0 0.032296 0.0389 0 1.3593 0.46628 0.14195 0.017337 10.7808 0.10793 0.00013781 0.78221 0.0083388 0.0092646 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.1566 0.94668 0.91951 0.0013963 0.99437 0.53815 0.0018812 0.42908 2.058 2.0574 16.003 144.9571 0.00015936 -85.6581 0.87294
5.977 0.9881 5.4848e-005 3.8183 0.011962 7.803e-005 0.0011636 0.23296 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3594 0.46633 0.14196 0.017338 10.7831 0.10794 0.00013782 0.7822 0.0083393 0.0092652 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.1566 0.9468 0.91956 0.0013963 0.99439 0.53831 0.0018812 0.42909 2.0583 2.0578 16.003 144.9572 0.0001593 -85.6581 0.87394
5.978 0.9881 5.4848e-005 3.8183 0.011962 7.8043e-005 0.0011636 0.23296 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3595 0.46637 0.14198 0.01734 10.7853 0.10795 0.00013783 0.78219 0.0083398 0.0092658 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15661 0.94691 0.9196 0.0013963 0.9944 0.53847 0.0018812 0.4291 2.0587 2.0582 16.003 144.9572 0.00015923 -85.6582 0.87494
5.979 0.9881 5.4848e-005 3.8183 0.011962 7.8056e-005 0.0011636 0.23296 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3596 0.46642 0.14199 0.017341 10.7876 0.10796 0.00013785 0.78218 0.0083404 0.0092663 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15661 0.94703 0.91965 0.0013963 0.99442 0.53863 0.0018812 0.42911 2.0591 2.0586 16.0029 144.9572 0.00015916 -85.6582 0.87594
5.98 0.9881 5.4848e-005 3.8183 0.011962 7.8069e-005 0.0011636 0.23296 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3597 0.46646 0.14201 0.017343 10.7898 0.10797 0.00013786 0.78217 0.0083409 0.0092669 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15661 0.94714 0.91969 0.0013963 0.99444 0.53879 0.0018812 0.42913 2.0595 2.0589 16.0029 144.9572 0.00015909 -85.6583 0.87694
5.981 0.9881 5.4848e-005 3.8183 0.011962 7.8082e-005 0.0011636 0.23296 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3598 0.46651 0.14202 0.017344 10.7921 0.10797 0.00013787 0.78216 0.0083415 0.0092675 0.0013848 0.98696 0.99172 2.9856e-006 1.1943e-005 0.15662 0.94726 0.91974 0.0013963 0.99446 0.53895 0.0018812 0.42914 2.0598 2.0593 16.0029 144.9572 0.00015902 -85.6583 0.87794
5.982 0.9881 5.4848e-005 3.8183 0.011962 7.8095e-005 0.0011636 0.23297 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3599 0.46656 0.14204 0.017345 10.7943 0.10798 0.00013788 0.78216 0.008342 0.0092681 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15662 0.94737 0.91978 0.0013963 0.99447 0.53912 0.0018812 0.42915 2.0602 2.0597 16.0028 144.9573 0.00015895 -85.6584 0.87894
5.983 0.9881 5.4848e-005 3.8183 0.011962 7.8107e-005 0.0011636 0.23297 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.36 0.4666 0.14205 0.017347 10.7966 0.10799 0.00013789 0.78215 0.0083425 0.0092687 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15663 0.94748 0.91982 0.0013963 0.99449 0.53928 0.0018812 0.42916 2.0606 2.0601 16.0028 144.9573 0.00015888 -85.6584 0.87994
5.984 0.9881 5.4848e-005 3.8183 0.011962 7.812e-005 0.0011636 0.23297 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3601 0.46665 0.14207 0.017348 10.7989 0.108 0.00013791 0.78214 0.0083431 0.0092692 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15663 0.9476 0.91987 0.0013963 0.99451 0.53944 0.0018812 0.42918 2.061 2.0604 16.0028 144.9573 0.00015881 -85.6585 0.88094
5.985 0.9881 5.4848e-005 3.8183 0.011962 7.8133e-005 0.0011636 0.23297 0.0006593 0.23362 0.21556 0 0.032296 0.0389 0 1.3602 0.4667 0.14208 0.017349 10.8011 0.10801 0.00013792 0.78213 0.0083436 0.0092698 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15664 0.94771 0.91991 0.0013963 0.99453 0.5396 0.0018812 0.42919 2.0613 2.0608 16.0028 144.9573 0.00015875 -85.6585 0.88194
5.986 0.9881 5.4848e-005 3.8183 0.011962 7.8146e-005 0.0011636 0.23297 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3603 0.46674 0.1421 0.017351 10.8034 0.10802 0.00013793 0.78212 0.0083442 0.0092704 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.15664 0.94782 0.91995 0.0013963 0.99454 0.53976 0.0018811 0.4292 2.0617 2.0612 16.0027 144.9573 0.00015868 -85.6586 0.88294
5.987 0.9881 5.4847e-005 3.8183 0.011962 7.8159e-005 0.0011636 0.23297 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3603 0.46679 0.14211 0.017352 10.8056 0.10802 0.00013794 0.78211 0.0083447 0.009271 0.0013847 0.98696 0.99172 2.9857e-006 1.1942e-005 0.15664 0.94793 0.92 0.0013963 0.99456 0.53992 0.0018811 0.42921 2.0621 2.0615 16.0027 144.9574 0.00015861 -85.6587 0.88394
5.988 0.9881 5.4847e-005 3.8183 0.011962 7.8172e-005 0.0011636 0.23297 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3604 0.46683 0.14213 0.017354 10.8079 0.10803 0.00013795 0.7821 0.0083452 0.0092716 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.15665 0.94804 0.92004 0.0013963 0.99458 0.54008 0.0018811 0.42923 2.0624 2.0619 16.0027 144.9574 0.00015854 -85.6587 0.88494
5.989 0.9881 5.4847e-005 3.8183 0.011962 7.8185e-005 0.0011637 0.23297 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3605 0.46688 0.14214 0.017355 10.8101 0.10804 0.00013797 0.7821 0.0083458 0.0092721 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.15665 0.94815 0.92008 0.0013962 0.9946 0.54024 0.0018811 0.42924 2.0628 2.0623 16.0026 144.9574 0.00015848 -85.6588 0.88594
5.99 0.9881 5.4847e-005 3.8183 0.011962 7.8198e-005 0.0011637 0.23297 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3606 0.46693 0.14216 0.017356 10.8124 0.10805 0.00013798 0.78209 0.0083463 0.0092727 0.0013847 0.98696 0.99172 2.9854e-006 1.1942e-005 0.15666 0.94826 0.92013 0.0013962 0.99461 0.5404 0.0018811 0.42925 2.0632 2.0626 16.0026 144.9574 0.00015841 -85.6588 0.88694
5.991 0.9881 5.4847e-005 3.8183 0.011962 7.8211e-005 0.0011637 0.23298 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3607 0.46697 0.14217 0.017358 10.8146 0.10806 0.00013799 0.78208 0.0083469 0.0092733 0.0013847 0.98696 0.99172 2.9853e-006 1.1942e-005 0.15666 0.94838 0.92017 0.0013962 0.99463 0.54056 0.0018811 0.42926 2.0635 2.063 16.0026 144.9574 0.00015834 -85.6589 0.88794
5.992 0.9881 5.4847e-005 3.8183 0.011962 7.8224e-005 0.0011637 0.23298 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3608 0.46702 0.14219 0.017359 10.8169 0.10807 0.000138 0.78207 0.0083474 0.0092739 0.0013847 0.98696 0.99172 2.9854e-006 1.1942e-005 0.15667 0.94848 0.92021 0.0013962 0.99465 0.54072 0.0018811 0.42928 2.0639 2.0634 16.0025 144.9575 0.00015828 -85.6589 0.88894
5.993 0.9881 5.4847e-005 3.8183 0.011962 7.8237e-005 0.0011637 0.23298 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.3609 0.46706 0.1422 0.01736 10.8191 0.10807 0.00013802 0.78206 0.0083479 0.0092745 0.0013847 0.98696 0.99172 2.9854e-006 1.1942e-005 0.15667 0.94859 0.92025 0.0013962 0.99466 0.54088 0.0018811 0.42929 2.0643 2.0637 16.0025 144.9575 0.00015821 -85.659 0.88994
5.994 0.9881 5.4847e-005 3.8183 0.011962 7.825e-005 0.0011637 0.23298 0.0006593 0.23363 0.21557 0 0.032295 0.0389 0 1.361 0.46711 0.14222 0.017362 10.8214 0.10808 0.00013803 0.78205 0.0083485 0.0092751 0.0013846 0.98696 0.99172 2.9855e-006 1.1942e-005 0.15667 0.9487 0.92029 0.0013962 0.99468 0.54104 0.0018811 0.4293 2.0646 2.0641 16.0025 144.9575 0.00015815 -85.659 0.89094
5.995 0.9881 5.4847e-005 3.8183 0.011962 7.8262e-005 0.0011637 0.23298 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3611 0.46716 0.14223 0.017363 10.8236 0.10809 0.00013804 0.78205 0.008349 0.0092756 0.0013846 0.98696 0.99172 2.9857e-006 1.1942e-005 0.15668 0.94881 0.92034 0.0013962 0.99469 0.5412 0.0018811 0.42931 2.065 2.0645 16.0024 144.9575 0.00015808 -85.659 0.89194
5.996 0.9881 5.4847e-005 3.8183 0.011962 7.8275e-005 0.0011637 0.23298 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3612 0.4672 0.14225 0.017365 10.8259 0.1081 0.00013805 0.78204 0.0083496 0.0092762 0.0013846 0.98697 0.99172 2.9857e-006 1.1942e-005 0.15668 0.94892 0.92038 0.0013962 0.99471 0.54136 0.0018811 0.42933 2.0653 2.0648 16.0024 144.9576 0.00015802 -85.6591 0.89294
5.997 0.9881 5.4847e-005 3.8183 0.011962 7.8288e-005 0.0011637 0.23298 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3613 0.46725 0.14226 0.017366 10.8282 0.10811 0.00013806 0.78203 0.0083501 0.0092768 0.0013846 0.98697 0.99172 2.9857e-006 1.1942e-005 0.15669 0.94903 0.92042 0.0013962 0.99473 0.54152 0.0018811 0.42934 2.0657 2.0652 16.0024 144.9576 0.00015795 -85.6591 0.89394
5.998 0.9881 5.4847e-005 3.8183 0.011962 7.8301e-005 0.0011637 0.23298 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3614 0.4673 0.14228 0.017367 10.8304 0.10812 0.00013808 0.78202 0.0083506 0.0092774 0.0013846 0.98697 0.99172 2.9856e-006 1.1941e-005 0.15669 0.94914 0.92046 0.0013962 0.99474 0.54168 0.0018811 0.42935 2.0661 2.0656 16.0023 144.9576 0.00015789 -85.6592 0.89494
5.999 0.9881 5.4847e-005 3.8183 0.011962 7.8314e-005 0.0011637 0.23298 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3615 0.46734 0.14229 0.017369 10.8327 0.10813 0.00013809 0.78201 0.0083512 0.009278 0.0013846 0.98697 0.99172 2.9855e-006 1.1941e-005 0.1567 0.94924 0.9205 0.0013962 0.99476 0.54184 0.001881 0.42936 2.0664 2.0659 16.0023 144.9576 0.00015782 -85.6592 0.89594
6 0.9881 5.4846e-005 3.8183 0.011962 7.8327e-005 0.0011637 0.23299 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3616 0.46739 0.14231 0.01737 10.8349 0.10813 0.0001381 0.782 0.0083517 0.0092785 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.1567 0.94935 0.92054 0.0013962 0.99477 0.542 0.001881 0.42937 2.0668 2.0663 16.0023 144.9576 0.00015776 -85.6593 0.89694
6.001 0.9881 5.4846e-005 3.8183 0.011962 7.834e-005 0.0011637 0.23299 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3617 0.46743 0.14232 0.017371 10.8372 0.10814 0.00013811 0.782 0.0083522 0.0092791 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.1567 0.94946 0.92059 0.0013962 0.99479 0.54216 0.001881 0.42939 2.0671 2.0666 16.0022 144.9577 0.00015769 -85.6593 0.89794
6.002 0.9881 5.4846e-005 3.8183 0.011962 7.8353e-005 0.0011637 0.23299 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3617 0.46748 0.14234 0.017373 10.8394 0.10815 0.00013812 0.78199 0.0083528 0.0092797 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.15671 0.94957 0.92063 0.0013962 0.99481 0.54232 0.001881 0.4294 2.0675 2.067 16.0022 144.9577 0.00015763 -85.6594 0.89894
6.003 0.9881 5.4846e-005 3.8183 0.011962 7.8366e-005 0.0011637 0.23299 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3618 0.46753 0.14235 0.017374 10.8417 0.10816 0.00013814 0.78198 0.0083533 0.0092803 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.15671 0.94967 0.92067 0.0013962 0.99482 0.54247 0.001881 0.42941 2.0679 2.0674 16.0022 144.9577 0.00015756 -85.6594 0.89994
6.004 0.9881 5.4846e-005 3.8183 0.011962 7.8379e-005 0.0011637 0.23299 0.0006593 0.23364 0.21558 0 0.032295 0.0389 0 1.3619 0.46757 0.14237 0.017375 10.844 0.10817 0.00013815 0.78197 0.0083539 0.0092809 0.0013845 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15672 0.94978 0.92071 0.0013962 0.99484 0.54263 0.001881 0.42942 2.0682 2.0677 16.0021 144.9577 0.0001575 -85.6595 0.90094
6.005 0.9881 5.4846e-005 3.8183 0.011962 7.8392e-005 0.0011637 0.23299 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.362 0.46762 0.14238 0.017377 10.8462 0.10818 0.00013816 0.78196 0.0083544 0.0092814 0.0013845 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15672 0.94988 0.92075 0.0013962 0.99485 0.54279 0.001881 0.42944 2.0686 2.0681 16.0021 144.9577 0.00015744 -85.6595 0.90194
6.006 0.9881 5.4846e-005 3.8183 0.011962 7.8405e-005 0.0011637 0.23299 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3621 0.46767 0.1424 0.017378 10.8485 0.10818 0.00013817 0.78195 0.0083549 0.009282 0.0013845 0.98697 0.99172 2.9853e-006 1.1941e-005 0.15672 0.94999 0.92079 0.0013961 0.99487 0.54295 0.001881 0.42945 2.0689 2.0684 16.0021 144.9578 0.00015737 -85.6596 0.90294
6.007 0.9881 5.4846e-005 3.8183 0.011962 7.8418e-005 0.0011637 0.23299 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3622 0.46771 0.14241 0.01738 10.8507 0.10819 0.00013819 0.78195 0.0083555 0.0092826 0.0013845 0.98697 0.99172 2.9852e-006 1.194e-005 0.15673 0.95009 0.92083 0.0013961 0.99488 0.54311 0.001881 0.42946 2.0693 2.0688 16.002 144.9578 0.00015731 -85.6596 0.90394
6.008 0.9881 5.4846e-005 3.8183 0.011962 7.843e-005 0.0011637 0.23299 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3623 0.46776 0.14243 0.017381 10.853 0.1082 0.0001382 0.78194 0.008356 0.0092832 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.15673 0.9502 0.92087 0.0013961 0.9949 0.54327 0.001881 0.42947 2.0696 2.0691 16.002 144.9578 0.00015725 -85.6596 0.90494
6.009 0.9881 5.4846e-005 3.8183 0.011962 7.8443e-005 0.0011637 0.233 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3624 0.4678 0.14244 0.017382 10.8552 0.10821 0.00013821 0.78193 0.0083566 0.0092837 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.15674 0.9503 0.92091 0.0013961 0.99491 0.54343 0.001881 0.42949 2.07 2.0695 16.002 144.9578 0.00015719 -85.6597 0.90594
6.01 0.9881 5.4846e-005 3.8183 0.011962 7.8456e-005 0.0011637 0.233 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3625 0.46785 0.14246 0.017384 10.8575 0.10822 0.00013822 0.78192 0.0083571 0.0092843 0.0013845 0.98697 0.99172 2.9849e-006 1.194e-005 0.15674 0.95041 0.92095 0.0013961 0.99493 0.54359 0.001881 0.4295 2.0704 2.0699 16.002 144.9578 0.00015712 -85.6597 0.90694
6.011 0.9881 5.4846e-005 3.8183 0.011962 7.8469e-005 0.0011637 0.233 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3626 0.4679 0.14247 0.017385 10.8598 0.10823 0.00013823 0.78191 0.0083576 0.0092849 0.0013845 0.98697 0.99172 2.9849e-006 1.194e-005 0.15675 0.95051 0.92099 0.0013961 0.99494 0.54375 0.001881 0.42951 2.0707 2.0702 16.0019 144.9579 0.00015706 -85.6598 0.90794
6.012 0.9881 5.4846e-005 3.8183 0.011962 7.8482e-005 0.0011637 0.233 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3627 0.46794 0.14248 0.017386 10.862 0.10823 0.00013825 0.7819 0.0083582 0.0092855 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.15675 0.95061 0.92103 0.0013961 0.99495 0.54391 0.001881 0.42952 2.0711 2.0706 16.0019 144.9579 0.000157 -85.6598 0.90894
6.013 0.9881 5.4845e-005 3.8183 0.011962 7.8495e-005 0.0011637 0.233 0.0006593 0.23365 0.21559 0 0.032294 0.0389 0 1.3628 0.46799 0.1425 0.017388 10.8643 0.10824 0.00013826 0.7819 0.0083587 0.0092861 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.15675 0.95072 0.92107 0.0013961 0.99497 0.54407 0.0018809 0.42954 2.0714 2.0709 16.0019 144.9579 0.00015694 -85.6599 0.90994
6.014 0.9881 5.4845e-005 3.8183 0.011962 7.8508e-005 0.0011637 0.233 0.0006593 0.23366 0.21559 0 0.032294 0.0389 0 1.3629 0.46804 0.14251 0.017389 10.8666 0.10825 0.00013827 0.78189 0.0083592 0.0092866 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.15676 0.95082 0.92111 0.0013961 0.99498 0.54422 0.0018809 0.42955 2.0718 2.0713 16.0018 144.9579 0.00015688 -85.6599 0.91094
6.015 0.9881 5.4845e-005 3.8183 0.011962 7.8521e-005 0.0011637 0.233 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.363 0.46808 0.14253 0.017391 10.8688 0.10826 0.00013828 0.78188 0.0083598 0.0092872 0.0013844 0.98697 0.99172 2.9851e-006 1.194e-005 0.15676 0.95092 0.92115 0.0013961 0.995 0.54438 0.0018809 0.42956 2.0721 2.0716 16.0018 144.9579 0.00015681 -85.6599 0.91194
6.016 0.9881 5.4845e-005 3.8183 0.011962 7.8534e-005 0.0011637 0.233 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.363 0.46813 0.14254 0.017392 10.8711 0.10827 0.00013829 0.78187 0.0083603 0.0092878 0.0013844 0.98697 0.99172 2.9852e-006 1.194e-005 0.15677 0.95102 0.92119 0.0013961 0.99501 0.54454 0.0018809 0.42957 2.0725 2.072 16.0018 144.958 0.00015675 -85.66 0.91294
6.017 0.9881 5.4845e-005 3.8183 0.011962 7.8547e-005 0.0011638 0.233 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.3631 0.46817 0.14256 0.017393 10.8733 0.10828 0.00013831 0.78186 0.0083609 0.0092884 0.0013844 0.98697 0.99172 2.9851e-006 1.194e-005 0.15677 0.95112 0.92122 0.0013961 0.99503 0.5447 0.0018809 0.42959 2.0728 2.0723 16.0017 144.958 0.00015669 -85.66 0.91394
6.018 0.9881 5.4845e-005 3.8183 0.011962 7.856e-005 0.0011638 0.23301 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.3632 0.46822 0.14257 0.017395 10.8756 0.10828 0.00013832 0.78185 0.0083614 0.009289 0.0013844 0.98697 0.99172 2.9851e-006 1.194e-005 0.15678 0.95122 0.92126 0.0013961 0.99504 0.54486 0.0018809 0.4296 2.0732 2.0727 16.0017 144.958 0.00015663 -85.6601 0.91494
6.019 0.9881 5.4845e-005 3.8183 0.011962 7.8573e-005 0.0011638 0.23301 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.3633 0.46827 0.14259 0.017396 10.8779 0.10829 0.00013833 0.78185 0.0083619 0.0092895 0.0013844 0.98697 0.99172 2.985e-006 1.1939e-005 0.15678 0.95133 0.9213 0.0013961 0.99505 0.54502 0.0018809 0.42961 2.0735 2.073 16.0017 144.958 0.00015657 -85.6601 0.91594
6.02 0.9881 5.4845e-005 3.8183 0.011962 7.8585e-005 0.0011638 0.23301 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.3634 0.46831 0.1426 0.017397 10.8801 0.1083 0.00013834 0.78184 0.0083625 0.0092901 0.0013844 0.98697 0.99172 2.985e-006 1.1939e-005 0.15678 0.95143 0.92134 0.0013961 0.99507 0.54518 0.0018809 0.42962 2.0739 2.0734 16.0016 144.958 0.00015651 -85.6601 0.91694
6.021 0.9881 5.4845e-005 3.8183 0.011962 7.8598e-005 0.0011638 0.23301 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.3635 0.46836 0.14262 0.017399 10.8824 0.10831 0.00013836 0.78183 0.008363 0.0092907 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.15679 0.95153 0.92138 0.0013961 0.99508 0.54534 0.0018809 0.42963 2.0742 2.0737 16.0016 144.9581 0.00015645 -85.6602 0.91794
6.022 0.9881 5.4845e-005 3.8183 0.011962 7.8611e-005 0.0011638 0.23301 0.0006593 0.23366 0.2156 0 0.032294 0.0389 0 1.3636 0.4684 0.14263 0.0174 10.8847 0.10832 0.00013837 0.78182 0.0083635 0.0092913 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.15679 0.95163 0.92142 0.0013961 0.99509 0.54549 0.0018809 0.42965 2.0746 2.0741 16.0016 144.9581 0.00015639 -85.6602 0.91894
6.023 0.9881 5.4845e-005 3.8183 0.011962 7.8624e-005 0.0011638 0.23301 0.0006593 0.23367 0.2156 0 0.032293 0.0389 0 1.3637 0.46845 0.14265 0.017402 10.8869 0.10833 0.00013838 0.78181 0.0083641 0.0092918 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.1568 0.95173 0.92146 0.0013961 0.99511 0.54565 0.0018809 0.42966 2.0749 2.0744 16.0015 144.9581 0.00015633 -85.6603 0.91994
6.024 0.9881 5.4845e-005 3.8183 0.011962 7.8637e-005 0.0011638 0.23301 0.0006593 0.23367 0.2156 0 0.032293 0.0389 0 1.3638 0.4685 0.14266 0.017403 10.8892 0.10833 0.00013839 0.7818 0.0083646 0.0092924 0.0013843 0.98697 0.99172 2.9849e-006 1.1939e-005 0.1568 0.95183 0.92149 0.0013961 0.99512 0.54581 0.0018809 0.42967 2.0752 2.0748 16.0015 144.9581 0.00015627 -85.6603 0.92094
6.025 0.9881 5.4845e-005 3.8183 0.011962 7.865e-005 0.0011638 0.23301 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3639 0.46854 0.14268 0.017404 10.8915 0.10834 0.0001384 0.7818 0.0083651 0.009293 0.0013843 0.98697 0.99172 2.9849e-006 1.1939e-005 0.1568 0.95193 0.92153 0.0013961 0.99514 0.54597 0.0018809 0.42968 2.0756 2.0751 16.0015 144.9581 0.00015621 -85.6603 0.92194
6.026 0.9881 5.4844e-005 3.8183 0.011962 7.8663e-005 0.0011638 0.23301 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.364 0.46859 0.14269 0.017406 10.8937 0.10835 0.00013842 0.78179 0.0083657 0.0092936 0.0013843 0.98697 0.99172 2.9848e-006 1.1939e-005 0.15681 0.95202 0.92157 0.0013961 0.99515 0.54613 0.0018809 0.4297 2.0759 2.0755 16.0014 144.9582 0.00015615 -85.6604 0.92294
6.027 0.9881 5.4844e-005 3.8183 0.011962 7.8676e-005 0.0011638 0.23301 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3641 0.46864 0.14271 0.017407 10.896 0.10836 0.00013843 0.78178 0.0083662 0.0092942 0.0013843 0.98697 0.99172 2.9848e-006 1.1939e-005 0.15681 0.95212 0.92161 0.001396 0.99516 0.54628 0.0018809 0.42971 2.0763 2.0758 16.0014 144.9582 0.00015609 -85.6604 0.92394
6.028 0.9881 5.4844e-005 3.8183 0.011962 7.8689e-005 0.0011638 0.23302 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3642 0.46868 0.14272 0.017408 10.8983 0.10837 0.00013844 0.78177 0.0083668 0.0092947 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.15682 0.95222 0.92165 0.001396 0.99517 0.54644 0.0018809 0.42972 2.0766 2.0761 16.0014 144.9582 0.00015604 -85.6604 0.92494
6.029 0.9881 5.4844e-005 3.8183 0.011962 7.8702e-005 0.0011638 0.23302 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3643 0.46873 0.14274 0.01741 10.9005 0.10838 0.00013845 0.78176 0.0083673 0.0092953 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.15682 0.95232 0.92168 0.001396 0.99519 0.5466 0.0018808 0.42973 2.077 2.0765 16.0013 144.9582 0.00015598 -85.6605 0.92594
6.03 0.9881 5.4844e-005 3.8183 0.011961 7.8715e-005 0.0011638 0.23302 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3643 0.46877 0.14275 0.017411 10.9028 0.10838 0.00013846 0.78175 0.0083678 0.0092959 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15683 0.95242 0.92172 0.001396 0.9952 0.54676 0.0018808 0.42974 2.0773 2.0768 16.0013 144.9583 0.00015592 -85.6605 0.92694
6.031 0.9881 5.4844e-005 3.8183 0.011961 7.8728e-005 0.0011638 0.23302 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3644 0.46882 0.14277 0.017412 10.9051 0.10839 0.00013848 0.78175 0.0083684 0.0092965 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15683 0.95251 0.92176 0.001396 0.99521 0.54692 0.0018808 0.42976 2.0777 2.0772 16.0013 144.9583 0.00015586 -85.6605 0.92794
6.032 0.9881 5.4844e-005 3.8183 0.011961 7.874e-005 0.0011638 0.23302 0.0006593 0.23367 0.21561 0 0.032293 0.0389 0 1.3645 0.46887 0.14278 0.017414 10.9073 0.1084 0.00013849 0.78174 0.0083689 0.009297 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15683 0.95261 0.92179 0.001396 0.99523 0.54707 0.0018808 0.42977 2.078 2.0775 16.0012 144.9583 0.0001558 -85.6606 0.92894
6.033 0.9881 5.4844e-005 3.8183 0.011961 7.8753e-005 0.0011638 0.23302 0.0006593 0.23368 0.21561 0 0.032293 0.0389 0 1.3646 0.46891 0.1428 0.017415 10.9096 0.10841 0.0001385 0.78173 0.0083694 0.0092976 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.15684 0.95271 0.92183 0.001396 0.99524 0.54723 0.0018808 0.42978 2.0783 2.0779 16.0012 144.9583 0.00015574 -85.6606 0.92994
6.034 0.9881 5.4844e-005 3.8183 0.011961 7.8766e-005 0.0011638 0.23302 0.0006593 0.23368 0.21561 0 0.032293 0.0389 0 1.3647 0.46896 0.14281 0.017417 10.9119 0.10842 0.00013851 0.78172 0.00837 0.0092982 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.15684 0.9528 0.92187 0.001396 0.99525 0.54739 0.0018808 0.42979 2.0787 2.0782 16.0012 144.9583 0.00015569 -85.6607 0.93094
6.035 0.9881 5.4844e-005 3.8183 0.011961 7.8779e-005 0.0011638 0.23302 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3648 0.46901 0.14283 0.017418 10.9141 0.10843 0.00013852 0.78171 0.0083705 0.0092988 0.0013843 0.98697 0.99172 2.9847e-006 1.1938e-005 0.15685 0.9529 0.9219 0.001396 0.99526 0.54755 0.0018808 0.42981 2.079 2.0785 16.0011 144.9584 0.00015563 -85.6607 0.93194
6.036 0.9881 5.4844e-005 3.8183 0.011961 7.8792e-005 0.0011638 0.23302 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3649 0.46905 0.14284 0.017419 10.9164 0.10843 0.00013854 0.7817 0.008371 0.0092993 0.0013842 0.98697 0.99172 2.9847e-006 1.1938e-005 0.15685 0.953 0.92194 0.001396 0.99528 0.5477 0.0018808 0.42982 2.0794 2.0789 16.0011 144.9584 0.00015557 -85.6607 0.93294
6.037 0.9881 5.4844e-005 3.8183 0.011961 7.8805e-005 0.0011638 0.23303 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.365 0.4691 0.14286 0.017421 10.9187 0.10844 0.00013855 0.7817 0.0083716 0.0092999 0.0013842 0.98697 0.99172 2.9846e-006 1.1938e-005 0.15686 0.95309 0.92198 0.001396 0.99529 0.54786 0.0018808 0.42983 2.0797 2.0792 16.0011 144.9584 0.00015552 -85.6608 0.93394
6.038 0.9881 5.4844e-005 3.8183 0.011961 7.8818e-005 0.0011638 0.23303 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3651 0.46914 0.14287 0.017422 10.9209 0.10845 0.00013856 0.78169 0.0083721 0.0093005 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.15686 0.95319 0.92201 0.001396 0.9953 0.54802 0.0018808 0.42984 2.08 2.0796 16.001 144.9584 0.00015546 -85.6608 0.93494
6.039 0.9881 5.4843e-005 3.8183 0.011961 7.8831e-005 0.0011638 0.23303 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3652 0.46919 0.14289 0.017423 10.9232 0.10846 0.00013857 0.78168 0.0083726 0.0093011 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.15686 0.95328 0.92205 0.001396 0.99531 0.54818 0.0018808 0.42985 2.0804 2.0799 16.001 144.9584 0.0001554 -85.6608 0.93594
6.04 0.9881 5.4843e-005 3.8183 0.011961 7.8844e-005 0.0011638 0.23303 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3653 0.46924 0.1429 0.017425 10.9255 0.10847 0.00013859 0.78167 0.0083732 0.0093017 0.0013842 0.98697 0.99172 2.9842e-006 1.1937e-005 0.15687 0.95338 0.92209 0.001396 0.99533 0.54833 0.0018808 0.42987 2.0807 2.0802 16.001 144.9585 0.00015535 -85.6609 0.93694
6.041 0.9881 5.4843e-005 3.8183 0.011961 7.8857e-005 0.0011638 0.23303 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3654 0.46928 0.14292 0.017426 10.9278 0.10848 0.0001386 0.78166 0.0083737 0.0093022 0.0013842 0.98697 0.99172 2.9842e-006 1.1937e-005 0.15687 0.95347 0.92212 0.001396 0.99534 0.54849 0.0018808 0.42988 2.081 2.0806 16.0009 144.9585 0.00015529 -85.6609 0.93794
6.042 0.9881 5.4843e-005 3.8183 0.011961 7.887e-005 0.0011638 0.23303 0.0006593 0.23368 0.21562 0 0.032293 0.0389 0 1.3655 0.46933 0.14293 0.017427 10.93 0.10848 0.00013861 0.78166 0.0083743 0.0093028 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15688 0.95356 0.92216 0.001396 0.99535 0.54865 0.0018808 0.42989 2.0814 2.0809 16.0009 144.9585 0.00015523 -85.6609 0.93894
6.043 0.9881 5.4843e-005 3.8183 0.011961 7.8883e-005 0.0011638 0.23303 0.0006593 0.23369 0.21562 0 0.032292 0.0389 0 1.3656 0.46938 0.14295 0.017429 10.9323 0.10849 0.00013862 0.78165 0.0083748 0.0093034 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.15688 0.95366 0.92219 0.001396 0.99536 0.54881 0.0018808 0.4299 2.0817 2.0812 16.0009 144.9585 0.00015518 -85.661 0.93994
6.044 0.9881 5.4843e-005 3.8183 0.011961 7.8895e-005 0.0011638 0.23303 0.0006593 0.23369 0.21562 0 0.032292 0.0389 0 1.3657 0.46942 0.14296 0.01743 10.9346 0.1085 0.00013863 0.78164 0.0083753 0.009304 0.0013842 0.98697 0.99172 2.9845e-006 1.1937e-005 0.15688 0.95375 0.92223 0.001396 0.99537 0.54896 0.0018808 0.42992 2.082 2.0816 16.0008 144.9585 0.00015512 -85.661 0.94094
6.045 0.9881 5.4843e-005 3.8183 0.011961 7.8908e-005 0.0011639 0.23303 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.3657 0.46947 0.14298 0.017432 10.9368 0.10851 0.00013865 0.78163 0.0083759 0.0093045 0.0013842 0.98697 0.99172 2.9847e-006 1.1938e-005 0.15689 0.95384 0.92227 0.001396 0.99538 0.54912 0.0018808 0.42993 2.0824 2.0819 16.0008 144.9586 0.00015507 -85.661 0.94194
6.046 0.9881 5.4843e-005 3.8183 0.011961 7.8921e-005 0.0011639 0.23303 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.3658 0.46951 0.14299 0.017433 10.9391 0.10852 0.00013866 0.78162 0.0083764 0.0093051 0.0013842 0.98697 0.99172 2.9848e-006 1.1938e-005 0.15689 0.95394 0.9223 0.001396 0.9954 0.54928 0.0018808 0.42994 2.0827 2.0822 16.0008 144.9586 0.00015501 -85.6611 0.94294
6.047 0.9881 5.4843e-005 3.8183 0.011961 7.8934e-005 0.0011639 0.23304 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.3659 0.46956 0.14301 0.017434 10.9414 0.10853 0.00013867 0.78161 0.0083769 0.0093057 0.0013842 0.98697 0.99172 2.9848e-006 1.1938e-005 0.1569 0.95403 0.92234 0.001396 0.99541 0.54943 0.0018808 0.42995 2.083 2.0826 16.0007 144.9586 0.00015496 -85.6611 0.94394
6.048 0.9881 5.4843e-005 3.8183 0.011961 7.8947e-005 0.0011639 0.23304 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.366 0.46961 0.14302 0.017436 10.9437 0.10853 0.00013868 0.78161 0.0083775 0.0093063 0.0013842 0.98697 0.99172 2.9847e-006 1.1937e-005 0.1569 0.95412 0.92237 0.001396 0.99542 0.54959 0.0018807 0.42996 2.0834 2.0829 16.0007 144.9586 0.0001549 -85.6611 0.94494
6.049 0.9881 5.4843e-005 3.8183 0.011961 7.896e-005 0.0011639 0.23304 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.3661 0.46965 0.14304 0.017437 10.9459 0.10854 0.00013869 0.7816 0.008378 0.0093068 0.0013842 0.98697 0.99172 2.9846e-006 1.1937e-005 0.15691 0.95421 0.92241 0.001396 0.99543 0.54975 0.0018807 0.42998 2.0837 2.0832 16.0007 144.9586 0.00015485 -85.6611 0.94594
6.05 0.9881 5.4843e-005 3.8183 0.011961 7.8973e-005 0.0011639 0.23304 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.3662 0.4697 0.14305 0.017438 10.9482 0.10855 0.00013871 0.78159 0.0083785 0.0093074 0.0013841 0.98697 0.99172 2.9845e-006 1.1937e-005 0.15691 0.9543 0.92244 0.001396 0.99544 0.54991 0.0018807 0.42999 2.084 2.0836 16.0006 144.9587 0.00015479 -85.6612 0.94694
6.051 0.9881 5.4843e-005 3.8183 0.011961 7.8986e-005 0.0011639 0.23304 0.0006593 0.23369 0.21563 0 0.032292 0.0389 0 1.3663 0.46974 0.14307 0.01744 10.9505 0.10856 0.00013872 0.78158 0.0083791 0.009308 0.0013841 0.98697 0.99172 2.9845e-006 1.1937e-005 0.15691 0.9544 0.92248 0.0013959 0.99545 0.55006 0.0018807 0.43 2.0844 2.0839 16.0006 144.9587 0.00015474 -85.6612 0.94794
6.052 0.9881 5.4842e-005 3.8183 0.011961 7.8999e-005 0.0011639 0.23304 0.0006593 0.2337 0.21563 0 0.032292 0.0389 0 1.3664 0.46979 0.14308 0.017441 10.9528 0.10857 0.00013873 0.78157 0.0083796 0.0093086 0.0013841 0.98697 0.99172 2.9845e-006 1.1937e-005 0.15692 0.95449 0.92251 0.0013959 0.99546 0.55022 0.0018807 0.43001 2.0847 2.0842 16.0006 144.9587 0.00015468 -85.6612 0.94894
6.053 0.9881 5.4842e-005 3.8183 0.011961 7.9012e-005 0.0011639 0.23304 0.0006593 0.2337 0.21563 0 0.032292 0.0389 0 1.3665 0.46984 0.1431 0.017442 10.955 0.10857 0.00013874 0.78156 0.0083801 0.0093091 0.0013841 0.98697 0.99172 2.9844e-006 1.1937e-005 0.15692 0.95458 0.92254 0.0013959 0.99548 0.55038 0.0018807 0.43003 2.085 2.0846 16.0005 144.9587 0.00015463 -85.6613 0.94994
6.054 0.9881 5.4842e-005 3.8183 0.011961 7.9025e-005 0.0011639 0.23304 0.0006593 0.2337 0.21563 0 0.032292 0.0389 0 1.3666 0.46988 0.14311 0.017444 10.9573 0.10858 0.00013875 0.78156 0.0083807 0.0093097 0.0013841 0.98697 0.99172 2.9845e-006 1.1937e-005 0.15693 0.95467 0.92258 0.0013959 0.99549 0.55053 0.0018807 0.43004 2.0854 2.0849 16.0005 144.9587 0.00015457 -85.6613 0.95094
6.055 0.9881 5.4842e-005 3.8183 0.011961 7.9038e-005 0.0011639 0.23304 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.3667 0.46993 0.14313 0.017445 10.9596 0.10859 0.00013877 0.78155 0.0083812 0.0093103 0.0013841 0.98697 0.99172 2.9845e-006 1.1937e-005 0.15693 0.95476 0.92261 0.0013959 0.9955 0.55069 0.0018807 0.43005 2.0857 2.0852 16.0005 144.9588 0.00015452 -85.6613 0.95194
6.056 0.9881 5.4842e-005 3.8183 0.011961 7.905e-005 0.0011639 0.23304 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.3668 0.46998 0.14314 0.017447 10.9619 0.1086 0.00013878 0.78154 0.0083817 0.0093109 0.0013841 0.98697 0.99172 2.9844e-006 1.1937e-005 0.15693 0.95485 0.92265 0.0013959 0.99551 0.55085 0.0018807 0.43006 2.086 2.0856 16.0004 144.9588 0.00015447 -85.6614 0.95294
6.057 0.9881 5.4842e-005 3.8183 0.011961 7.9063e-005 0.0011639 0.23305 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.3669 0.47002 0.14316 0.017448 10.9641 0.10861 0.00013879 0.78153 0.0083823 0.0093114 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.15694 0.95494 0.92268 0.0013959 0.99552 0.551 0.0018807 0.43007 2.0863 2.0859 16.0004 144.9588 0.00015441 -85.6614 0.95394
6.058 0.9881 5.4842e-005 3.8183 0.011961 7.9076e-005 0.0011639 0.23305 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.367 0.47007 0.14317 0.017449 10.9664 0.10862 0.0001388 0.78152 0.0083828 0.009312 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.15694 0.95503 0.92272 0.0013959 0.99553 0.55116 0.0018807 0.43009 2.0867 2.0862 16.0004 144.9588 0.00015436 -85.6614 0.95494
6.059 0.9881 5.4842e-005 3.8183 0.011961 7.9089e-005 0.0011639 0.23305 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.367 0.47011 0.14319 0.017451 10.9687 0.10862 0.00013882 0.78151 0.0083833 0.0093126 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15695 0.95512 0.92275 0.0013959 0.99554 0.55131 0.0018807 0.4301 2.087 2.0865 16.0003 144.9588 0.00015431 -85.6614 0.95594
6.06 0.9881 5.4842e-005 3.8183 0.011961 7.9102e-005 0.0011639 0.23305 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.3671 0.47016 0.1432 0.017452 10.971 0.10863 0.00013883 0.78151 0.0083839 0.0093132 0.0013841 0.98697 0.99172 2.984e-006 1.1936e-005 0.15695 0.95521 0.92278 0.0013959 0.99555 0.55147 0.0018807 0.43011 2.0873 2.0869 16.0003 144.9589 0.00015425 -85.6615 0.95694
6.061 0.9881 5.4842e-005 3.8183 0.011961 7.9115e-005 0.0011639 0.23305 0.0006593 0.2337 0.21564 0 0.032292 0.0389 0 1.3672 0.47021 0.14322 0.017453 10.9733 0.10864 0.00013884 0.7815 0.0083844 0.0093137 0.0013841 0.98697 0.99172 2.9839e-006 1.1936e-005 0.15696 0.95529 0.92282 0.0013959 0.99556 0.55163 0.0018807 0.43012 2.0877 2.0872 16.0003 144.9589 0.0001542 -85.6615 0.95794
6.062 0.9881 5.4842e-005 3.8183 0.011961 7.9128e-005 0.0011639 0.23305 0.0006593 0.23371 0.21564 0 0.032291 0.0389 0 1.3673 0.47025 0.14323 0.017455 10.9755 0.10865 0.00013885 0.78149 0.0083849 0.0093143 0.0013841 0.98697 0.99172 2.984e-006 1.1936e-005 0.15696 0.95538 0.92285 0.0013959 0.99557 0.55178 0.0018807 0.43013 2.088 2.0875 16.0002 144.9589 0.00015415 -85.6615 0.95894
6.063 0.9881 5.4842e-005 3.8183 0.011961 7.9141e-005 0.0011639 0.23305 0.0006593 0.23371 0.21564 0 0.032291 0.0389 0 1.3674 0.4703 0.14325 0.017456 10.9778 0.10866 0.00013886 0.78148 0.0083855 0.0093149 0.0013841 0.98697 0.99172 2.9841e-006 1.1936e-005 0.15696 0.95547 0.92288 0.0013959 0.99558 0.55194 0.0018807 0.43015 2.0883 2.0879 16.0002 144.9589 0.0001541 -85.6616 0.95994
6.064 0.9881 5.4842e-005 3.8183 0.011961 7.9154e-005 0.0011639 0.23305 0.0006593 0.23371 0.21564 0 0.032291 0.0389 0 1.3675 0.47034 0.14326 0.017457 10.9801 0.10867 0.00013888 0.78147 0.008386 0.0093155 0.001384 0.98697 0.99172 2.9842e-006 1.1936e-005 0.15697 0.95556 0.92292 0.0013959 0.99559 0.5521 0.0018807 0.43016 2.0886 2.0882 16.0002 144.9589 0.00015404 -85.6616 0.96094
6.065 0.9881 5.4841e-005 3.8183 0.011961 7.9167e-005 0.0011639 0.23305 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.3676 0.47039 0.14328 0.017459 10.9824 0.10867 0.00013889 0.78146 0.0083865 0.009316 0.001384 0.98697 0.99172 2.9844e-006 1.1936e-005 0.15697 0.95565 0.92295 0.0013959 0.9956 0.55225 0.0018807 0.43017 2.089 2.0885 16.0001 144.959 0.00015399 -85.6616 0.96194
6.066 0.9881 5.4841e-005 3.8183 0.011961 7.918e-005 0.0011639 0.23305 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.3677 0.47044 0.14329 0.01746 10.9847 0.10868 0.0001389 0.78146 0.0083871 0.0093166 0.001384 0.98697 0.99172 2.9843e-006 1.1936e-005 0.15698 0.95573 0.92298 0.0013959 0.99561 0.55241 0.0018807 0.43018 2.0893 2.0888 16.0001 144.959 0.00015394 -85.6616 0.96294
6.067 0.9881 5.4841e-005 3.8183 0.011961 7.9193e-005 0.0011639 0.23306 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.3678 0.47048 0.14331 0.017462 10.9869 0.10869 0.00013891 0.78145 0.0083876 0.0093172 0.001384 0.98697 0.99172 2.9842e-006 1.1936e-005 0.15698 0.95582 0.92302 0.0013959 0.99562 0.55256 0.0018807 0.43019 2.0896 2.0891 16.0001 144.959 0.00015389 -85.6617 0.96394
6.068 0.9881 5.4841e-005 3.8183 0.011961 7.9205e-005 0.0011639 0.23306 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.3679 0.47053 0.14332 0.017463 10.9892 0.1087 0.00013892 0.78144 0.0083881 0.0093177 0.001384 0.98697 0.99172 2.984e-006 1.1936e-005 0.15698 0.95591 0.92305 0.0013959 0.99563 0.55272 0.0018807 0.43021 2.0899 2.0895 16 144.959 0.00015384 -85.6617 0.96494
6.069 0.9881 5.4841e-005 3.8183 0.011961 7.9218e-005 0.0011639 0.23306 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.368 0.47058 0.14334 0.017464 10.9915 0.10871 0.00013894 0.78143 0.0083887 0.0093183 0.001384 0.98697 0.99172 2.9838e-006 1.1936e-005 0.15699 0.95599 0.92308 0.0013959 0.99564 0.55287 0.0018807 0.43022 2.0902 2.0898 16 144.9591 0.00015379 -85.6617 0.96594
6.07 0.9881 5.4841e-005 3.8183 0.011961 7.9231e-005 0.0011639 0.23306 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.3681 0.47062 0.14335 0.017466 10.9938 0.10872 0.00013895 0.78142 0.0083892 0.0093189 0.001384 0.98697 0.99172 2.9835e-006 1.1935e-005 0.15699 0.95608 0.92312 0.0013959 0.99565 0.55303 0.0018806 0.43023 2.0906 2.0901 16 144.9591 0.00015374 -85.6617 0.96694
6.071 0.9881 5.4841e-005 3.8183 0.011961 7.9244e-005 0.0011639 0.23306 0.0006593 0.23371 0.21565 0 0.032291 0.0389 0 1.3682 0.47067 0.14337 0.017467 10.9961 0.10872 0.00013896 0.78141 0.0083897 0.0093195 0.001384 0.98697 0.99172 2.9834e-006 1.1935e-005 0.157 0.95616 0.92315 0.0013959 0.99566 0.55319 0.0018806 0.43024 2.0909 2.0904 15.9999 144.9591 0.00015368 -85.6618 0.96794
6.072 0.9881 5.4841e-005 3.8183 0.011961 7.9257e-005 0.0011639 0.23306 0.0006593 0.23372 0.21565 0 0.032291 0.0389 0 1.3683 0.47071 0.14338 0.017468 10.9983 0.10873 0.00013897 0.78141 0.0083903 0.00932 0.001384 0.98697 0.99172 2.9834e-006 1.1935e-005 0.157 0.95625 0.92318 0.0013959 0.99567 0.55334 0.0018806 0.43025 2.0912 2.0908 15.9999 144.9591 0.00015363 -85.6618 0.96894
6.073 0.9881 5.4841e-005 3.8183 0.011961 7.927e-005 0.001164 0.23306 0.0006593 0.23372 0.21565 0 0.032291 0.0389 0 1.3683 0.47076 0.1434 0.01747 11.0006 0.10874 0.00013898 0.7814 0.0083908 0.0093206 0.001384 0.98697 0.99172 2.9834e-006 1.1935e-005 0.15701 0.95634 0.92321 0.0013959 0.99568 0.5535 0.0018806 0.43027 2.0915 2.0911 15.9999 144.9591 0.00015358 -85.6618 0.96994
6.074 0.9881 5.4841e-005 3.8183 0.011961 7.9283e-005 0.001164 0.23306 0.0006593 0.23372 0.21565 0 0.032291 0.0389 0 1.3684 0.47081 0.14341 0.017471 11.0029 0.10875 0.000139 0.78139 0.0083913 0.0093212 0.001384 0.98697 0.99172 2.9835e-006 1.1935e-005 0.15701 0.95642 0.92325 0.0013959 0.99569 0.55365 0.0018806 0.43028 2.0918 2.0914 15.9998 144.9592 0.00015353 -85.6618 0.97094
6.075 0.9881 5.4841e-005 3.8183 0.011961 7.9296e-005 0.001164 0.23306 0.0006593 0.23372 0.21565 0 0.032291 0.0389 0 1.3685 0.47085 0.14343 0.017472 11.0052 0.10876 0.00013901 0.78138 0.0083919 0.0093218 0.001384 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15701 0.9565 0.92328 0.0013959 0.9957 0.55381 0.0018806 0.43029 2.0922 2.0917 15.9998 144.9592 0.00015348 -85.6619 0.97194
6.076 0.9881 5.4841e-005 3.8183 0.011961 7.9309e-005 0.001164 0.23306 0.0006593 0.23372 0.21566 0 0.032291 0.0389 0 1.3686 0.4709 0.14344 0.017474 11.0075 0.10877 0.00013902 0.78137 0.0083924 0.0093223 0.001384 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15702 0.95659 0.92331 0.0013959 0.99571 0.55396 0.0018806 0.4303 2.0925 2.092 15.9998 144.9592 0.00015343 -85.6619 0.97294
6.077 0.9881 5.4841e-005 3.8183 0.011961 7.9322e-005 0.001164 0.23307 0.0006593 0.23372 0.21566 0 0.032291 0.0389 0 1.3687 0.47095 0.14346 0.017475 11.0098 0.10877 0.00013903 0.78136 0.0083929 0.0093229 0.001384 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15702 0.95667 0.92334 0.0013959 0.99572 0.55412 0.0018806 0.43031 2.0928 2.0924 15.9997 144.9592 0.00015338 -85.6619 0.97394
6.078 0.9881 5.484e-005 3.8183 0.011961 7.9335e-005 0.001164 0.23307 0.0006593 0.23372 0.21566 0 0.032291 0.0389 0 1.3688 0.47099 0.14347 0.017477 11.012 0.10878 0.00013904 0.78136 0.0083935 0.0093235 0.001384 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15703 0.95676 0.92337 0.0013959 0.99573 0.55427 0.0018806 0.43033 2.0931 2.0927 15.9997 144.9592 0.00015333 -85.6619 0.97494
6.079 0.9881 5.484e-005 3.8183 0.011961 7.9348e-005 0.001164 0.23307 0.0006593 0.23372 0.21566 0 0.032291 0.0389 0 1.3689 0.47104 0.14349 0.017478 11.0143 0.10879 0.00013906 0.78135 0.008394 0.009324 0.0013839 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15703 0.95684 0.9234 0.0013959 0.99574 0.55443 0.0018806 0.43034 2.0934 2.093 15.9997 144.9593 0.00015328 -85.662 0.97594
6.08 0.9881 5.484e-005 3.8183 0.011961 7.936e-005 0.001164 0.23307 0.0006593 0.23372 0.21566 0 0.032291 0.0389 0 1.369 0.47108 0.1435 0.017479 11.0166 0.1088 0.00013907 0.78134 0.0083945 0.0093246 0.0013839 0.98697 0.99172 2.9835e-006 1.1935e-005 0.15704 0.95692 0.92344 0.0013959 0.99575 0.55458 0.0018806 0.43035 2.0937 2.0933 15.9996 144.9593 0.00015323 -85.662 0.97694
6.081 0.9881 5.484e-005 3.8183 0.011961 7.9373e-005 0.001164 0.23307 0.0006593 0.23372 0.21566 0 0.032291 0.0389 0 1.3691 0.47113 0.14352 0.017481 11.0189 0.10881 0.00013908 0.78133 0.0083951 0.0093252 0.0013839 0.98697 0.99172 2.9835e-006 1.1935e-005 0.15704 0.95701 0.92347 0.0013959 0.99576 0.55474 0.0018806 0.43036 2.0941 2.0936 15.9996 144.9593 0.00015318 -85.662 0.97794
6.082 0.9881 5.484e-005 3.8183 0.011961 7.9386e-005 0.001164 0.23307 0.0006593 0.23373 0.21566 0 0.03229 0.0389 0 1.3692 0.47118 0.14353 0.017482 11.0212 0.10882 0.00013909 0.78132 0.0083956 0.0093258 0.0013839 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15704 0.95709 0.9235 0.0013958 0.99577 0.5549 0.0018806 0.43037 2.0944 2.0939 15.9996 144.9593 0.00015313 -85.662 0.97894
6.083 0.9881 5.484e-005 3.8183 0.011961 7.9399e-005 0.001164 0.23307 0.0006593 0.23373 0.21566 0 0.03229 0.0389 0 1.3693 0.47122 0.14355 0.017483 11.0235 0.10882 0.0001391 0.78132 0.0083961 0.0093263 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15705 0.95717 0.92353 0.0013958 0.99578 0.55505 0.0018806 0.43039 2.0947 2.0943 15.9995 144.9593 0.00015309 -85.662 0.97994
6.084 0.9881 5.484e-005 3.8183 0.011961 7.9412e-005 0.001164 0.23307 0.0006593 0.23373 0.21566 0 0.03229 0.0389 0 1.3694 0.47127 0.14356 0.017485 11.0257 0.10883 0.00013912 0.78131 0.0083967 0.0093269 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.15705 0.95726 0.92356 0.0013958 0.99579 0.55521 0.0018806 0.4304 2.095 2.0946 15.9995 144.9594 0.00015304 -85.6621 0.98094
6.085 0.9881 5.484e-005 3.8183 0.011961 7.9425e-005 0.001164 0.23307 0.00065931 0.23373 0.21566 0 0.03229 0.0389 0 1.3695 0.47131 0.14358 0.017486 11.028 0.10884 0.00013913 0.7813 0.0083972 0.0093275 0.0013839 0.98697 0.99172 2.984e-006 1.1935e-005 0.15706 0.95734 0.92359 0.0013958 0.9958 0.55536 0.0018806 0.43041 2.0953 2.0949 15.9995 144.9594 0.00015299 -85.6621 0.98194
6.086 0.9881 5.484e-005 3.8183 0.011961 7.9438e-005 0.001164 0.23307 0.00065931 0.23373 0.21567 0 0.03229 0.0389 0 1.3696 0.47136 0.14359 0.017487 11.0303 0.10885 0.00013914 0.78129 0.0083977 0.0093281 0.0013839 0.98697 0.99172 2.984e-006 1.1935e-005 0.15706 0.95742 0.92362 0.0013958 0.9958 0.55551 0.0018806 0.43042 2.0956 2.0952 15.9994 144.9594 0.00015294 -85.6621 0.98294
6.087 0.9881 5.484e-005 3.8183 0.011961 7.9451e-005 0.001164 0.23308 0.00065931 0.23373 0.21567 0 0.03229 0.0389 0 1.3696 0.47141 0.14361 0.017489 11.0326 0.10886 0.00013915 0.78128 0.0083983 0.0093286 0.0013839 0.98697 0.99172 2.9839e-006 1.1935e-005 0.15706 0.9575 0.92366 0.0013958 0.99581 0.55567 0.0018806 0.43043 2.096 2.0955 15.9994 144.9594 0.00015289 -85.6621 0.98394
6.088 0.9881 5.484e-005 3.8183 0.011961 7.9464e-005 0.001164 0.23308 0.00065931 0.23373 0.21567 0 0.03229 0.0389 0 1.3697 0.47145 0.14362 0.01749 11.0349 0.10887 0.00013917 0.78127 0.0083988 0.0093292 0.0013839 0.98697 0.99172 2.9838e-006 1.1935e-005 0.15707 0.95758 0.92369 0.0013958 0.99582 0.55582 0.0018806 0.43045 2.0963 2.0958 15.9994 144.9594 0.00015284 -85.6622 0.98494
6.089 0.9881 5.484e-005 3.8183 0.011961 7.9477e-005 0.001164 0.23308 0.00065931 0.23373 0.21567 0 0.03229 0.0389 0 1.3698 0.4715 0.14363 0.017491 11.0372 0.10887 0.00013918 0.78127 0.0083993 0.0093298 0.0013839 0.98697 0.99172 2.9836e-006 1.1935e-005 0.15707 0.95766 0.92372 0.0013958 0.99583 0.55598 0.0018806 0.43046 2.0966 2.0961 15.9993 144.9595 0.0001528 -85.6622 0.98594
6.09 0.9881 5.484e-005 3.8183 0.01196 7.949e-005 0.001164 0.23308 0.00065931 0.23373 0.21567 0 0.03229 0.0389 0 1.3699 0.47155 0.14365 0.017493 11.0395 0.10888 0.00013919 0.78126 0.0083998 0.0093303 0.0013839 0.98697 0.99172 2.9833e-006 1.1935e-005 0.15708 0.95774 0.92375 0.0013958 0.99584 0.55613 0.0018806 0.43047 2.0969 2.0965 15.9993 144.9595 0.00015275 -85.6622 0.98694
6.091 0.9881 5.4839e-005 3.8183 0.01196 7.9502e-005 0.001164 0.23308 0.00065931 0.23373 0.21567 0 0.03229 0.0389 0 1.37 0.47159 0.14366 0.017494 11.0418 0.10889 0.0001392 0.78125 0.0084004 0.0093309 0.0013839 0.98697 0.99172 2.9832e-006 1.1934e-005 0.15708 0.95783 0.92378 0.0013958 0.99585 0.55629 0.0018806 0.43048 2.0972 2.0968 15.9993 144.9595 0.0001527 -85.6622 0.98794
6.092 0.9881 5.4839e-005 3.8183 0.01196 7.9515e-005 0.001164 0.23308 0.00065931 0.23374 0.21567 0 0.03229 0.0389 0 1.3701 0.47164 0.14368 0.017496 11.0441 0.1089 0.00013921 0.78124 0.0084009 0.0093315 0.0013839 0.98697 0.99172 2.9832e-006 1.1934e-005 0.15708 0.95791 0.92381 0.0013958 0.99586 0.55644 0.0018806 0.43049 2.0975 2.0971 15.9992 144.9595 0.00015265 -85.6622 0.98894
6.093 0.9881 5.4839e-005 3.8183 0.01196 7.9528e-005 0.001164 0.23308 0.00065931 0.23374 0.21567 0 0.03229 0.0389 0 1.3702 0.47168 0.14369 0.017497 11.0463 0.10891 0.00013923 0.78123 0.0084014 0.0093321 0.0013839 0.98697 0.99172 2.9833e-006 1.1934e-005 0.15709 0.95799 0.92384 0.0013958 0.99587 0.5566 0.0018806 0.43051 2.0978 2.0974 15.9992 144.9595 0.0001526 -85.6623 0.98994
6.094 0.9881 5.4839e-005 3.8183 0.01196 7.9541e-005 0.001164 0.23308 0.00065931 0.23374 0.21567 0 0.03229 0.0389 0 1.3703 0.47173 0.14371 0.017498 11.0486 0.10891 0.00013924 0.78122 0.008402 0.0093326 0.0013839 0.98697 0.99172 2.9833e-006 1.1934e-005 0.15709 0.95807 0.92387 0.0013958 0.99587 0.55675 0.0018806 0.43052 2.0981 2.0977 15.9992 144.9596 0.00015256 -85.6623 0.99094
6.095 0.9881 5.4839e-005 3.8183 0.01196 7.9554e-005 0.001164 0.23308 0.00065931 0.23374 0.21567 0 0.03229 0.0389 0 1.3704 0.47178 0.14372 0.0175 11.0509 0.10892 0.00013925 0.78122 0.0084025 0.0093332 0.0013839 0.98697 0.99172 2.9834e-006 1.1934e-005 0.1571 0.95815 0.9239 0.0013958 0.99588 0.55691 0.0018806 0.43053 2.0984 2.098 15.9991 144.9596 0.00015251 -85.6623 0.99194
6.096 0.9881 5.4839e-005 3.8183 0.01196 7.9567e-005 0.001164 0.23308 0.00065931 0.23374 0.21567 0 0.03229 0.0389 0 1.3705 0.47182 0.14374 0.017501 11.0532 0.10893 0.00013926 0.78121 0.008403 0.0093338 0.0013839 0.98697 0.99172 2.9835e-006 1.1934e-005 0.1571 0.95822 0.92393 0.0013958 0.99589 0.55706 0.0018806 0.43054 2.0987 2.0983 15.9991 144.9596 0.00015246 -85.6623 0.99294
6.097 0.9881 5.4839e-005 3.8183 0.01196 7.958e-005 0.001164 0.23309 0.00065931 0.23374 0.21568 0 0.03229 0.0389 0 1.3706 0.47187 0.14375 0.017502 11.0555 0.10894 0.00013927 0.7812 0.0084036 0.0093343 0.0013839 0.98697 0.99172 2.9837e-006 1.1935e-005 0.15711 0.9583 0.92396 0.0013958 0.9959 0.55721 0.0018806 0.43055 2.0991 2.0986 15.9991 144.9596 0.00015242 -85.6623 0.99394
6.098 0.9881 5.4839e-005 3.8183 0.01196 7.9593e-005 0.001164 0.23309 0.00065931 0.23374 0.21568 0 0.03229 0.0389 0 1.3707 0.47191 0.14377 0.017504 11.0578 0.10895 0.00013929 0.78119 0.0084041 0.0093349 0.0013839 0.98697 0.99172 2.9837e-006 1.1934e-005 0.15711 0.95838 0.92399 0.0013958 0.99591 0.55737 0.0018805 0.43057 2.0994 2.0989 15.999 144.9596 0.00015237 -85.6624 0.99494
6.099 0.9881 5.4839e-005 3.8183 0.01196 7.9606e-005 0.001164 0.23309 0.00065931 0.23374 0.21568 0 0.03229 0.0389 0 1.3708 0.47196 0.14378 0.017505 11.0601 0.10896 0.0001393 0.78118 0.0084046 0.0093355 0.0013839 0.98697 0.99172 2.9836e-006 1.1934e-005 0.15711 0.95846 0.92402 0.0013958 0.99592 0.55752 0.0018805 0.43058 2.0997 2.0992 15.999 144.9597 0.00015232 -85.6624 0.99594
6.1 0.9881 5.4839e-005 3.8183 0.01196 7.9619e-005 0.0011641 0.23309 0.00065931 0.23374 0.21568 0 0.03229 0.0389 0 1.3709 0.47201 0.1438 0.017506 11.0624 0.10896 0.00013931 0.78117 0.0084052 0.0093361 0.001384 0.98697 0.99172 2.9837e-006 1.1934e-005 0.15712 0.95854 0.92405 0.0013958 0.99592 0.55768 0.0018805 0.43059 2.1 2.0996 15.999 144.9597 0.00015228 -85.6575 0.99694
6.101 0.9881 5.4839e-005 3.8183 0.01196 7.9632e-005 0.0011641 0.23309 0.00065931 0.23374 0.21568 0 0.03229 0.0389 0 1.3709 0.47205 0.14381 0.017508 11.0647 0.10897 0.00013932 0.78117 0.0084057 0.0093366 0.0064793 0.98322 0.99099 1.4532e-005 5.3384e-005 0.15712 0.95857 0.92408 0.0027744 0.99592 0.55781 0.002396 0.43055 2.1003 2.0999 15.9989 144.9597 0.00015224 -76.1548 0.99794
6.102 0.9881 5.4839e-005 3.8183 0.01196 7.9645e-005 0.0011641 0.23309 0.00065931 0.23375 0.21568 0 0.03229 0.0389 0 1.371 0.4721 0.14383 0.017509 11.067 0.10898 0.00013933 0.78116 0.0084062 0.0093372 0.026243 0.9717 0.98766 6.6038e-005 0.0002297 0.15713 0.95837 0.92411 0.0053028 0.99587 0.55793 0.0033369 0.43043 2.1006 2.1002 15.9988 144.9597 0.00015223 -67.141 0.99894
6.103 0.9881 5.4839e-005 3.8183 0.01196 7.9657e-005 0.0011641 0.23309 0.00065931 0.23375 0.21568 0 0.032289 0.0389 0 1.3711 0.47215 0.14384 0.01751 11.0693 0.10899 0.00013935 0.78115 0.0084067 0.0093378 0.094951 0.9472 0.97731 0.00028467 0.00091393 0.15713 0.95763 0.92413 0.0092506 0.9956 0.55803 0.0044258 0.43026 2.1009 2.1005 15.9988 144.9596 0.00015223 -58.009 0.99994
6.104 0.9881 5.4838e-005 3.8183 0.01196 7.967e-005 0.0011641 0.23309 0.00065931 0.23375 0.21568 0 0.032289 0.0389 0 1.3712 0.47219 0.14386 0.017512 11.0715 0.109 0.00013936 0.78114 0.0084073 0.0093383 0.48898 0.8559 0.93866 0.0021859 0.0054898 0.15713 0.95563 0.92416 0.01576 0.99148 0.55806 0.005625 0.43007 2.1012 2.1008 15.9995 144.9596 0.00015227 -37.1648 0.15505
6.105 0.9881 5.4838e-005 3.8183 0.01196 7.9683e-005 0.0011641 0.23309 0.00065931 0.23375 0.21568 0 0.032289 0.0389 0 1.3713 0.47224 0.14387 0.017513 11.0738 0.10901 0.00013937 0.78113 0.0084078 0.0093389 0.99962 0.0021566 0.71197 0.94202 0.99646 0.15714 0.92226 0.92112 0.33515 0.96406 0.5458 0.044434 0.42987 2.0494 0.95759 16.0034 144.9593 0.00024402 24.9076 0.0019467
6.106 0.9881 5.4838e-005 3.8183 0.01196 7.9696e-005 0.0011641 0.23309 0.00065931 0.23375 0.21568 0 0.032289 0.0389 0 1.3714 0.47228 0.14389 0.017515 11.0761 0.10901 0.00013938 0.78113 0.0084083 0.0093395 0.99949 1.3175e-006 0.52806 0.99801 0.99955 0.15714 0.88231 0.90289 0.62235 0.93691 0.53053 0.099568 0.42967 1.8474 0.60432 16.003 144.9579 0.00035822 21.3772 0.0029467
6.107 0.9881 5.4838e-005 3.8183 0.01196 7.9709e-005 0.0011641 0.2331 0.00065931 0.23375 0.21568 0 0.032289 0.0389 0 1.3715 0.47233 0.1439 0.017516 11.0784 0.10902 0.00013939 0.78112 0.0084089 0.00934 0.99913 9.0761e-010 0.39193 0.99623 0.99894 0.15715 0.84455 0.87929 0.7478 0.91052 0.51584 0.14228 0.42946 1.6577 0.58566 16.0026 144.9562 0.00043194 16.3202 0.0039467
6.108 0.9881 5.4838e-005 3.8183 0.01196 7.9722e-005 0.0011641 0.2331 0.00065931 0.23375 0.21569 0 0.032289 0.0389 0 1.3716 0.47238 0.14392 0.017517 11.0807 0.10903 0.00013941 0.78111 0.0084094 0.0093406 0.99873 -9.3803e-011 0.29119 0.99301 0.99802 0.15715 0.80936 0.85289 0.80279 0.88488 0.50185 0.17587 0.42926 1.5002 0.62942 16.0023 144.9543 0.00048778 12.827 0.0049467
6.109 0.9881 5.4838e-005 3.8183 0.01196 7.9735e-005 0.0011641 0.2331 0.00065931 0.23375 0.21569 0 0.032289 0.0389 0 1.3717 0.47242 0.14393 0.017519 11.083 0.10904 0.00013942 0.7811 0.0084099 0.0093412 0.99836 -2.7891e-011 0.21654 0.98927 0.99698 0.15716 0.77667 0.82494 0.82676 0.85996 0.48857 0.20398 0.42905 1.3754 0.69297 16.002 144.9525 0.00053111 10.5181 0.0059467
6.11 0.9881 5.4838e-005 3.8183 0.01196 7.9748e-005 0.0011641 0.2331 0.00065931 0.23375 0.21569 0 0.032289 0.0389 0 1.3718 0.47247 0.14395 0.01752 11.0853 0.10905 0.00013943 0.78109 0.0084105 0.0093418 0.99802 -1.6775e-010 0.16115 0.98528 0.99588 0.15716 0.74621 0.79631 0.83543 0.83575 0.47597 0.22844 0.42885 1.2798 0.76076 16.0016 144.9507 0.00056456 8.8036 0.0069467
6.111 0.9881 5.4838e-005 3.8183 0.01196 7.9761e-005 0.0011641 0.2331 0.00065931 0.23375 0.21569 0 0.032289 0.0389 0 1.3719 0.47251 0.14396 0.017521 11.0876 0.10906 0.00013944 0.78108 0.008411 0.0093423 0.99769 1.4094e-011 0.12003 0.98101 0.99469 0.15716 0.71777 0.76763 0.83571 0.81222 0.464 0.25014 0.42864 1.209 0.8247 16.0013 144.949 0.00059022 7.3739 0.0079467
6.112 0.9881 5.4838e-005 3.8183 0.01196 7.9774e-005 0.0011641 0.2331 0.00065931 0.23375 0.21569 0 0.032289 0.0389 0 1.372 0.47256 0.14398 0.017523 11.0899 0.10906 0.00013945 0.78108 0.0084115 0.0093429 0.99734 -1.8915e-011 0.089464 0.97632 0.99336 0.15717 0.69118 0.73938 0.83101 0.78936 0.45266 0.26957 0.42844 1.1582 0.8804 16.001 144.9474 0.00060993 6.0833 0.0089467
6.113 0.9881 5.4838e-005 3.8183 0.01196 7.9787e-005 0.0011641 0.2331 0.00065931 0.23376 0.21569 0 0.032289 0.0389 0 1.3721 0.47261 0.14399 0.017524 11.0922 0.10907 0.00013947 0.78107 0.008412 0.0093435 0.99696 3.4949e-011 0.066737 0.97103 0.99183 0.15717 0.66632 0.71188 0.8231 0.76714 0.44192 0.28702 0.42824 1.1228 0.92609 16.0007 144.9458 0.00062526 4.8589 0.0099467
6.114 0.9881 5.4838e-005 3.8183 0.01196 7.98e-005 0.0011641 0.2331 0.00065931 0.23376 0.21569 0 0.032289 0.0389 0 1.3721 0.47265 0.14401 0.017525 11.0945 0.10908 0.00013948 0.78106 0.0084126 0.009344 0.99653 1.1393e-011 0.049826 0.96496 0.99003 0.15718 0.6431 0.68536 0.81293 0.74555 0.4318 0.30271 0.42803 1.0991 0.96189 16.0005 144.9444 0.00063743 3.6596 0.010947
6.115 0.9881 5.4838e-005 3.8183 0.01196 7.9812e-005 0.0011641 0.2331 0.00065931 0.23376 0.21569 0 0.032289 0.0389 0 1.3722 0.4727 0.14402 0.017527 11.0968 0.10909 0.00013949 0.78105 0.0084131 0.0093446 0.99605 6.5799e-011 0.037236 0.95788 0.98787 0.15718 0.62146 0.65999 0.80103 0.72458 0.4223 0.31678 0.42783 1.0837 0.989 16.0002 144.943 0.00064734 2.4587 0.011947
6.116 0.9881 5.4838e-005 3.8183 0.01196 7.9825e-005 0.0011641 0.2331 0.00065931 0.23376 0.21569 0 0.032289 0.0389 0 1.3723 0.47275 0.14404 0.017528 11.0991 0.1091 0.0001395 0.78104 0.0084136 0.0093452 0.99548 1.6872e-011 0.027857 0.94952 0.98525 0.15718 0.60133 0.6359 0.78765 0.7042 0.41342 0.32934 0.42762 1.0743 1.0091 15.9999 144.9417 0.00065563 1.2352 0.012947
6.117 0.9881 5.4837e-005 3.8183 0.01196 7.9838e-005 0.0011641 0.2331 0.00065931 0.23376 0.21569 0 0.032289 0.0389 0 1.3724 0.47279 0.14405 0.017529 11.1014 0.1091 0.00013951 0.78103 0.0084142 0.0093457 0.9948 8.8652e-011 0.020867 0.93954 0.98201 0.15719 0.58266 0.61317 0.7729 0.6844 0.40519 0.34049 0.42742 1.0689 1.0238 15.9996 144.9404 0.00066271 -0.030989 0.013947
6.118 0.9881 5.4837e-005 3.8183 0.01196 7.9851e-005 0.0011641 0.23311 0.00065931 0.23376 0.21569 0 0.032289 0.0389 0 1.3725 0.47284 0.14407 0.017531 11.1037 0.10911 0.00013953 0.78103 0.0084147 0.0093463 0.99398 1.0805e-010 0.015654 0.9275 0.978 0.15719 0.56543 0.59189 0.75676 0.66517 0.39761 0.35029 0.42722 1.0663 1.0347 15.9994 144.9393 0.00066887 -1.3621 0.014947
6.119 0.9881 5.4837e-005 3.8183 0.01196 7.9864e-005 0.0011641 0.23311 0.00065931 0.23376 0.2157 0 0.032289 0.0389 0 1.3726 0.47288 0.14408 0.017532 11.106 0.10912 0.00013954 0.78102 0.0084152 0.0093469 0.99295 7.4633e-012 0.011764 0.91282 0.97285 0.1572 0.54961 0.57214 0.73914 0.64648 0.39072 0.35878 0.42701 1.0655 1.0428 15.9991 144.9382 0.00067426 -2.7861 0.015947
6.12 0.9881 5.4837e-005 3.8183 0.01196 7.9877e-005 0.0011641 0.23311 0.00065931 0.23376 0.2157 0 0.032289 0.0389 0 1.3727 0.47293 0.1441 0.017534 11.1083 0.10913 0.00013955 0.78101 0.0084157 0.0093474 0.99163 2.0427e-011 0.00886 0.89468 0.96625 0.1572 0.5352 0.55403 0.71985 0.62834 0.38455 0.36601 0.42681 1.0659 1.049 15.9989 144.9372 0.00067897 -4.34 0.016947
6.121 0.9881 5.4837e-005 3.8183 0.01196 7.989e-005 0.0011641 0.23311 0.00065931 0.23376 0.2157 0 0.032289 0.0389 0 1.3728 0.47298 0.14411 0.017535 11.1106 0.10914 0.00013956 0.781 0.0084163 0.009348 0.98986 -1.1237e-011 0.0066912 0.87192 0.95749 0.15721 0.52222 0.53766 0.69861 0.61072 0.37912 0.37197 0.42661 1.0671 1.0539 15.9986 144.9363 0.00068305 -6.0757 0.017947
6.122 0.9881 5.4837e-005 3.8183 0.01196 7.9903e-005 0.0011641 0.23311 0.00065931 0.23376 0.2157 0 0.032289 0.0389 0 1.3729 0.47302 0.14413 0.017536 11.1129 0.10915 0.00013957 0.78099 0.0084168 0.0093486 0.98735 5.6314e-012 0.0050716 0.84287 0.94558 0.15721 0.51069 0.52315 0.67506 0.59363 0.37447 0.37666 0.42641 1.0688 1.0581 15.9984 144.9354 0.00068649 -8.0666 0.018947
6.123 0.9881 5.4837e-005 3.8183 0.01196 7.9916e-005 0.0011641 0.23311 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.373 0.47307 0.14414 0.017538 11.1152 0.10915 0.00013959 0.78099 0.0084173 0.0093492 0.98356 -2.7351e-012 0.0038634 0.80505 0.92888 0.15721 0.50068 0.51068 0.64876 0.57706 0.37063 0.38007 0.4262 1.0708 1.0616 15.9982 144.9346 0.00068925 -10.4171 0.019947
6.124 0.9881 5.4837e-005 3.8183 0.01196 7.9929e-005 0.0011641 0.23311 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.3731 0.47311 0.14416 0.017539 11.1175 0.10916 0.0001396 0.78098 0.0084179 0.0093497 0.97741 2.3966e-012 0.0029646 0.75481 0.90474 0.15722 0.49224 0.5004 0.61923 0.56102 0.36763 0.38215 0.426 1.0731 1.0649 15.998 144.9339 0.00069125 -13.2703 0.020947
6.125 0.9881 5.4837e-005 3.8183 0.01196 7.9942e-005 0.0011641 0.23311 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.3732 0.47316 0.14417 0.01754 11.1198 0.10917 0.00013961 0.78097 0.0084184 0.0093503 0.9665 -1.5836e-012 0.0023004 0.68697 0.86877 0.15722 0.48543 0.49248 0.5861 0.54556 0.36545 0.38291 0.4258 1.0754 1.0679 15.9978 144.9333 0.00069238 -16.804 0.021947
6.126 0.9881 5.4837e-005 3.8183 0.01196 7.9954e-005 0.0011641 0.23311 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.3733 0.47321 0.14419 0.017542 11.1221 0.10918 0.00013962 0.78096 0.0084189 0.0093509 0.94548 -4.2926e-014 0.0018169 0.59498 0.81407 0.15723 0.48021 0.48694 0.54933 0.53081 0.364 0.3824 0.4256 1.0779 1.0707 15.9976 144.9328 0.00069254 -21.1754 0.022947
6.127 0.9881 5.4837e-005 3.8183 0.01196 7.9967e-005 0.0011641 0.23311 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.3734 0.47325 0.1442 0.017543 11.1244 0.10919 0.00013963 0.78095 0.0084194 0.0093514 0.90323 1.7746e-013 0.0014749 0.47367 0.73118 0.15723 0.4764 0.48357 0.50913 0.51707 0.36313 0.38075 0.42539 1.0804 1.0735 15.9974 144.9323 0.00069173 -26.3596 0.023947
6.128 0.9881 5.4837e-005 3.8183 0.01196 7.998e-005 0.0011642 0.23312 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.3734 0.4733 0.14422 0.017544 11.1267 0.1092 0.00013965 0.78094 0.00842 0.009352 0.82356 -6.2334e-014 0.0012429 0.32817 0.61209 0.15723 0.47366 0.4818 0.46512 0.5051 0.36268 0.37808 0.42519 1.083 1.0762 15.9973 144.9319 0.00069015 -31.9307 0.024947
6.129 0.9881 5.4837e-005 3.8183 0.01196 7.9993e-005 0.0011642 0.23312 0.00065931 0.23377 0.2157 0 0.032288 0.0389 0 1.3735 0.47335 0.14423 0.017546 11.129 0.1092 0.00013966 0.78094 0.0084205 0.0093526 0.70133 3.5247e-014 0.0010906 0.18507 0.46128 0.15724 0.47166 0.48091 0.41553 0.49621 0.36248 0.37431 0.42499 1.0855 1.0789 15.9972 144.9316 0.00068817 -37.1744 0.025947
6.13 0.9881 5.4836e-005 3.8183 0.01196 8.0006e-005 0.0011642 0.23312 0.00065931 0.23377 0.21571 0 0.032288 0.0389 0 1.3736 0.47339 0.14425 0.017547 11.1313 0.10921 0.00013967 0.78093 0.008421 0.0093531 0.55895 0.00015918 0.0010358 0.08055 0.30357 0.15724 0.47016 0.48062 0.35872 0.49146 0.36243 0.36911 0.4248 1.0881 1.0815 15.9971 144.9314 0.00068605 -41.6602 0.026947
6.131 0.9881 5.4836e-005 3.8183 0.01196 8.0019e-005 0.0011642 0.23312 0.00065931 0.23377 0.21571 0 0.032288 0.0389 0 1.3737 0.47344 0.14426 0.017548 11.1336 0.10922 0.00013968 0.78092 0.0084216 0.0093537 0.42769 0.00072882 0.0012253 0.026816 0.17124 0.15725 0.46905 0.48119 0.29562 0.49037 0.36247 0.36211 0.4246 1.0907 1.0842 15.9971 144.9312 0.00068388 -45.3697 0.027947
6.132 0.9881 5.4836e-005 3.8183 0.01196 8.0032e-005 0.0011642 0.23312 0.00065931 0.23377 0.21571 0 0.032288 0.0389 0 1.3738 0.47348 0.14428 0.01755 11.1359 0.10923 0.00013969 0.78091 0.0084221 0.0093543 0.32443 0.0016552 0.001677 0.0075415 0.082614 0.15725 0.46828 0.48284 0.23055 0.49134 0.36257 0.35302 0.42441 1.0933 1.0868 15.997 144.9311 0.00068166 -48.405 0.028947
6.133 0.9881 5.4836e-005 3.8183 0.01196 8.0045e-005 0.0011642 0.23312 0.00065931 0.23377 0.21571 0 0.032288 0.0389 0 1.3739 0.47353 0.14429 0.017551 11.1382 0.10924 0.00013971 0.7809 0.0084226 0.0093548 0.24994 0.0030432 0.0024157 0.0024496 0.034948 0.15725 0.4678 0.48538 0.16968 0.4931 0.36269 0.34174 0.42422 1.0958 1.0894 15.997 144.931 0.00067942 -50.8797 0.029947
6.134 0.9881 5.4836e-005 3.8183 0.01196 8.0058e-005 0.0011642 0.23312 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.374 0.47358 0.14431 0.017552 11.1405 0.10924 0.00013972 0.78089 0.0084231 0.0093554 0.19759 0.0049701 0.0034528 0.0012248 0.013939 0.15726 0.46756 0.4884 0.11841 0.49505 0.36283 0.32836 0.42403 1.0984 1.092 15.997 144.9309 0.00067715 -52.9115 0.030947
6.135 0.9881 5.4836e-005 3.8183 0.01196 8.0071e-005 0.0011642 0.23312 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.3741 0.47362 0.14432 0.017554 11.1428 0.10925 0.00013973 0.78089 0.0084237 0.009356 0.16028 0.0074925 0.004791 0.00081927 0.0060187 0.15726 0.46754 0.49163 0.079396 0.49699 0.36297 0.31311 0.42385 1.101 1.0946 15.997 144.9308 0.00067487 -54.6146 0.031947
6.136 0.9881 5.4836e-005 3.8183 0.01196 8.0084e-005 0.0011642 0.23312 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.3742 0.47367 0.14433 0.017555 11.1451 0.10926 0.00013974 0.78088 0.0084242 0.0093565 0.1327 0.010659 0.0064309 0.00060927 0.0032328 0.15727 0.46768 0.49489 0.052309 0.49883 0.36313 0.29628 0.42366 1.1036 1.0972 15.997 144.9308 0.00067257 -56.0881 0.032947
6.137 0.9881 5.4836e-005 3.8183 0.01196 8.0096e-005 0.0011642 0.23312 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.3743 0.47371 0.14435 0.017557 11.1474 0.10927 0.00013975 0.78087 0.0084247 0.0093571 0.11144 0.014524 0.0083771 0.00047373 0.002162 0.15727 0.46798 0.49816 0.034933 0.50057 0.36328 0.27816 0.42348 1.1061 1.0998 15.997 144.9308 0.00067027 -57.4083 0.033947
6.138 0.9881 5.4836e-005 3.8183 0.01196 8.0109e-005 0.0011642 0.23312 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.3744 0.47376 0.14436 0.017558 11.1497 0.10928 0.00013977 0.78086 0.0084252 0.0093577 0.094446 0.019157 0.010641 0.00037762 0.0016321 0.15728 0.46841 0.50139 0.024453 0.50222 0.36344 0.25904 0.42331 1.1087 1.1023 15.997 144.9307 0.00066796 -58.6284 0.034947
6.139 0.9881 5.4836e-005 3.8183 0.01196 8.0122e-005 0.0011642 0.23313 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.3745 0.47381 0.14438 0.017559 11.152 0.10929 0.00013978 0.78085 0.0084258 0.0093582 0.080495 0.024643 0.013239 0.0003052 0.0012942 0.15728 0.46896 0.5046 0.018357 0.50378 0.3636 0.23917 0.42314 1.1113 1.1049 15.997 144.9307 0.00066565 -59.7821 0.035947
6.14 0.9881 5.4836e-005 3.8183 0.01196 8.0135e-005 0.0011642 0.23313 0.00065931 0.23378 0.21571 0 0.032288 0.0389 0 1.3746 0.47385 0.14439 0.017561 11.1543 0.10929 0.00013979 0.78085 0.0084263 0.0093588 0.068854 0.031089 0.016194 0.00024963 0.0010475 0.15728 0.46961 0.50777 0.014799 0.50526 0.36376 0.21882 0.42297 1.1139 1.1075 15.997 144.9307 0.00066333 -60.8889 0.036947
6.141 0.9881 5.4836e-005 3.8183 0.01196 8.0148e-005 0.0011642 0.23313 0.00065931 0.23378 0.21572 0 0.032288 0.0389 0 1.3747 0.4739 0.14441 0.017562 11.1566 0.1093 0.0001398 0.78084 0.0084268 0.0093594 0.059052 0.038615 0.019534 0.00020541 0.00085696 0.15729 0.47036 0.51091 0.012602 0.50668 0.36391 0.19827 0.4228 1.1164 1.1101 15.997 144.9307 0.00066101 -61.9597 0.037947
6.142 0.9881 5.4836e-005 3.8183 0.01196 8.0161e-005 0.0011642 0.23313 0.00065931 0.23378 0.21572 0 0.032288 0.0389 0 1.3747 0.47395 0.14442 0.017563 11.1589 0.10931 0.00013981 0.78083 0.0084274 0.0093599 0.050759 0.047352 0.023289 0.00017021 0.00070652 0.15729 0.4712 0.51402 0.011104 0.50803 0.36407 0.17777 0.42264 1.119 1.1127 15.9971 144.9306 0.00065868 -62.9999 0.038947
6.143 0.9881 5.4835e-005 3.8183 0.01196 8.0174e-005 0.0011642 0.23313 0.00065931 0.23378 0.21572 0 0.032288 0.0389 0 1.3748 0.47399 0.14444 0.017565 11.1613 0.10932 0.00013983 0.78082 0.0084279 0.0093605 0.043725 0.057444 0.027492 0.0001418 0.00058615 0.1573 0.47211 0.5171 0.0099675 0.50934 0.36423 0.15764 0.42248 1.1215 1.1153 15.9971 144.9306 0.00065636 -64.0126 0.039947
6.144 0.9881 5.4835e-005 3.8183 0.01196 8.0187e-005 0.0011642 0.23313 0.00065931 0.23379 0.21572 0 0.032288 0.0389 0 1.3749 0.47404 0.14445 0.017566 11.1636 0.10933 0.00013984 0.78081 0.0084284 0.0093611 0.037749 0.069036 0.032178 0.00011871 0.00048906 0.1573 0.4731 0.52014 0.0090357 0.51061 0.36439 0.13814 0.42232 1.1241 1.1178 15.9972 144.9306 0.00065403 -64.9992 0.040947
6.145 0.9881 5.4835e-005 3.8183 0.01196 8.02e-005 0.0011642 0.23313 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.375 0.47408 0.14447 0.017567 11.1659 0.10934 0.00013985 0.7808 0.0084289 0.0093616 0.032666 0.082279 0.037385 9.9878e-005 0.0004102 0.1573 0.47415 0.52315 0.0082375 0.51184 0.36455 0.11955 0.42217 1.1267 1.1204 15.9972 144.9306 0.0006517 -65.9606 0.041947
6.146 0.9881 5.4835e-005 3.8183 0.01196 8.0213e-005 0.0011642 0.23313 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.3751 0.47413 0.14448 0.017569 11.1682 0.10934 0.00013986 0.7808 0.0084295 0.0093622 0.028337 0.097318 0.043155 8.442e-005 0.0003458 0.15731 0.47525 0.52613 0.0075395 0.51306 0.36471 0.10212 0.42203 1.1292 1.123 15.9973 144.9305 0.00064937 -66.8974 0.042947
6.147 0.9881 5.4835e-005 3.8183 0.01196 8.0226e-005 0.0011642 0.23313 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.3752 0.47418 0.1445 0.01757 11.1705 0.10935 0.00013987 0.78079 0.00843 0.0093628 0.024645 0.1143 0.049534 7.1682e-005 0.00029294 0.15731 0.47641 0.52907 0.0069233 0.51425 0.36488 0.086065 0.42188 1.1318 1.1256 15.9973 144.9305 0.00064704 -67.8098 0.043947
6.148 0.9881 5.4835e-005 3.8183 0.01196 8.0239e-005 0.0011642 0.23313 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.3753 0.47422 0.14451 0.017571 11.1728 0.10936 0.00013989 0.78078 0.0084305 0.0093633 0.021494 0.13334 0.05657 6.1146e-005 0.00024936 0.15732 0.4776 0.53198 0.006376 0.51544 0.36504 0.071544 0.42175 1.1343 1.1281 15.9974 144.9305 0.00064472 -68.6976 0.044947
6.149 0.9881 5.4835e-005 3.8183 0.01196 8.0251e-005 0.0011642 0.23314 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.3754 0.47427 0.14453 0.017573 11.1751 0.10937 0.0001399 0.78077 0.008431 0.0093639 0.018801 0.15455 0.064318 5.2396e-005 0.00021329 0.15732 0.47884 0.53487 0.0058886 0.51662 0.3652 0.058663 0.42161 1.1369 1.1307 15.9974 144.9304 0.00064239 -69.5606 0.045947
6.15 0.9881 5.4835e-005 3.8183 0.01196 8.0264e-005 0.0011642 0.23314 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.3755 0.47431 0.14454 0.017574 11.1774 0.10938 0.00013991 0.78076 0.0084316 0.0093645 0.016498 0.17801 0.072837 4.5111e-005 0.00018332 0.15733 0.48011 0.53772 0.0054534 0.5178 0.36536 0.047467 0.42149 1.1394 1.1333 15.9975 144.9304 0.00064006 -70.3982 0.046947
6.151 0.9881 5.4835e-005 3.8183 0.011959 8.0277e-005 0.0011642 0.23314 0.00065931 0.23379 0.21572 0 0.032287 0.0389 0 1.3756 0.47436 0.14456 0.017575 11.1797 0.10938 0.00013992 0.78076 0.0084321 0.009365 0.014526 0.20376 0.08219 3.9021e-005 0.00015834 0.15733 0.48141 0.54054 0.0050641 0.519 0.36552 0.037939 0.42137 1.142 1.1358 15.9976 144.9304 0.00063774 -71.2098 0.047947
6.152 0.9881 5.4835e-005 3.8183 0.011959 8.029e-005 0.0011642 0.23314 0.00065931 0.23379 0.21573 0 0.032287 0.0389 0 1.3757 0.47441 0.14457 0.017577 11.182 0.10939 0.00013993 0.78075 0.0084326 0.0093656 0.012836 0.23179 0.092442 3.3919e-005 0.00013745 0.15733 0.48274 0.54332 0.0047154 0.5202 0.36569 0.030006 0.42125 1.1445 1.1384 15.9976 144.9303 0.00063542 -71.9944 0.048947
6.153 0.9881 5.4835e-005 3.8183 0.011959 8.0303e-005 0.0011642 0.23314 0.00065931 0.23379 0.21573 0 0.032287 0.0389 0 1.3758 0.47445 0.14459 0.017578 11.1843 0.1094 0.00013995 0.78074 0.0084331 0.0093662 0.011387 0.26204 0.10366 2.9636e-005 0.00011995 0.15734 0.48409 0.54608 0.0044028 0.52142 0.36586 0.023546 0.42114 1.147 1.1409 15.9977 144.9303 0.0006331 -72.7511 0.049947
6.154 0.9881 5.4835e-005 3.8183 0.011959 8.0316e-005 0.0011642 0.23314 0.00065931 0.23379 0.21573 0 0.032287 0.0389 0 1.3759 0.4745 0.1446 0.01758 11.1866 0.10941 0.00013996 0.78073 0.0084337 0.0093667 0.010142 0.2944 0.1159 2.6027e-005 0.00010523 0.15734 0.48545 0.54881 0.0041226 0.52267 0.36602 0.018404 0.42103 1.1496 1.1435 15.9978 144.9303 0.00063078 -73.4787 0.050947
6.155 0.9881 5.4835e-005 3.8183 0.011959 8.0329e-005 0.0011643 0.23314 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3759 0.47455 0.14462 0.017581 11.189 0.10942 0.00013997 0.78072 0.0084342 0.0093673 0.0090739 0.32867 0.12923 2.2983e-005 9.2824e-005 0.15735 0.48684 0.55151 0.0038712 0.52394 0.36619 0.014399 0.42093 1.1521 1.146 15.9979 144.9303 0.00062847 -74.1763 0.051947
6.156 0.9881 5.4834e-005 3.8183 0.011959 8.0342e-005 0.0011643 0.23314 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.376 0.47459 0.14463 0.017582 11.1913 0.10943 0.00013998 0.78071 0.0084347 0.0093679 0.0081554 0.36461 0.14369 2.0409e-005 8.2349e-005 0.15735 0.48824 0.55418 0.0036458 0.52524 0.36636 0.011348 0.42084 1.1546 1.1486 15.998 144.9302 0.00062616 -74.8429 0.052947
6.157 0.9881 5.4834e-005 3.8183 0.011959 8.0355e-005 0.0011643 0.23314 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3761 0.47464 0.14465 0.017584 11.1936 0.10943 0.00013999 0.78071 0.0084352 0.0093684 0.0073643 0.40189 0.15929 1.8225e-005 7.3479e-005 0.15735 0.48964 0.55683 0.0034438 0.52657 0.36653 0.0090685 0.42075 1.1572 1.1511 15.9981 144.9302 0.00062386 -75.4777 0.053947
6.158 0.9881 5.4834e-005 3.8183 0.011959 8.0368e-005 0.0011643 0.23314 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3762 0.47468 0.14466 0.017585 11.1959 0.10944 0.00014001 0.7807 0.0084358 0.009369 0.0066834 0.44016 0.17605 1.6371e-005 6.5952e-005 0.15736 0.49106 0.55944 0.0032627 0.52794 0.3667 0.0073948 0.42066 1.1597 1.1537 15.9982 144.9302 0.00062157 -76.0799 0.054947
6.159 0.9881 5.4834e-005 3.8183 0.011959 8.0381e-005 0.0011643 0.23314 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3763 0.47473 0.14468 0.017586 11.1982 0.10945 0.00014002 0.78069 0.0084363 0.0093696 0.0060961 0.47899 0.19393 1.4792e-005 5.955e-005 0.15736 0.49249 0.56203 0.0031004 0.52935 0.36688 0.0061829 0.42058 1.1622 1.1562 15.9983 144.9302 0.00061927 -76.6493 0.055947
6.16 0.9881 5.4834e-005 3.8183 0.011959 8.0393e-005 0.0011643 0.23315 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3764 0.47478 0.14469 0.017588 11.2005 0.10946 0.00014003 0.78068 0.0084368 0.0093701 0.0055889 0.51795 0.21289 1.3445e-005 5.4091e-005 0.15737 0.49392 0.56459 0.0029552 0.5308 0.36705 0.0053128 0.42051 1.1647 1.1588 15.9984 144.9301 0.00061699 -77.1856 0.056947
6.161 0.9881 5.4834e-005 3.8183 0.011959 8.0406e-005 0.0011643 0.23315 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3765 0.47482 0.14471 0.017589 11.2028 0.10947 0.00014004 0.78067 0.0084373 0.0093707 0.0051505 0.55659 0.23284 1.2292e-005 4.9425e-005 0.15737 0.49536 0.56712 0.0028252 0.53228 0.36723 0.0046887 0.42044 1.1672 1.1613 15.9985 144.9301 0.00061471 -77.689 0.057947
6.162 0.9881 5.4834e-005 3.8183 0.011959 8.0419e-005 0.0011643 0.23315 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3766 0.47487 0.14472 0.01759 11.2051 0.10948 0.00014005 0.78067 0.0084379 0.0093713 0.0047706 0.59448 0.25368 1.1304e-005 4.5427e-005 0.15737 0.49681 0.56963 0.0027089 0.53381 0.36741 0.0042379 0.42037 1.1698 1.1638 15.9986 144.9301 0.00061244 -78.16 0.058947
6.163 0.9881 5.4834e-005 3.8183 0.011959 8.0432e-005 0.0011643 0.23315 0.00065931 0.2338 0.21573 0 0.032287 0.0389 0 1.3767 0.47491 0.14474 0.017592 11.2075 0.10948 0.00014007 0.78066 0.0084384 0.0093718 0.0044413 0.63119 0.27529 1.0454e-005 4.1992e-005 0.15738 0.49825 0.57211 0.0026048 0.53538 0.36759 0.0039071 0.42031 1.1723 1.1664 15.9987 144.9301 0.00061018 -78.5991 0.059947
6.164 0.9881 5.4834e-005 3.8183 0.011959 8.0445e-005 0.0011643 0.23315 0.00065931 0.2338 0.21574 0 0.032287 0.0389 0 1.3768 0.47496 0.14475 0.017593 11.2098 0.10949 0.00014008 0.78065 0.0084389 0.0093724 0.0041553 0.66637 0.29754 9.7215e-006 3.9033e-005 0.15738 0.4997 0.57456 0.0025118 0.537 0.36777 0.0036586 0.42025 1.1748 1.1689 15.9988 144.93 0.00060792 -79.0072 0.060947
6.165 0.9881 5.4834e-005 3.8183 0.011959 8.0458e-005 0.0011643 0.23315 0.00065931 0.2338 0.21574 0 0.032287 0.0389 0 1.3769 0.47501 0.14477 0.017594 11.2121 0.1095 0.00014009 0.78064 0.0084394 0.0093729 0.003906 0.69971 0.32027 9.0888e-006 3.6478e-005 0.15739 0.50115 0.57699 0.0024286 0.53865 0.36796 0.0034668 0.4202 1.1773 1.1714 15.9989 144.93 0.00060568 -79.3855 0.061947
6.166 0.9881 5.4834e-005 3.8183 0.011959 8.0471e-005 0.0011643 0.23315 0.00065931 0.23381 0.21574 0 0.032287 0.0389 0 1.377 0.47505 0.14478 0.017596 11.2144 0.10951 0.0001401 0.78063 0.00844 0.0093735 0.0036884 0.73096 0.34335 8.5404e-006 3.4266e-005 0.15739 0.5026 0.5794 0.0023542 0.54034 0.36814 0.0033141 0.42015 1.1798 1.1739 15.999 144.93 0.00060344 -79.7353 0.062947
6.167 0.9881 5.4834e-005 3.8183 0.011959 8.0484e-005 0.0011643 0.23315 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3771 0.4751 0.1448 0.017597 11.2167 0.10952 0.00014011 0.78062 0.0084405 0.0093741 0.0034987 0.75996 0.36663 8.0641e-006 3.2345e-005 0.15739 0.50405 0.58178 0.0022876 0.54207 0.36833 0.0031891 0.4201 1.1823 1.1764 15.9991 144.93 0.00060121 -80.0578 0.063947
6.168 0.9881 5.4834e-005 3.8183 0.011959 8.0497e-005 0.0011643 0.23315 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3772 0.47514 0.14481 0.017598 11.219 0.10952 0.00014013 0.78062 0.008441 0.0093746 0.0033326 0.78661 0.38997 7.6496e-006 3.0673e-005 0.1574 0.5055 0.58413 0.002228 0.54384 0.36852 0.0030842 0.42006 1.1848 1.1789 15.9992 144.93 0.00059899 -80.3546 0.064947
6.169 0.9881 5.4833e-005 3.8183 0.011959 8.051e-005 0.0011643 0.23315 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3772 0.47519 0.14483 0.0176 11.2213 0.10953 0.00014014 0.78061 0.0084415 0.0093752 0.0031864 0.81086 0.41325 7.2877e-006 2.9215e-005 0.1574 0.50695 0.58646 0.0021747 0.54564 0.36871 0.0029945 0.42002 1.1873 1.1815 15.9993 144.93 0.00059678 -80.6273 0.065947
6.17 0.9881 5.4833e-005 3.8183 0.011959 8.0523e-005 0.0011643 0.23315 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3773 0.47524 0.14484 0.017601 11.2237 0.10954 0.00014015 0.7806 0.0084421 0.0093758 0.0030582 0.83273 0.43635 6.9706e-006 2.7938e-005 0.15741 0.5084 0.58877 0.002127 0.54747 0.3689 0.0029168 0.41998 1.1898 1.184 15.9994 144.93 0.00059458 -80.8773 0.066947
6.171 0.9881 5.4833e-005 3.8183 0.011959 8.0535e-005 0.0011643 0.23316 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3774 0.47528 0.14486 0.017602 11.226 0.10955 0.00014016 0.78059 0.0084426 0.0093763 0.0029452 0.85231 0.45917 6.6926e-006 2.6818e-005 0.15741 0.50984 0.59105 0.0020842 0.54933 0.36909 0.0028487 0.41995 1.1922 1.1865 15.9995 144.93 0.00059239 -81.1062 0.067947
6.172 0.9881 5.4833e-005 3.8183 0.011959 8.0548e-005 0.0011643 0.23316 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3775 0.47533 0.14487 0.017604 11.2283 0.10956 0.00014017 0.78058 0.0084431 0.0093769 0.0028453 0.86968 0.48161 6.4481e-006 2.5833e-005 0.15742 0.51129 0.59332 0.0020458 0.55122 0.36928 0.0027888 0.41992 1.1947 1.189 15.9996 144.9299 0.00059021 -81.3156 0.068947
6.173 0.9881 5.4833e-005 3.8183 0.011959 8.0561e-005 0.0011643 0.23316 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3776 0.47538 0.14488 0.017605 11.2306 0.10957 0.00014019 0.78057 0.0084436 0.0093775 0.002757 0.885 0.50361 6.2324e-006 2.4965e-005 0.15742 0.51273 0.59555 0.0020114 0.55314 0.36947 0.0027357 0.41989 1.1972 1.1915 15.9997 144.9299 0.00058805 -81.507 0.069947
6.174 0.9881 5.4833e-005 3.8183 0.011959 8.0574e-005 0.0011643 0.23316 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3777 0.47542 0.1449 0.017606 11.2329 0.10957 0.0001402 0.78057 0.0084442 0.009378 0.0026787 0.89842 0.5251 6.0417e-006 2.4198e-005 0.15742 0.51417 0.59777 0.0019805 0.55507 0.36967 0.0026885 0.41986 1.1997 1.194 15.9999 144.9299 0.00058589 -81.6818 0.070947
6.175 0.9881 5.4833e-005 3.8183 0.011959 8.0587e-005 0.0011643 0.23316 0.00065931 0.23381 0.21574 0 0.032286 0.0389 0 1.3778 0.47547 0.14491 0.017608 11.2352 0.10958 0.00014021 0.78056 0.0084447 0.0093786 0.0026091 0.9101 0.54602 5.8728e-006 2.3519e-005 0.15743 0.5156 0.59996 0.0019527 0.55703 0.36986 0.0026464 0.41983 1.2022 1.1965 16 144.9299 0.00058374 -81.8413 0.071947
6.176 0.9881 5.4833e-005 3.8183 0.011959 8.06e-005 0.0011643 0.23316 0.00065931 0.23381 0.21575 0 0.032286 0.0389 0 1.3779 0.47551 0.14493 0.017609 11.2376 0.10959 0.00014022 0.78055 0.0084452 0.0093792 0.0025471 0.92021 0.56634 5.7228e-006 2.2915e-005 0.15743 0.51703 0.60214 0.0019277 0.55901 0.37006 0.0026088 0.41981 1.2046 1.1989 16.0001 144.9299 0.00058161 -81.987 0.072947
6.177 0.9881 5.4833e-005 3.8183 0.011959 8.0613e-005 0.0011643 0.23316 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.378 0.47556 0.14494 0.017611 11.2399 0.1096 0.00014023 0.78054 0.0084457 0.0093797 0.0024918 0.92892 0.58602 5.5892e-006 2.2378e-005 0.15744 0.51846 0.60429 0.0019051 0.561 0.37025 0.0025751 0.41978 1.2071 1.2014 16.0002 144.9299 0.00057948 -82.1199 0.073947
6.178 0.9881 5.4833e-005 3.8183 0.011959 8.0626e-005 0.0011643 0.23316 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3781 0.47561 0.14496 0.017612 11.2422 0.10961 0.00014024 0.78053 0.0084463 0.0093803 0.0024424 0.9364 0.60504 5.47e-006 2.1899e-005 0.15744 0.51989 0.60642 0.0018848 0.563 0.37045 0.0025449 0.41976 1.2096 1.2039 16.0003 144.9299 0.00057737 -82.2413 0.074947
6.179 0.9881 5.4833e-005 3.8183 0.011959 8.0639e-005 0.0011643 0.23316 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3782 0.47565 0.14497 0.017613 11.2445 0.10961 0.00014026 0.78053 0.0084468 0.0093808 0.002398 0.9428 0.62339 5.3633e-006 2.147e-005 0.15744 0.52132 0.60853 0.0018664 0.56502 0.37065 0.0025177 0.41974 1.212 1.2064 16.0004 144.9299 0.00057527 -82.3522 0.075947
6.18 0.9881 5.4833e-005 3.8183 0.011959 8.0652e-005 0.0011643 0.23316 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3783 0.4757 0.14499 0.017615 11.2468 0.10962 0.00014027 0.78052 0.0084473 0.0093814 0.0023582 0.94824 0.64106 5.2675e-006 2.1085e-005 0.15745 0.52274 0.61061 0.0018497 0.56705 0.37085 0.0024932 0.41972 1.2145 1.2089 16.0005 144.9299 0.00057317 -82.4535 0.076947
6.181 0.9881 5.4833e-005 3.8183 0.011959 8.0665e-005 0.0011643 0.23316 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3784 0.47574 0.145 0.017616 11.2492 0.10963 0.00014028 0.78051 0.0084478 0.009382 0.0023223 0.95287 0.65804 5.1816e-006 2.0739e-005 0.15745 0.52415 0.61268 0.0018346 0.56909 0.37104 0.0024711 0.4197 1.2169 1.2113 16.0006 144.9299 0.0005711 -82.5462 0.077947
6.182 0.9881 5.4832e-005 3.8183 0.011959 8.0677e-005 0.0011643 0.23317 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3784 0.47579 0.14502 0.017617 11.2515 0.10964 0.00014029 0.7805 0.0084484 0.0093825 0.0022897 0.9568 0.67434 5.1043e-006 2.0428e-005 0.15746 0.52557 0.61473 0.0018209 0.57113 0.37124 0.0024511 0.41969 1.2194 1.2138 16.0007 144.9299 0.00056903 -82.6312 0.078947
6.183 0.9881 5.4832e-005 3.8183 0.011959 8.069e-005 0.0011644 0.23317 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3785 0.47584 0.14503 0.017619 11.2538 0.10965 0.0001403 0.78049 0.0084489 0.0093831 0.0022606 0.96012 0.68996 5.0338e-006 2.0146e-005 0.15746 0.52697 0.61676 0.0018084 0.57319 0.37144 0.002433 0.41967 1.2218 1.2163 16.0009 144.9299 0.00056697 -82.7091 0.079947
6.184 0.9881 5.4832e-005 3.8183 0.011959 8.0703e-005 0.0011644 0.23317 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3786 0.47588 0.14505 0.01762 11.2561 0.10966 0.00014032 0.78048 0.0084494 0.0093837 0.0022341 0.96293 0.70492 4.9701e-006 1.989e-005 0.15746 0.52838 0.61877 0.001797 0.57524 0.37164 0.0024165 0.41965 1.2243 1.2187 16.001 144.9299 0.00056492 -82.7806 0.080947
6.185 0.9881 5.4832e-005 3.8183 0.011959 8.0716e-005 0.0011644 0.23317 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3787 0.47593 0.14506 0.017621 11.2584 0.10966 0.00014033 0.78048 0.0084499 0.0093842 0.0022098 0.9653 0.71923 4.9125e-006 1.9658e-005 0.15747 0.52978 0.62076 0.0017866 0.5773 0.37184 0.0024015 0.41964 1.2267 1.2212 16.0011 144.9299 0.00056289 -82.8465 0.081947
6.186 0.9881 5.4832e-005 3.8183 0.011959 8.0729e-005 0.0011644 0.23317 0.00065931 0.23382 0.21575 0 0.032286 0.0389 0 1.3788 0.47597 0.14508 0.017623 11.2608 0.10967 0.00014034 0.78047 0.0084505 0.0093848 0.0021875 0.96731 0.7329 4.86e-006 1.9447e-005 0.15747 0.53118 0.62273 0.001777 0.57936 0.37204 0.0023878 0.41962 1.2292 1.2237 16.0012 144.9299 0.00056087 -82.9072 0.082947
6.187 0.9881 5.4832e-005 3.8183 0.011959 8.0742e-005 0.0011644 0.23317 0.00065931 0.23382 0.21576 0 0.032286 0.0389 0 1.3789 0.47602 0.14509 0.017624 11.2631 0.10968 0.00014035 0.78046 0.008451 0.0093854 0.0021672 0.96901 0.74596 4.8119e-006 1.9254e-005 0.15748 0.53257 0.62468 0.0017682 0.58142 0.37224 0.0023753 0.41961 1.2316 1.2261 16.0013 144.9299 0.00055886 -82.9633 0.083947
6.188 0.9881 5.4832e-005 3.8183 0.011959 8.0755e-005 0.0011644 0.23317 0.00065931 0.23383 0.21576 0 0.032286 0.0389 0 1.379 0.47607 0.14511 0.017625 11.2654 0.10969 0.00014036 0.78045 0.0084515 0.0093859 0.0021487 0.97044 0.75841 4.7677e-006 1.9077e-005 0.15748 0.53396 0.62661 0.0017602 0.58349 0.37244 0.0023638 0.4196 1.234 1.2286 16.0014 144.9299 0.00055685 -83.0152 0.084947
6.189 0.9881 5.4832e-005 3.8183 0.011959 8.0768e-005 0.0011644 0.23317 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3791 0.47611 0.14512 0.017627 11.2677 0.1097 0.00014038 0.78044 0.008452 0.0093865 0.0021319 0.97166 0.77027 4.727e-006 1.8914e-005 0.15749 0.53535 0.62852 0.0017527 0.58555 0.37265 0.0023532 0.41959 1.2364 1.231 16.0015 144.9299 0.00055487 -83.0633 0.085947
6.19 0.9881 5.4832e-005 3.8183 0.011959 8.0781e-005 0.0011644 0.23317 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3792 0.47616 0.14514 0.017628 11.2701 0.1097 0.00014039 0.78044 0.0084525 0.009387 0.0021162 0.97269 0.78158 4.6895e-006 1.8764e-005 0.15749 0.53673 0.63042 0.0017458 0.58761 0.37285 0.0023435 0.41957 1.2389 1.2334 16.0016 144.9299 0.00055289 -83.1081 0.086947
6.191 0.9881 5.4832e-005 3.8183 0.011959 8.0794e-005 0.0011644 0.23317 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3793 0.47621 0.14515 0.017629 11.2724 0.10971 0.0001404 0.78043 0.0084531 0.0093876 0.0021016 0.97356 0.79234 4.6549e-006 1.8625e-005 0.15749 0.53811 0.6323 0.0017394 0.58967 0.37305 0.0023345 0.41956 1.2413 1.2359 16.0017 144.9299 0.00055092 -83.1499 0.087947
6.192 0.9881 5.4832e-005 3.8183 0.011959 8.0807e-005 0.0011644 0.23317 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3794 0.47625 0.14517 0.017631 11.2747 0.10972 0.00014041 0.78042 0.0084536 0.0093882 0.0020879 0.97431 0.80259 4.6229e-006 1.8496e-005 0.1575 0.53949 0.63416 0.0017334 0.59173 0.37325 0.0023261 0.41955 1.2437 1.2383 16.0018 144.9299 0.00054896 -83.189 0.088947
6.193 0.9881 5.4832e-005 3.8183 0.011959 8.082e-005 0.0011644 0.23317 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3795 0.4763 0.14518 0.017632 11.277 0.10973 0.00014042 0.78041 0.0084541 0.0093887 0.0020751 0.97495 0.81233 4.593e-006 1.8376e-005 0.1575 0.54086 0.636 0.0017278 0.59379 0.37345 0.0023183 0.41954 1.2461 1.2407 16.0019 144.9299 0.00054702 -83.2256 0.089947
6.194 0.9881 5.4831e-005 3.8183 0.011959 8.0832e-005 0.0011644 0.23318 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3796 0.47634 0.1452 0.017633 11.2794 0.10974 0.00014044 0.7804 0.0084546 0.0093893 0.0020633 0.9755 0.82159 4.565e-006 1.8264e-005 0.15751 0.54222 0.63783 0.0017226 0.59584 0.37365 0.0023111 0.41953 1.2485 1.2432 16.002 144.9299 0.00054508 -83.2601 0.090947
6.195 0.9881 5.4831e-005 3.8183 0.011959 8.0845e-005 0.0011644 0.23318 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3796 0.47639 0.14521 0.017635 11.2817 0.10975 0.00014045 0.7804 0.0084552 0.0093898 0.0020524 0.97598 0.83039 4.5387e-006 1.8159e-005 0.15751 0.54359 0.63964 0.0017177 0.59789 0.37386 0.0023043 0.41952 1.2509 1.2456 16.0021 144.9299 0.00054316 -83.2925 0.091947
6.196 0.9881 5.4831e-005 3.8183 0.011959 8.0858e-005 0.0011644 0.23318 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3797 0.47644 0.14523 0.017636 11.284 0.10975 0.00014046 0.78039 0.0084557 0.0093904 0.0020421 0.97639 0.83875 4.514e-006 1.806e-005 0.15751 0.54495 0.64143 0.001713 0.59993 0.37406 0.0022979 0.41951 1.2533 1.248 16.0022 144.9299 0.00054125 -83.3232 0.092947
6.197 0.9881 5.4831e-005 3.8183 0.011959 8.0871e-005 0.0011644 0.23318 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3798 0.47648 0.14524 0.017637 11.2863 0.10976 0.00014047 0.78038 0.0084562 0.009391 0.0020323 0.97675 0.84669 4.4908e-006 1.7967e-005 0.15752 0.5463 0.64321 0.0017087 0.60197 0.37426 0.0022918 0.4195 1.2557 1.2504 16.0023 144.9299 0.00053935 -83.3523 0.093947
6.198 0.9881 5.4831e-005 3.8183 0.011959 8.0884e-005 0.0011644 0.23318 0.00065931 0.23383 0.21576 0 0.032285 0.0389 0 1.3799 0.47653 0.14526 0.017639 11.2887 0.10977 0.00014048 0.78037 0.0084567 0.0093915 0.002023 0.97707 0.85422 4.4688e-006 1.7878e-005 0.15752 0.54765 0.64497 0.0017045 0.604 0.37446 0.0022862 0.41949 1.2581 1.2529 16.0025 144.9299 0.00053746 -83.38 0.094947
6.199 0.9881 5.4831e-005 3.8183 0.011959 8.0897e-005 0.0011644 0.23318 0.00065931 0.23383 0.21577 0 0.032285 0.0389 0 1.38 0.47657 0.14527 0.01764 11.291 0.10978 0.0001405 0.78036 0.0084573 0.0093921 0.0020139 0.97735 0.86137 4.4481e-006 1.7795e-005 0.15753 0.549 0.64671 0.0017006 0.60603 0.37467 0.0022808 0.41948 1.2605 1.2553 16.0026 144.9299 0.00053558 -83.4064 0.095947
6.2 0.9881 5.4831e-005 3.8183 0.011959 8.091e-005 0.0011644 0.23318 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3801 0.47662 0.14529 0.017641 11.2933 0.10979 0.00014051 0.78035 0.0084578 0.0093927 0.0020054 0.97759 0.86816 4.4283e-006 1.7716e-005 0.15753 0.55034 0.64844 0.0016968 0.60806 0.37487 0.0022756 0.41948 1.2629 1.2577 16.0027 144.9299 0.00053371 -83.4316 0.096947
6.201 0.9881 5.4831e-005 3.8183 0.011959 8.0923e-005 0.0011644 0.23318 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3802 0.47667 0.1453 0.017643 11.2956 0.10979 0.00014052 0.78035 0.0084583 0.0093932 0.0019974 0.97782 0.8746 4.4094e-006 1.764e-005 0.15753 0.55168 0.65015 0.0016932 0.61007 0.37507 0.0022708 0.41947 1.2653 1.2601 16.0028 144.93 0.00053185 -83.4557 0.097947
6.202 0.9881 5.4831e-005 3.8183 0.011959 8.0936e-005 0.0011644 0.23318 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3803 0.47671 0.14532 0.017644 11.298 0.1098 0.00014053 0.78034 0.0084588 0.0093938 0.0019899 0.97802 0.8807 4.3912e-006 1.7567e-005 0.15754 0.55301 0.65185 0.0016898 0.61209 0.37528 0.0022661 0.41946 1.2677 1.2625 16.0029 144.93 0.00053 -83.4789 0.098947
6.203 0.9881 5.4831e-005 3.8183 0.011959 8.0949e-005 0.0011644 0.23318 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3804 0.47676 0.14533 0.017645 11.3003 0.10981 0.00014054 0.78033 0.0084593 0.0093943 0.0019827 0.9782 0.88649 4.3738e-006 1.7498e-005 0.15754 0.55434 0.65353 0.0016864 0.61409 0.37548 0.0022616 0.41945 1.2701 1.2649 16.003 144.93 0.00052816 -83.5013 0.099947
6.204 0.9881 5.4831e-005 3.8183 0.011959 8.0962e-005 0.0011644 0.23318 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3805 0.4768 0.14535 0.017647 11.3026 0.10982 0.00014056 0.78032 0.0084599 0.0093949 0.0019758 0.97836 0.89198 4.3571e-006 1.7431e-005 0.15755 0.55567 0.6552 0.0016833 0.61609 0.37568 0.0022573 0.41945 1.2724 1.2673 16.0031 144.93 0.00052633 -83.5228 0.10095
6.205 0.9881 5.4831e-005 3.8183 0.011959 8.0974e-005 0.0011644 0.23319 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3806 0.47685 0.14536 0.017648 11.3049 0.10983 0.00014057 0.78031 0.0084604 0.0093955 0.0019689 0.97851 0.89718 4.341e-006 1.7366e-005 0.15755 0.55699 0.65685 0.0016802 0.61809 0.37588 0.0022532 0.41944 1.2748 1.2696 16.0032 144.93 0.00052452 -83.5437 0.10195
6.206 0.9881 5.4831e-005 3.8183 0.011959 8.0987e-005 0.0011644 0.23319 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3807 0.4769 0.14537 0.01765 11.3073 0.10984 0.00014058 0.78031 0.0084609 0.009396 0.0019621 0.97865 0.90211 4.3256e-006 1.7304e-005 0.15755 0.55831 0.65849 0.0016772 0.62008 0.37609 0.0022492 0.41943 1.2772 1.272 16.0033 144.93 0.00052271 -83.5639 0.10295
6.207 0.9881 5.483e-005 3.8183 0.011959 8.1e-005 0.0011644 0.23319 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3808 0.47694 0.14539 0.017651 11.3096 0.10984 0.00014059 0.7803 0.0084614 0.0093966 0.0019555 0.97878 0.90678 4.3106e-006 1.7244e-005 0.15756 0.55963 0.66011 0.0016743 0.62206 0.37629 0.0022454 0.41943 1.2795 1.2744 16.0033 144.93 0.00052091 -83.5835 0.10395
6.208 0.9881 5.483e-005 3.8183 0.011959 8.1013e-005 0.0011644 0.23319 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3809 0.47699 0.1454 0.017652 11.3119 0.10985 0.0001406 0.78029 0.0084619 0.0093971 0.0019493 0.97891 0.9112 4.2961e-006 1.7186e-005 0.15756 0.56094 0.66172 0.0016715 0.62403 0.37649 0.0022416 0.41942 1.2819 1.2768 16.0034 144.93 0.00051912 -83.6026 0.10495
6.209 0.9881 5.483e-005 3.8183 0.011959 8.1026e-005 0.0011644 0.23319 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.3809 0.47704 0.14542 0.017654 11.3143 0.10986 0.00014061 0.78028 0.0084625 0.0093977 0.0019433 0.97902 0.91539 4.2819e-006 1.7129e-005 0.15757 0.56225 0.66331 0.0016688 0.626 0.3767 0.002238 0.41941 1.2843 1.2792 16.0035 144.93 0.00051735 -83.6212 0.10595
6.21 0.9881 5.483e-005 3.8183 0.011959 8.1039e-005 0.0011645 0.23319 0.00065931 0.23384 0.21577 0 0.032285 0.0389 0 1.381 0.47708 0.14543 0.017655 11.3166 0.10987 0.00014063 0.78027 0.008463 0.0093983 0.0019377 0.97913 0.91936 4.2681e-006 1.7074e-005 0.15757 0.56355 0.66489 0.0016661 0.62796 0.3769 0.0022345 0.41941 1.2866 1.2815 16.0036 144.93 0.00051558 -83.6394 0.10695
6.211 0.9881 5.483e-005 3.8183 0.011958 8.1052e-005 0.0011645 0.23319 0.00065931 0.23385 0.21578 0 0.032285 0.0389 0 1.3811 0.47713 0.14545 0.017656 11.3189 0.10988 0.00014064 0.78026 0.0084635 0.0093988 0.0019321 0.97923 0.92312 4.2546e-006 1.7021e-005 0.15758 0.56485 0.66645 0.0016636 0.62991 0.3771 0.002231 0.4194 1.289 1.2839 16.0037 144.93 0.00051382 -83.6572 0.10795
6.212 0.9881 5.483e-005 3.8183 0.011958 8.1065e-005 0.0011645 0.23319 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3812 0.47717 0.14546 0.017658 11.3213 0.10988 0.00014065 0.78026 0.008464 0.0093994 0.0019265 0.97933 0.92668 4.2416e-006 1.6968e-005 0.15758 0.56614 0.66801 0.001661 0.63186 0.37731 0.0022277 0.4194 1.2913 1.2863 16.0038 144.93 0.00051208 -83.6745 0.10895
6.213 0.9881 5.483e-005 3.8183 0.011958 8.1078e-005 0.0011645 0.23319 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3813 0.47722 0.14548 0.017659 11.3236 0.10989 0.00014066 0.78025 0.0084646 0.0094 0.0019209 0.97942 0.93005 4.2288e-006 1.6917e-005 0.15758 0.56743 0.66955 0.0016585 0.6338 0.37751 0.0022244 0.41939 1.2937 1.2886 16.0039 144.93 0.00051034 -83.6916 0.10995
6.214 0.9881 5.483e-005 3.8183 0.011958 8.1091e-005 0.0011645 0.23319 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3814 0.47727 0.14549 0.01766 11.3259 0.1099 0.00014067 0.78024 0.0084651 0.0094005 0.0019154 0.97952 0.93324 4.2164e-006 1.6867e-005 0.15759 0.56872 0.67107 0.0016561 0.63574 0.37772 0.0022212 0.41939 1.296 1.291 16.004 144.93 0.00050861 -83.7083 0.11095
6.215 0.9881 5.483e-005 3.8183 0.011958 8.1104e-005 0.0011645 0.23319 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3815 0.47731 0.14551 0.017662 11.3282 0.10991 0.00014069 0.78023 0.0084656 0.0094011 0.0019102 0.9796 0.93626 4.2042e-006 1.6818e-005 0.15759 0.57001 0.67258 0.0016537 0.63766 0.37792 0.002218 0.41938 1.2983 1.2933 16.0041 144.93 0.00050689 -83.7247 0.11195
6.216 0.9881 5.483e-005 3.8183 0.011958 8.1116e-005 0.0011645 0.23319 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3816 0.47736 0.14552 0.017663 11.3306 0.10992 0.0001407 0.78022 0.0084661 0.0094016 0.0019053 0.97969 0.93911 4.1922e-006 1.677e-005 0.1576 0.57128 0.67408 0.0016514 0.63958 0.37812 0.002215 0.41938 1.3007 1.2957 16.0042 144.93 0.00050518 -83.7408 0.11295
6.217 0.9881 5.483e-005 3.8183 0.011958 8.1129e-005 0.0011645 0.2332 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3817 0.4774 0.14554 0.017664 11.3329 0.10992 0.00014071 0.78022 0.0084666 0.0094022 0.0019005 0.97977 0.94182 4.1804e-006 1.6723e-005 0.1576 0.57256 0.67557 0.0016491 0.64149 0.37833 0.0022119 0.41937 1.303 1.298 16.0043 144.93 0.00050348 -83.7566 0.11395
6.218 0.9881 5.483e-005 3.8183 0.011958 8.1142e-005 0.0011645 0.2332 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3818 0.47745 0.14555 0.017666 11.3352 0.10993 0.00014072 0.78021 0.0084672 0.0094028 0.0018957 0.97985 0.94438 4.1689e-006 1.6677e-005 0.1576 0.57383 0.67704 0.0016469 0.6434 0.37853 0.002209 0.41937 1.3053 1.3003 16.0044 144.93 0.00050179 -83.7722 0.11495
6.219 0.9881 5.483e-005 3.8183 0.011958 8.1155e-005 0.0011645 0.2332 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3819 0.4775 0.14557 0.017667 11.3376 0.10994 0.00014073 0.7802 0.0084677 0.0094033 0.0018908 0.97992 0.9468 4.1575e-006 1.6632e-005 0.15761 0.5751 0.6785 0.0016446 0.64529 0.37873 0.0022061 0.41936 1.3076 1.3027 16.0045 144.9301 0.00050011 -83.7876 0.11595
6.22 0.9881 5.4829e-005 3.8183 0.011958 8.1168e-005 0.0011645 0.2332 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.382 0.47754 0.14558 0.017668 11.3399 0.10995 0.00014075 0.78019 0.0084682 0.0094039 0.0018857 0.98 0.94909 4.1464e-006 1.6587e-005 0.15761 0.57636 0.67995 0.0016425 0.64718 0.37894 0.0022032 0.41936 1.3099 1.305 16.0046 144.9301 0.00049844 -83.8028 0.11695
6.221 0.9881 5.4829e-005 3.8183 0.011958 8.1181e-005 0.0011645 0.2332 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3821 0.47759 0.1456 0.01767 11.3422 0.10996 0.00014076 0.78018 0.0084687 0.0094044 0.0018809 0.98007 0.95126 4.1355e-006 1.6543e-005 0.15762 0.57762 0.68139 0.0016403 0.64907 0.37914 0.0022004 0.41936 1.3122 1.3073 16.0047 144.9301 0.00049678 -83.8177 0.11795
6.222 0.9881 5.4829e-005 3.8183 0.011958 8.1194e-005 0.0011645 0.2332 0.00065931 0.23385 0.21578 0 0.032284 0.0389 0 1.3821 0.47763 0.14561 0.017671 11.3446 0.10997 0.00014077 0.78018 0.0084692 0.009405 0.0018763 0.98014 0.95332 4.1247e-006 1.65e-005 0.15762 0.57888 0.68281 0.0016382 0.65094 0.37935 0.0021976 0.41935 1.3146 1.3097 16.0047 144.9301 0.00049513 -83.8325 0.11895
6.223 0.9881 5.4829e-005 3.8183 0.011958 8.1207e-005 0.0011645 0.2332 0.00065931 0.23386 0.21578 0 0.032284 0.0389 0 1.3822 0.47768 0.14563 0.017672 11.3469 0.10997 0.00014078 0.78017 0.0084698 0.0094055 0.001872 0.98021 0.95526 4.114e-006 1.6457e-005 0.15762 0.58013 0.68422 0.0016361 0.65281 0.37955 0.0021948 0.41935 1.3169 1.312 16.0048 144.9301 0.00049348 -83.8471 0.11995
6.224 0.9881 5.4829e-005 3.8183 0.011958 8.122e-005 0.0011645 0.2332 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3823 0.47773 0.14564 0.017674 11.3492 0.10998 0.00014079 0.78016 0.0084703 0.0094061 0.0018678 0.98028 0.95709 4.1035e-006 1.6416e-005 0.15763 0.58138 0.68562 0.001634 0.65467 0.37975 0.0021921 0.41935 1.3192 1.3143 16.0049 144.9301 0.00049185 -83.8615 0.12095
6.225 0.9881 5.4829e-005 3.8183 0.011958 8.1233e-005 0.0011645 0.2332 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3824 0.47777 0.14566 0.017675 11.3516 0.10999 0.00014081 0.78015 0.0084708 0.0094067 0.0018634 0.98035 0.95883 4.0932e-006 1.6374e-005 0.15763 0.58263 0.68701 0.001632 0.65652 0.37996 0.0021895 0.41934 1.3214 1.3166 16.005 144.9301 0.00049022 -83.8757 0.12195
6.226 0.9881 5.4829e-005 3.8183 0.011958 8.1245e-005 0.0011645 0.2332 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3825 0.47782 0.14567 0.017676 11.3539 0.11 0.00014082 0.78014 0.0084713 0.0094072 0.0018589 0.98041 0.96048 4.083e-006 1.6333e-005 0.15764 0.58387 0.68839 0.00163 0.65837 0.38016 0.0021868 0.41934 1.3237 1.3189 16.0051 144.9301 0.0004886 -83.8898 0.12295
6.227 0.9881 5.4829e-005 3.8183 0.011958 8.1258e-005 0.0011645 0.2332 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3826 0.47787 0.14569 0.017678 11.3563 0.11001 0.00014083 0.78013 0.0084718 0.0094078 0.0018543 0.98048 0.96203 4.073e-006 1.6293e-005 0.15764 0.58511 0.68975 0.001628 0.66021 0.38037 0.0021842 0.41934 1.326 1.3212 16.0052 144.9301 0.000487 -83.9037 0.12395
6.228 0.9881 5.4829e-005 3.8183 0.011958 8.1271e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3827 0.47791 0.1457 0.017679 11.3586 0.11001 0.00014084 0.78013 0.0084724 0.0094083 0.0018499 0.98054 0.9635 4.0631e-006 1.6254e-005 0.15764 0.58634 0.69111 0.0016261 0.66204 0.38057 0.0021817 0.41933 1.3283 1.3235 16.0053 144.9301 0.0004854 -83.9175 0.12495
6.229 0.9881 5.4829e-005 3.8183 0.011958 8.1284e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3828 0.47796 0.14572 0.01768 11.3609 0.11002 0.00014085 0.78012 0.0084729 0.0094089 0.0018457 0.9806 0.96489 4.0533e-006 1.6214e-005 0.15765 0.58757 0.69245 0.0016241 0.66386 0.38077 0.0021791 0.41933 1.3306 1.3258 16.0053 144.9301 0.00048381 -83.9311 0.12595
6.23 0.9881 5.4829e-005 3.8183 0.011958 8.1297e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3829 0.478 0.14573 0.017682 11.3633 0.11003 0.00014086 0.78011 0.0084734 0.0094095 0.0018418 0.98066 0.96621 4.0436e-006 1.6176e-005 0.15765 0.5888 0.69378 0.0016222 0.66568 0.38098 0.0021766 0.41933 1.3329 1.3281 16.0054 144.9301 0.00048223 -83.9446 0.12695
6.231 0.9881 5.4829e-005 3.8183 0.011958 8.131e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.383 0.47805 0.14575 0.017683 11.3656 0.11004 0.00014088 0.7801 0.0084739 0.00941 0.0018379 0.98073 0.96745 4.0341e-006 1.6138e-005 0.15766 0.59002 0.6951 0.0016203 0.66748 0.38118 0.0021741 0.41933 1.3351 1.3304 16.0055 144.9301 0.00048065 -83.9579 0.12795
6.232 0.9881 5.4829e-005 3.8183 0.011958 8.1323e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3831 0.4781 0.14576 0.017684 11.3679 0.11005 0.00014089 0.78009 0.0084744 0.0094106 0.0018339 0.98078 0.96863 4.0247e-006 1.61e-005 0.15766 0.59124 0.69641 0.0016184 0.66929 0.38139 0.0021717 0.41933 1.3374 1.3327 16.0056 144.9301 0.00047909 -83.9712 0.12895
6.233 0.9881 5.4828e-005 3.8183 0.011958 8.1336e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3832 0.47814 0.14577 0.017686 11.3703 0.11006 0.0001409 0.78009 0.008475 0.0094111 0.0018298 0.98084 0.96974 4.0153e-006 1.6063e-005 0.15766 0.59245 0.69771 0.0016166 0.67108 0.38159 0.0021692 0.41932 1.3397 1.335 16.0057 144.9302 0.00047753 -83.9843 0.12995
6.234 0.9881 5.4828e-005 3.8183 0.011958 8.1349e-005 0.0011645 0.23321 0.00065931 0.23386 0.21579 0 0.032284 0.0389 0 1.3833 0.47819 0.14579 0.017687 11.3726 0.11006 0.00014091 0.78008 0.0084755 0.0094117 0.0018257 0.9809 0.97079 4.0061e-006 1.6026e-005 0.15767 0.59366 0.699 0.0016147 0.67287 0.38179 0.0021668 0.41932 1.3419 1.3372 16.0058 144.9302 0.00047598 -83.9972 0.13095
6.235 0.9881 5.4828e-005 3.8183 0.011958 8.1362e-005 0.0011645 0.23321 0.00065931 0.23387 0.21579 0 0.032283 0.0389 0 1.3833 0.47823 0.1458 0.017688 11.375 0.11007 0.00014092 0.78007 0.008476 0.0094123 0.0018218 0.98096 0.97179 3.997e-006 1.5989e-005 0.15767 0.59487 0.70028 0.0016129 0.67464 0.382 0.0021645 0.41932 1.3442 1.3395 16.0058 144.9302 0.00047445 -84.0101 0.13195
6.236 0.9881 5.4828e-005 3.8183 0.011958 8.1375e-005 0.0011645 0.23321 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3834 0.47828 0.14582 0.01769 11.3773 0.11008 0.00014094 0.78006 0.0084765 0.0094128 0.001818 0.98102 0.97273 3.988e-006 1.5953e-005 0.15768 0.59608 0.70155 0.0016111 0.67642 0.3822 0.0021621 0.41932 1.3464 1.3418 16.0059 144.9302 0.00047292 -84.0228 0.13295
6.237 0.9881 5.4828e-005 3.8183 0.011958 8.1387e-005 0.0011646 0.23321 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3835 0.47833 0.14583 0.017691 11.3796 0.11009 0.00014095 0.78005 0.008477 0.0094134 0.0018142 0.98107 0.97362 3.9791e-006 1.5918e-005 0.15768 0.59728 0.70281 0.0016094 0.67818 0.38241 0.0021598 0.41932 1.3487 1.344 16.006 144.9302 0.00047139 -84.0354 0.13395
6.238 0.9881 5.4828e-005 3.8183 0.011958 8.14e-005 0.0011646 0.23321 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3836 0.47837 0.14585 0.017692 11.382 0.1101 0.00014096 0.78004 0.0084776 0.0094139 0.0018105 0.98113 0.97446 3.9703e-006 1.5882e-005 0.15768 0.59847 0.70406 0.0016076 0.67993 0.38261 0.0021575 0.41932 1.3509 1.3463 16.0061 144.9302 0.00046988 -84.0479 0.13495
6.239 0.9881 5.4828e-005 3.8183 0.011958 8.1413e-005 0.0011646 0.23321 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3837 0.47842 0.14586 0.017694 11.3843 0.1101 0.00014097 0.78004 0.0084781 0.0094145 0.0018068 0.98118 0.97526 3.9616e-006 1.5848e-005 0.15769 0.59967 0.70529 0.0016059 0.68168 0.38281 0.0021552 0.41932 1.3532 1.3485 16.0062 144.9302 0.00046837 -84.0603 0.13595
6.24 0.9881 5.4828e-005 3.8183 0.011958 8.1426e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3838 0.47846 0.14588 0.017695 11.3867 0.11011 0.00014098 0.78003 0.0084786 0.009415 0.0018032 0.98123 0.97601 3.953e-006 1.5813e-005 0.15769 0.60086 0.70652 0.0016041 0.68342 0.38302 0.002153 0.41931 1.3554 1.3508 16.0062 144.9302 0.00046687 -84.0726 0.13695
6.241 0.9881 5.4828e-005 3.8183 0.011958 8.1439e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3839 0.47851 0.14589 0.017696 11.389 0.11012 0.000141 0.78002 0.0084791 0.0094156 0.0017997 0.98129 0.97673 3.9445e-006 1.5779e-005 0.1577 0.60204 0.70774 0.0016024 0.68516 0.38322 0.0021507 0.41931 1.3576 1.353 16.0063 144.9302 0.00046539 -84.0848 0.13795
6.242 0.9881 5.4828e-005 3.8183 0.011958 8.1452e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.384 0.47856 0.14591 0.017698 11.3913 0.11013 0.00014101 0.78001 0.0084796 0.0094162 0.0017961 0.98134 0.9774 3.9361e-006 1.5746e-005 0.1577 0.60322 0.70895 0.0016007 0.68688 0.38343 0.0021485 0.41931 1.3599 1.3553 16.0064 144.9302 0.0004639 -84.0968 0.13895
6.243 0.9881 5.4828e-005 3.8183 0.011958 8.1465e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3841 0.4786 0.14592 0.017699 11.3937 0.11014 0.00014102 0.78 0.0084801 0.0094167 0.0017925 0.98139 0.97804 3.9278e-006 1.5712e-005 0.15771 0.6044 0.71015 0.0015991 0.6886 0.38363 0.0021463 0.41931 1.3621 1.3575 16.0065 144.9302 0.00046243 -84.1088 0.13995
6.244 0.9881 5.4828e-005 3.8183 0.011958 8.1478e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3842 0.47865 0.14594 0.0177 11.396 0.11014 0.00014103 0.78 0.0084807 0.0094173 0.001789 0.98144 0.97864 3.9196e-006 1.5679e-005 0.15771 0.60558 0.71134 0.0015974 0.69031 0.38384 0.0021441 0.41931 1.3643 1.3598 16.0066 144.9302 0.00046096 -84.1207 0.14095
6.245 0.9881 5.4828e-005 3.8183 0.011958 8.1491e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3843 0.47869 0.14595 0.017702 11.3984 0.11015 0.00014104 0.77999 0.0084812 0.0094178 0.0017854 0.98149 0.97921 3.9114e-006 1.5647e-005 0.15771 0.60675 0.71252 0.0015957 0.69202 0.38404 0.002142 0.41931 1.3665 1.362 16.0066 144.9303 0.00045951 -84.1324 0.14195
6.246 0.9881 5.4827e-005 3.8183 0.011958 8.1504e-005 0.0011646 0.23322 0.00065931 0.23387 0.2158 0 0.032283 0.0389 0 1.3844 0.47874 0.14597 0.017703 11.4007 0.11016 0.00014105 0.77998 0.0084817 0.0094184 0.0017819 0.98154 0.97975 3.9034e-006 1.5614e-005 0.15772 0.60792 0.71369 0.0015941 0.69372 0.38424 0.0021399 0.41931 1.3687 1.3642 16.0067 144.9303 0.00045806 -84.1441 0.14295
6.247 0.9881 5.4827e-005 3.8183 0.011958 8.1517e-005 0.0011646 0.23322 0.00065931 0.23388 0.2158 0 0.032283 0.0389 0 1.3845 0.47879 0.14598 0.017704 11.403 0.11017 0.00014107 0.77997 0.0084822 0.0094189 0.0017785 0.98159 0.98026 3.8954e-006 1.5582e-005 0.15772 0.60908 0.71485 0.0015925 0.6954 0.38445 0.0021378 0.41931 1.3709 1.3664 16.0068 144.9303 0.00045661 -84.1557 0.14395
6.248 0.9881 5.4827e-005 3.8183 0.011958 8.1529e-005 0.0011646 0.23322 0.00065931 0.23388 0.2158 0 0.032283 0.0389 0 1.3845 0.47883 0.146 0.017706 11.4054 0.11018 0.00014108 0.77996 0.0084827 0.0094195 0.001775 0.98164 0.98075 3.8875e-006 1.5551e-005 0.15773 0.61024 0.71601 0.0015909 0.69709 0.38465 0.0021357 0.41931 1.3731 1.3686 16.0069 144.9303 0.00045518 -84.1671 0.14495
6.249 0.9881 5.4827e-005 3.8183 0.011958 8.1542e-005 0.0011646 0.23322 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3846 0.47888 0.14601 0.017707 11.4077 0.11019 0.00014109 0.77996 0.0084833 0.0094201 0.0017717 0.98169 0.9812 3.8797e-006 1.552e-005 0.15773 0.6114 0.71715 0.0015893 0.69876 0.38486 0.0021336 0.41931 1.3753 1.3709 16.0069 144.9303 0.00045375 -84.1785 0.14595
6.25 0.9881 5.4827e-005 3.8183 0.011958 8.1555e-005 0.0011646 0.23322 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3847 0.47893 0.14603 0.017708 11.4101 0.11019 0.0001411 0.77995 0.0084838 0.0094206 0.0017684 0.98174 0.98164 3.8719e-006 1.5489e-005 0.15773 0.61255 0.71829 0.0015878 0.70043 0.38506 0.0021316 0.41931 1.3775 1.3731 16.007 144.9303 0.00045233 -84.1898 0.14695
6.251 0.9881 5.4827e-005 3.8183 0.011958 8.1568e-005 0.0011646 0.23322 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3848 0.47897 0.14604 0.01771 11.4124 0.1102 0.00014111 0.77994 0.0084843 0.0094212 0.0017651 0.98178 0.98205 3.8643e-006 1.5458e-005 0.15774 0.6137 0.71942 0.0015862 0.70209 0.38526 0.0021295 0.41931 1.3797 1.3753 16.0071 144.9303 0.00045092 -84.201 0.14795
6.252 0.9881 5.4827e-005 3.8183 0.011958 8.1581e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3849 0.47902 0.14606 0.017711 11.4148 0.11021 0.00014113 0.77993 0.0084848 0.0094217 0.0017619 0.98183 0.98244 3.8567e-006 1.5428e-005 0.15774 0.61485 0.72053 0.0015847 0.70374 0.38547 0.0021275 0.41931 1.3819 1.3775 16.0072 144.9303 0.00044952 -84.2121 0.14895
6.253 0.9881 5.4827e-005 3.8183 0.011958 8.1594e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.385 0.47906 0.14607 0.017712 11.4171 0.11022 0.00014114 0.77992 0.0084853 0.0094223 0.0017586 0.98188 0.9828 3.8492e-006 1.5398e-005 0.15775 0.61599 0.72164 0.0015831 0.70538 0.38567 0.0021255 0.41931 1.3841 1.3797 16.0072 144.9303 0.00044812 -84.2231 0.14995
6.254 0.9881 5.4827e-005 3.8183 0.011958 8.1607e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3851 0.47911 0.14609 0.017714 11.4195 0.11023 0.00014115 0.77992 0.0084858 0.0094228 0.0017554 0.98192 0.98315 3.8418e-006 1.5368e-005 0.15775 0.61713 0.72275 0.0015816 0.70702 0.38588 0.0021235 0.41932 1.3863 1.3819 16.0073 144.9303 0.00044673 -84.234 0.15095
6.255 0.9881 5.4827e-005 3.8183 0.011958 8.162e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3852 0.47916 0.1461 0.017715 11.4218 0.11023 0.00014116 0.77991 0.0084864 0.0094234 0.0017523 0.98197 0.98348 3.8344e-006 1.5338e-005 0.15775 0.61827 0.72384 0.0015801 0.70865 0.38608 0.0021216 0.41932 1.3884 1.384 16.0074 144.9304 0.00044535 -84.2448 0.15195
6.256 0.9881 5.4827e-005 3.8183 0.011958 8.1633e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3853 0.4792 0.14612 0.017716 11.4241 0.11024 0.00014117 0.7799 0.0084869 0.009424 0.0017491 0.98201 0.98379 3.8271e-006 1.5309e-005 0.15776 0.6194 0.72492 0.0015787 0.71027 0.38629 0.0021196 0.41932 1.3906 1.3862 16.0074 144.9304 0.00044398 -84.2555 0.15295
6.257 0.9881 5.4827e-005 3.8183 0.011958 8.1646e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3854 0.47925 0.14613 0.017718 11.4265 0.11025 0.00014119 0.77989 0.0084874 0.0094245 0.001746 0.98206 0.98409 3.8199e-006 1.5281e-005 0.15776 0.62053 0.726 0.0015772 0.71189 0.38649 0.0021177 0.41932 1.3928 1.3884 16.0075 144.9304 0.00044261 -84.2662 0.15395
6.258 0.9881 5.4827e-005 3.8183 0.011958 8.1659e-005 0.0011646 0.23323 0.00065931 0.23388 0.21581 0 0.032283 0.0389 0 1.3855 0.47929 0.14615 0.017719 11.4288 0.11026 0.0001412 0.77988 0.0084879 0.0094251 0.001743 0.9821 0.98437 3.8128e-006 1.5252e-005 0.15777 0.62166 0.72707 0.0015757 0.71349 0.38669 0.0021158 0.41932 1.3949 1.3906 16.0076 144.9304 0.00044125 -84.2767 0.15495
6.259 0.9881 5.4826e-005 3.8183 0.011958 8.1671e-005 0.0011646 0.23323 0.00065931 0.23389 0.21581 0 0.032283 0.0389 0 1.3856 0.47934 0.14616 0.01772 11.4312 0.11027 0.00014121 0.77987 0.0084884 0.0094256 0.00174 0.98214 0.98464 3.8057e-006 1.5224e-005 0.15777 0.62278 0.72813 0.0015743 0.71509 0.3869 0.0021139 0.41932 1.3971 1.3928 16.0077 144.9304 0.0004399 -84.2872 0.15595
6.26 0.9881 5.4826e-005 3.8183 0.011958 8.1684e-005 0.0011646 0.23323 0.00065931 0.23389 0.21581 0 0.032282 0.0389 0 1.3857 0.47939 0.14617 0.017722 11.4335 0.11027 0.00014122 0.77987 0.008489 0.0094262 0.001737 0.98219 0.98489 3.7988e-006 1.5196e-005 0.15777 0.6239 0.72918 0.0015729 0.71669 0.3871 0.0021121 0.41932 1.3992 1.3949 16.0077 144.9304 0.00043855 -84.2976 0.15695
6.261 0.9881 5.4826e-005 3.8183 0.011958 8.1697e-005 0.0011646 0.23323 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3857 0.47943 0.14619 0.017723 11.4359 0.11028 0.00014123 0.77986 0.0084895 0.0094267 0.001734 0.98223 0.98513 3.7918e-006 1.5168e-005 0.15778 0.62501 0.73023 0.0015714 0.71827 0.38731 0.0021102 0.41933 1.4014 1.3971 16.0078 144.9304 0.00043721 -84.3079 0.15795
6.262 0.9881 5.4826e-005 3.8183 0.011958 8.171e-005 0.0011646 0.23323 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3858 0.47948 0.1462 0.017724 11.4382 0.11029 0.00014124 0.77985 0.00849 0.0094273 0.0017311 0.98227 0.98535 3.785e-006 1.5141e-005 0.15778 0.62612 0.73127 0.00157 0.71985 0.38751 0.0021084 0.41933 1.4035 1.3992 16.0079 144.9304 0.00043588 -84.3181 0.15895
6.263 0.9881 5.4826e-005 3.8183 0.011958 8.1723e-005 0.0011647 0.23323 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3859 0.47952 0.14622 0.017726 11.4406 0.1103 0.00014126 0.77984 0.0084905 0.0094279 0.0017282 0.98231 0.98557 3.7782e-006 1.5114e-005 0.15779 0.62723 0.7323 0.0015686 0.72142 0.38772 0.0021065 0.41933 1.4057 1.4014 16.0079 144.9304 0.00043456 -84.3283 0.15995
6.264 0.9881 5.4826e-005 3.8183 0.011958 8.1736e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.386 0.47957 0.14623 0.017727 11.4429 0.11031 0.00014127 0.77983 0.008491 0.0094284 0.0017253 0.98235 0.98577 3.7715e-006 1.5087e-005 0.15779 0.62834 0.73332 0.0015673 0.72299 0.38792 0.0021047 0.41933 1.4078 1.4035 16.008 144.9304 0.00043324 -84.3383 0.16095
6.265 0.9881 5.4826e-005 3.8183 0.011958 8.1749e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3861 0.47962 0.14625 0.017728 11.4453 0.11032 0.00014128 0.77983 0.0084915 0.009429 0.0017225 0.98239 0.98597 3.7648e-006 1.506e-005 0.15779 0.62944 0.73433 0.0015659 0.72454 0.38812 0.002103 0.41933 1.4099 1.4057 16.0081 144.9305 0.00043193 -84.3483 0.16195
6.266 0.9881 5.4826e-005 3.8183 0.011958 8.1762e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3862 0.47966 0.14626 0.01773 11.4476 0.11032 0.00014129 0.77982 0.0084921 0.0094295 0.0017197 0.98243 0.98615 3.7582e-006 1.5034e-005 0.1578 0.63054 0.73534 0.0015645 0.72609 0.38833 0.0021012 0.41934 1.412 1.4078 16.0081 144.9305 0.00043062 -84.3582 0.16295
6.267 0.9881 5.4826e-005 3.8183 0.011958 8.1775e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3863 0.47971 0.14628 0.017731 11.45 0.11033 0.0001413 0.77981 0.0084926 0.0094301 0.0017169 0.98247 0.98632 3.7517e-006 1.5008e-005 0.1578 0.63163 0.73634 0.0015632 0.72763 0.38853 0.0020994 0.41934 1.4142 1.41 16.0082 144.9305 0.00042933 -84.368 0.16395
6.268 0.9881 5.4826e-005 3.8183 0.011958 8.1788e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3864 0.47975 0.14629 0.017732 11.4523 0.11034 0.00014132 0.7798 0.0084931 0.0094306 0.0017141 0.98251 0.98649 3.7452e-006 1.4982e-005 0.15781 0.63273 0.73734 0.0015619 0.72917 0.38874 0.0020977 0.41934 1.4163 1.4121 16.0083 144.9305 0.00042804 -84.3778 0.16495
6.269 0.9881 5.4826e-005 3.8183 0.011958 8.18e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3865 0.4798 0.14631 0.017734 11.4547 0.11035 0.00014133 0.77979 0.0084936 0.0094312 0.0017114 0.98255 0.98665 3.7388e-006 1.4956e-005 0.15781 0.63381 0.73832 0.0015605 0.7307 0.38894 0.002096 0.41934 1.4184 1.4142 16.0083 144.9305 0.00042675 -84.3874 0.16595
6.27 0.9881 5.4826e-005 3.8183 0.011958 8.1813e-005 0.0011647 0.23324 0.00065931 0.23389 0.21582 0 0.032282 0.0389 0 1.3866 0.47985 0.14632 0.017735 11.457 0.11036 0.00014134 0.77979 0.0084941 0.0094317 0.0017086 0.98259 0.98679 3.7325e-006 1.4931e-005 0.15781 0.6349 0.7393 0.0015592 0.73222 0.38915 0.0020942 0.41935 1.4205 1.4163 16.0084 144.9305 0.00042548 -84.397 0.16695
6.271 0.9881 5.4826e-005 3.8183 0.011957 8.1826e-005 0.0011647 0.23324 0.00065931 0.2339 0.21582 0 0.032282 0.0389 0 1.3867 0.47989 0.14634 0.017736 11.4594 0.11036 0.00014135 0.77978 0.0084946 0.0094323 0.0017059 0.98263 0.98694 3.7262e-006 1.4906e-005 0.15782 0.63598 0.74027 0.0015579 0.73373 0.38935 0.0020926 0.41935 1.4226 1.4185 16.0085 144.9305 0.00042421 -84.4065 0.16795
6.272 0.9881 5.4825e-005 3.8183 0.011957 8.1839e-005 0.0011647 0.23324 0.00065931 0.2339 0.21582 0 0.032282 0.0389 0 1.3868 0.47994 0.14635 0.017738 11.4617 0.11037 0.00014136 0.77977 0.0084952 0.0094329 0.0017032 0.98267 0.98707 3.72e-006 1.4881e-005 0.15782 0.63706 0.74124 0.0015566 0.73524 0.38955 0.0020909 0.41935 1.4247 1.4206 16.0085 144.9305 0.00042294 -84.4159 0.16895
6.273 0.9881 5.4825e-005 3.8183 0.011957 8.1852e-005 0.0011647 0.23324 0.00065931 0.2339 0.21582 0 0.032282 0.0389 0 1.3868 0.47998 0.14637 0.017739 11.4641 0.11038 0.00014138 0.77976 0.0084957 0.0094334 0.0017005 0.9827 0.9872 3.7138e-006 1.4856e-005 0.15783 0.63813 0.74219 0.0015554 0.73673 0.38976 0.0020892 0.41936 1.4268 1.4227 16.0086 144.9305 0.00042169 -84.4253 0.16995
6.274 0.9881 5.4825e-005 3.8183 0.011957 8.1865e-005 0.0011647 0.23324 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3869 0.48003 0.14638 0.01774 11.4664 0.11039 0.00014139 0.77975 0.0084962 0.009434 0.0016979 0.98274 0.98732 3.7078e-006 1.4832e-005 0.15783 0.63921 0.74314 0.0015541 0.73823 0.38996 0.0020876 0.41936 1.4289 1.4248 16.0087 144.9306 0.00042044 -84.4346 0.17095
6.275 0.9881 5.4825e-005 3.8183 0.011957 8.1878e-005 0.0011647 0.23324 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.387 0.48008 0.1464 0.017742 11.4688 0.1104 0.0001414 0.77974 0.0084967 0.0094345 0.0016953 0.98278 0.98744 3.7017e-006 1.4808e-005 0.15783 0.64027 0.74409 0.0015529 0.73971 0.39017 0.0020859 0.41936 1.431 1.4269 16.0087 144.9306 0.00041919 -84.4438 0.17195
6.276 0.9881 5.4825e-005 3.8183 0.011957 8.1891e-005 0.0011647 0.23324 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3871 0.48012 0.14641 0.017743 11.4711 0.1104 0.00014141 0.77974 0.0084972 0.0094351 0.0016927 0.98281 0.98755 3.6957e-006 1.4784e-005 0.15784 0.64134 0.74503 0.0015516 0.74119 0.39037 0.0020843 0.41936 1.4331 1.429 16.0088 144.9306 0.00041796 -84.4529 0.17295
6.277 0.9881 5.4825e-005 3.8183 0.011957 8.1904e-005 0.0011647 0.23325 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3872 0.48017 0.14643 0.017744 11.4735 0.11041 0.00014142 0.77973 0.0084977 0.0094356 0.0016901 0.98285 0.98765 3.6898e-006 1.476e-005 0.15784 0.6424 0.74596 0.0015504 0.74266 0.39058 0.0020827 0.41937 1.4351 1.4311 16.0088 144.9306 0.00041673 -84.462 0.17395
6.278 0.9881 5.4825e-005 3.8183 0.011957 8.1917e-005 0.0011647 0.23325 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3873 0.48022 0.14644 0.017746 11.4758 0.11042 0.00014143 0.77972 0.0084982 0.0094362 0.0016876 0.98288 0.98775 3.684e-006 1.4736e-005 0.15785 0.64346 0.74688 0.0015492 0.74412 0.39078 0.0020811 0.41937 1.4372 1.4332 16.0089 144.9306 0.0004155 -84.471 0.17495
6.279 0.9881 5.4825e-005 3.8183 0.011957 8.193e-005 0.0011647 0.23325 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3874 0.48026 0.14646 0.017747 11.4782 0.11043 0.00014145 0.77971 0.0084988 0.0094367 0.0016852 0.98292 0.98785 3.6781e-006 1.4713e-005 0.15785 0.64452 0.7478 0.001548 0.74558 0.39098 0.0020795 0.41938 1.4393 1.4353 16.009 144.9306 0.00041428 -84.4799 0.17595
6.28 0.9881 5.4825e-005 3.8183 0.011957 8.1942e-005 0.0011647 0.23325 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3875 0.48031 0.14647 0.017748 11.4806 0.11044 0.00014146 0.7797 0.0084993 0.0094373 0.0016827 0.98295 0.98794 3.6724e-006 1.469e-005 0.15785 0.64557 0.74871 0.0015468 0.74703 0.39119 0.0020779 0.41938 1.4414 1.4373 16.009 144.9306 0.00041307 -84.4887 0.17695
6.281 0.9881 5.4825e-005 3.8183 0.011957 8.1955e-005 0.0011647 0.23325 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3876 0.48035 0.14649 0.01775 11.4829 0.11045 0.00014147 0.7797 0.0084998 0.0094378 0.0016803 0.98299 0.98803 3.6667e-006 1.4667e-005 0.15786 0.64662 0.74962 0.0015456 0.74847 0.39139 0.0020764 0.41938 1.4434 1.4394 16.0091 144.9306 0.00041187 -84.4975 0.17795
6.282 0.9881 5.4825e-005 3.8183 0.011957 8.1968e-005 0.0011647 0.23325 0.00065931 0.2339 0.21583 0 0.032282 0.0389 0 1.3877 0.4804 0.1465 0.017751 11.4853 0.11045 0.00014148 0.77969 0.0085003 0.0094384 0.0016779 0.98302 0.98811 3.661e-006 1.4645e-005 0.15786 0.64766 0.75052 0.0015444 0.7499 0.3916 0.0020749 0.41939 1.4455 1.4415 16.0092 144.9306 0.00041067 -84.5062 0.17895
6.283 0.9881 5.4825e-005 3.8183 0.011957 8.1981e-005 0.0011647 0.23325 0.00065931 0.23391 0.21583 0 0.032282 0.0389 0 1.3878 0.48045 0.14651 0.017752 11.4876 0.11046 0.00014149 0.77968 0.0085008 0.009439 0.0016755 0.98306 0.98819 3.6554e-006 1.4622e-005 0.15787 0.64871 0.75141 0.0015432 0.75133 0.3918 0.0020733 0.41939 1.4475 1.4435 16.0092 144.9307 0.00040948 -84.5149 0.17995
6.284 0.9881 5.4825e-005 3.8183 0.011957 8.1994e-005 0.0011647 0.23325 0.00065931 0.23391 0.21583 0 0.032281 0.0389 0 1.3879 0.48049 0.14653 0.017754 11.49 0.11047 0.00014151 0.77967 0.0085013 0.0094395 0.0016732 0.98309 0.98827 3.6499e-006 1.46e-005 0.15787 0.64975 0.7523 0.0015421 0.75275 0.39201 0.0020718 0.4194 1.4496 1.4456 16.0093 144.9307 0.00040829 -84.5235 0.18095
6.285 0.9881 5.4824e-005 3.8183 0.011957 8.2007e-005 0.0011647 0.23325 0.00065931 0.23391 0.21583 0 0.032281 0.0389 0 1.388 0.48054 0.14654 0.017755 11.4923 0.11048 0.00014152 0.77966 0.0085019 0.0094401 0.0016708 0.98312 0.98834 3.6444e-006 1.4578e-005 0.15787 0.65078 0.75318 0.0015409 0.75417 0.39221 0.0020703 0.4194 1.4516 1.4477 16.0093 144.9307 0.00040711 -84.532 0.18195
6.286 0.9881 5.4824e-005 3.8183 0.011957 8.202e-005 0.0011647 0.23325 0.00065931 0.23391 0.21583 0 0.032281 0.0389 0 1.388 0.48058 0.14656 0.017756 11.4947 0.11049 0.00014153 0.77966 0.0085024 0.0094406 0.0016685 0.98316 0.98841 3.6389e-006 1.4556e-005 0.15788 0.65181 0.75405 0.0015398 0.75557 0.39241 0.0020688 0.4194 1.4537 1.4497 16.0094 144.9307 0.00040593 -84.5404 0.18295
6.287 0.9881 5.4824e-005 3.8183 0.011957 8.2033e-005 0.0011647 0.23325 0.00065931 0.23391 0.21583 0 0.032281 0.0389 0 1.3881 0.48063 0.14657 0.017758 11.497 0.11049 0.00014154 0.77965 0.0085029 0.0094412 0.0016661 0.98319 0.98847 3.6336e-006 1.4535e-005 0.15788 0.65284 0.75492 0.0015387 0.75697 0.39262 0.0020674 0.41941 1.4557 1.4518 16.0094 144.9307 0.00040477 -84.5488 0.18395
6.288 0.9881 5.4824e-005 3.8183 0.011957 8.2046e-005 0.0011647 0.23325 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3882 0.48068 0.14659 0.017759 11.4994 0.1105 0.00014155 0.77964 0.0085034 0.0094417 0.0016638 0.98322 0.98854 3.6282e-006 1.4513e-005 0.15789 0.65387 0.75578 0.0015375 0.75837 0.39282 0.0020659 0.41941 1.4577 1.4538 16.0095 144.9307 0.0004036 -84.5571 0.18495
6.289 0.9881 5.4824e-005 3.8183 0.011957 8.2059e-005 0.0011647 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3883 0.48072 0.1466 0.01776 11.5018 0.11051 0.00014156 0.77963 0.0085039 0.0094423 0.0016615 0.98325 0.9886 3.6229e-006 1.4492e-005 0.15789 0.65489 0.75664 0.0015364 0.75975 0.39303 0.0020644 0.41942 1.4597 1.4558 16.0096 144.9307 0.00040245 -84.5653 0.18595
6.29 0.9881 5.4824e-005 3.8183 0.011957 8.2072e-005 0.0011648 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3884 0.48077 0.14662 0.017762 11.5041 0.11052 0.00014158 0.77962 0.0085044 0.0094428 0.0016592 0.98328 0.98866 3.6177e-006 1.4471e-005 0.1579 0.65592 0.75749 0.0015353 0.76113 0.39323 0.002063 0.41942 1.4618 1.4579 16.0096 144.9307 0.0004013 -84.5735 0.18695
6.291 0.9881 5.4824e-005 3.8183 0.011957 8.2084e-005 0.0011648 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3885 0.48081 0.14663 0.017763 11.5065 0.11053 0.00014159 0.77962 0.0085049 0.0094434 0.0016569 0.98331 0.98871 3.6125e-006 1.4451e-005 0.1579 0.65693 0.75833 0.0015342 0.76251 0.39343 0.0020616 0.41943 1.4638 1.4599 16.0097 144.9308 0.00040015 -84.5816 0.18795
6.292 0.9881 5.4824e-005 3.8183 0.011957 8.2097e-005 0.0011648 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3886 0.48086 0.14665 0.017764 11.5088 0.11053 0.0001416 0.77961 0.0085055 0.0094439 0.0016547 0.98335 0.98877 3.6074e-006 1.443e-005 0.1579 0.65795 0.75917 0.0015332 0.76387 0.39364 0.0020602 0.41943 1.4658 1.4619 16.0097 144.9308 0.00039901 -84.5897 0.18895
6.293 0.9881 5.4824e-005 3.8183 0.011957 8.211e-005 0.0011648 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3887 0.48091 0.14666 0.017766 11.5112 0.11054 0.00014161 0.7796 0.008506 0.0094445 0.0016525 0.98338 0.98882 3.6023e-006 1.441e-005 0.15791 0.65896 0.76001 0.0015321 0.76523 0.39384 0.0020588 0.41944 1.4678 1.464 16.0098 144.9308 0.00039788 -84.5977 0.18995
6.294 0.9881 5.4824e-005 3.8183 0.011957 8.2123e-005 0.0011648 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3888 0.48095 0.14668 0.017767 11.5135 0.11055 0.00014162 0.77959 0.0085065 0.009445 0.0016504 0.98341 0.98887 3.5972e-006 1.4389e-005 0.15791 0.65997 0.76084 0.001531 0.76658 0.39405 0.0020574 0.41944 1.4698 1.466 16.0098 144.9308 0.00039675 -84.6056 0.19095
6.295 0.9881 5.4824e-005 3.8183 0.011957 8.2136e-005 0.0011648 0.23326 0.00065931 0.23391 0.21584 0 0.032281 0.0389 0 1.3889 0.481 0.14669 0.017768 11.5159 0.11056 0.00014164 0.77958 0.008507 0.0094456 0.0016483 0.98344 0.98892 3.5922e-006 1.4369e-005 0.15792 0.66097 0.76166 0.00153 0.76793 0.39425 0.002056 0.41945 1.4718 1.468 16.0099 144.9308 0.00039563 -84.6134 0.19195
6.296 0.9881 5.4824e-005 3.8183 0.011957 8.2149e-005 0.0011648 0.23326 0.00065931 0.23392 0.21584 0 0.032281 0.0389 0 1.389 0.48104 0.14671 0.01777 11.5183 0.11057 0.00014165 0.77958 0.0085075 0.0094461 0.0016461 0.98347 0.98896 3.5873e-006 1.435e-005 0.15792 0.66197 0.76248 0.0015289 0.76927 0.39445 0.0020546 0.41945 1.4738 1.47 16.01 144.9308 0.00039452 -84.6212 0.19295
6.297 0.9881 5.4824e-005 3.8183 0.011957 8.2162e-005 0.0011648 0.23326 0.00065931 0.23392 0.21584 0 0.032281 0.0389 0 1.3891 0.48109 0.14672 0.017771 11.5206 0.11057 0.00014166 0.77957 0.008508 0.0094467 0.001644 0.9835 0.98901 3.5824e-006 1.433e-005 0.15792 0.66297 0.76329 0.0015279 0.7706 0.39466 0.0020533 0.41946 1.4758 1.472 16.01 144.9308 0.00039341 -84.629 0.19395
6.298 0.9881 5.4823e-005 3.8183 0.011957 8.2175e-005 0.0011648 0.23326 0.00065931 0.23392 0.21584 0 0.032281 0.0389 0 1.3892 0.48114 0.14674 0.017772 11.523 0.11058 0.00014167 0.77956 0.0085085 0.0094473 0.0016418 0.98352 0.98905 3.5775e-006 1.431e-005 0.15793 0.66397 0.7641 0.0015269 0.77192 0.39486 0.0020519 0.41946 1.4778 1.474 16.0101 144.9308 0.0003923 -84.6367 0.19495
6.299 0.9881 5.4823e-005 3.8183 0.011957 8.2188e-005 0.0011648 0.23326 0.00065931 0.23392 0.21584 0 0.032281 0.0389 0 1.3892 0.48118 0.14675 0.017774 11.5253 0.11059 0.00014168 0.77955 0.0085091 0.0094478 0.0016396 0.98355 0.98909 3.5727e-006 1.4291e-005 0.15793 0.66496 0.7649 0.0015258 0.77324 0.39507 0.0020506 0.41947 1.4798 1.476 16.0101 144.9309 0.0003912 -84.6443 0.19595
6.3 0.9881 5.4823e-005 3.8183 0.011957 8.2201e-005 0.0011648 0.23326 0.00065931 0.23392 0.21584 0 0.032281 0.0389 0 1.3893 0.48123 0.14677 0.017775 11.5277 0.1106 0.00014169 0.77954 0.0085096 0.0094484 0.0016375 0.98358 0.98913 3.5679e-006 1.4272e-005 0.15794 0.66595 0.76569 0.0015248 0.77455 0.39527 0.0020493 0.41947 1.4817 1.478 16.0102 144.9309 0.00039011 -84.6518 0.19695
6.301 0.9881 5.4823e-005 3.8183 0.011957 8.2213e-005 0.0011648 0.23326 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3894 0.48127 0.14678 0.017776 11.5301 0.11061 0.00014171 0.77953 0.0085101 0.0094489 0.0016354 0.98361 0.98917 3.5632e-006 1.4253e-005 0.15794 0.66694 0.76648 0.0015238 0.77586 0.39547 0.002048 0.41948 1.4837 1.48 16.0102 144.9309 0.00038902 -84.6593 0.19795
6.302 0.9881 5.4823e-005 3.8183 0.011957 8.2226e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3895 0.48132 0.1468 0.017778 11.5324 0.11061 0.00014172 0.77953 0.0085106 0.0094495 0.0016334 0.98364 0.98921 3.5585e-006 1.4234e-005 0.15794 0.66792 0.76727 0.0015228 0.77716 0.39568 0.0020467 0.41949 1.4857 1.482 16.0103 144.9309 0.00038794 -84.6668 0.19895
6.303 0.9881 5.4823e-005 3.8183 0.011957 8.2239e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3896 0.48137 0.14681 0.017779 11.5348 0.11062 0.00014173 0.77952 0.0085111 0.00945 0.0016314 0.98367 0.98924 3.5538e-006 1.4216e-005 0.15795 0.6689 0.76805 0.0015219 0.77845 0.39588 0.0020454 0.41949 1.4877 1.4839 16.0103 144.9309 0.00038686 -84.6742 0.19995
6.304 0.9881 5.4823e-005 3.8183 0.011957 8.2252e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3897 0.48141 0.14682 0.01778 11.5372 0.11063 0.00014174 0.77951 0.0085116 0.0094506 0.0016295 0.98369 0.98928 3.5492e-006 1.4197e-005 0.15795 0.66988 0.76883 0.0015209 0.77973 0.39609 0.0020441 0.4195 1.4896 1.4859 16.0104 144.9309 0.00038579 -84.6815 0.20095
6.305 0.9881 5.4823e-005 3.8183 0.011957 8.2265e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3898 0.48146 0.14684 0.017782 11.5395 0.11064 0.00014175 0.7795 0.0085121 0.0094511 0.0016276 0.98372 0.98931 3.5447e-006 1.4179e-005 0.15796 0.67085 0.7696 0.0015199 0.78101 0.39629 0.0020429 0.4195 1.4916 1.4879 16.0104 144.9309 0.00038473 -84.6888 0.20195
6.306 0.9881 5.4823e-005 3.8183 0.011957 8.2278e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3899 0.4815 0.14685 0.017783 11.5419 0.11065 0.00014177 0.77949 0.0085127 0.0094517 0.0016257 0.98375 0.98934 3.5401e-006 1.4161e-005 0.15796 0.67182 0.77036 0.001519 0.78228 0.39649 0.0020416 0.41951 1.4935 1.4898 16.0105 144.9309 0.00038367 -84.696 0.20295
6.307 0.9881 5.4823e-005 3.8183 0.011957 8.2291e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.39 0.48155 0.14687 0.017784 11.5442 0.11066 0.00014178 0.77949 0.0085132 0.0094522 0.0016238 0.98377 0.98937 3.5356e-006 1.4143e-005 0.15796 0.67279 0.77112 0.001518 0.78355 0.3967 0.0020404 0.41952 1.4955 1.4918 16.0105 144.931 0.00038261 -84.7031 0.20395
6.308 0.9881 5.4823e-005 3.8183 0.011957 8.2304e-005 0.0011648 0.23327 0.00065931 0.23392 0.21585 0 0.032281 0.0389 0 1.3901 0.4816 0.14688 0.017786 11.5466 0.11066 0.00014179 0.77948 0.0085137 0.0094528 0.0016219 0.9838 0.9894 3.5312e-006 1.4125e-005 0.15797 0.67376 0.77188 0.0015171 0.78481 0.3969 0.0020391 0.41952 1.4974 1.4938 16.0106 144.931 0.00038156 -84.7103 0.20495
6.309 0.9881 5.4823e-005 3.8183 0.011957 8.2317e-005 0.0011648 0.23327 0.00065931 0.23393 0.21585 0 0.032281 0.0389 0 1.3902 0.48164 0.1469 0.017787 11.549 0.11067 0.0001418 0.77947 0.0085142 0.0094533 0.00162 0.98383 0.98943 3.5268e-006 1.4108e-005 0.15797 0.67472 0.77263 0.0015161 0.78606 0.3971 0.0020379 0.41953 1.4993 1.4957 16.0106 144.931 0.00038052 -84.7173 0.20595
6.31 0.9881 5.4823e-005 3.8183 0.011957 8.233e-005 0.0011648 0.23327 0.00065931 0.23393 0.21585 0 0.03228 0.0389 0 1.3903 0.48169 0.14691 0.017788 11.5513 0.11068 0.00014181 0.77946 0.0085147 0.0094539 0.0016182 0.98385 0.98946 3.5224e-006 1.409e-005 0.15798 0.67568 0.77337 0.0015152 0.78731 0.39731 0.0020367 0.41954 1.5013 1.4977 16.0107 144.931 0.00037948 -84.7243 0.20695
6.311 0.9881 5.4822e-005 3.8183 0.011957 8.2343e-005 0.0011648 0.23327 0.00065931 0.23393 0.21585 0 0.03228 0.0389 0 1.3904 0.48173 0.14693 0.01779 11.5537 0.11069 0.00014182 0.77945 0.0085152 0.0094544 0.0016163 0.98388 0.98949 3.5181e-006 1.4073e-005 0.15798 0.67664 0.77412 0.0015143 0.78855 0.39751 0.0020355 0.41954 1.5032 1.4996 16.0107 144.931 0.00037844 -84.7312 0.20795
6.312 0.9881 5.4822e-005 3.8183 0.011957 8.2355e-005 0.0011648 0.23327 0.00065931 0.23393 0.21585 0 0.03228 0.0389 0 1.3904 0.48178 0.14694 0.017791 11.5561 0.1107 0.00014184 0.77945 0.0085157 0.009455 0.0016145 0.9839 0.98952 3.5138e-006 1.4056e-005 0.15798 0.67759 0.77485 0.0015134 0.78978 0.39771 0.0020343 0.41955 1.5051 1.5015 16.0108 144.931 0.00037742 -84.7381 0.20895
6.313 0.9881 5.4822e-005 3.8183 0.011957 8.2368e-005 0.0011648 0.23327 0.00065931 0.23393 0.21585 0 0.03228 0.0389 0 1.3905 0.48183 0.14696 0.017792 11.5584 0.1107 0.00014185 0.77944 0.0085162 0.0094555 0.0016126 0.98393 0.98954 3.5096e-006 1.4039e-005 0.15799 0.67854 0.77558 0.0015125 0.79101 0.39792 0.0020331 0.41955 1.5071 1.5035 16.0108 144.931 0.00037639 -84.745 0.20995
6.314 0.9881 5.4822e-005 3.8183 0.011957 8.2381e-005 0.0011648 0.23327 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3906 0.48187 0.14697 0.017794 11.5608 0.11071 0.00014186 0.77943 0.0085168 0.0094561 0.0016107 0.98396 0.98957 3.5054e-006 1.4022e-005 0.15799 0.67949 0.77631 0.0015116 0.79223 0.39812 0.0020319 0.41956 1.509 1.5054 16.0109 144.931 0.00037537 -84.7517 0.21095
6.315 0.9881 5.4822e-005 3.8183 0.011957 8.2394e-005 0.0011648 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3907 0.48192 0.14699 0.017795 11.5632 0.11072 0.00014187 0.77942 0.0085173 0.0094566 0.0016089 0.98398 0.98959 3.5012e-006 1.4005e-005 0.158 0.68043 0.77703 0.0015107 0.79344 0.39833 0.0020308 0.41957 1.5109 1.5073 16.0109 144.9311 0.00037436 -84.7585 0.21195
6.316 0.9881 5.4822e-005 3.8183 0.011957 8.2407e-005 0.0011648 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3908 0.48197 0.147 0.017796 11.5655 0.11073 0.00014188 0.77941 0.0085178 0.0094572 0.0016071 0.984 0.98962 3.4971e-006 1.3989e-005 0.158 0.68137 0.77775 0.0015098 0.79465 0.39853 0.0020296 0.41957 1.5128 1.5092 16.011 144.9311 0.00037335 -84.7651 0.21295
6.317 0.9881 5.4822e-005 3.8183 0.011957 8.242e-005 0.0011649 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3909 0.48201 0.14702 0.017798 11.5679 0.11074 0.0001419 0.77941 0.0085183 0.0094577 0.0016053 0.98403 0.98964 3.493e-006 1.3972e-005 0.158 0.68231 0.77847 0.0015089 0.79585 0.39873 0.0020285 0.41958 1.5147 1.5112 16.011 144.9311 0.00037235 -84.7718 0.21395
6.318 0.9881 5.4822e-005 3.8183 0.011957 8.2433e-005 0.0011649 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.391 0.48206 0.14703 0.017799 11.5703 0.11074 0.00014191 0.7794 0.0085188 0.0094583 0.0016035 0.98405 0.98967 3.4889e-006 1.3956e-005 0.15801 0.68325 0.77918 0.0015081 0.79704 0.39894 0.0020274 0.41959 1.5166 1.5131 16.0111 144.9311 0.00037135 -84.7783 0.21495
6.319 0.9881 5.4822e-005 3.8183 0.011957 8.2446e-005 0.0011649 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3911 0.4821 0.14705 0.0178 11.5726 0.11075 0.00014192 0.77939 0.0085193 0.0094588 0.0016017 0.98408 0.98969 3.4849e-006 1.394e-005 0.15801 0.68418 0.77988 0.0015072 0.79823 0.39914 0.0020262 0.4196 1.5185 1.515 16.0111 144.9311 0.00037036 -84.7849 0.21595
6.32 0.9881 5.4822e-005 3.8183 0.011957 8.2459e-005 0.0011649 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3912 0.48215 0.14706 0.017802 11.575 0.11076 0.00014193 0.77938 0.0085198 0.0094594 0.0016 0.9841 0.98971 3.4809e-006 1.3924e-005 0.15802 0.68511 0.78058 0.0015063 0.79942 0.39934 0.0020251 0.4196 1.5204 1.5169 16.0111 144.9311 0.00036937 -84.7913 0.21695
6.321 0.9881 5.4822e-005 3.8183 0.011957 8.2472e-005 0.0011649 0.23328 0.00065931 0.23393 0.21586 0 0.03228 0.0389 0 1.3913 0.4822 0.14708 0.017803 11.5774 0.11077 0.00014194 0.77937 0.0085203 0.0094599 0.0015982 0.98412 0.98973 3.4769e-006 1.3908e-005 0.15802 0.68604 0.78128 0.0015055 0.80059 0.39955 0.002024 0.41961 1.5223 1.5188 16.0112 144.9311 0.00036839 -84.7977 0.21795
6.322 0.9881 5.4822e-005 3.8183 0.011957 8.2484e-005 0.0011649 0.23328 0.00065931 0.23394 0.21586 0 0.03228 0.0389 0 1.3914 0.48224 0.14709 0.017804 11.5797 0.11078 0.00014195 0.77937 0.0085209 0.0094605 0.0015965 0.98415 0.98975 3.473e-006 1.3893e-005 0.15802 0.68697 0.78197 0.0015046 0.80176 0.39975 0.0020229 0.41962 1.5241 1.5207 16.0112 144.9312 0.00036741 -84.8041 0.21895
6.323 0.9881 5.4822e-005 3.8183 0.011957 8.2497e-005 0.0011649 0.23328 0.00065931 0.23394 0.21586 0 0.03228 0.0389 0 1.3915 0.48229 0.14711 0.017806 11.5821 0.11078 0.00014197 0.77936 0.0085214 0.009461 0.0015949 0.98417 0.98977 3.4691e-006 1.3877e-005 0.15803 0.68789 0.78266 0.0015038 0.80293 0.39995 0.0020218 0.41962 1.526 1.5225 16.0113 144.9312 0.00036644 -84.8104 0.21995
6.324 0.9881 5.4821e-005 3.8183 0.011957 8.251e-005 0.0011649 0.23328 0.00065931 0.23394 0.21586 0 0.03228 0.0389 0 1.3915 0.48233 0.14712 0.017807 11.5845 0.11079 0.00014198 0.77935 0.0085219 0.0094616 0.0015933 0.98419 0.98979 3.4653e-006 1.3862e-005 0.15803 0.68881 0.78334 0.001503 0.80408 0.40016 0.0020207 0.41963 1.5279 1.5244 16.0113 144.9312 0.00036547 -84.8167 0.22095
6.325 0.9881 5.4821e-005 3.8183 0.011957 8.2523e-005 0.0011649 0.23328 0.00065931 0.23394 0.21586 0 0.03228 0.0389 0 1.3916 0.48238 0.14713 0.017808 11.5869 0.1108 0.00014199 0.77934 0.0085224 0.0094621 0.0015916 0.98422 0.98981 3.4615e-006 1.3846e-005 0.15804 0.68972 0.78402 0.0015022 0.80523 0.40036 0.0020197 0.41964 1.5298 1.5263 16.0114 144.9312 0.0003645 -84.8229 0.22195
6.326 0.9881 5.4821e-005 3.8183 0.011957 8.2536e-005 0.0011649 0.23328 0.00065931 0.23394 0.21586 0 0.03228 0.0389 0 1.3917 0.48243 0.14715 0.01781 11.5892 0.11081 0.000142 0.77933 0.0085229 0.0094627 0.00159 0.98424 0.98983 3.4577e-006 1.3831e-005 0.15804 0.69064 0.7847 0.0015014 0.80638 0.40056 0.0020186 0.41965 1.5316 1.5282 16.0114 144.9312 0.00036354 -84.8291 0.22295
6.327 0.9881 5.4821e-005 3.8183 0.011957 8.2549e-005 0.0011649 0.23328 0.00065931 0.23394 0.21586 0 0.03228 0.0389 0 1.3918 0.48247 0.14716 0.017811 11.5916 0.11082 0.00014201 0.77933 0.0085234 0.0094632 0.0015885 0.98426 0.98985 3.4539e-006 1.3816e-005 0.15804 0.69155 0.78537 0.0015006 0.80752 0.40077 0.0020176 0.41965 1.5335 1.5301 16.0115 144.9312 0.00036259 -84.8353 0.22395
6.328 0.9881 5.4821e-005 3.8183 0.011957 8.2562e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.3919 0.48252 0.14718 0.017812 11.594 0.11082 0.00014203 0.77932 0.0085239 0.0094638 0.0015869 0.98428 0.98987 3.4502e-006 1.3801e-005 0.15805 0.69245 0.78603 0.0014998 0.80865 0.40097 0.0020165 0.41966 1.5353 1.5319 16.0115 144.9312 0.00036164 -84.8413 0.22495
6.329 0.9881 5.4821e-005 3.8183 0.011957 8.2575e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.392 0.48256 0.14719 0.017814 11.5963 0.11083 0.00014204 0.77931 0.0085244 0.0094643 0.0015853 0.9843 0.98989 3.4465e-006 1.3787e-005 0.15805 0.69336 0.7867 0.001499 0.80978 0.40117 0.0020155 0.41967 1.5372 1.5338 16.0115 144.9313 0.0003607 -84.8474 0.22595
6.33 0.9881 5.4821e-005 3.8183 0.011957 8.2588e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.3921 0.48261 0.14721 0.017815 11.5987 0.11084 0.00014205 0.7793 0.008525 0.0094649 0.0015838 0.98433 0.98991 3.4429e-006 1.3772e-005 0.15806 0.69426 0.78736 0.0014982 0.8109 0.40138 0.0020144 0.41968 1.539 1.5356 16.0116 144.9313 0.00035976 -84.8534 0.22695
6.331 0.9881 5.4821e-005 3.8183 0.011956 8.2601e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.3922 0.48266 0.14722 0.017816 11.6011 0.11085 0.00014206 0.77929 0.0085255 0.0094654 0.0015822 0.98435 0.98992 3.4393e-006 1.3757e-005 0.15806 0.69516 0.78801 0.0014974 0.81201 0.40158 0.0020134 0.41969 1.5409 1.5375 16.0116 144.9313 0.00035882 -84.8593 0.22795
6.332 0.9881 5.4821e-005 3.8183 0.011956 8.2613e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.3923 0.4827 0.14724 0.017818 11.6034 0.11086 0.00014207 0.77929 0.008526 0.009466 0.0015807 0.98437 0.98994 3.4357e-006 1.3743e-005 0.15806 0.69606 0.78866 0.0014967 0.81312 0.40178 0.0020124 0.41969 1.5427 1.5393 16.0117 144.9313 0.00035789 -84.8652 0.22895
6.333 0.9881 5.4821e-005 3.8183 0.011956 8.2626e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.3924 0.48275 0.14725 0.017819 11.6058 0.11086 0.00014208 0.77928 0.0085265 0.0094665 0.0015791 0.98439 0.98996 3.4321e-006 1.3729e-005 0.15807 0.69695 0.78931 0.0014959 0.81423 0.40199 0.0020114 0.4197 1.5445 1.5412 16.0117 144.9313 0.00035696 -84.8711 0.22995
6.334 0.9881 5.4821e-005 3.8183 0.011956 8.2639e-005 0.0011649 0.23329 0.00065931 0.23394 0.21587 0 0.03228 0.0389 0 1.3925 0.48279 0.14727 0.01782 11.6082 0.11087 0.0001421 0.77927 0.008527 0.0094671 0.0015776 0.98441 0.98998 3.4286e-006 1.3715e-005 0.15807 0.69784 0.78995 0.0014951 0.81532 0.40219 0.0020104 0.41971 1.5464 1.543 16.0117 144.9313 0.00035604 -84.8769 0.23095
6.335 0.9881 5.4821e-005 3.8183 0.011956 8.2652e-005 0.0011649 0.23329 0.00065931 0.23395 0.21587 0 0.03228 0.0389 0 1.3926 0.48284 0.14728 0.017822 11.6106 0.11088 0.00014211 0.77926 0.0085275 0.0094676 0.001576 0.98443 0.98999 3.4251e-006 1.3701e-005 0.15808 0.69873 0.79059 0.0014944 0.81642 0.40239 0.0020094 0.41972 1.5482 1.5449 16.0118 144.9313 0.00035512 -84.8827 0.23195
6.336 0.9881 5.4821e-005 3.8183 0.011956 8.2665e-005 0.0011649 0.23329 0.00065931 0.23395 0.21587 0 0.032279 0.0389 0 1.3927 0.48289 0.1473 0.017823 11.6129 0.11089 0.00014212 0.77925 0.008528 0.0094682 0.0015745 0.98445 0.99001 3.4216e-006 1.3687e-005 0.15808 0.69962 0.79123 0.0014936 0.8175 0.4026 0.0020085 0.41973 1.55 1.5467 16.0118 144.9314 0.00035421 -84.8884 0.23295
6.337 0.9881 5.482e-005 3.8183 0.011956 8.2678e-005 0.0011649 0.23329 0.00065931 0.23395 0.21587 0 0.032279 0.0389 0 1.3927 0.48293 0.14731 0.017824 11.6153 0.1109 0.00014213 0.77925 0.0085285 0.0094687 0.001573 0.98447 0.99002 3.4182e-006 1.3673e-005 0.15808 0.7005 0.79186 0.0014929 0.81858 0.4028 0.0020075 0.41973 1.5518 1.5485 16.0119 144.9314 0.0003533 -84.8941 0.23395
6.338 0.9881 5.482e-005 3.8183 0.011956 8.2691e-005 0.0011649 0.23329 0.00065931 0.23395 0.21587 0 0.032279 0.0389 0 1.3928 0.48298 0.14733 0.017826 11.6177 0.11091 0.00014214 0.77924 0.008529 0.0094693 0.0015714 0.98449 0.99004 3.4148e-006 1.3659e-005 0.15809 0.70138 0.79249 0.0014921 0.81965 0.403 0.0020065 0.41974 1.5536 1.5503 16.0119 144.9314 0.0003524 -84.8997 0.23495
6.339 0.9881 5.482e-005 3.8183 0.011956 8.2704e-005 0.0011649 0.23329 0.00065931 0.23395 0.21587 0 0.032279 0.0389 0 1.3929 0.48302 0.14734 0.017827 11.6201 0.11091 0.00014215 0.77923 0.0085296 0.0094698 0.0015699 0.98451 0.99005 3.4114e-006 1.3646e-005 0.15809 0.70226 0.79311 0.0014914 0.82072 0.4032 0.0020056 0.41975 1.5554 1.5522 16.0119 144.9314 0.0003515 -84.9053 0.23595
6.34 0.9881 5.482e-005 3.8183 0.011956 8.2717e-005 0.0011649 0.23329 0.00065931 0.23395 0.21587 0 0.032279 0.0389 0 1.393 0.48307 0.14736 0.017828 11.6224 0.11092 0.00014217 0.77922 0.0085301 0.0094704 0.0015684 0.98453 0.99007 3.4081e-006 1.3633e-005 0.1581 0.70313 0.79373 0.0014907 0.82178 0.40341 0.0020046 0.41976 1.5572 1.554 16.012 144.9314 0.00035061 -84.9108 0.23695
6.341 0.9881 5.482e-005 3.8183 0.011956 8.273e-005 0.0011649 0.2333 0.00065931 0.23395 0.21587 0 0.032279 0.0389 0 1.3931 0.48312 0.14737 0.017829 11.6248 0.11093 0.00014218 0.77921 0.0085306 0.0094709 0.001567 0.98455 0.99008 3.4047e-006 1.3619e-005 0.1581 0.704 0.79435 0.00149 0.82284 0.40361 0.0020037 0.41977 1.559 1.5558 16.012 144.9314 0.00034972 -84.9163 0.23795
6.342 0.9881 5.482e-005 3.8183 0.011956 8.2743e-005 0.0011649 0.2333 0.00065931 0.23395 0.21588 0 0.032279 0.0389 0 1.3932 0.48316 0.14739 0.017831 11.6272 0.11094 0.00014219 0.7792 0.0085311 0.0094715 0.0015655 0.98457 0.9901 3.4014e-006 1.3606e-005 0.1581 0.70487 0.79496 0.0014892 0.82389 0.40381 0.0020028 0.41978 1.5608 1.5576 16.0121 144.9314 0.00034883 -84.9218 0.23895
6.343 0.9881 5.482e-005 3.8183 0.011956 8.2755e-005 0.001165 0.2333 0.00065931 0.23395 0.21588 0 0.032279 0.0389 0 1.3933 0.48321 0.1474 0.017832 11.6296 0.11095 0.0001422 0.7792 0.0085316 0.009472 0.0015641 0.98459 0.99011 3.3982e-006 1.3593e-005 0.15811 0.70574 0.79557 0.0014885 0.82493 0.40402 0.0020018 0.41978 1.5626 1.5594 16.0121 144.9315 0.00034795 -84.9272 0.23995
6.344 0.9881 5.482e-005 3.8183 0.011956 8.2768e-005 0.001165 0.2333 0.00065931 0.23395 0.21588 0 0.032279 0.0389 0 1.3934 0.48325 0.14742 0.017833 11.6319 0.11095 0.00014221 0.77919 0.0085321 0.0094726 0.0015628 0.98461 0.99013 3.3949e-006 1.358e-005 0.15811 0.7066 0.79618 0.0014878 0.82597 0.40422 0.0020009 0.41979 1.5644 1.5612 16.0121 144.9315 0.00034707 -84.9326 0.24095
6.345 0.9881 5.482e-005 3.8183 0.011956 8.2781e-005 0.001165 0.2333 0.00065931 0.23395 0.21588 0 0.032279 0.0389 0 1.3935 0.4833 0.14743 0.017835 11.6343 0.11096 0.00014223 0.77918 0.0085326 0.0094731 0.0015614 0.98463 0.99014 3.3917e-006 1.3567e-005 0.15812 0.70746 0.79678 0.0014871 0.82701 0.40442 0.002 0.4198 1.5662 1.563 16.0122 144.9315 0.0003462 -84.938 0.24195
6.346 0.9881 5.482e-005 3.8183 0.011956 8.2794e-005 0.001165 0.2333 0.00065931 0.23395 0.21588 0 0.032279 0.0389 0 1.3936 0.48335 0.14744 0.017836 11.6367 0.11097 0.00014224 0.77917 0.0085331 0.0094737 0.00156 0.98465 0.99016 3.3886e-006 1.3555e-005 0.15812 0.70832 0.79738 0.0014864 0.82803 0.40462 0.0019991 0.41981 1.568 1.5648 16.0122 144.9315 0.00034533 -84.9433 0.24295
6.347 0.9881 5.482e-005 3.8183 0.011956 8.2807e-005 0.001165 0.2333 0.00065931 0.23395 0.21588 0 0.032279 0.0389 0 1.3937 0.48339 0.14746 0.017837 11.6391 0.11098 0.00014225 0.77916 0.0085336 0.0094742 0.0015587 0.98466 0.99017 3.3854e-006 1.3542e-005 0.15812 0.70918 0.79798 0.0014857 0.82906 0.40483 0.0019982 0.41982 1.5697 1.5665 16.0122 144.9315 0.00034446 -84.9485 0.24395
6.348 0.9881 5.482e-005 3.8183 0.011956 8.282e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3938 0.48344 0.14747 0.017839 11.6415 0.11099 0.00014226 0.77916 0.0085341 0.0094748 0.0015573 0.98468 0.99018 3.3823e-006 1.3529e-005 0.15813 0.71003 0.79857 0.0014851 0.83007 0.40503 0.0019973 0.41983 1.5715 1.5683 16.0123 144.9315 0.0003436 -84.9537 0.24495
6.349 0.9881 5.4819e-005 3.8183 0.011956 8.2833e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3938 0.48348 0.14749 0.01784 11.6438 0.11099 0.00014227 0.77915 0.0085347 0.0094753 0.001556 0.9847 0.9902 3.3792e-006 1.3517e-005 0.15813 0.71088 0.79916 0.0014844 0.83108 0.40523 0.0019964 0.41984 1.5732 1.5701 16.0123 144.9315 0.00034275 -84.9589 0.24595
6.35 0.9881 5.4819e-005 3.8183 0.011956 8.2846e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3939 0.48353 0.1475 0.017841 11.6462 0.111 0.00014228 0.77914 0.0085352 0.0094759 0.0015546 0.98472 0.99021 3.3761e-006 1.3505e-005 0.15814 0.71173 0.79975 0.0014837 0.83209 0.40543 0.0019956 0.41985 1.575 1.5719 16.0124 144.9316 0.0003419 -84.9641 0.24695
6.351 0.98811 5.4819e-005 3.8183 0.011956 8.2859e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.394 0.48358 0.14752 0.017843 11.6486 0.11101 0.0001423 0.77913 0.0085357 0.0094764 0.0015533 0.98474 0.99022 3.3731e-006 1.3492e-005 0.15814 0.71258 0.80033 0.0014831 0.83309 0.40564 0.0019947 0.41986 1.5768 1.5736 16.0124 144.9316 0.00034105 -84.9692 0.24795
6.352 0.98811 5.4819e-005 3.8183 0.011956 8.2872e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3941 0.48362 0.14753 0.017844 11.651 0.11102 0.00014231 0.77912 0.0085362 0.009477 0.0015521 0.98475 0.99024 3.37e-006 1.348e-005 0.15814 0.71342 0.80091 0.0014824 0.83408 0.40584 0.0019938 0.41986 1.5785 1.5754 16.0124 144.9316 0.0003402 -84.9742 0.24895
6.353 0.98811 5.4819e-005 3.8183 0.011956 8.2884e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3942 0.48367 0.14755 0.017845 11.6533 0.11103 0.00014232 0.77912 0.0085367 0.0094775 0.0015508 0.98477 0.99025 3.367e-006 1.3468e-005 0.15815 0.71426 0.80148 0.0014818 0.83507 0.40604 0.001993 0.41987 1.5803 1.5771 16.0125 144.9316 0.00033936 -84.9793 0.24995
6.354 0.98811 5.4819e-005 3.8183 0.011956 8.2897e-005 0.001165 0.2333 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3943 0.48371 0.14756 0.017847 11.6557 0.11103 0.00014233 0.77911 0.0085372 0.0094781 0.0015496 0.98479 0.99026 3.3641e-006 1.3457e-005 0.15815 0.7151 0.80205 0.0014811 0.83605 0.40624 0.0019921 0.41988 1.582 1.5789 16.0125 144.9316 0.00033853 -84.9842 0.25095
6.355 0.98811 5.4819e-005 3.8183 0.011956 8.291e-005 0.001165 0.23331 0.00065931 0.23396 0.21588 0 0.032279 0.0389 0 1.3944 0.48376 0.14758 0.017848 11.6581 0.11104 0.00014234 0.7791 0.0085377 0.0094786 0.0015484 0.98481 0.99027 3.3611e-006 1.3445e-005 0.15816 0.71593 0.80262 0.0014805 0.83703 0.40645 0.0019913 0.41989 1.5837 1.5806 16.0125 144.9316 0.0003377 -84.9892 0.25195
6.356 0.98811 5.4819e-005 3.8183 0.011956 8.2923e-005 0.001165 0.23331 0.00065931 0.23396 0.21589 0 0.032279 0.0389 0 1.3945 0.48381 0.14759 0.017849 11.6605 0.11105 0.00014235 0.77909 0.0085382 0.0094792 0.0015471 0.98482 0.99029 3.3582e-006 1.3433e-005 0.15816 0.71676 0.80319 0.0014798 0.838 0.40665 0.0019905 0.4199 1.5855 1.5824 16.0126 144.9317 0.00033687 -84.9941 0.25295
6.357 0.98811 5.4819e-005 3.8183 0.011956 8.2936e-005 0.001165 0.23331 0.00065931 0.23396 0.21589 0 0.032279 0.0389 0 1.3946 0.48385 0.14761 0.017851 11.6629 0.11106 0.00014237 0.77908 0.0085387 0.0094797 0.0015458 0.98484 0.9903 3.3553e-006 1.3421e-005 0.15816 0.71759 0.80375 0.0014792 0.83897 0.40685 0.0019896 0.41991 1.5872 1.5841 16.0126 144.9317 0.00033605 -84.999 0.25395
6.358 0.98811 5.4819e-005 3.8183 0.011956 8.2949e-005 0.001165 0.23331 0.00065931 0.23396 0.21589 0 0.032279 0.0389 0 1.3947 0.4839 0.14762 0.017852 11.6652 0.11107 0.00014238 0.77908 0.0085392 0.0094803 0.0015445 0.98486 0.99031 3.3524e-006 1.341e-005 0.15817 0.71842 0.80431 0.0014786 0.83993 0.40705 0.0019888 0.41992 1.5889 1.5858 16.0126 144.9317 0.00033523 -85.0038 0.25495
6.359 0.98811 5.4819e-005 3.8183 0.011956 8.2962e-005 0.001165 0.23331 0.00065931 0.23396 0.21589 0 0.032279 0.0389 0 1.3948 0.48394 0.14764 0.017853 11.6676 0.11107 0.00014239 0.77907 0.0085398 0.0094808 0.0015431 0.98487 0.99032 3.3496e-006 1.3399e-005 0.15817 0.71925 0.80487 0.001478 0.84089 0.40726 0.001988 0.41993 1.5906 1.5876 16.0127 144.9317 0.00033441 -85.0086 0.25595
6.36 0.98811 5.4819e-005 3.8183 0.011956 8.2975e-005 0.001165 0.23331 0.00065931 0.23396 0.21589 0 0.032279 0.0389 0 1.3949 0.48399 0.14765 0.017855 11.67 0.11108 0.0001424 0.77906 0.0085403 0.0094813 0.0015418 0.98489 0.99033 3.3468e-006 1.3387e-005 0.15818 0.72007 0.80542 0.0014774 0.84184 0.40746 0.0019872 0.41994 1.5923 1.5893 16.0127 144.9317 0.0003336 -85.0134 0.25695
6.361 0.98811 5.4819e-005 3.8183 0.011956 8.2988e-005 0.001165 0.23331 0.00065931 0.23396 0.21589 0 0.032279 0.0389 0 1.3949 0.48404 0.14767 0.017856 11.6724 0.11109 0.00014241 0.77905 0.0085408 0.0094819 0.0015406 0.98491 0.99035 3.344e-006 1.3376e-005 0.15818 0.72089 0.80597 0.0014768 0.84279 0.40766 0.0019864 0.41995 1.5941 1.591 16.0127 144.9317 0.00033279 -85.0181 0.25795
6.362 0.98811 5.4818e-005 3.8183 0.011956 8.3001e-005 0.001165 0.23331 0.00065931 0.23397 0.21589 0 0.032279 0.0389 0 1.395 0.48408 0.14768 0.017857 11.6748 0.1111 0.00014243 0.77904 0.0085413 0.0094824 0.0015393 0.98492 0.99036 3.3412e-006 1.3365e-005 0.15818 0.72171 0.80652 0.0014762 0.84373 0.40786 0.0019856 0.41996 1.5958 1.5927 16.0128 144.9317 0.00033199 -85.0228 0.25895
6.363 0.98811 5.4818e-005 3.8183 0.011956 8.3013e-005 0.001165 0.23331 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3951 0.48413 0.14769 0.017859 11.6772 0.11111 0.00014244 0.77904 0.0085418 0.009483 0.0015381 0.98494 0.99037 3.3384e-006 1.3354e-005 0.15819 0.72252 0.80706 0.0014756 0.84466 0.40806 0.0019848 0.41997 1.5975 1.5944 16.0128 144.9318 0.00033119 -85.0275 0.25995
6.364 0.98811 5.4818e-005 3.8183 0.011956 8.3026e-005 0.001165 0.23331 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3952 0.48417 0.14771 0.01786 11.6795 0.11111 0.00014245 0.77903 0.0085423 0.0094835 0.001537 0.98496 0.99038 3.3357e-006 1.3343e-005 0.15819 0.72333 0.80761 0.001475 0.84559 0.40827 0.001984 0.41998 1.5992 1.5962 16.0128 144.9318 0.00033039 -85.0321 0.26095
6.365 0.98811 5.4818e-005 3.8183 0.011956 8.3039e-005 0.001165 0.23331 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3953 0.48422 0.14772 0.017861 11.6819 0.11112 0.00014246 0.77902 0.0085428 0.0094841 0.0015359 0.98497 0.99039 3.333e-006 1.3332e-005 0.1582 0.72414 0.80814 0.0014744 0.84651 0.40847 0.0019833 0.41999 1.6009 1.5979 16.0129 144.9318 0.0003296 -85.0367 0.26195
6.366 0.98811 5.4818e-005 3.8183 0.011956 8.3052e-005 0.001165 0.23331 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3954 0.48427 0.14774 0.017863 11.6843 0.11113 0.00014247 0.77901 0.0085433 0.0094846 0.0015348 0.98499 0.9904 3.3303e-006 1.3321e-005 0.1582 0.72495 0.80868 0.0014738 0.84743 0.40867 0.0019825 0.42 1.6025 1.5996 16.0129 144.9318 0.00032881 -85.0412 0.26295
6.367 0.98811 5.4818e-005 3.8183 0.011956 8.3065e-005 0.001165 0.23331 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3955 0.48431 0.14775 0.017864 11.6867 0.11114 0.00014248 0.779 0.0085438 0.0094852 0.0015337 0.985 0.99041 3.3276e-006 1.3311e-005 0.1582 0.72575 0.80921 0.0014732 0.84835 0.40887 0.0019817 0.42001 1.6042 1.6013 16.0129 144.9318 0.00032803 -85.0458 0.26395
6.368 0.98811 5.4818e-005 3.8183 0.011956 8.3078e-005 0.001165 0.23332 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3956 0.48436 0.14777 0.017865 11.6891 0.11115 0.0001425 0.779 0.0085443 0.0094857 0.0015326 0.98502 0.99042 3.325e-006 1.33e-005 0.15821 0.72656 0.80974 0.0014726 0.84926 0.40907 0.001981 0.42002 1.6059 1.6029 16.013 144.9318 0.00032725 -85.0503 0.26495
6.369 0.98811 5.4818e-005 3.8183 0.011956 8.3091e-005 0.001165 0.23332 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3957 0.4844 0.14778 0.017867 11.6915 0.11115 0.00014251 0.77899 0.0085448 0.0094863 0.0015316 0.98503 0.99043 3.3224e-006 1.329e-005 0.15821 0.72736 0.81027 0.001472 0.85016 0.40928 0.0019802 0.42003 1.6076 1.6046 16.013 144.9319 0.00032647 -85.0547 0.26595
6.37 0.98811 5.4818e-005 3.8183 0.011956 8.3104e-005 0.0011651 0.23332 0.00065931 0.23397 0.21589 0 0.032278 0.0389 0 1.3958 0.48445 0.1478 0.017868 11.6939 0.11116 0.00014252 0.77898 0.0085454 0.0094868 0.0015305 0.98505 0.99044 3.3198e-006 1.3279e-005 0.15821 0.72815 0.81079 0.0014714 0.85106 0.40948 0.0019795 0.42004 1.6093 1.6063 16.013 144.9319 0.0003257 -85.0591 0.26695
6.371 0.98811 5.4818e-005 3.8183 0.011956 8.3117e-005 0.0011651 0.23332 0.00065931 0.23397 0.2159 0 0.032278 0.0389 0 1.3959 0.4845 0.14781 0.017869 11.6962 0.11117 0.00014253 0.77897 0.0085459 0.0094874 0.0015294 0.98506 0.99045 3.3172e-006 1.3269e-005 0.15822 0.72895 0.81131 0.0014709 0.85195 0.40968 0.0019788 0.42005 1.6109 1.608 16.013 144.9319 0.00032493 -85.0635 0.26795
6.372 0.98811 5.4818e-005 3.8183 0.011956 8.313e-005 0.0011651 0.23332 0.00065931 0.23397 0.2159 0 0.032278 0.0389 0 1.396 0.48454 0.14783 0.01787 11.6986 0.11118 0.00014254 0.77896 0.0085464 0.0094879 0.0015283 0.98508 0.99047 3.3147e-006 1.3259e-005 0.15822 0.72974 0.81183 0.0014703 0.85284 0.40988 0.001978 0.42006 1.6126 1.6097 16.0131 144.9319 0.00032416 -85.0679 0.26895
6.373 0.98811 5.4818e-005 3.8183 0.011956 8.3142e-005 0.0011651 0.23332 0.00065931 0.23397 0.2159 0 0.032278 0.0389 0 1.3961 0.48459 0.14784 0.017872 11.701 0.11119 0.00014255 0.77896 0.0085469 0.0094885 0.0015272 0.98509 0.99048 3.3121e-006 1.3249e-005 0.15823 0.73053 0.81234 0.0014697 0.85373 0.41008 0.0019773 0.42007 1.6142 1.6113 16.0131 144.9319 0.0003234 -85.0722 0.26995
6.374 0.98811 5.4818e-005 3.8183 0.011956 8.3155e-005 0.0011651 0.23332 0.00065931 0.23397 0.2159 0 0.032278 0.0389 0 1.3961 0.48463 0.14786 0.017873 11.7034 0.11119 0.00014257 0.77895 0.0085474 0.009489 0.001526 0.98511 0.99049 3.3096e-006 1.3239e-005 0.15823 0.73132 0.81286 0.0014692 0.8546 0.41028 0.0019766 0.42008 1.6159 1.613 16.0131 144.9319 0.00032264 -85.0765 0.27095
6.375 0.98811 5.4817e-005 3.8183 0.011956 8.3168e-005 0.0011651 0.23332 0.00065931 0.23397 0.2159 0 0.032278 0.0389 0 1.3962 0.48468 0.14787 0.017874 11.7058 0.1112 0.00014258 0.77894 0.0085479 0.0094895 0.0015248 0.98512 0.9905 3.3071e-006 1.3229e-005 0.15823 0.7321 0.81337 0.0014687 0.85548 0.41049 0.0019759 0.42009 1.6175 1.6147 16.0132 144.932 0.00032188 -85.0807 0.27195
6.376 0.98811 5.4817e-005 3.8183 0.011956 8.3181e-005 0.0011651 0.23332 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3963 0.48473 0.14789 0.017876 11.7082 0.11121 0.00014259 0.77893 0.0085484 0.0094901 0.0015237 0.98514 0.99051 3.3046e-006 1.3219e-005 0.15824 0.73289 0.81387 0.0014681 0.85635 0.41069 0.0019751 0.4201 1.6192 1.6163 16.0132 144.932 0.00032113 -85.0849 0.27295
6.377 0.98811 5.4817e-005 3.8183 0.011956 8.3194e-005 0.0011651 0.23332 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3964 0.48477 0.1479 0.017877 11.7106 0.11122 0.0001426 0.77892 0.0085489 0.0094906 0.0015226 0.98515 0.99052 3.3022e-006 1.3209e-005 0.15824 0.73367 0.81438 0.0014676 0.85721 0.41089 0.0019744 0.42011 1.6208 1.618 16.0132 144.932 0.00032038 -85.0891 0.27395
6.378 0.98811 5.4817e-005 3.8183 0.011956 8.3207e-005 0.0011651 0.23332 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3965 0.48482 0.14792 0.017878 11.7129 0.11123 0.00014261 0.77892 0.0085494 0.0094912 0.0015215 0.98516 0.99052 3.2998e-006 1.3199e-005 0.15825 0.73444 0.81488 0.0014671 0.85807 0.41109 0.0019737 0.42012 1.6225 1.6196 16.0132 144.932 0.00031964 -85.0933 0.27495
6.379 0.98811 5.4817e-005 3.8183 0.011956 8.322e-005 0.0011651 0.23332 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3966 0.48486 0.14793 0.01788 11.7153 0.11123 0.00014262 0.77891 0.0085499 0.0094917 0.0015204 0.98518 0.99053 3.2974e-006 1.319e-005 0.15825 0.73522 0.81538 0.0014666 0.85892 0.41129 0.0019731 0.42013 1.6241 1.6213 16.0133 144.932 0.0003189 -85.0974 0.27595
6.38 0.98811 5.4817e-005 3.8183 0.011956 8.3233e-005 0.0011651 0.23332 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3967 0.48491 0.14795 0.017881 11.7177 0.11124 0.00014264 0.7789 0.0085504 0.0094923 0.0015194 0.98519 0.99054 3.295e-006 1.318e-005 0.15825 0.73599 0.81587 0.001466 0.85977 0.41149 0.0019724 0.42014 1.6257 1.6229 16.0133 144.932 0.00031816 -85.1015 0.27695
6.381 0.98811 5.4817e-005 3.8183 0.011956 8.3246e-005 0.0011651 0.23332 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3968 0.48496 0.14796 0.017882 11.7201 0.11125 0.00014265 0.77889 0.0085509 0.0094928 0.0015184 0.98521 0.99055 3.2926e-006 1.3171e-005 0.15826 0.73676 0.81637 0.0014655 0.86062 0.41169 0.0019717 0.42015 1.6274 1.6245 16.0133 144.9321 0.00031743 -85.1056 0.27795
6.382 0.98811 5.4817e-005 3.8183 0.011956 8.3259e-005 0.0011651 0.23333 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3969 0.485 0.14797 0.017884 11.7225 0.11126 0.00014266 0.77888 0.0085514 0.0094934 0.0015173 0.98522 0.99056 3.2902e-006 1.3161e-005 0.15826 0.73753 0.81686 0.001465 0.86145 0.4119 0.001971 0.42016 1.629 1.6262 16.0134 144.9321 0.0003167 -85.1096 0.27895
6.383 0.98811 5.4817e-005 3.8183 0.011956 8.3271e-005 0.0011651 0.23333 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.397 0.48505 0.14799 0.017885 11.7249 0.11127 0.00014267 0.77888 0.008552 0.0094939 0.0015164 0.98523 0.99057 3.2879e-006 1.3152e-005 0.15827 0.7383 0.81734 0.0014645 0.86229 0.4121 0.0019703 0.42017 1.6306 1.6278 16.0134 144.9321 0.00031597 -85.1136 0.27995
6.384 0.98811 5.4817e-005 3.8183 0.011956 8.3284e-005 0.0011651 0.23333 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3971 0.48509 0.148 0.017886 11.7273 0.11127 0.00014268 0.77887 0.0085525 0.0094945 0.0015154 0.98525 0.99058 3.2856e-006 1.3143e-005 0.15827 0.73906 0.81783 0.001464 0.86312 0.4123 0.0019697 0.42018 1.6322 1.6294 16.0134 144.9321 0.00031525 -85.1176 0.28095
6.385 0.98811 5.4817e-005 3.8183 0.011956 8.3297e-005 0.0011651 0.23333 0.00065931 0.23398 0.2159 0 0.032278 0.0389 0 1.3972 0.48514 0.14802 0.017888 11.7297 0.11128 0.0001427 0.77886 0.008553 0.009495 0.0015144 0.98526 0.99059 3.2833e-006 1.3133e-005 0.15827 0.73982 0.81831 0.0014635 0.86394 0.4125 0.001969 0.42019 1.6338 1.631 16.0134 144.9321 0.00031453 -85.1216 0.28195
6.386 0.98811 5.4817e-005 3.8183 0.011956 8.331e-005 0.0011651 0.23333 0.00065931 0.23398 0.21591 0 0.032278 0.0389 0 1.3972 0.48519 0.14803 0.017889 11.7321 0.11129 0.00014271 0.77885 0.0085535 0.0094955 0.0015135 0.98527 0.9906 3.281e-006 1.3124e-005 0.15828 0.74058 0.81879 0.001463 0.86476 0.4127 0.0019684 0.4202 1.6354 1.6326 16.0135 144.9321 0.00031381 -85.1255 0.28295
6.387 0.98811 5.4817e-005 3.8183 0.011956 8.3323e-005 0.0011651 0.23333 0.00065931 0.23398 0.21591 0 0.032278 0.0389 0 1.3973 0.48523 0.14805 0.01789 11.7345 0.1113 0.00014272 0.77884 0.008554 0.0094961 0.0015125 0.98529 0.99061 3.2788e-006 1.3115e-005 0.15828 0.74134 0.81927 0.0014625 0.86558 0.4129 0.0019677 0.42021 1.637 1.6343 16.0135 144.9321 0.0003131 -85.1294 0.28395
6.388 0.98811 5.4816e-005 3.8183 0.011956 8.3336e-005 0.0011651 0.23333 0.00065931 0.23398 0.21591 0 0.032278 0.0389 0 1.3974 0.48528 0.14806 0.017892 11.7368 0.11131 0.00014273 0.77884 0.0085545 0.0094966 0.0015115 0.9853 0.99062 3.2765e-006 1.3106e-005 0.15829 0.74209 0.81975 0.001462 0.86639 0.4131 0.0019671 0.42022 1.6386 1.6359 16.0135 144.9322 0.00031239 -85.1332 0.28495
6.389 0.98811 5.4816e-005 3.8183 0.011956 8.3349e-005 0.0011651 0.23333 0.00065931 0.23398 0.21591 0 0.032278 0.0389 0 1.3975 0.48532 0.14808 0.017893 11.7392 0.11131 0.00014274 0.77883 0.008555 0.0094972 0.0015105 0.98531 0.99063 3.2743e-006 1.3097e-005 0.15829 0.74284 0.82022 0.0014615 0.8672 0.4133 0.0019664 0.42023 1.6402 1.6375 16.0135 144.9322 0.00031168 -85.1371 0.28595
6.39 0.98811 5.4816e-005 3.8183 0.011956 8.3362e-005 0.0011651 0.23333 0.00065931 0.23399 0.21591 0 0.032278 0.0389 0 1.3976 0.48537 0.14809 0.017894 11.7416 0.11132 0.00014275 0.77882 0.0085555 0.0094977 0.0015095 0.98533 0.99063 3.2721e-006 1.3089e-005 0.15829 0.74359 0.82069 0.001461 0.868 0.41351 0.0019658 0.42025 1.6418 1.6391 16.0136 144.9322 0.00031098 -85.1409 0.28695
6.391 0.98811 5.4816e-005 3.8183 0.011955 8.3375e-005 0.0011651 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3977 0.48542 0.14811 0.017896 11.744 0.11133 0.00014277 0.77881 0.008556 0.0094983 0.0015086 0.98534 0.99064 3.2699e-006 1.308e-005 0.1583 0.74434 0.82116 0.0014605 0.86879 0.41371 0.0019651 0.42026 1.6434 1.6406 16.0136 144.9322 0.00031028 -85.1446 0.28795
6.392 0.98811 5.4816e-005 3.8183 0.011955 8.3388e-005 0.0011651 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3978 0.48546 0.14812 0.017897 11.7464 0.11134 0.00014278 0.7788 0.0085565 0.0094988 0.0015077 0.98535 0.99065 3.2678e-006 1.3071e-005 0.1583 0.74508 0.82162 0.00146 0.86959 0.41391 0.0019645 0.42027 1.645 1.6422 16.0136 144.9322 0.00030958 -85.1484 0.28895
6.393 0.98811 5.4816e-005 3.8183 0.011955 8.34e-005 0.0011651 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3979 0.48551 0.14814 0.017898 11.7488 0.11135 0.00014279 0.7788 0.008557 0.0094994 0.0015068 0.98536 0.99066 3.2656e-006 1.3063e-005 0.15831 0.74583 0.82209 0.0014595 0.87037 0.41411 0.0019639 0.42028 1.6465 1.6438 16.0136 144.9322 0.00030889 -85.1521 0.28995
6.394 0.98811 5.4816e-005 3.8183 0.011955 8.3413e-005 0.0011651 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.398 0.48555 0.14815 0.017899 11.7512 0.11135 0.0001428 0.77879 0.0085575 0.0094999 0.0015059 0.98538 0.99067 3.2635e-006 1.3054e-005 0.15831 0.74657 0.82255 0.0014591 0.87116 0.41431 0.0019633 0.42029 1.6481 1.6454 16.0137 144.9323 0.0003082 -85.1558 0.29095
6.395 0.98811 5.4816e-005 3.8183 0.011955 8.3426e-005 0.0011651 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3981 0.4856 0.14817 0.017901 11.7536 0.11136 0.00014281 0.77878 0.008558 0.0095004 0.0015051 0.98539 0.99068 3.2614e-006 1.3046e-005 0.15831 0.7473 0.823 0.0014586 0.87194 0.41451 0.0019627 0.4203 1.6497 1.647 16.0137 144.9323 0.00030751 -85.1595 0.29195
6.396 0.98811 5.4816e-005 3.8183 0.011955 8.3439e-005 0.0011652 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3982 0.48565 0.14818 0.017902 11.756 0.11137 0.00014282 0.77877 0.0085585 0.009501 0.0015041 0.9854 0.99069 3.2593e-006 1.3037e-005 0.15832 0.74804 0.82346 0.0014581 0.87271 0.41471 0.0019621 0.42031 1.6512 1.6485 16.0137 144.9323 0.00030683 -85.1631 0.29295
6.397 0.98811 5.4816e-005 3.8183 0.011955 8.3452e-005 0.0011652 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3983 0.48569 0.1482 0.017903 11.7584 0.11138 0.00014284 0.77876 0.008559 0.0095015 0.0015032 0.98541 0.99069 3.2572e-006 1.3029e-005 0.15832 0.74877 0.82391 0.0014577 0.87348 0.41491 0.0019615 0.42032 1.6528 1.6501 16.0137 144.9323 0.00030615 -85.1667 0.29395
6.398 0.98811 5.4816e-005 3.8183 0.011955 8.3465e-005 0.0011652 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3983 0.48574 0.14821 0.017905 11.7608 0.11139 0.00014285 0.77876 0.0085596 0.0095021 0.0015022 0.98542 0.9907 3.2551e-006 1.3021e-005 0.15833 0.7495 0.82437 0.0014572 0.87424 0.41511 0.0019609 0.42033 1.6543 1.6517 16.0137 144.9323 0.00030547 -85.1703 0.29495
6.399 0.98811 5.4816e-005 3.8183 0.011955 8.3478e-005 0.0011652 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3984 0.48578 0.14822 0.017906 11.7632 0.11139 0.00014286 0.77875 0.0085601 0.0095026 0.0015012 0.98544 0.99071 3.2531e-006 1.3012e-005 0.15833 0.75023 0.82481 0.0014568 0.87501 0.41531 0.0019603 0.42034 1.6559 1.6532 16.0138 144.9323 0.0003048 -85.1738 0.29595
6.4 0.98811 5.4816e-005 3.8183 0.011955 8.3491e-005 0.0011652 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.3985 0.48583 0.14824 0.017907 11.7656 0.1114 0.00014287 0.77874 0.0085606 0.0095032 0.0015003 0.98545 0.99072 3.251e-006 1.3004e-005 0.15833 0.75096 0.82526 0.0014563 0.87576 0.41551 0.0019597 0.42036 1.6574 1.6548 16.0138 144.9324 0.00030413 -85.1774 0.29695
6.401 0.98811 5.4815e-005 3.8183 0.011955 8.3504e-005 0.0011652 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.3986 0.48588 0.14825 0.017909 11.768 0.11141 0.00014288 0.77873 0.0085611 0.0095037 0.0014994 0.98546 0.99073 3.249e-006 1.2996e-005 0.15834 0.75168 0.8257 0.0014559 0.87651 0.41571 0.0019591 0.42037 1.659 1.6563 16.0138 144.9324 0.00030346 -85.1809 0.29795
6.402 0.98811 5.4815e-005 3.8183 0.011955 8.3517e-005 0.0011652 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.3987 0.48592 0.14827 0.01791 11.7704 0.11142 0.00014289 0.77872 0.0085616 0.0095042 0.0014985 0.98547 0.99073 3.247e-006 1.2988e-005 0.15834 0.7524 0.82615 0.0014554 0.87726 0.41591 0.0019585 0.42038 1.6605 1.6579 16.0138 144.9324 0.00030279 -85.1844 0.29895
6.403 0.98811 5.4815e-005 3.8183 0.011955 8.3529e-005 0.0011652 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.3988 0.48597 0.14828 0.017911 11.7728 0.11143 0.00014291 0.77872 0.0085621 0.0095048 0.0014977 0.98548 0.99074 3.245e-006 1.298e-005 0.15835 0.75312 0.82659 0.001455 0.878 0.41611 0.0019579 0.42039 1.6621 1.6594 16.0139 144.9324 0.00030213 -85.1878 0.29995
6.404 0.98811 5.4815e-005 3.8183 0.011955 8.3542e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3989 0.48601 0.1483 0.017913 11.7752 0.11143 0.00014292 0.77871 0.0085626 0.0095053 0.0014968 0.98549 0.99075 3.2431e-006 1.2972e-005 0.15835 0.75384 0.82702 0.0014545 0.87874 0.41631 0.0019574 0.4204 1.6636 1.661 16.0139 144.9324 0.00030147 -85.1912 0.30095
6.405 0.98811 5.4815e-005 3.8183 0.011955 8.3555e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.399 0.48606 0.14831 0.017914 11.7776 0.11144 0.00014293 0.7787 0.0085631 0.0095059 0.001496 0.98551 0.99076 3.2411e-006 1.2965e-005 0.15835 0.75456 0.82746 0.0014541 0.87948 0.41652 0.0019568 0.42041 1.6651 1.6625 16.0139 144.9324 0.00030082 -85.1946 0.30195
6.406 0.98811 5.4815e-005 3.8183 0.011955 8.3568e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3991 0.48611 0.14833 0.017915 11.78 0.11145 0.00014294 0.77869 0.0085636 0.0095064 0.0014952 0.98552 0.99076 3.2392e-006 1.2957e-005 0.15836 0.75527 0.82789 0.0014537 0.88021 0.41672 0.0019563 0.42042 1.6666 1.664 16.0139 144.9325 0.00030017 -85.198 0.30295
6.407 0.98811 5.4815e-005 3.8183 0.011955 8.3581e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3992 0.48615 0.14834 0.017917 11.7824 0.11146 0.00014295 0.77868 0.0085641 0.009507 0.0014944 0.98553 0.99077 3.2373e-006 1.2949e-005 0.15836 0.75598 0.82832 0.0014533 0.88093 0.41692 0.0019557 0.42043 1.6682 1.6656 16.0139 144.9325 0.00029952 -85.2014 0.30395
6.408 0.98811 5.4815e-005 3.8183 0.011955 8.3594e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3993 0.4862 0.14836 0.017918 11.7848 0.11147 0.00014296 0.77868 0.0085646 0.0095075 0.0014936 0.98554 0.99078 3.2354e-006 1.2942e-005 0.15837 0.75669 0.82875 0.0014528 0.88166 0.41712 0.0019551 0.42045 1.6697 1.6671 16.014 144.9325 0.00029887 -85.2047 0.30495
6.409 0.98811 5.4815e-005 3.8183 0.011955 8.3607e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3994 0.48624 0.14837 0.017919 11.7872 0.11147 0.00014298 0.77867 0.0085651 0.009508 0.0014929 0.98555 0.99079 3.2335e-006 1.2934e-005 0.15837 0.7574 0.82918 0.0014524 0.88237 0.41732 0.0019546 0.42046 1.6712 1.6686 16.014 144.9325 0.00029823 -85.208 0.30595
6.41 0.98811 5.4815e-005 3.8183 0.011955 8.362e-005 0.0011652 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3994 0.48629 0.14839 0.017921 11.7896 0.11148 0.00014299 0.77866 0.0085656 0.0095086 0.0014921 0.98556 0.99079 3.2316e-006 1.2927e-005 0.15837 0.7581 0.8296 0.001452 0.88309 0.41752 0.001954 0.42047 1.6727 1.6701 16.014 144.9325 0.00029759 -85.2113 0.30695
6.411 0.98811 5.4815e-005 3.8183 0.011955 8.3633e-005 0.0011652 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3995 0.48634 0.1484 0.017922 11.792 0.11149 0.000143 0.77865 0.0085661 0.0095091 0.0014913 0.98557 0.9908 3.2298e-006 1.2919e-005 0.15838 0.7588 0.83002 0.0014516 0.8838 0.41772 0.0019535 0.42048 1.6742 1.6716 16.014 144.9326 0.00029695 -85.2145 0.30795
6.412 0.98811 5.4815e-005 3.8183 0.011955 8.3646e-005 0.0011652 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3996 0.48638 0.14842 0.017923 11.7944 0.1115 0.00014301 0.77864 0.0085666 0.0095097 0.0014905 0.98558 0.99081 3.2279e-006 1.2912e-005 0.15838 0.7595 0.83044 0.0014512 0.8845 0.41792 0.001953 0.42049 1.6757 1.6731 16.014 144.9326 0.00029631 -85.2177 0.30895
6.413 0.98811 5.4815e-005 3.8183 0.011955 8.3658e-005 0.0011652 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3997 0.48643 0.14843 0.017924 11.7968 0.11151 0.00014302 0.77864 0.0085671 0.0095102 0.0014897 0.98559 0.99081 3.2261e-006 1.2904e-005 0.15839 0.7602 0.83086 0.0014508 0.8852 0.41812 0.0019524 0.4205 1.6772 1.6746 16.0141 144.9326 0.00029568 -85.2209 0.30995
6.414 0.98811 5.4814e-005 3.8183 0.011955 8.3671e-005 0.0011652 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3998 0.48647 0.14845 0.017926 11.7992 0.11151 0.00014303 0.77863 0.0085676 0.0095108 0.0014889 0.9856 0.99082 3.2243e-006 1.2897e-005 0.15839 0.7609 0.83128 0.0014504 0.8859 0.41832 0.0019519 0.42052 1.6787 1.6761 16.0141 144.9326 0.00029505 -85.2241 0.31095
6.415 0.98811 5.4814e-005 3.8183 0.011955 8.3684e-005 0.0011652 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.3999 0.48652 0.14846 0.017927 11.8016 0.11152 0.00014305 0.77862 0.0085681 0.0095113 0.0014881 0.98561 0.99083 3.2225e-006 1.289e-005 0.15839 0.76159 0.83169 0.00145 0.88659 0.41852 0.0019514 0.42053 1.6802 1.6776 16.0141 144.9326 0.00029443 -85.2273 0.31195
6.416 0.98811 5.4814e-005 3.8183 0.011955 8.3697e-005 0.0011652 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.4 0.48657 0.14847 0.017928 11.804 0.11153 0.00014306 0.77861 0.0085686 0.0095118 0.0014873 0.98562 0.99084 3.2207e-006 1.2883e-005 0.1584 0.76228 0.8321 0.0014496 0.88728 0.41872 0.0019509 0.42054 1.6816 1.6791 16.0141 144.9326 0.00029381 -85.2304 0.31295
6.417 0.98811 5.4814e-005 3.8183 0.011955 8.371e-005 0.0011652 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.4001 0.48661 0.14849 0.01793 11.8064 0.11154 0.00014307 0.77861 0.0085692 0.0095124 0.0014866 0.98563 0.99084 3.2189e-006 1.2876e-005 0.1584 0.76297 0.83251 0.0014492 0.88796 0.41892 0.0019504 0.42055 1.6831 1.6806 16.0141 144.9327 0.00029319 -85.2335 0.31395
6.418 0.98811 5.4814e-005 3.8183 0.011955 8.3723e-005 0.0011652 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.4002 0.48666 0.1485 0.017931 11.8088 0.11155 0.00014308 0.7786 0.0085697 0.0095129 0.0014858 0.98564 0.99085 3.2171e-006 1.2869e-005 0.1584 0.76366 0.83292 0.0014488 0.88864 0.41912 0.0019498 0.42056 1.6846 1.6821 16.0142 144.9327 0.00029257 -85.2366 0.31495
6.419 0.98811 5.4814e-005 3.8183 0.011955 8.3736e-005 0.0011652 0.23335 0.00065931 0.23401 0.21593 0 0.032277 0.0389 0 1.4003 0.4867 0.14852 0.017932 11.8112 0.11155 0.00014309 0.77859 0.0085702 0.0095135 0.001485 0.98565 0.99086 3.2154e-006 1.2862e-005 0.15841 0.76434 0.83333 0.0014484 0.88932 0.41931 0.0019493 0.42057 1.6861 1.6836 16.0142 144.9327 0.00029195 -85.2397 0.31595
6.42 0.98811 5.4814e-005 3.8183 0.011955 8.3749e-005 0.0011652 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4004 0.48675 0.14853 0.017934 11.8136 0.11156 0.0001431 0.77858 0.0085707 0.009514 0.0014842 0.98566 0.99086 3.2137e-006 1.2855e-005 0.15841 0.76503 0.83373 0.001448 0.88999 0.41951 0.0019488 0.42059 1.6875 1.6851 16.0142 144.9327 0.00029134 -85.2427 0.31695
6.421 0.98811 5.4814e-005 3.8183 0.011955 8.3762e-005 0.0011652 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4005 0.4868 0.14855 0.017935 11.816 0.11157 0.00014312 0.77857 0.0085712 0.0095146 0.0014834 0.98567 0.99087 3.212e-006 1.2848e-005 0.15842 0.76571 0.83413 0.0014476 0.89066 0.41971 0.0019483 0.4206 1.689 1.6865 16.0142 144.9327 0.00029073 -85.2457 0.31795
6.422 0.98811 5.4814e-005 3.8183 0.011955 8.3775e-005 0.0011653 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4005 0.48684 0.14856 0.017936 11.8184 0.11158 0.00014313 0.77857 0.0085717 0.0095151 0.0014827 0.98568 0.99088 3.2102e-006 1.2841e-005 0.15842 0.76638 0.83453 0.0014472 0.89133 0.41991 0.0019478 0.42061 1.6904 1.688 16.0142 144.9327 0.00029013 -85.2487 0.31895
6.423 0.98811 5.4814e-005 3.8183 0.011955 8.3787e-005 0.0011653 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4006 0.48689 0.14858 0.017938 11.8208 0.11159 0.00014314 0.77856 0.0085722 0.0095156 0.0014819 0.98569 0.99088 3.2086e-006 1.2834e-005 0.15842 0.76706 0.83493 0.0014469 0.89199 0.42011 0.0019473 0.42062 1.6919 1.6895 16.0142 144.9328 0.00028953 -85.2517 0.31995
6.424 0.98811 5.4814e-005 3.8183 0.011955 8.38e-005 0.0011653 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4007 0.48693 0.14859 0.017939 11.8232 0.11159 0.00014315 0.77855 0.0085727 0.0095162 0.0014812 0.9857 0.99089 3.2069e-006 1.2828e-005 0.15843 0.76774 0.83533 0.0014465 0.89264 0.42031 0.0019468 0.42063 1.6934 1.6909 16.0143 144.9328 0.00028893 -85.2547 0.32095
6.425 0.98811 5.4814e-005 3.8183 0.011955 8.3813e-005 0.0011653 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4008 0.48698 0.14861 0.01794 11.8256 0.1116 0.00014316 0.77854 0.0085732 0.0095167 0.0014805 0.98571 0.9909 3.2052e-006 1.2821e-005 0.15843 0.76841 0.83572 0.0014461 0.89329 0.42051 0.0019464 0.42065 1.6948 1.6924 16.0143 144.9328 0.00028833 -85.2576 0.32195
6.426 0.98811 5.4814e-005 3.8183 0.011955 8.3826e-005 0.0011653 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4009 0.48703 0.14862 0.017942 11.828 0.11161 0.00014317 0.77853 0.0085737 0.0095173 0.0014797 0.98572 0.9909 3.2036e-006 1.2814e-005 0.15844 0.76908 0.83611 0.0014458 0.89394 0.42071 0.0019459 0.42066 1.6962 1.6938 16.0143 144.9328 0.00028773 -85.2605 0.32295
6.427 0.98811 5.4813e-005 3.8183 0.011955 8.3839e-005 0.0011653 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.401 0.48707 0.14864 0.017943 11.8304 0.11162 0.00014319 0.77853 0.0085742 0.0095178 0.001479 0.98573 0.99091 3.2019e-006 1.2808e-005 0.15844 0.76975 0.8365 0.0014454 0.89459 0.42091 0.0019454 0.42067 1.6977 1.6953 16.0143 144.9328 0.00028714 -85.2634 0.32395
6.428 0.98811 5.4813e-005 3.8183 0.011955 8.3852e-005 0.0011653 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4011 0.48712 0.14865 0.017944 11.8328 0.11163 0.0001432 0.77852 0.0085747 0.0095183 0.0014783 0.98574 0.99091 3.2003e-006 1.2801e-005 0.15844 0.77041 0.83689 0.001445 0.89523 0.42111 0.0019449 0.42068 1.6991 1.6967 16.0143 144.9328 0.00028655 -85.2663 0.32495
6.429 0.98811 5.4813e-005 3.8183 0.011955 8.3865e-005 0.0011653 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4012 0.48716 0.14867 0.017945 11.8352 0.11163 0.00014321 0.77851 0.0085752 0.0095189 0.0014776 0.98575 0.99092 3.1987e-006 1.2795e-005 0.15845 0.77108 0.83728 0.0014447 0.89587 0.42131 0.0019445 0.42069 1.7005 1.6982 16.0143 144.9329 0.00028597 -85.2691 0.32595
6.43 0.98811 5.4813e-005 3.8183 0.011955 8.3878e-005 0.0011653 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.4013 0.48721 0.14868 0.017947 11.8376 0.11164 0.00014322 0.7785 0.0085757 0.0095194 0.001477 0.98576 0.99093 3.1971e-006 1.2788e-005 0.15845 0.77174 0.83766 0.0014443 0.8965 0.42151 0.001944 0.42071 1.702 1.6996 16.0144 144.9329 0.00028538 -85.2719 0.32695
6.431 0.98811 5.4813e-005 3.8183 0.011955 8.3891e-005 0.0011653 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.4014 0.48726 0.14869 0.017948 11.84 0.11165 0.00014323 0.77849 0.0085762 0.00952 0.0014763 0.98577 0.99093 3.1955e-006 1.2782e-005 0.15846 0.7724 0.83804 0.001444 0.89713 0.42171 0.0019435 0.42072 1.7034 1.701 16.0144 144.9329 0.0002848 -85.2747 0.32795
6.432 0.98811 5.4813e-005 3.8183 0.011955 8.3904e-005 0.0011653 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.4015 0.4873 0.14871 0.017949 11.8424 0.11166 0.00014325 0.77849 0.0085767 0.0095205 0.0014756 0.98578 0.99094 3.1939e-006 1.2776e-005 0.15846 0.77306 0.83842 0.0014436 0.89776 0.42191 0.0019431 0.42073 1.7048 1.7025 16.0144 144.9329 0.00028422 -85.2775 0.32895
6.433 0.98811 5.4813e-005 3.8183 0.011955 8.3916e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4016 0.48735 0.14872 0.017951 11.8448 0.11167 0.00014326 0.77848 0.0085772 0.009521 0.001475 0.98579 0.99094 3.1924e-006 1.277e-005 0.15846 0.77371 0.8388 0.0014433 0.89838 0.42211 0.0019426 0.42074 1.7062 1.7039 16.0144 144.9329 0.00028365 -85.2803 0.32995
6.434 0.98811 5.4813e-005 3.8183 0.011955 8.3929e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4016 0.48739 0.14874 0.017952 11.8472 0.11167 0.00014327 0.77847 0.0085777 0.0095216 0.0014743 0.9858 0.99095 3.1908e-006 1.2763e-005 0.15847 0.77437 0.83918 0.0014429 0.899 0.4223 0.0019422 0.42075 1.7076 1.7053 16.0144 144.9329 0.00028307 -85.283 0.33095
6.435 0.98811 5.4813e-005 3.8183 0.011955 8.3942e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4017 0.48744 0.14875 0.017953 11.8496 0.11168 0.00014328 0.77846 0.0085782 0.0095221 0.0014737 0.9858 0.99096 3.1893e-006 1.2757e-005 0.15847 0.77502 0.83955 0.0014426 0.89961 0.4225 0.0019417 0.42077 1.7091 1.7067 16.0144 144.933 0.0002825 -85.2857 0.33195
6.436 0.98811 5.4813e-005 3.8183 0.011955 8.3955e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4018 0.48749 0.14877 0.017955 11.8521 0.11169 0.00014329 0.77845 0.0085787 0.0095227 0.001473 0.98581 0.99096 3.1877e-006 1.2751e-005 0.15848 0.77567 0.83993 0.0014422 0.90022 0.4227 0.0019413 0.42078 1.7105 1.7081 16.0144 144.933 0.00028193 -85.2885 0.33295
6.437 0.98811 5.4813e-005 3.8183 0.011955 8.3968e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4019 0.48753 0.14878 0.017956 11.8545 0.1117 0.0001433 0.77845 0.0085792 0.0095232 0.0014723 0.98582 0.99097 3.1862e-006 1.2745e-005 0.15848 0.77632 0.8403 0.0014419 0.90083 0.4229 0.0019408 0.42079 1.7119 1.7095 16.0145 144.933 0.00028137 -85.2911 0.33395
6.438 0.98811 5.4813e-005 3.8183 0.011955 8.3981e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.402 0.48758 0.1488 0.017957 11.8569 0.11171 0.00014332 0.77844 0.0085797 0.0095238 0.0014717 0.98583 0.99097 3.1847e-006 1.2739e-005 0.15848 0.77696 0.84067 0.0014416 0.90143 0.4231 0.0019404 0.4208 1.7133 1.7109 16.0145 144.933 0.00028081 -85.2938 0.33495
6.439 0.98811 5.4812e-005 3.8183 0.011955 8.3994e-005 0.0011653 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4021 0.48762 0.14881 0.017959 11.8593 0.11171 0.00014333 0.77843 0.0085802 0.0095243 0.001471 0.98584 0.99098 3.1832e-006 1.2733e-005 0.15849 0.7776 0.84103 0.0014412 0.90203 0.4233 0.0019399 0.42082 1.7147 1.7123 16.0145 144.933 0.00028024 -85.2964 0.33595
6.44 0.98811 5.4812e-005 3.8183 0.011955 8.4007e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4022 0.48767 0.14883 0.01796 11.8617 0.11172 0.00014334 0.77842 0.0085807 0.0095248 0.0014704 0.98585 0.99099 3.1818e-006 1.2727e-005 0.15849 0.77825 0.8414 0.0014409 0.90263 0.4235 0.0019395 0.42083 1.716 1.7137 16.0145 144.9331 0.00027969 -85.2991 0.33695
6.441 0.98811 5.4812e-005 3.8183 0.011955 8.402e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4023 0.48772 0.14884 0.017961 11.8641 0.11173 0.00014335 0.77841 0.0085812 0.0095254 0.0014697 0.98586 0.99099 3.1803e-006 1.2721e-005 0.1585 0.77889 0.84176 0.0014406 0.90322 0.4237 0.0019391 0.42084 1.7174 1.7151 16.0145 144.9331 0.00027913 -85.3017 0.33795
6.442 0.98811 5.4812e-005 3.8183 0.011955 8.4033e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4024 0.48776 0.14886 0.017963 11.8665 0.11174 0.00014336 0.77841 0.0085817 0.0095259 0.001469 0.98586 0.991 3.1788e-006 1.2715e-005 0.1585 0.77952 0.84213 0.0014402 0.90381 0.42389 0.0019387 0.42085 1.7188 1.7165 16.0145 144.9331 0.00027858 -85.3043 0.33895
6.443 0.98811 5.4812e-005 3.8183 0.011955 8.4045e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4025 0.48781 0.14887 0.017964 11.8689 0.11174 0.00014337 0.7784 0.0085822 0.0095265 0.0014684 0.98587 0.991 3.1774e-006 1.271e-005 0.1585 0.78016 0.84249 0.0014399 0.9044 0.42409 0.0019382 0.42087 1.7202 1.7179 16.0145 144.9331 0.00027803 -85.3068 0.33995
6.444 0.98811 5.4812e-005 3.8183 0.011955 8.4058e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4026 0.48785 0.14889 0.017965 11.8713 0.11175 0.00014339 0.77839 0.0085827 0.009527 0.0014677 0.98588 0.99101 3.176e-006 1.2704e-005 0.15851 0.78079 0.84285 0.0014396 0.90498 0.42429 0.0019378 0.42088 1.7216 1.7193 16.0145 144.9331 0.00027748 -85.3094 0.34095
6.445 0.98811 5.4812e-005 3.8183 0.011955 8.4071e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4027 0.4879 0.1489 0.017966 11.8737 0.11176 0.0001434 0.77838 0.0085833 0.0095275 0.0014671 0.98589 0.99101 3.1745e-006 1.2698e-005 0.15851 0.78143 0.8432 0.0014393 0.90556 0.42449 0.0019374 0.42089 1.7229 1.7207 16.0146 144.9331 0.00027694 -85.3119 0.34195
6.446 0.98811 5.4812e-005 3.8183 0.011955 8.4084e-005 0.0011653 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.4027 0.48795 0.14891 0.017968 11.8762 0.11177 0.00014341 0.77837 0.0085838 0.0095281 0.0014665 0.9859 0.99102 3.1731e-006 1.2693e-005 0.15851 0.78205 0.84356 0.0014389 0.90614 0.42469 0.001937 0.4209 1.7243 1.722 16.0146 144.9332 0.00027639 -85.3144 0.34295
6.447 0.98811 5.4812e-005 3.8183 0.011955 8.4097e-005 0.0011653 0.23337 0.00065931 0.23402 0.21595 0 0.032276 0.0389 0 1.4028 0.48799 0.14893 0.017969 11.8786 0.11178 0.00014342 0.77837 0.0085843 0.0095286 0.0014659 0.98591 0.99102 3.1717e-006 1.2687e-005 0.15852 0.78268 0.84391 0.0014386 0.90671 0.42489 0.0019366 0.42092 1.7257 1.7234 16.0146 144.9332 0.00027585 -85.3169 0.34395
6.448 0.98811 5.4812e-005 3.8183 0.011955 8.411e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.4029 0.48804 0.14894 0.01797 11.881 0.11178 0.00014343 0.77836 0.0085848 0.0095291 0.0014653 0.98591 0.99103 3.1704e-006 1.2681e-005 0.15852 0.78331 0.84427 0.0014383 0.90728 0.42508 0.0019362 0.42093 1.727 1.7248 16.0146 144.9332 0.00027531 -85.3194 0.34495
6.449 0.98811 5.4812e-005 3.8183 0.011955 8.4123e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.403 0.48808 0.14896 0.017972 11.8834 0.11179 0.00014344 0.77835 0.0085853 0.0095297 0.0014647 0.98592 0.99103 3.169e-006 1.2676e-005 0.15853 0.78393 0.84462 0.001438 0.90784 0.42528 0.0019358 0.42094 1.7284 1.7261 16.0146 144.9332 0.00027478 -85.3218 0.34595
6.45 0.98811 5.4812e-005 3.8183 0.011955 8.4136e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4031 0.48813 0.14897 0.017973 11.8858 0.1118 0.00014345 0.77834 0.0085858 0.0095302 0.0014641 0.98593 0.99104 3.1676e-006 1.267e-005 0.15853 0.78455 0.84497 0.0014377 0.9084 0.42548 0.0019354 0.42095 1.7297 1.7275 16.0146 144.9332 0.00027425 -85.3243 0.34695
6.451 0.98811 5.4812e-005 3.8183 0.011954 8.4149e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4032 0.48818 0.14899 0.017974 11.8882 0.11181 0.00014347 0.77833 0.0085863 0.0095308 0.0014635 0.98594 0.99104 3.1663e-006 1.2665e-005 0.15853 0.78518 0.84531 0.0014374 0.90896 0.42568 0.001935 0.42097 1.7311 1.7289 16.0146 144.9333 0.00027371 -85.3267 0.34795
6.452 0.98811 5.4811e-005 3.8183 0.011954 8.4162e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4033 0.48822 0.149 0.017976 11.8906 0.11182 0.00014348 0.77833 0.0085868 0.0095313 0.0014629 0.98594 0.99105 3.1649e-006 1.266e-005 0.15854 0.78579 0.84566 0.0014371 0.90952 0.42588 0.0019346 0.42098 1.7324 1.7302 16.0146 144.9333 0.00027319 -85.3291 0.34895
6.453 0.98811 5.4811e-005 3.8183 0.011954 8.4174e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4034 0.48827 0.14902 0.017977 11.893 0.11182 0.00014349 0.77832 0.0085873 0.0095318 0.0014624 0.98595 0.99105 3.1636e-006 1.2654e-005 0.15854 0.78641 0.846 0.0014368 0.91007 0.42607 0.0019342 0.42099 1.7338 1.7316 16.0147 144.9333 0.00027266 -85.3315 0.34995
6.454 0.98811 5.4811e-005 3.8183 0.011954 8.4187e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4035 0.48831 0.14903 0.017978 11.8955 0.11183 0.0001435 0.77831 0.0085878 0.0095324 0.0014619 0.98596 0.99106 3.1622e-006 1.2649e-005 0.15855 0.78702 0.84635 0.0014365 0.91062 0.42627 0.0019338 0.421 1.7351 1.7329 16.0147 144.9333 0.00027214 -85.3339 0.35095
6.455 0.98811 5.4811e-005 3.8183 0.011954 8.42e-005 0.0011654 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4036 0.48836 0.14905 0.01798 11.8979 0.11184 0.00014351 0.7783 0.0085883 0.0095329 0.0014613 0.98597 0.99106 3.1609e-006 1.2644e-005 0.15855 0.78764 0.84669 0.0014362 0.91116 0.42647 0.0019334 0.42102 1.7364 1.7342 16.0147 144.9333 0.00027161 -85.3362 0.35195
6.456 0.98811 5.4811e-005 3.8183 0.011954 8.4213e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4037 0.48841 0.14906 0.017981 11.9003 0.11185 0.00014352 0.7783 0.0085888 0.0095335 0.0014608 0.98597 0.99107 3.1596e-006 1.2639e-005 0.15855 0.78825 0.84703 0.0014359 0.9117 0.42667 0.001933 0.42103 1.7378 1.7356 16.0147 144.9333 0.0002711 -85.3385 0.35295
6.457 0.98811 5.4811e-005 3.8183 0.011954 8.4226e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4038 0.48845 0.14908 0.017982 11.9027 0.11186 0.00014354 0.77829 0.0085893 0.009534 0.0014602 0.98598 0.99107 3.1583e-006 1.2633e-005 0.15856 0.78886 0.84736 0.0014356 0.91224 0.42687 0.0019326 0.42104 1.7391 1.7369 16.0147 144.9334 0.00027058 -85.3409 0.35395
6.458 0.98811 5.4811e-005 3.8183 0.011954 8.4239e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4038 0.4885 0.14909 0.017983 11.9051 0.11186 0.00014355 0.77828 0.0085898 0.0095345 0.0014597 0.98599 0.99108 3.157e-006 1.2628e-005 0.15856 0.78946 0.8477 0.0014353 0.91278 0.42706 0.0019323 0.42105 1.7404 1.7382 16.0147 144.9334 0.00027006 -85.3432 0.35495
6.459 0.98811 5.4811e-005 3.8183 0.011954 8.4252e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4039 0.48854 0.14911 0.017985 11.9075 0.11187 0.00014356 0.77827 0.0085903 0.0095351 0.0014591 0.986 0.99108 3.1558e-006 1.2623e-005 0.15857 0.79007 0.84803 0.0014351 0.91331 0.42726 0.0019319 0.42107 1.7417 1.7396 16.0147 144.9334 0.00026955 -85.3454 0.35595
6.46 0.98811 5.4811e-005 3.8183 0.011954 8.4265e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.404 0.48859 0.14912 0.017986 11.91 0.11188 0.00014357 0.77826 0.0085908 0.0095356 0.0014586 0.986 0.99109 3.1545e-006 1.2618e-005 0.15857 0.79067 0.84837 0.0014348 0.91384 0.42746 0.0019315 0.42108 1.7431 1.7409 16.0147 144.9334 0.00026904 -85.3477 0.35695
6.461 0.98811 5.4811e-005 3.8183 0.011954 8.4278e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4041 0.48864 0.14913 0.017987 11.9124 0.11189 0.00014358 0.77826 0.0085913 0.0095362 0.001458 0.98601 0.99109 3.1532e-006 1.2613e-005 0.15857 0.79127 0.8487 0.0014345 0.91436 0.42766 0.0019311 0.42109 1.7444 1.7422 16.0147 144.9334 0.00026854 -85.35 0.35795
6.462 0.98811 5.4811e-005 3.8183 0.011954 8.429e-005 0.0011654 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.4042 0.48868 0.14915 0.017989 11.9148 0.1119 0.00014359 0.77825 0.0085918 0.0095367 0.0014574 0.98602 0.9911 3.152e-006 1.2608e-005 0.15858 0.79187 0.84903 0.0014342 0.91488 0.42785 0.0019308 0.42111 1.7457 1.7435 16.0147 144.9334 0.00026803 -85.3522 0.35895
6.463 0.98811 5.4811e-005 3.8183 0.011954 8.4303e-005 0.0011654 0.23338 0.00065931 0.23403 0.21596 0 0.032275 0.0389 0 1.4043 0.48873 0.14916 0.01799 11.9172 0.1119 0.00014361 0.77824 0.0085923 0.0095372 0.0014569 0.98603 0.9911 3.1508e-006 1.2603e-005 0.15858 0.79247 0.84936 0.0014339 0.9154 0.42805 0.0019304 0.42112 1.747 1.7448 16.0147 144.9335 0.00026753 -85.3544 0.35995
6.464 0.98811 5.4811e-005 3.8183 0.011954 8.4316e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4044 0.48877 0.14918 0.017991 11.9196 0.11191 0.00014362 0.77823 0.0085928 0.0095378 0.0014563 0.98603 0.99111 3.1495e-006 1.2598e-005 0.15859 0.79306 0.84968 0.0014337 0.91592 0.42825 0.00193 0.42113 1.7483 1.7462 16.0148 144.9335 0.00026703 -85.3566 0.36095
6.465 0.98811 5.481e-005 3.8183 0.011954 8.4329e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4045 0.48882 0.14919 0.017993 11.922 0.11192 0.00014363 0.77822 0.0085933 0.0095383 0.0014558 0.98604 0.99111 3.1483e-006 1.2593e-005 0.15859 0.79366 0.85001 0.0014334 0.91643 0.42845 0.0019297 0.42114 1.7496 1.7475 16.0148 144.9335 0.00026653 -85.3588 0.36195
6.466 0.98811 5.481e-005 3.8183 0.011954 8.4342e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4046 0.48886 0.14921 0.017994 11.9245 0.11193 0.00014364 0.77822 0.0085938 0.0095388 0.0014552 0.98605 0.99112 3.1471e-006 1.2588e-005 0.15859 0.79425 0.85033 0.0014331 0.91694 0.42864 0.0019293 0.42116 1.7509 1.7488 16.0148 144.9335 0.00026603 -85.361 0.36295
6.467 0.98811 5.481e-005 3.8183 0.011954 8.4355e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4047 0.48891 0.14922 0.017995 11.9269 0.11194 0.00014365 0.77821 0.0085943 0.0095394 0.0014547 0.98605 0.99112 3.1459e-006 1.2584e-005 0.1586 0.79484 0.85066 0.0014328 0.91745 0.42884 0.001929 0.42117 1.7522 1.7501 16.0148 144.9335 0.00026554 -85.3631 0.36395
6.468 0.98811 5.481e-005 3.8183 0.011954 8.4368e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4048 0.48896 0.14924 0.017997 11.9293 0.11194 0.00014366 0.7782 0.0085948 0.0095399 0.0014542 0.98606 0.99113 3.1447e-006 1.2579e-005 0.1586 0.79543 0.85098 0.0014326 0.91795 0.42904 0.0019286 0.42118 1.7535 1.7514 16.0148 144.9336 0.00026504 -85.3653 0.36495
6.469 0.98811 5.481e-005 3.8183 0.011954 8.4381e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4049 0.489 0.14925 0.017998 11.9317 0.11195 0.00014368 0.77819 0.0085953 0.0095405 0.0014536 0.98607 0.99113 3.1435e-006 1.2574e-005 0.1586 0.79601 0.8513 0.0014323 0.91845 0.42923 0.0019283 0.4212 1.7547 1.7526 16.0148 144.9336 0.00026455 -85.3674 0.36595
6.47 0.98811 5.481e-005 3.8183 0.011954 8.4394e-005 0.0011654 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4049 0.48905 0.14927 0.017999 11.9341 0.11196 0.00014369 0.77818 0.0085958 0.009541 0.0014531 0.98607 0.99114 3.1424e-006 1.257e-005 0.15861 0.7966 0.85161 0.001432 0.91895 0.42943 0.0019279 0.42121 1.756 1.7539 16.0148 144.9336 0.00026407 -85.3695 0.36695
6.471 0.98811 5.481e-005 3.8183 0.011954 8.4407e-005 0.0011654 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.405 0.48909 0.14928 0.018 11.9366 0.11197 0.0001437 0.77818 0.0085963 0.0095415 0.0014526 0.98608 0.99114 3.1412e-006 1.2565e-005 0.15861 0.79718 0.85193 0.0014318 0.91944 0.42963 0.0019276 0.42122 1.7573 1.7552 16.0148 144.9336 0.00026358 -85.3716 0.36795
6.472 0.98811 5.481e-005 3.8183 0.011954 8.4419e-005 0.0011654 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4051 0.48914 0.1493 0.018002 11.939 0.11198 0.00014371 0.77817 0.0085968 0.0095421 0.0014521 0.98609 0.99114 3.1401e-006 1.256e-005 0.15862 0.79776 0.85225 0.0014315 0.91994 0.42983 0.0019273 0.42123 1.7586 1.7565 16.0148 144.9336 0.0002631 -85.3737 0.36895
6.473 0.98811 5.481e-005 3.8183 0.011954 8.4432e-005 0.0011654 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4052 0.48919 0.14931 0.018003 11.9414 0.11198 0.00014372 0.77816 0.0085973 0.0095426 0.0014516 0.98609 0.99115 3.1389e-006 1.2556e-005 0.15862 0.79834 0.85256 0.0014313 0.92042 0.43002 0.0019269 0.42125 1.7598 1.7578 16.0148 144.9336 0.00026262 -85.3757 0.36995
6.474 0.98811 5.481e-005 3.8183 0.011954 8.4445e-005 0.0011655 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4053 0.48923 0.14933 0.018004 11.9438 0.11199 0.00014373 0.77815 0.0085978 0.0095431 0.0014511 0.9861 0.99115 3.1378e-006 1.2551e-005 0.15862 0.79892 0.85287 0.001431 0.92091 0.43022 0.0019266 0.42126 1.7611 1.759 16.0148 144.9337 0.00026214 -85.3778 0.37095
6.475 0.98811 5.481e-005 3.8183 0.011954 8.4458e-005 0.0011655 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4054 0.48928 0.14934 0.018006 11.9462 0.112 0.00014375 0.77814 0.0085983 0.0095437 0.0014506 0.98611 0.99116 3.1366e-006 1.2547e-005 0.15863 0.7995 0.85318 0.0014307 0.92139 0.43042 0.0019262 0.42127 1.7624 1.7603 16.0148 144.9337 0.00026166 -85.3798 0.37195
6.476 0.98811 5.481e-005 3.8183 0.011954 8.4471e-005 0.0011655 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4055 0.48932 0.14935 0.018007 11.9487 0.11201 0.00014376 0.77814 0.0085988 0.0095442 0.0014501 0.98611 0.99116 3.1355e-006 1.2542e-005 0.15863 0.80007 0.85349 0.0014305 0.92187 0.43061 0.0019259 0.42129 1.7636 1.7616 16.0148 144.9337 0.00026119 -85.3818 0.37295
6.477 0.98811 5.481e-005 3.8183 0.011954 8.4484e-005 0.0011655 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4056 0.48937 0.14937 0.018008 11.9511 0.11201 0.00014377 0.77813 0.0085993 0.0095448 0.0014497 0.98612 0.99117 3.1344e-006 1.2538e-005 0.15864 0.80064 0.8538 0.0014302 0.92235 0.43081 0.0019256 0.4213 1.7649 1.7628 16.0149 144.9337 0.00026071 -85.3838 0.37395
6.478 0.98811 5.4809e-005 3.8183 0.011954 8.4497e-005 0.0011655 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.4057 0.48942 0.14938 0.01801 11.9535 0.11202 0.00014378 0.77812 0.0085998 0.0095453 0.0014492 0.98613 0.99117 3.1333e-006 1.2533e-005 0.15864 0.80121 0.85411 0.00143 0.92282 0.43101 0.0019253 0.42131 1.7661 1.7641 16.0149 144.9337 0.00026024 -85.3858 0.37495
6.479 0.98811 5.4809e-005 3.8183 0.011954 8.451e-005 0.0011655 0.23339 0.00065931 0.23405 0.21596 0 0.032275 0.0389 0 1.4058 0.48946 0.1494 0.018011 11.9559 0.11203 0.00014379 0.77811 0.0086003 0.0095458 0.0014487 0.98613 0.99117 3.1322e-006 1.2529e-005 0.15864 0.80178 0.85441 0.0014297 0.92329 0.4312 0.0019249 0.42133 1.7674 1.7654 16.0149 144.9338 0.00025977 -85.3878 0.37595
6.48 0.98811 5.4809e-005 3.8183 0.011954 8.4523e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032275 0.0389 0 1.4059 0.48951 0.14941 0.018012 11.9584 0.11204 0.0001438 0.77811 0.0086008 0.0095464 0.0014483 0.98614 0.99118 3.1311e-006 1.2524e-005 0.15865 0.80235 0.85472 0.0014295 0.92376 0.4314 0.0019246 0.42134 1.7686 1.7666 16.0149 144.9338 0.00025931 -85.3898 0.37695
6.481 0.98811 5.4809e-005 3.8183 0.011954 8.4536e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032275 0.0389 0 1.406 0.48955 0.14943 0.018014 11.9608 0.11205 0.00014382 0.7781 0.0086013 0.0095469 0.0014478 0.98614 0.99118 3.13e-006 1.252e-005 0.15865 0.80291 0.85502 0.0014293 0.92423 0.4316 0.0019243 0.42135 1.7699 1.7679 16.0149 144.9338 0.00025884 -85.3917 0.37795
6.482 0.98811 5.4809e-005 3.8183 0.011954 8.4548e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.406 0.4896 0.14944 0.018015 11.9632 0.11205 0.00014383 0.77809 0.0086018 0.0095474 0.0014474 0.98615 0.99119 3.129e-006 1.2516e-005 0.15866 0.80347 0.85532 0.001429 0.92469 0.43179 0.001924 0.42137 1.7711 1.7691 16.0149 144.9338 0.00025838 -85.3936 0.37895
6.483 0.98811 5.4809e-005 3.8183 0.011954 8.4561e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4061 0.48965 0.14946 0.018016 11.9656 0.11206 0.00014384 0.77808 0.0086023 0.009548 0.0014469 0.98616 0.99119 3.1279e-006 1.2512e-005 0.15866 0.80404 0.85562 0.0014288 0.92515 0.43199 0.0019237 0.42138 1.7723 1.7704 16.0149 144.9338 0.00025792 -85.3956 0.37995
6.484 0.98811 5.4809e-005 3.8183 0.011954 8.4574e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4062 0.48969 0.14947 0.018017 11.9681 0.11207 0.00014385 0.77807 0.0086028 0.0095485 0.0014464 0.98616 0.99119 3.1269e-006 1.2507e-005 0.15866 0.8046 0.85592 0.0014285 0.9256 0.43218 0.0019234 0.42139 1.7736 1.7716 16.0149 144.9339 0.00025746 -85.3975 0.38095
6.485 0.98811 5.4809e-005 3.8183 0.011954 8.4587e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4063 0.48974 0.14949 0.018019 11.9705 0.11208 0.00014386 0.77807 0.0086033 0.009549 0.001446 0.98617 0.9912 3.1258e-006 1.2503e-005 0.15867 0.80515 0.85621 0.0014283 0.92606 0.43238 0.001923 0.42141 1.7748 1.7728 16.0149 144.9339 0.00025701 -85.3993 0.38195
6.486 0.98811 5.4809e-005 3.8183 0.011954 8.46e-005 0.0011655 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4064 0.48978 0.1495 0.01802 11.9729 0.11209 0.00014387 0.77806 0.0086038 0.0095496 0.0014455 0.98617 0.9912 3.1248e-006 1.2499e-005 0.15867 0.80571 0.85651 0.0014281 0.92651 0.43258 0.0019227 0.42142 1.776 1.7741 16.0149 144.9339 0.00025655 -85.4012 0.38295
6.487 0.98811 5.4809e-005 3.8183 0.011954 8.4613e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4065 0.48983 0.14952 0.018021 11.9753 0.11209 0.00014389 0.77805 0.0086043 0.0095501 0.0014451 0.98618 0.99121 3.1237e-006 1.2495e-005 0.15868 0.80626 0.8568 0.0014278 0.92696 0.43277 0.0019224 0.42143 1.7773 1.7753 16.0149 144.9339 0.0002561 -85.4031 0.38395
6.488 0.98811 5.4809e-005 3.8183 0.011954 8.4626e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4066 0.48988 0.14953 0.018023 11.9778 0.1121 0.0001439 0.77804 0.0086048 0.0095507 0.0014446 0.98619 0.99121 3.1227e-006 1.2491e-005 0.15868 0.80682 0.8571 0.0014276 0.9274 0.43297 0.0019221 0.42145 1.7785 1.7765 16.0149 144.9339 0.00025565 -85.4049 0.38495
6.489 0.98811 5.4809e-005 3.8183 0.011954 8.4639e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4067 0.48992 0.14954 0.018024 11.9802 0.11211 0.00014391 0.77803 0.0086053 0.0095512 0.0014441 0.98619 0.99121 3.1217e-006 1.2487e-005 0.15868 0.80737 0.85739 0.0014274 0.92784 0.43317 0.0019218 0.42146 1.7797 1.7777 16.0149 144.9339 0.0002552 -85.4068 0.38595
6.49 0.98811 5.4809e-005 3.8183 0.011954 8.4652e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4068 0.48997 0.14956 0.018025 11.9826 0.11212 0.00014392 0.77803 0.0086058 0.0095517 0.0014437 0.9862 0.99122 3.1207e-006 1.2483e-005 0.15869 0.80792 0.85768 0.0014271 0.92828 0.43336 0.0019215 0.42147 1.7809 1.779 16.0149 144.934 0.00025475 -85.4086 0.38695
6.491 0.98811 5.4808e-005 3.8183 0.011954 8.4664e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4069 0.49001 0.14957 0.018027 11.985 0.11213 0.00014393 0.77802 0.0086063 0.0095523 0.0014432 0.9862 0.99122 3.1197e-006 1.2479e-005 0.15869 0.80847 0.85797 0.0014269 0.92872 0.43356 0.0019212 0.42148 1.7821 1.7802 16.0149 144.934 0.00025431 -85.4104 0.38795
6.492 0.98811 5.4808e-005 3.8183 0.011954 8.4677e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.407 0.49006 0.14959 0.018028 11.9875 0.11213 0.00014394 0.77801 0.0086068 0.0095528 0.0014428 0.98621 0.99122 3.1187e-006 1.2475e-005 0.15869 0.80901 0.85826 0.0014267 0.92916 0.43375 0.0019209 0.4215 1.7833 1.7814 16.0149 144.934 0.00025387 -85.4122 0.38895
6.493 0.98811 5.4808e-005 3.8183 0.011954 8.469e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.407 0.49011 0.1496 0.018029 11.9899 0.11214 0.00014396 0.778 0.0086073 0.0095533 0.0014423 0.98621 0.99123 3.1177e-006 1.2471e-005 0.1587 0.80956 0.85854 0.0014265 0.92959 0.43395 0.0019207 0.42151 1.7845 1.7826 16.0149 144.934 0.00025342 -85.414 0.38995
6.494 0.98811 5.4808e-005 3.8183 0.011954 8.4703e-005 0.0011655 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.4071 0.49015 0.14962 0.01803 11.9923 0.11215 0.00014397 0.77799 0.0086078 0.0095539 0.0014419 0.98622 0.99123 3.1167e-006 1.2467e-005 0.1587 0.8101 0.85883 0.0014262 0.93002 0.43414 0.0019204 0.42152 1.7857 1.7838 16.0149 144.934 0.00025299 -85.4158 0.39095
6.495 0.98811 5.4808e-005 3.8183 0.011954 8.4716e-005 0.0011655 0.2334 0.00065931 0.23406 0.21597 0 0.032274 0.0389 0 1.4072 0.4902 0.14963 0.018032 11.9948 0.11216 0.00014398 0.77799 0.0086083 0.0095544 0.0014415 0.98623 0.99124 3.1158e-006 1.2463e-005 0.15871 0.81064 0.85911 0.001426 0.93044 0.43434 0.0019201 0.42154 1.7869 1.785 16.0149 144.9341 0.00025255 -85.4175 0.39195
6.496 0.98811 5.4808e-005 3.8183 0.011954 8.4729e-005 0.0011655 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4073 0.49024 0.14965 0.018033 11.9972 0.11217 0.00014399 0.77798 0.0086088 0.0095549 0.0014411 0.98623 0.99124 3.1148e-006 1.2459e-005 0.15871 0.81118 0.85939 0.0014258 0.93087 0.43454 0.0019198 0.42155 1.7881 1.7862 16.0149 144.9341 0.00025211 -85.4193 0.39295
6.497 0.98811 5.4808e-005 3.8183 0.011954 8.4742e-005 0.0011655 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4074 0.49029 0.14966 0.018034 11.9996 0.11217 0.000144 0.77797 0.0086093 0.0095555 0.0014407 0.98624 0.99124 3.1138e-006 1.2455e-005 0.15871 0.81172 0.85968 0.0014256 0.93129 0.43473 0.0019195 0.42157 1.7893 1.7874 16.0149 144.9341 0.00025168 -85.421 0.39395
6.498 0.98811 5.4808e-005 3.8183 0.011954 8.4755e-005 0.0011655 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4075 0.49034 0.14968 0.018036 12.002 0.11218 0.00014401 0.77796 0.0086098 0.009556 0.0014403 0.98624 0.99125 3.1129e-006 1.2452e-005 0.15872 0.81225 0.85996 0.0014254 0.93171 0.43493 0.0019192 0.42158 1.7905 1.7886 16.0149 144.9341 0.00025125 -85.4227 0.39495
6.499 0.98811 5.4808e-005 3.8183 0.011954 8.4768e-005 0.0011655 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4076 0.49038 0.14969 0.018037 12.0045 0.11219 0.00014402 0.77796 0.0086103 0.0095565 0.0014399 0.98625 0.99125 3.112e-006 1.2448e-005 0.15872 0.81279 0.86023 0.0014252 0.93212 0.43512 0.001919 0.42159 1.7917 1.7898 16.015 144.9341 0.00025082 -85.4244 0.39595
6.5 0.98811 5.4808e-005 3.8183 0.011954 8.4781e-005 0.0011656 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4077 0.49043 0.14971 0.018038 12.0069 0.1122 0.00014404 0.77795 0.0086108 0.0095571 0.0014395 0.98625 0.99125 3.111e-006 1.2444e-005 0.15873 0.81332 0.86051 0.001425 0.93254 0.43532 0.0019187 0.42161 1.7928 1.791 16.015 144.9342 0.00025039 -85.4261 0.39695
6.501 0.98811 5.4808e-005 3.8183 0.011954 8.4793e-005 0.0011656 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4078 0.49047 0.14972 0.01804 12.0093 0.1122 0.00014405 0.77794 0.0086113 0.0095576 0.0014391 0.98626 0.99126 3.1101e-006 1.244e-005 0.15873 0.81385 0.86079 0.0014248 0.93295 0.43551 0.0019184 0.42162 1.794 1.7921 16.015 144.9342 0.00024997 -85.4278 0.39795
6.502 0.98811 5.4808e-005 3.8183 0.011954 8.4806e-005 0.0011656 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4079 0.49052 0.14974 0.018041 12.0118 0.11221 0.00014406 0.77793 0.0086118 0.0095581 0.0014387 0.98626 0.99126 3.1092e-006 1.2437e-005 0.15873 0.81438 0.86106 0.0014246 0.93336 0.43571 0.0019181 0.42163 1.7952 1.7933 16.015 144.9342 0.00024954 -85.4295 0.39895
6.503 0.98811 5.4808e-005 3.8183 0.011954 8.4819e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.408 0.49056 0.14975 0.018042 12.0142 0.11222 0.00014407 0.77792 0.0086123 0.0095587 0.0014384 0.98627 0.99126 3.1083e-006 1.2433e-005 0.15874 0.81491 0.86134 0.0014243 0.93376 0.4359 0.0019179 0.42165 1.7964 1.7945 16.015 144.9342 0.00024912 -85.4311 0.39995
6.504 0.98811 5.4807e-005 3.8183 0.011954 8.4832e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4081 0.49061 0.14976 0.018044 12.0166 0.11223 0.00014408 0.77792 0.0086128 0.0095592 0.001438 0.98627 0.99127 3.1074e-006 1.2429e-005 0.15874 0.81543 0.86161 0.0014241 0.93417 0.4361 0.0019176 0.42166 1.7975 1.7957 16.015 144.9342 0.0002487 -85.4328 0.40095
6.505 0.98811 5.4807e-005 3.8183 0.011954 8.4845e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4081 0.49066 0.14978 0.018045 12.0191 0.11224 0.00014409 0.77791 0.0086132 0.0095597 0.0014376 0.98628 0.99127 3.1065e-006 1.2426e-005 0.15874 0.81596 0.86188 0.0014239 0.93457 0.43629 0.0019173 0.42167 1.7987 1.7968 16.015 144.9342 0.00024828 -85.4344 0.40195
6.506 0.98811 5.4807e-005 3.8183 0.011954 8.4858e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4082 0.4907 0.14979 0.018046 12.0215 0.11224 0.00014411 0.7779 0.0086137 0.0095603 0.0014372 0.98628 0.99127 3.1056e-006 1.2422e-005 0.15875 0.81648 0.86215 0.0014237 0.93496 0.43649 0.0019171 0.42169 1.7998 1.798 16.015 144.9343 0.00024787 -85.436 0.40295
6.507 0.98811 5.4807e-005 3.8183 0.011954 8.4871e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4083 0.49075 0.14981 0.018047 12.0239 0.11225 0.00014412 0.77789 0.0086142 0.0095608 0.0014368 0.98629 0.99128 3.1047e-006 1.2419e-005 0.15875 0.817 0.86242 0.0014235 0.93536 0.43668 0.0019168 0.4217 1.801 1.7992 16.015 144.9343 0.00024745 -85.4377 0.40395
6.508 0.98811 5.4807e-005 3.8183 0.011954 8.4884e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4084 0.49079 0.14982 0.018049 12.0264 0.11226 0.00014413 0.77788 0.0086147 0.0095614 0.0014364 0.98629 0.99128 3.1038e-006 1.2415e-005 0.15876 0.81752 0.86269 0.0014233 0.93575 0.43688 0.0019165 0.42171 1.8022 1.8003 16.015 144.9343 0.00024704 -85.4393 0.40495
6.509 0.98811 5.4807e-005 3.8183 0.011954 8.4897e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4085 0.49084 0.14984 0.01805 12.0288 0.11227 0.00014414 0.77788 0.0086152 0.0095619 0.001436 0.9863 0.99128 3.1029e-006 1.2412e-005 0.15876 0.81804 0.86296 0.0014231 0.93614 0.43707 0.0019163 0.42173 1.8033 1.8015 16.015 144.9343 0.00024663 -85.4409 0.40595
6.51 0.98811 5.4807e-005 3.8183 0.011953 8.4909e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4086 0.49089 0.14985 0.018051 12.0312 0.11228 0.00014415 0.77787 0.0086157 0.0095624 0.0014356 0.9863 0.99129 3.1021e-006 1.2408e-005 0.15876 0.81855 0.86322 0.0014229 0.93653 0.43727 0.001916 0.42174 1.8045 1.8026 16.015 144.9343 0.00024622 -85.4424 0.40695
6.511 0.98811 5.4807e-005 3.8183 0.011953 8.4922e-005 0.0011656 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.4087 0.49093 0.14987 0.018053 12.0337 0.11228 0.00014416 0.77786 0.0086162 0.009563 0.0014352 0.98631 0.99129 3.1012e-006 1.2405e-005 0.15877 0.81907 0.86349 0.0014227 0.93692 0.43746 0.0019158 0.42175 1.8056 1.8038 16.015 144.9344 0.00024581 -85.444 0.40795
6.512 0.98811 5.4807e-005 3.8183 0.011953 8.4935e-005 0.0011656 0.23341 0.00065931 0.23407 0.21598 0 0.032274 0.0389 0 1.4088 0.49098 0.14988 0.018054 12.0361 0.11229 0.00014418 0.77785 0.0086167 0.0095635 0.0014348 0.98631 0.99129 3.1003e-006 1.2401e-005 0.15877 0.81958 0.86375 0.0014225 0.9373 0.43766 0.0019155 0.42177 1.8067 1.8049 16.015 144.9344 0.0002454 -85.4456 0.40895
6.513 0.98811 5.4807e-005 3.8183 0.011953 8.4948e-005 0.0011656 0.23341 0.00065931 0.23407 0.21599 0 0.032274 0.0389 0 1.4089 0.49102 0.1499 0.018055 12.0385 0.1123 0.00014419 0.77784 0.0086172 0.009564 0.0014344 0.98632 0.9913 3.0995e-006 1.2398e-005 0.15878 0.82009 0.86401 0.0014223 0.93768 0.43785 0.0019153 0.42178 1.8079 1.8061 16.015 144.9344 0.000245 -85.4471 0.40995
6.514 0.98811 5.4807e-005 3.8183 0.011953 8.4961e-005 0.0011656 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.409 0.49107 0.14991 0.018057 12.041 0.11231 0.0001442 0.77784 0.0086177 0.0095646 0.001434 0.98632 0.9913 3.0987e-006 1.2395e-005 0.15878 0.8206 0.86427 0.0014221 0.93806 0.43805 0.001915 0.42179 1.809 1.8072 16.015 144.9344 0.0002446 -85.4486 0.41095
6.515 0.98811 5.4807e-005 3.8183 0.011953 8.4974e-005 0.0011656 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4091 0.49112 0.14993 0.018058 12.0434 0.11232 0.00014421 0.77783 0.0086182 0.0095651 0.0014336 0.98633 0.9913 3.0978e-006 1.2391e-005 0.15878 0.82111 0.86453 0.0014219 0.93844 0.43824 0.0019148 0.42181 1.8101 1.8084 16.015 144.9344 0.0002442 -85.4502 0.41195
6.516 0.98811 5.4806e-005 3.8183 0.011953 8.4987e-005 0.0011656 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4092 0.49116 0.14994 0.018059 12.0458 0.11232 0.00014422 0.77782 0.0086187 0.0095656 0.0014332 0.98633 0.99131 3.097e-006 1.2388e-005 0.15879 0.82162 0.86479 0.0014218 0.93881 0.43844 0.0019145 0.42182 1.8113 1.8095 16.015 144.9345 0.0002438 -85.4517 0.41295
6.517 0.98811 5.4806e-005 3.8183 0.011953 8.5e-005 0.0011656 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4092 0.49121 0.14995 0.01806 12.0483 0.11233 0.00014423 0.77781 0.0086192 0.0095662 0.0014329 0.98634 0.99131 3.0962e-006 1.2385e-005 0.15879 0.82212 0.86505 0.0014216 0.93919 0.43863 0.0019143 0.42184 1.8124 1.8106 16.015 144.9345 0.0002434 -85.4532 0.41395
6.518 0.98811 5.4806e-005 3.8183 0.011953 8.5013e-005 0.0011656 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4093 0.49125 0.14997 0.018062 12.0507 0.11234 0.00014424 0.77781 0.0086197 0.0095667 0.0014325 0.98634 0.99131 3.0954e-006 1.2381e-005 0.1588 0.82263 0.86531 0.0014214 0.93956 0.43882 0.001914 0.42185 1.8135 1.8117 16.015 144.9345 0.000243 -85.4547 0.41495
6.519 0.98811 5.4806e-005 3.8183 0.011953 8.5026e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4094 0.4913 0.14998 0.018063 12.0531 0.11235 0.00014426 0.7778 0.0086202 0.0095672 0.0014322 0.98635 0.99132 3.0946e-006 1.2378e-005 0.1588 0.82313 0.86556 0.0014212 0.93992 0.43902 0.0019138 0.42186 1.8146 1.8129 16.015 144.9345 0.00024261 -85.4561 0.41595
6.52 0.98811 5.4806e-005 3.8183 0.011953 8.5038e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4095 0.49135 0.15 0.018064 12.0556 0.11235 0.00014427 0.77779 0.0086207 0.0095678 0.0014319 0.98635 0.99132 3.0937e-006 1.2375e-005 0.1588 0.82363 0.86582 0.001421 0.94029 0.43921 0.0019136 0.42188 1.8158 1.814 16.015 144.9345 0.00024222 -85.4576 0.41695
6.521 0.98811 5.4806e-005 3.8183 0.011953 8.5051e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4096 0.49139 0.15001 0.018066 12.058 0.11236 0.00014428 0.77778 0.0086212 0.0095683 0.0014315 0.98636 0.99132 3.093e-006 1.2372e-005 0.15881 0.82413 0.86607 0.0014208 0.94065 0.43941 0.0019133 0.42189 1.8169 1.8151 16.015 144.9345 0.00024183 -85.4591 0.41795
6.522 0.98811 5.4806e-005 3.8183 0.011953 8.5064e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4097 0.49144 0.15003 0.018067 12.0605 0.11237 0.00014429 0.77777 0.0086217 0.0095688 0.0014312 0.98636 0.99132 3.0922e-006 1.2369e-005 0.15881 0.82462 0.86632 0.0014207 0.94101 0.4396 0.0019131 0.4219 1.818 1.8162 16.015 144.9346 0.00024144 -85.4605 0.41895
6.523 0.98811 5.4806e-005 3.8183 0.011953 8.5077e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4098 0.49148 0.15004 0.018068 12.0629 0.11238 0.0001443 0.77777 0.0086222 0.0095694 0.0014309 0.98636 0.99133 3.0914e-006 1.2365e-005 0.15881 0.82512 0.86657 0.0014205 0.94137 0.4398 0.0019128 0.42192 1.8191 1.8173 16.015 144.9346 0.00024105 -85.4619 0.41995
6.524 0.98811 5.4806e-005 3.8183 0.011953 8.509e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4099 0.49153 0.15006 0.01807 12.0653 0.11239 0.00014431 0.77776 0.0086227 0.0095699 0.0014306 0.98637 0.99133 3.0906e-006 1.2362e-005 0.15882 0.82561 0.86682 0.0014203 0.94173 0.43999 0.0019126 0.42193 1.8202 1.8185 16.015 144.9346 0.00024067 -85.4634 0.42095
6.525 0.98811 5.4806e-005 3.8183 0.011953 8.5103e-005 0.0011656 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.41 0.49158 0.15007 0.018071 12.0678 0.11239 0.00014433 0.77775 0.0086232 0.0095704 0.0014303 0.98637 0.99133 3.0898e-006 1.2359e-005 0.15882 0.82611 0.86707 0.0014201 0.94208 0.44018 0.0019124 0.42195 1.8213 1.8196 16.015 144.9346 0.00024028 -85.4648 0.42195
6.526 0.98811 5.4806e-005 3.8183 0.011953 8.5116e-005 0.0011657 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4101 0.49162 0.15009 0.018072 12.0702 0.1124 0.00014434 0.77774 0.0086237 0.0095709 0.00143 0.98638 0.99134 3.0891e-006 1.2356e-005 0.15883 0.8266 0.86732 0.00142 0.94243 0.44038 0.0019122 0.42196 1.8224 1.8207 16.015 144.9346 0.0002399 -85.4662 0.42295
6.527 0.98811 5.4806e-005 3.8183 0.011953 8.5129e-005 0.0011657 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.4102 0.49167 0.1501 0.018073 12.0727 0.11241 0.00014435 0.77773 0.0086242 0.0095715 0.0014296 0.98638 0.99134 3.0883e-006 1.2353e-005 0.15883 0.82709 0.86757 0.0014198 0.94278 0.44057 0.0019119 0.42197 1.8235 1.8218 16.015 144.9347 0.00023952 -85.4676 0.42395
6.528 0.98811 5.4806e-005 3.8183 0.011953 8.5142e-005 0.0011657 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.4102 0.49171 0.15012 0.018075 12.0751 0.11242 0.00014436 0.77773 0.0086247 0.009572 0.0014293 0.98639 0.99134 3.0875e-006 1.235e-005 0.15883 0.82757 0.86781 0.0014196 0.94313 0.44077 0.0019117 0.42199 1.8246 1.8229 16.015 144.9347 0.00023914 -85.469 0.42495
6.529 0.98811 5.4805e-005 3.8183 0.011953 8.5154e-005 0.0011657 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.4103 0.49176 0.15013 0.018076 12.0775 0.11243 0.00014437 0.77772 0.0086252 0.0095725 0.001429 0.98639 0.99134 3.0868e-006 1.2347e-005 0.15884 0.82806 0.86806 0.0014195 0.94348 0.44096 0.0019115 0.422 1.8257 1.824 16.015 144.9347 0.00023876 -85.4704 0.42595
6.53 0.98811 5.4805e-005 3.8183 0.011953 8.5167e-005 0.0011657 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.4104 0.4918 0.15014 0.018077 12.08 0.11243 0.00014438 0.77771 0.0086257 0.0095731 0.0014287 0.9864 0.99135 3.086e-006 1.2344e-005 0.15884 0.82855 0.8683 0.0014193 0.94382 0.44115 0.0019113 0.42201 1.8268 1.825 16.015 144.9347 0.00023839 -85.4717 0.42695
6.531 0.98811 5.4805e-005 3.8183 0.011953 8.518e-005 0.0011657 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4105 0.49185 0.15016 0.018079 12.0824 0.11244 0.0001444 0.7777 0.0086262 0.0095736 0.0014283 0.9864 0.99135 3.0853e-006 1.2341e-005 0.15885 0.82903 0.86855 0.0014191 0.94416 0.44135 0.001911 0.42203 1.8278 1.8261 16.015 144.9347 0.00023801 -85.4731 0.42795
6.532 0.98811 5.4805e-005 3.8183 0.011953 8.5193e-005 0.0011657 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4106 0.4919 0.15017 0.01808 12.0849 0.11245 0.00014441 0.7777 0.0086267 0.0095741 0.001428 0.9864 0.99135 3.0845e-006 1.2338e-005 0.15885 0.82951 0.86879 0.001419 0.9445 0.44154 0.0019108 0.42204 1.8289 1.8272 16.015 144.9348 0.00023764 -85.4744 0.42895
6.533 0.98811 5.4805e-005 3.8183 0.011953 8.5206e-005 0.0011657 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4107 0.49194 0.15019 0.018081 12.0873 0.11246 0.00014442 0.77769 0.0086271 0.0095747 0.0014277 0.98641 0.99136 3.0838e-006 1.2335e-005 0.15885 0.82999 0.86903 0.0014188 0.94483 0.44173 0.0019106 0.42206 1.83 1.8283 16.015 144.9348 0.00023727 -85.4758 0.42995
6.534 0.98811 5.4805e-005 3.8183 0.011953 8.5219e-005 0.0011657 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4108 0.49199 0.1502 0.018083 12.0897 0.11246 0.00014443 0.77768 0.0086276 0.0095752 0.0014273 0.98641 0.99136 3.0831e-006 1.2332e-005 0.15886 0.83047 0.86927 0.0014186 0.94517 0.44193 0.0019104 0.42207 1.8311 1.8294 16.015 144.9348 0.0002369 -85.4771 0.43095
6.535 0.98811 5.4805e-005 3.8183 0.011953 8.5232e-005 0.0011657 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4109 0.49203 0.15022 0.018084 12.0922 0.11247 0.00014444 0.77767 0.0086281 0.0095757 0.001427 0.98642 0.99136 3.0824e-006 1.2329e-005 0.15886 0.83095 0.86951 0.0014185 0.9455 0.44212 0.0019102 0.42208 1.8321 1.8305 16.015 144.9348 0.00023653 -85.4784 0.43195
6.536 0.98811 5.4805e-005 3.8183 0.011953 8.5245e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.411 0.49208 0.15023 0.018085 12.0946 0.11248 0.00014445 0.77766 0.0086286 0.0095763 0.0014267 0.98642 0.99136 3.0817e-006 1.2327e-005 0.15887 0.83143 0.86974 0.0014183 0.94583 0.44231 0.00191 0.4221 1.8332 1.8315 16.0149 144.9348 0.00023616 -85.4797 0.43295
6.537 0.98811 5.4805e-005 3.8183 0.011953 8.5258e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4111 0.49213 0.15025 0.018086 12.0971 0.11249 0.00014446 0.77766 0.0086291 0.0095768 0.0014264 0.98642 0.99137 3.0809e-006 1.2324e-005 0.15887 0.8319 0.86998 0.0014181 0.94616 0.44251 0.0019097 0.42211 1.8343 1.8326 16.0149 144.9349 0.0002358 -85.481 0.43395
6.538 0.98811 5.4805e-005 3.8183 0.011953 8.5271e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4112 0.49217 0.15026 0.018088 12.0995 0.1125 0.00014448 0.77765 0.0086296 0.0095773 0.001426 0.98643 0.99137 3.0802e-006 1.2321e-005 0.15887 0.83237 0.87022 0.001418 0.94649 0.4427 0.0019095 0.42212 1.8353 1.8337 16.0149 144.9349 0.00023543 -85.4823 0.43495
6.539 0.98811 5.4805e-005 3.8183 0.011953 8.5283e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4113 0.49222 0.15028 0.018089 12.102 0.1125 0.00014449 0.77764 0.0086301 0.0095779 0.0014257 0.98643 0.99137 3.0795e-006 1.2318e-005 0.15888 0.83284 0.87045 0.0014178 0.94681 0.44289 0.0019093 0.42214 1.8364 1.8347 16.0149 144.9349 0.00023507 -85.4836 0.43595
6.54 0.98811 5.4805e-005 3.8183 0.011953 8.5296e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4113 0.49226 0.15029 0.01809 12.1044 0.11251 0.0001445 0.77763 0.0086306 0.0095784 0.0014254 0.98644 0.99137 3.0788e-006 1.2315e-005 0.15888 0.83331 0.87068 0.0014176 0.94713 0.44309 0.0019091 0.42215 1.8375 1.8358 16.0149 144.9349 0.00023471 -85.4849 0.43695
6.541 0.98811 5.4805e-005 3.8183 0.011953 8.5309e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4114 0.49231 0.15031 0.018092 12.1068 0.11252 0.00014451 0.77762 0.0086311 0.0095789 0.0014251 0.98644 0.99138 3.0782e-006 1.2313e-005 0.15888 0.83378 0.87092 0.0014175 0.94745 0.44328 0.0019089 0.42217 1.8385 1.8369 16.0149 144.9349 0.00023435 -85.4861 0.43795
6.542 0.98811 5.4804e-005 3.8183 0.011953 8.5322e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4115 0.49236 0.15032 0.018093 12.1093 0.11253 0.00014452 0.77762 0.0086316 0.0095795 0.0014248 0.98644 0.99138 3.0775e-006 1.231e-005 0.15889 0.83425 0.87115 0.0014173 0.94777 0.44347 0.0019087 0.42218 1.8396 1.8379 16.0149 144.9349 0.000234 -85.4874 0.43895
6.543 0.98811 5.4804e-005 3.8183 0.011953 8.5335e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4116 0.4924 0.15033 0.018094 12.1117 0.11254 0.00014453 0.77761 0.0086321 0.00958 0.0014245 0.98645 0.99138 3.0768e-006 1.2307e-005 0.15889 0.83472 0.87138 0.0014172 0.94809 0.44367 0.0019085 0.42219 1.8406 1.839 16.0149 144.935 0.00023364 -85.4886 0.43995
6.544 0.98811 5.4804e-005 3.8183 0.011953 8.5348e-005 0.0011657 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.4117 0.49245 0.15035 0.018095 12.1142 0.11254 0.00014455 0.7776 0.0086326 0.0095805 0.0014242 0.98645 0.99138 3.0761e-006 1.2304e-005 0.1589 0.83518 0.87161 0.001417 0.9484 0.44386 0.0019083 0.42221 1.8416 1.84 16.0149 144.935 0.00023329 -85.4899 0.44095
6.545 0.98811 5.4804e-005 3.8183 0.011953 8.5361e-005 0.0011657 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.4118 0.49249 0.15036 0.018097 12.1166 0.11255 0.00014456 0.77759 0.0086331 0.0095811 0.0014239 0.98646 0.99139 3.0755e-006 1.2302e-005 0.1589 0.83564 0.87184 0.0014169 0.94871 0.44405 0.0019081 0.42222 1.8427 1.8411 16.0149 144.935 0.00023293 -85.4911 0.44195
6.546 0.98811 5.4804e-005 3.8183 0.011953 8.5374e-005 0.0011657 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.4119 0.49254 0.15038 0.018098 12.1191 0.11256 0.00014457 0.77759 0.0086336 0.0095816 0.0014237 0.98646 0.99139 3.0748e-006 1.2299e-005 0.1589 0.83611 0.87206 0.0014167 0.94902 0.44424 0.0019079 0.42224 1.8437 1.8421 16.0149 144.935 0.00023258 -85.4923 0.44295
6.547 0.98811 5.4804e-005 3.8183 0.011953 8.5387e-005 0.0011657 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.412 0.49259 0.15039 0.018099 12.1215 0.11257 0.00014458 0.77758 0.0086341 0.0095821 0.0014234 0.98646 0.99139 3.0741e-006 1.2297e-005 0.15891 0.83657 0.87229 0.0014166 0.94933 0.44444 0.0019077 0.42225 1.8448 1.8432 16.0149 144.935 0.00023223 -85.4935 0.44395
6.548 0.98811 5.4804e-005 3.8183 0.011953 8.5399e-005 0.0011657 0.23343 0.00065931 0.23409 0.216 0 0.032272 0.0389 0 1.4121 0.49263 0.15041 0.018101 12.124 0.11257 0.00014459 0.77757 0.0086346 0.0095826 0.0014231 0.98647 0.99139 3.0735e-006 1.2294e-005 0.15891 0.83702 0.87252 0.0014164 0.94964 0.44463 0.0019075 0.42226 1.8458 1.8442 16.0149 144.9351 0.00023188 -85.4947 0.44495
6.549 0.98811 5.4804e-005 3.8183 0.011953 8.5412e-005 0.0011657 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4122 0.49268 0.15042 0.018102 12.1264 0.11258 0.0001446 0.77756 0.0086351 0.0095832 0.0014229 0.98647 0.9914 3.0728e-006 1.2291e-005 0.15892 0.83748 0.87274 0.0014163 0.94994 0.44482 0.0019073 0.42228 1.8468 1.8452 16.0149 144.9351 0.00023154 -85.4959 0.44595
6.55 0.98811 5.4804e-005 3.8183 0.011953 8.5425e-005 0.0011657 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4123 0.49272 0.15044 0.018103 12.1289 0.11259 0.00014462 0.77755 0.0086356 0.0095837 0.0014226 0.98647 0.9914 3.0722e-006 1.2289e-005 0.15892 0.83794 0.87296 0.0014161 0.95025 0.44501 0.0019071 0.42229 1.8479 1.8463 16.0149 144.9351 0.00023119 -85.4971 0.44695
6.551 0.98811 5.4804e-005 3.8183 0.011953 8.5438e-005 0.0011658 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4123 0.49277 0.15045 0.018105 12.1313 0.1126 0.00014463 0.77755 0.0086361 0.0095842 0.0014223 0.98648 0.9914 3.0715e-006 1.2286e-005 0.15892 0.83839 0.87319 0.001416 0.95055 0.44521 0.0019069 0.4223 1.8489 1.8473 16.0149 144.9351 0.00023085 -85.4983 0.44795
6.552 0.98811 5.4804e-005 3.8183 0.011953 8.5451e-005 0.0011658 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4124 0.49282 0.15047 0.018106 12.1338 0.11261 0.00014464 0.77754 0.0086365 0.0095848 0.0014221 0.98648 0.9914 3.0709e-006 1.2284e-005 0.15893 0.83884 0.87341 0.0014159 0.95085 0.4454 0.0019068 0.42232 1.8499 1.8483 16.0149 144.9351 0.0002305 -85.4995 0.44895
6.553 0.98811 5.4804e-005 3.8183 0.011953 8.5464e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4125 0.49286 0.15048 0.018107 12.1362 0.11261 0.00014465 0.77753 0.008637 0.0095853 0.0014218 0.98648 0.99141 3.0703e-006 1.2281e-005 0.15893 0.8393 0.87363 0.0014157 0.95114 0.44559 0.0019066 0.42233 1.8509 1.8493 16.0149 144.9352 0.00023016 -85.5006 0.44995
6.554 0.98811 5.4804e-005 3.8183 0.011953 8.5477e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4126 0.49291 0.1505 0.018108 12.1387 0.11262 0.00014466 0.77752 0.0086375 0.0095858 0.0014215 0.98649 0.99141 3.0696e-006 1.2279e-005 0.15893 0.83975 0.87385 0.0014156 0.95144 0.44578 0.0019064 0.42235 1.8519 1.8504 16.0149 144.9352 0.00022982 -85.5018 0.45095
6.555 0.98811 5.4803e-005 3.8183 0.011953 8.549e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4127 0.49295 0.15051 0.01811 12.1411 0.11263 0.00014467 0.77751 0.008638 0.0095864 0.0014212 0.98649 0.99141 3.069e-006 1.2276e-005 0.15894 0.84019 0.87407 0.0014154 0.95173 0.44598 0.0019062 0.42236 1.853 1.8514 16.0149 144.9352 0.00022948 -85.5029 0.45195
6.556 0.98811 5.4803e-005 3.8183 0.011953 8.5503e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4128 0.493 0.15052 0.018111 12.1436 0.11264 0.00014468 0.77751 0.0086385 0.0095869 0.001421 0.9865 0.99141 3.0684e-006 1.2274e-005 0.15894 0.84064 0.87429 0.0014153 0.95202 0.44617 0.001906 0.42237 1.854 1.8524 16.0149 144.9352 0.00022915 -85.5041 0.45295
6.557 0.98811 5.4803e-005 3.8183 0.011953 8.5516e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4129 0.49304 0.15054 0.018112 12.146 0.11265 0.0001447 0.7775 0.008639 0.0095874 0.0014207 0.9865 0.99142 3.0678e-006 1.2271e-005 0.15895 0.84109 0.87451 0.0014152 0.95231 0.44636 0.0019058 0.42239 1.855 1.8534 16.0149 144.9352 0.00022881 -85.5052 0.45395
6.558 0.98811 5.4803e-005 3.8183 0.011953 8.5528e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.413 0.49309 0.15055 0.018114 12.1485 0.11265 0.00014471 0.77749 0.0086395 0.0095879 0.0014204 0.9865 0.99142 3.0672e-006 1.2269e-005 0.15895 0.84153 0.87472 0.001415 0.9526 0.44655 0.0019056 0.4224 1.856 1.8544 16.0149 144.9353 0.00022848 -85.5063 0.45495
6.559 0.98811 5.4803e-005 3.8183 0.011953 8.5541e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4131 0.49314 0.15057 0.018115 12.1509 0.11266 0.00014472 0.77748 0.00864 0.0095885 0.0014201 0.98651 0.99142 3.0666e-006 1.2266e-005 0.15895 0.84198 0.87494 0.0014149 0.95288 0.44674 0.0019055 0.42242 1.857 1.8554 16.0149 144.9353 0.00022814 -85.5074 0.45595
6.56 0.98811 5.4803e-005 3.8183 0.011953 8.5554e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4132 0.49318 0.15058 0.018116 12.1534 0.11267 0.00014473 0.77748 0.0086405 0.009589 0.0014198 0.98651 0.99142 3.066e-006 1.2264e-005 0.15896 0.84242 0.87515 0.0014147 0.95317 0.44694 0.0019053 0.42243 1.858 1.8564 16.0148 144.9353 0.00022781 -85.5085 0.45695
6.561 0.98811 5.4803e-005 3.8183 0.011953 8.5567e-005 0.0011658 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.4133 0.49323 0.1506 0.018118 12.1558 0.11268 0.00014474 0.77747 0.008641 0.0095895 0.0014195 0.98651 0.99142 3.0654e-006 1.2262e-005 0.15896 0.84286 0.87537 0.0014146 0.95345 0.44713 0.0019051 0.42244 1.859 1.8575 16.0148 144.9353 0.00022748 -85.5096 0.45795
6.562 0.98811 5.4803e-005 3.8183 0.011953 8.558e-005 0.0011658 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.4134 0.49327 0.15061 0.018119 12.1583 0.11268 0.00014475 0.77746 0.0086415 0.0095901 0.0014192 0.98652 0.99143 3.0648e-006 1.2259e-005 0.15897 0.8433 0.87558 0.0014144 0.95373 0.44732 0.0019049 0.42246 1.86 1.8585 16.0148 144.9353 0.00022715 -85.5107 0.45895
6.563 0.98811 5.4803e-005 3.8183 0.011953 8.5593e-005 0.0011658 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.4134 0.49332 0.15063 0.01812 12.1607 0.11269 0.00014477 0.77745 0.008642 0.0095906 0.001419 0.98652 0.99143 3.0642e-006 1.2257e-005 0.15897 0.84373 0.87579 0.0014143 0.95401 0.44751 0.0019048 0.42247 1.861 1.8594 16.0148 144.9354 0.00022683 -85.5118 0.45995
6.564 0.98811 5.4803e-005 3.8183 0.011953 8.5606e-005 0.0011658 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.4135 0.49337 0.15064 0.018121 12.1632 0.1127 0.00014478 0.77744 0.0086425 0.0095911 0.0014187 0.98652 0.99143 3.0636e-006 1.2255e-005 0.15897 0.84417 0.876 0.0014142 0.95429 0.4477 0.0019046 0.42249 1.862 1.8604 16.0148 144.9354 0.0002265 -85.5129 0.46095
6.565 0.98811 5.4803e-005 3.8183 0.011953 8.5619e-005 0.0011658 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.4136 0.49341 0.15066 0.018123 12.1656 0.11271 0.00014479 0.77744 0.008643 0.0095916 0.0014184 0.98653 0.99143 3.0631e-006 1.2252e-005 0.15898 0.84461 0.87621 0.001414 0.95456 0.44789 0.0019044 0.4225 1.863 1.8614 16.0148 144.9354 0.00022618 -85.5139 0.46195
6.566 0.98811 5.4803e-005 3.8183 0.011953 8.5632e-005 0.0011658 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.4137 0.49346 0.15067 0.018124 12.1681 0.11272 0.0001448 0.77743 0.0086435 0.0095922 0.0014182 0.98653 0.99143 3.0625e-006 1.225e-005 0.15898 0.84504 0.87642 0.0014139 0.95484 0.44809 0.0019042 0.42251 1.8639 1.8624 16.0148 144.9354 0.00022585 -85.515 0.46295
6.567 0.98811 5.4803e-005 3.8183 0.011953 8.5644e-005 0.0011658 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4138 0.4935 0.15068 0.018125 12.1705 0.11272 0.00014481 0.77742 0.0086439 0.0095927 0.001418 0.98653 0.99144 3.0619e-006 1.2248e-005 0.15898 0.84547 0.87663 0.0014137 0.95511 0.44828 0.0019041 0.42253 1.8649 1.8634 16.0148 144.9354 0.00022553 -85.516 0.46395
6.568 0.98811 5.4802e-005 3.8183 0.011953 8.5657e-005 0.0011658 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4139 0.49355 0.1507 0.018127 12.173 0.11273 0.00014482 0.77741 0.0086444 0.0095932 0.0014178 0.98654 0.99144 3.0613e-006 1.2245e-005 0.15899 0.8459 0.87684 0.0014136 0.95538 0.44847 0.0019039 0.42254 1.8659 1.8644 16.0148 144.9355 0.00022521 -85.5171 0.46495
6.569 0.98811 5.4802e-005 3.8183 0.011953 8.567e-005 0.0011658 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.414 0.4936 0.15071 0.018128 12.1754 0.11274 0.00014483 0.77741 0.0086449 0.0095938 0.0014176 0.98654 0.99144 3.0608e-006 1.2243e-005 0.15899 0.84633 0.87704 0.0014135 0.95565 0.44866 0.0019037 0.42256 1.8669 1.8654 16.0148 144.9355 0.00022489 -85.5181 0.46595
6.57 0.98811 5.4802e-005 3.8183 0.011952 8.5683e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4141 0.49364 0.15073 0.018129 12.1779 0.11275 0.00014485 0.7774 0.0086454 0.0095943 0.0014173 0.98654 0.99144 3.0602e-006 1.2241e-005 0.159 0.84676 0.87725 0.0014134 0.95591 0.44885 0.0019036 0.42257 1.8679 1.8664 16.0148 144.9355 0.00022457 -85.5192 0.46695
6.571 0.98811 5.4802e-005 3.8183 0.011952 8.5696e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4142 0.49369 0.15074 0.01813 12.1803 0.11276 0.00014486 0.77739 0.0086459 0.0095948 0.0014171 0.98655 0.99145 3.0597e-006 1.2239e-005 0.159 0.84719 0.87746 0.0014133 0.95618 0.44904 0.0019034 0.42258 1.8688 1.8673 16.0148 144.9355 0.00022425 -85.5202 0.46795
6.572 0.98811 5.4802e-005 3.8183 0.011952 8.5709e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4143 0.49373 0.15076 0.018132 12.1828 0.11276 0.00014487 0.77738 0.0086464 0.0095954 0.0014168 0.98655 0.99145 3.0591e-006 1.2236e-005 0.159 0.84761 0.87766 0.0014131 0.95644 0.44923 0.0019032 0.4226 1.8698 1.8683 16.0148 144.9355 0.00022394 -85.5212 0.46895
6.573 0.98811 5.4802e-005 3.8183 0.011952 8.5722e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4144 0.49378 0.15077 0.018133 12.1853 0.11277 0.00014488 0.77737 0.0086469 0.0095959 0.0014166 0.98655 0.99145 3.0586e-006 1.2234e-005 0.15901 0.84804 0.87786 0.001413 0.9567 0.44943 0.0019031 0.42261 1.8708 1.8693 16.0148 144.9355 0.00022363 -85.5222 0.46995
6.574 0.98811 5.4802e-005 3.8183 0.011952 8.5735e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4144 0.49382 0.15079 0.018134 12.1877 0.11278 0.00014489 0.77737 0.0086474 0.0095964 0.0014163 0.98655 0.99145 3.058e-006 1.2232e-005 0.15901 0.84846 0.87807 0.0014129 0.95696 0.44962 0.0019029 0.42263 1.8717 1.8702 16.0148 144.9356 0.00022331 -85.5232 0.47095
6.575 0.98811 5.4802e-005 3.8183 0.011952 8.5748e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4145 0.49387 0.1508 0.018136 12.1902 0.11279 0.0001449 0.77736 0.0086479 0.0095969 0.001416 0.98656 0.99145 3.0575e-006 1.223e-005 0.15902 0.84888 0.87827 0.0014128 0.95722 0.44981 0.0019028 0.42264 1.8727 1.8712 16.0147 144.9356 0.000223 -85.5242 0.47195
6.576 0.98811 5.4802e-005 3.8183 0.011952 8.576e-005 0.0011658 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4146 0.49392 0.15082 0.018137 12.1926 0.11279 0.00014491 0.77735 0.0086484 0.0095975 0.0014158 0.98656 0.99146 3.057e-006 1.2228e-005 0.15902 0.8493 0.87847 0.0014127 0.95748 0.45 0.0019026 0.42266 1.8736 1.8722 16.0147 144.9356 0.00022269 -85.5252 0.47295
6.577 0.98811 5.4802e-005 3.8183 0.011952 8.5773e-005 0.0011659 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4147 0.49396 0.15083 0.018138 12.1951 0.1128 0.00014493 0.77734 0.0086489 0.009598 0.0014156 0.98656 0.99146 3.0564e-006 1.2226e-005 0.15902 0.84972 0.87867 0.0014125 0.95773 0.45019 0.0019024 0.42267 1.8746 1.8731 16.0147 144.9356 0.00022238 -85.5262 0.47395
6.578 0.98811 5.4802e-005 3.8183 0.011952 8.5786e-005 0.0011659 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4148 0.49401 0.15085 0.018139 12.1975 0.11281 0.00014494 0.77733 0.0086494 0.0095985 0.0014153 0.98657 0.99146 3.0559e-006 1.2224e-005 0.15903 0.85014 0.87887 0.0014124 0.95799 0.45038 0.0019023 0.42268 1.8756 1.8741 16.0147 144.9356 0.00022207 -85.5271 0.47495
6.579 0.98811 5.4802e-005 3.8183 0.011952 8.5799e-005 0.0011659 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.4149 0.49405 0.15086 0.018141 12.2 0.11282 0.00014495 0.77733 0.0086499 0.009599 0.0014151 0.98657 0.99146 3.0554e-006 1.2222e-005 0.15903 0.85055 0.87907 0.0014123 0.95824 0.45057 0.0019021 0.4227 1.8765 1.875 16.0147 144.9357 0.00022177 -85.5281 0.47595
6.58 0.98811 5.4801e-005 3.8183 0.011952 8.5812e-005 0.0011659 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.415 0.4941 0.15087 0.018142 12.2025 0.11283 0.00014496 0.77732 0.0086503 0.0095996 0.0014149 0.98657 0.99146 3.0549e-006 1.2219e-005 0.15903 0.85097 0.87926 0.0014122 0.95849 0.45076 0.001902 0.42271 1.8775 1.876 16.0147 144.9357 0.00022146 -85.5291 0.47695
6.581 0.98811 5.4801e-005 3.8183 0.011952 8.5825e-005 0.0011659 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.4151 0.49415 0.15089 0.018143 12.2049 0.11283 0.00014497 0.77731 0.0086508 0.0096001 0.0014147 0.98658 0.99146 3.0544e-006 1.2217e-005 0.15904 0.85138 0.87946 0.0014121 0.95874 0.45095 0.0019018 0.42273 1.8784 1.877 16.0147 144.9357 0.00022116 -85.53 0.47795
6.582 0.98811 5.4801e-005 3.8183 0.011952 8.5838e-005 0.0011659 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.4152 0.49419 0.1509 0.018145 12.2074 0.11284 0.00014498 0.7773 0.0086513 0.0096006 0.0014145 0.98658 0.99147 3.0539e-006 1.2215e-005 0.15904 0.85179 0.87966 0.001412 0.95898 0.45114 0.0019017 0.42274 1.8793 1.8779 16.0147 144.9357 0.00022085 -85.531 0.47895
6.583 0.98811 5.4801e-005 3.8183 0.011952 8.5851e-005 0.0011659 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.4153 0.49424 0.15092 0.018146 12.2098 0.11285 0.000145 0.7773 0.0086518 0.0096012 0.0014143 0.98658 0.99147 3.0533e-006 1.2213e-005 0.15905 0.85221 0.87985 0.0014118 0.95923 0.45133 0.0019015 0.42275 1.8803 1.8788 16.0147 144.9357 0.00022055 -85.5319 0.47995
6.584 0.98811 5.4801e-005 3.8183 0.011952 8.5864e-005 0.0011659 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.4154 0.49428 0.15093 0.018147 12.2123 0.11286 0.00014501 0.77729 0.0086523 0.0096017 0.0014141 0.98658 0.99147 3.0528e-006 1.2211e-005 0.15905 0.85262 0.88005 0.0014117 0.95947 0.45152 0.0019014 0.42277 1.8812 1.8798 16.0147 144.9358 0.00022025 -85.5328 0.48095
6.585 0.98811 5.4801e-005 3.8183 0.011952 8.5876e-005 0.0011659 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.4154 0.49433 0.15095 0.018149 12.2148 0.11286 0.00014502 0.77728 0.0086528 0.0096022 0.0014139 0.98659 0.99147 3.0523e-006 1.2209e-005 0.15905 0.85302 0.88024 0.0014116 0.95971 0.45171 0.0019012 0.42278 1.8822 1.8807 16.0147 144.9358 0.00021995 -85.5337 0.48195
6.586 0.98811 5.4801e-005 3.8183 0.011952 8.5889e-005 0.0011659 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4155 0.49438 0.15096 0.01815 12.2172 0.11287 0.00014503 0.77727 0.0086533 0.0096027 0.0014137 0.98659 0.99147 3.0518e-006 1.2207e-005 0.15906 0.85343 0.88043 0.0014115 0.95996 0.4519 0.0019011 0.4228 1.8831 1.8817 16.0147 144.9358 0.00021966 -85.5347 0.48295
6.587 0.98811 5.4801e-005 3.8183 0.011952 8.5902e-005 0.0011659 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4156 0.49442 0.15098 0.018151 12.2197 0.11288 0.00014504 0.77726 0.0086538 0.0096033 0.0014135 0.98659 0.99148 3.0513e-006 1.2205e-005 0.15906 0.85384 0.88062 0.0014114 0.9602 0.45209 0.0019009 0.42281 1.884 1.8826 16.0146 144.9358 0.00021936 -85.5356 0.48395
6.588 0.98811 5.4801e-005 3.8183 0.011952 8.5915e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4157 0.49447 0.15099 0.018152 12.2221 0.11289 0.00014505 0.77726 0.0086543 0.0096038 0.0014133 0.9866 0.99148 3.0509e-006 1.2203e-005 0.15906 0.85424 0.88082 0.0014113 0.96043 0.45228 0.0019008 0.42282 1.8849 1.8835 16.0146 144.9358 0.00021906 -85.5365 0.48495
6.589 0.98811 5.4801e-005 3.8183 0.011952 8.5928e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4158 0.49451 0.15101 0.018154 12.2246 0.1129 0.00014506 0.77725 0.0086548 0.0096043 0.0014131 0.9866 0.99148 3.0504e-006 1.2201e-005 0.15907 0.85465 0.88101 0.0014112 0.96067 0.45247 0.0019006 0.42284 1.8859 1.8845 16.0146 144.9359 0.00021877 -85.5374 0.48595
6.59 0.98811 5.4801e-005 3.8183 0.011952 8.5941e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4159 0.49456 0.15102 0.018155 12.2271 0.1129 0.00014508 0.77724 0.0086553 0.0096048 0.0014129 0.9866 0.99148 3.0499e-006 1.22e-005 0.15907 0.85505 0.8812 0.001411 0.9609 0.45267 0.0019005 0.42285 1.8868 1.8854 16.0146 144.9359 0.00021848 -85.5383 0.48695
6.591 0.98811 5.4801e-005 3.8183 0.011952 8.5954e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.416 0.4946 0.15103 0.018156 12.2295 0.11291 0.00014509 0.77723 0.0086557 0.0096054 0.0014127 0.9866 0.99148 3.0494e-006 1.2198e-005 0.15908 0.85545 0.88138 0.0014109 0.96114 0.45286 0.0019003 0.42287 1.8877 1.8863 16.0146 144.9359 0.00021818 -85.5392 0.48795
6.592 0.98811 5.4801e-005 3.8183 0.011952 8.5967e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4161 0.49465 0.15105 0.018158 12.232 0.11292 0.0001451 0.77723 0.0086562 0.0096059 0.0014125 0.98661 0.99148 3.0489e-006 1.2196e-005 0.15908 0.85585 0.88157 0.0014108 0.96137 0.45305 0.0019002 0.42288 1.8886 1.8872 16.0146 144.9359 0.00021789 -85.54 0.48895
6.593 0.98811 5.48e-005 3.8183 0.011952 8.598e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4162 0.4947 0.15106 0.018159 12.2344 0.11293 0.00014511 0.77722 0.0086567 0.0096064 0.0014123 0.98661 0.99149 3.0485e-006 1.2194e-005 0.15908 0.85625 0.88176 0.0014107 0.9616 0.45323 0.0019001 0.42289 1.8896 1.8882 16.0146 144.9359 0.0002176 -85.5409 0.48995
6.594 0.98811 5.48e-005 3.8183 0.011952 8.5992e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4163 0.49474 0.15108 0.01816 12.2369 0.11294 0.00014512 0.77721 0.0086572 0.009607 0.001412 0.98661 0.99149 3.048e-006 1.2192e-005 0.15909 0.85665 0.88195 0.0014106 0.96183 0.45342 0.0018999 0.42291 1.8905 1.8891 16.0146 144.936 0.00021732 -85.5418 0.49095
6.595 0.98811 5.48e-005 3.8183 0.011952 8.6005e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4164 0.49479 0.15109 0.018161 12.2394 0.11294 0.00014513 0.7772 0.0086577 0.0096075 0.0014118 0.98661 0.99149 3.0475e-006 1.219e-005 0.15909 0.85704 0.88213 0.0014105 0.96206 0.45361 0.0018998 0.42292 1.8914 1.89 16.0146 144.936 0.00021703 -85.5427 0.49195
6.596 0.98811 5.48e-005 3.8183 0.011952 8.6018e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4164 0.49483 0.15111 0.018163 12.2418 0.11295 0.00014515 0.77719 0.0086582 0.009608 0.0014116 0.98662 0.99149 3.0471e-006 1.2188e-005 0.1591 0.85744 0.88232 0.0014104 0.96228 0.4538 0.0018996 0.42294 1.8923 1.8909 16.0146 144.936 0.00021674 -85.5435 0.49295
6.597 0.98811 5.48e-005 3.8183 0.011952 8.6031e-005 0.0011659 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.4165 0.49488 0.15112 0.018164 12.2443 0.11296 0.00014516 0.77719 0.0086587 0.0096085 0.0014114 0.98662 0.99149 3.0466e-006 1.2186e-005 0.1591 0.85783 0.8825 0.0014103 0.96251 0.45399 0.0018995 0.42295 1.8932 1.8918 16.0146 144.936 0.00021646 -85.5444 0.49395
6.598 0.98811 5.48e-005 3.8183 0.011952 8.6044e-005 0.0011659 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.4166 0.49493 0.15114 0.018165 12.2468 0.11297 0.00014517 0.77718 0.0086592 0.0096091 0.0014112 0.98662 0.9915 3.0462e-006 1.2185e-005 0.1591 0.85822 0.88269 0.0014102 0.96273 0.45418 0.0018994 0.42297 1.8941 1.8927 16.0145 144.936 0.00021617 -85.5452 0.49495
6.599 0.98811 5.48e-005 3.8183 0.011952 8.6057e-005 0.0011659 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.4167 0.49497 0.15115 0.018167 12.2492 0.11297 0.00014518 0.77717 0.0086597 0.0096096 0.0014109 0.98662 0.9915 3.0457e-006 1.2183e-005 0.15911 0.85861 0.88287 0.0014101 0.96295 0.45437 0.0018992 0.42298 1.895 1.8936 16.0145 144.9361 0.00021589 -85.546 0.49595
6.6 0.98811 5.48e-005 3.8183 0.011952 8.607e-005 0.0011659 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.4168 0.49502 0.15117 0.018168 12.2517 0.11298 0.00014519 0.77716 0.0086602 0.0096101 0.0014107 0.98663 0.9915 3.0453e-006 1.2181e-005 0.15911 0.859 0.88305 0.00141 0.96317 0.45456 0.0018991 0.42299 1.8959 1.8945 16.0145 144.9361 0.00021561 -85.5469 0.49695
6.601 0.98811 5.48e-005 3.8183 0.011952 8.6083e-005 0.0011659 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.4169 0.49506 0.15118 0.018169 12.2542 0.11299 0.0001452 0.77716 0.0086607 0.0096106 0.0014105 0.98663 0.9915 3.0448e-006 1.2179e-005 0.15911 0.85939 0.88323 0.0014099 0.96339 0.45475 0.001899 0.42301 1.8968 1.8954 16.0145 144.9361 0.00021533 -85.5477 0.49795
6.602 0.98811 5.48e-005 3.8183 0.011952 8.6096e-005 0.001166 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.417 0.49511 0.15119 0.01817 12.2566 0.113 0.00014521 0.77715 0.0086611 0.0096112 0.0014103 0.98663 0.9915 3.0444e-006 1.2177e-005 0.15912 0.85978 0.88341 0.0014098 0.96361 0.45494 0.0018988 0.42302 1.8977 1.8963 16.0145 144.9361 0.00021505 -85.5485 0.49895
6.603 0.98811 5.48e-005 3.8183 0.011952 8.6109e-005 0.001166 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.4171 0.49516 0.15121 0.018172 12.2591 0.11301 0.00014523 0.77714 0.0086616 0.0096117 0.0014101 0.98663 0.9915 3.0439e-006 1.2176e-005 0.15912 0.86017 0.88359 0.0014097 0.96383 0.45513 0.0018987 0.42304 1.8986 1.8972 16.0145 144.9361 0.00021477 -85.5493 0.49995
6.604 0.98811 5.48e-005 3.8183 0.011952 8.6121e-005 0.001166 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.4172 0.4952 0.15122 0.018173 12.2616 0.11301 0.00014524 0.77713 0.0086621 0.0096122 0.0014099 0.98664 0.99151 3.0435e-006 1.2174e-005 0.15913 0.86055 0.88377 0.0014096 0.96404 0.45532 0.0018986 0.42305 1.8995 1.8981 16.0145 144.9362 0.00021449 -85.5501 0.50095
6.605 0.98811 5.48e-005 3.8183 0.011952 8.6134e-005 0.001166 0.23346 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4173 0.49525 0.15124 0.018174 12.264 0.11302 0.00014525 0.77712 0.0086626 0.0096127 0.0014098 0.98664 0.99151 3.0431e-006 1.2172e-005 0.15913 0.86094 0.88395 0.0014095 0.96425 0.45551 0.0018984 0.42306 1.9004 1.899 16.0145 144.9362 0.00021422 -85.551 0.50195
6.606 0.98811 5.4799e-005 3.8183 0.011952 8.6147e-005 0.001166 0.23346 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4174 0.49529 0.15125 0.018176 12.2665 0.11303 0.00014526 0.77712 0.0086631 0.0096133 0.0014096 0.98664 0.99151 3.0426e-006 1.217e-005 0.15913 0.86132 0.88413 0.0014094 0.96447 0.4557 0.0018983 0.42308 1.9012 1.8999 16.0145 144.9362 0.00021394 -85.5518 0.50295
6.607 0.98811 5.4799e-005 3.8183 0.011952 8.616e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4175 0.49534 0.15127 0.018177 12.269 0.11304 0.00014527 0.77711 0.0086636 0.0096138 0.0014094 0.98664 0.99151 3.0422e-006 1.2169e-005 0.15914 0.8617 0.88431 0.0014093 0.96468 0.45589 0.0018982 0.42309 1.9021 1.9008 16.0144 144.9362 0.00021367 -85.5525 0.50395
6.608 0.98811 5.4799e-005 3.8183 0.011952 8.6173e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4175 0.49538 0.15128 0.018178 12.2714 0.11304 0.00014528 0.7771 0.0086641 0.0096143 0.0014093 0.98665 0.99151 3.0418e-006 1.2167e-005 0.15914 0.86208 0.88448 0.0014092 0.96489 0.45608 0.001898 0.42311 1.903 1.9017 16.0144 144.9362 0.0002134 -85.5533 0.50495
6.609 0.98811 5.4799e-005 3.8183 0.011952 8.6186e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4176 0.49543 0.1513 0.018179 12.2739 0.11305 0.00014529 0.77709 0.0086646 0.0096148 0.0014091 0.98665 0.99151 3.0414e-006 1.2165e-005 0.15915 0.86246 0.88466 0.0014091 0.96509 0.45627 0.0018979 0.42312 1.9039 1.9025 16.0144 144.9363 0.00021313 -85.5541 0.50595
6.61 0.98811 5.4799e-005 3.8183 0.011952 8.6199e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4177 0.49548 0.15131 0.018181 12.2764 0.11306 0.00014531 0.77708 0.0086651 0.0096154 0.001409 0.98665 0.99151 3.0409e-006 1.2164e-005 0.15915 0.86284 0.88483 0.001409 0.9653 0.45645 0.0018978 0.42314 1.9047 1.9034 16.0144 144.9363 0.00021286 -85.5549 0.50695
6.611 0.98811 5.4799e-005 3.8183 0.011952 8.6212e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4178 0.49552 0.15133 0.018182 12.2788 0.11307 0.00014532 0.77708 0.0086656 0.0096159 0.0014088 0.98665 0.99152 3.0405e-006 1.2162e-005 0.15915 0.86321 0.88501 0.0014089 0.96551 0.45664 0.0018977 0.42315 1.9056 1.9043 16.0144 144.9363 0.00021259 -85.5557 0.50795
6.612 0.98811 5.4799e-005 3.8183 0.011952 8.6225e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4179 0.49557 0.15134 0.018183 12.2813 0.11308 0.00014533 0.77707 0.008666 0.0096164 0.0014087 0.98666 0.99152 3.0401e-006 1.216e-005 0.15916 0.86359 0.88518 0.0014088 0.96571 0.45683 0.0018975 0.42316 1.9065 1.9052 16.0144 144.9363 0.00021232 -85.5564 0.50895
6.613 0.98811 5.4799e-005 3.8183 0.011952 8.6237e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.418 0.49561 0.15136 0.018185 12.2838 0.11308 0.00014534 0.77706 0.0086665 0.0096169 0.0014085 0.98666 0.99152 3.0397e-006 1.2159e-005 0.15916 0.86396 0.88535 0.0014087 0.96591 0.45702 0.0018974 0.42318 1.9074 1.9061 16.0144 144.9363 0.00021205 -85.5572 0.50995
6.614 0.98811 5.4799e-005 3.8183 0.011952 8.625e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4181 0.49566 0.15137 0.018186 12.2862 0.11309 0.00014535 0.77705 0.008667 0.0096175 0.0014083 0.98666 0.99152 3.0393e-006 1.2157e-005 0.15916 0.86434 0.88553 0.0014086 0.96611 0.45721 0.0018973 0.42319 1.9082 1.9069 16.0144 144.9364 0.00021178 -85.5579 0.51095
6.615 0.98811 5.4799e-005 3.8183 0.011952 8.6263e-005 0.001166 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.4182 0.49571 0.15138 0.018187 12.2887 0.1131 0.00014536 0.77705 0.0086675 0.009618 0.0014081 0.98666 0.99152 3.0389e-006 1.2156e-005 0.15917 0.86471 0.8857 0.0014085 0.96631 0.4574 0.0018972 0.42321 1.9091 1.9078 16.0144 144.9364 0.00021152 -85.5587 0.51195
6.616 0.98811 5.4799e-005 3.8183 0.011952 8.6276e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.4183 0.49575 0.1514 0.018188 12.2912 0.11311 0.00014537 0.77704 0.008668 0.0096185 0.001408 0.98667 0.99152 3.0385e-006 1.2154e-005 0.15917 0.86508 0.88587 0.0014084 0.96651 0.45759 0.0018971 0.42322 1.91 1.9087 16.0143 144.9364 0.00021126 -85.5594 0.51295
6.617 0.98811 5.4799e-005 3.8183 0.011952 8.6289e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.4184 0.4958 0.15141 0.01819 12.2936 0.11311 0.00014539 0.77703 0.0086685 0.009619 0.0014078 0.98667 0.99153 3.0381e-006 1.2152e-005 0.15918 0.86545 0.88604 0.0014083 0.96671 0.45777 0.0018969 0.42324 1.9108 1.9095 16.0143 144.9364 0.00021099 -85.5602 0.51395
6.618 0.98811 5.4799e-005 3.8183 0.011952 8.6302e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.4185 0.49584 0.15143 0.018191 12.2961 0.11312 0.0001454 0.77702 0.008669 0.0096196 0.0014076 0.98667 0.99153 3.0377e-006 1.2151e-005 0.15918 0.86582 0.88621 0.0014082 0.96691 0.45796 0.0018968 0.42325 1.9117 1.9104 16.0143 144.9364 0.00021073 -85.5609 0.51495
6.619 0.98811 5.4798e-005 3.8183 0.011952 8.6315e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.4185 0.49589 0.15144 0.018192 12.2986 0.11313 0.00014541 0.77701 0.0086695 0.0096201 0.0014073 0.98667 0.99153 3.0373e-006 1.2149e-005 0.15918 0.86619 0.88638 0.0014081 0.9671 0.45815 0.0018967 0.42326 1.9125 1.9112 16.0143 144.9365 0.00021047 -85.5616 0.51595
6.62 0.98811 5.4798e-005 3.8183 0.011952 8.6328e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.4186 0.49594 0.15146 0.018194 12.3011 0.11314 0.00014542 0.77701 0.00867 0.0096206 0.0014071 0.98667 0.99153 3.0369e-006 1.2148e-005 0.15919 0.86655 0.88654 0.001408 0.9673 0.45834 0.0018966 0.42328 1.9134 1.9121 16.0143 144.9365 0.00021021 -85.5624 0.51695
6.621 0.98811 5.4798e-005 3.8183 0.011952 8.6341e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.4187 0.49598 0.15147 0.018195 12.3035 0.11315 0.00014543 0.777 0.0086704 0.0096211 0.001407 0.98668 0.99153 3.0365e-006 1.2146e-005 0.15919 0.86692 0.88671 0.0014079 0.96749 0.45853 0.0018965 0.42329 1.9142 1.9129 16.0143 144.9365 0.00020995 -85.5631 0.51795
6.622 0.98811 5.4798e-005 3.8183 0.011952 8.6353e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.4188 0.49603 0.15149 0.018196 12.306 0.11315 0.00014544 0.77699 0.0086709 0.0096217 0.0014068 0.98668 0.99153 3.0362e-006 1.2145e-005 0.15919 0.86728 0.88688 0.0014079 0.96768 0.45872 0.0018964 0.42331 1.9151 1.9138 16.0143 144.9365 0.00020969 -85.5638 0.51895
6.623 0.98811 5.4798e-005 3.8183 0.011952 8.6366e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.4189 0.49607 0.1515 0.018197 12.3085 0.11316 0.00014546 0.77698 0.0086714 0.0096222 0.0014067 0.98668 0.99153 3.0358e-006 1.2143e-005 0.1592 0.86765 0.88704 0.0014078 0.96787 0.4589 0.0018962 0.42332 1.9159 1.9146 16.0143 144.9365 0.00020944 -85.5645 0.51995
6.624 0.98811 5.4798e-005 3.8183 0.011952 8.6379e-005 0.001166 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.419 0.49612 0.15152 0.018199 12.311 0.11317 0.00014547 0.77698 0.0086719 0.0096227 0.0014066 0.98668 0.99153 3.0354e-006 1.2142e-005 0.1592 0.86801 0.88721 0.0014077 0.96806 0.45909 0.0018961 0.42333 1.9168 1.9155 16.0142 144.9366 0.00020918 -85.5652 0.52095
6.625 0.98811 5.4798e-005 3.8183 0.011952 8.6392e-005 0.001166 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4191 0.49616 0.15153 0.0182 12.3134 0.11318 0.00014548 0.77697 0.0086724 0.0096232 0.0014064 0.98668 0.99154 3.035e-006 1.214e-005 0.15921 0.86837 0.88737 0.0014076 0.96825 0.45928 0.001896 0.42335 1.9176 1.9163 16.0142 144.9366 0.00020893 -85.5659 0.52195
6.626 0.98811 5.4798e-005 3.8183 0.011952 8.6405e-005 0.001166 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4192 0.49621 0.15154 0.018201 12.3159 0.11319 0.00014549 0.77696 0.0086729 0.0096238 0.0014062 0.98669 0.99154 3.0346e-006 1.2139e-005 0.15921 0.86873 0.88754 0.0014075 0.96843 0.45947 0.0018959 0.42336 1.9184 1.9172 16.0142 144.9366 0.00020867 -85.5666 0.52295
6.627 0.98811 5.4798e-005 3.8183 0.011952 8.6418e-005 0.001166 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4193 0.49626 0.15156 0.018203 12.3184 0.11319 0.0001455 0.77695 0.0086734 0.0096243 0.001406 0.98669 0.99154 3.0343e-006 1.2137e-005 0.15921 0.86909 0.8877 0.0014075 0.96862 0.45966 0.0018958 0.42338 1.9193 1.918 16.0142 144.9366 0.00020842 -85.5673 0.52395
6.628 0.98811 5.4798e-005 3.8183 0.011952 8.6431e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4194 0.4963 0.15157 0.018204 12.3208 0.1132 0.00014551 0.77694 0.0086739 0.0096248 0.0014058 0.98669 0.99154 3.0339e-006 1.2136e-005 0.15922 0.86944 0.88787 0.0014074 0.9688 0.45984 0.0018957 0.42339 1.9201 1.9189 16.0142 144.9366 0.00020817 -85.568 0.52495
6.629 0.98811 5.4798e-005 3.8183 0.011951 8.6444e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4195 0.49635 0.15159 0.018205 12.3233 0.11321 0.00014552 0.77694 0.0086743 0.0096253 0.0014056 0.98669 0.99154 3.0335e-006 1.2134e-005 0.15922 0.8698 0.88803 0.0014073 0.96899 0.46003 0.0018956 0.42341 1.9209 1.9197 16.0142 144.9367 0.00020792 -85.5686 0.52595
6.63 0.98811 5.4798e-005 3.8183 0.011951 8.6457e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4195 0.49639 0.1516 0.018206 12.3258 0.11322 0.00014554 0.77693 0.0086748 0.0096259 0.0014054 0.9867 0.99154 3.0332e-006 1.2133e-005 0.15923 0.87015 0.88819 0.0014072 0.96917 0.46022 0.0018955 0.42342 1.9218 1.9205 16.0142 144.9367 0.00020767 -85.5693 0.52695
6.631 0.98811 5.4797e-005 3.8183 0.011951 8.6469e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4196 0.49644 0.15162 0.018208 12.3283 0.11322 0.00014555 0.77692 0.0086753 0.0096264 0.0014053 0.9867 0.99154 3.0328e-006 1.2131e-005 0.15923 0.87051 0.88835 0.0014071 0.96935 0.46041 0.0018954 0.42343 1.9226 1.9214 16.0142 144.9367 0.00020742 -85.57 0.52795
6.632 0.98811 5.4797e-005 3.8183 0.011951 8.6482e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4197 0.49649 0.15163 0.018209 12.3307 0.11323 0.00014556 0.77691 0.0086758 0.0096269 0.0014052 0.9867 0.99155 3.0325e-006 1.213e-005 0.15923 0.87086 0.88851 0.001407 0.96953 0.46059 0.0018953 0.42345 1.9234 1.9222 16.0141 144.9367 0.00020717 -85.5707 0.52895
6.633 0.98811 5.4797e-005 3.8183 0.011951 8.6495e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4198 0.49653 0.15165 0.01821 12.3332 0.11324 0.00014557 0.77691 0.0086763 0.0096274 0.0014051 0.9867 0.99155 3.0321e-006 1.2128e-005 0.15924 0.87121 0.88867 0.001407 0.96971 0.46078 0.0018951 0.42346 1.9243 1.923 16.0141 144.9367 0.00020692 -85.5713 0.52995
6.634 0.98811 5.4797e-005 3.8183 0.011951 8.6508e-005 0.0011661 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.4199 0.49658 0.15166 0.018212 12.3357 0.11325 0.00014558 0.7769 0.0086768 0.009628 0.001405 0.9867 0.99155 3.0318e-006 1.2127e-005 0.15924 0.87156 0.88883 0.0014069 0.96989 0.46097 0.001895 0.42348 1.9251 1.9238 16.0141 144.9368 0.00020668 -85.572 0.53095
6.635 0.98811 5.4797e-005 3.8183 0.011951 8.6521e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.42 0.49662 0.15168 0.018213 12.3382 0.11326 0.00014559 0.77689 0.0086773 0.0096285 0.0014048 0.98671 0.99155 3.0314e-006 1.2126e-005 0.15924 0.87191 0.88899 0.0014068 0.97006 0.46116 0.0018949 0.42349 1.9259 1.9247 16.0141 144.9368 0.00020643 -85.5726 0.53195
6.636 0.98811 5.4797e-005 3.8183 0.011951 8.6534e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4201 0.49667 0.15169 0.018214 12.3407 0.11326 0.0001456 0.77688 0.0086778 0.009629 0.0014047 0.98671 0.99155 3.0311e-006 1.2124e-005 0.15925 0.87226 0.88915 0.0014067 0.97024 0.46134 0.0018948 0.42351 1.9267 1.9255 16.0141 144.9368 0.00020619 -85.5733 0.53295
6.637 0.98811 5.4797e-005 3.8183 0.011951 8.6547e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4202 0.49671 0.1517 0.018215 12.3431 0.11327 0.00014562 0.77687 0.0086782 0.0096295 0.0014045 0.98671 0.99155 3.0307e-006 1.2123e-005 0.15925 0.87261 0.8893 0.0014067 0.97041 0.46153 0.0018947 0.42352 1.9275 1.9263 16.0141 144.9368 0.00020595 -85.5739 0.53395
6.638 0.98811 5.4797e-005 3.8183 0.011951 8.656e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4203 0.49676 0.15172 0.018217 12.3456 0.11328 0.00014563 0.77687 0.0086787 0.00963 0.0014043 0.98671 0.99155 3.0304e-006 1.2121e-005 0.15926 0.87296 0.88946 0.0014066 0.97058 0.46172 0.0018946 0.42353 1.9283 1.9271 16.0141 144.9368 0.00020571 -85.5746 0.53495
6.639 0.98811 5.4797e-005 3.8183 0.011951 8.6573e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4204 0.49681 0.15173 0.018218 12.3481 0.11329 0.00014564 0.77686 0.0086792 0.0096306 0.001404 0.98671 0.99155 3.03e-006 1.212e-005 0.15926 0.8733 0.88961 0.0014065 0.97076 0.46191 0.0018945 0.42355 1.9292 1.9279 16.014 144.9368 0.00020546 -85.5752 0.53595
6.64 0.98811 5.4797e-005 3.8183 0.011951 8.6585e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4205 0.49685 0.15175 0.018219 12.3506 0.11329 0.00014565 0.77685 0.0086797 0.0096311 0.0014039 0.98672 0.99156 3.0297e-006 1.2119e-005 0.15926 0.87365 0.88977 0.0014064 0.97093 0.46209 0.0018944 0.42356 1.93 1.9288 16.014 144.9369 0.00020522 -85.5758 0.53695
6.641 0.98811 5.4797e-005 3.8183 0.011951 8.6598e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4205 0.4969 0.15176 0.018221 12.353 0.1133 0.00014566 0.77684 0.0086802 0.0096316 0.0014037 0.98672 0.99156 3.0294e-006 1.2117e-005 0.15927 0.87399 0.88992 0.0014063 0.9711 0.46228 0.0018943 0.42358 1.9308 1.9296 16.014 144.9369 0.00020499 -85.5764 0.53795
6.642 0.98811 5.4797e-005 3.8183 0.011951 8.6611e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4206 0.49694 0.15178 0.018222 12.3555 0.11331 0.00014567 0.77684 0.0086807 0.0096321 0.0014036 0.98672 0.99156 3.029e-006 1.2116e-005 0.15927 0.87433 0.89008 0.0014062 0.97126 0.46247 0.0018942 0.42359 1.9316 1.9304 16.014 144.9369 0.00020475 -85.5771 0.53895
6.643 0.98811 5.4797e-005 3.8183 0.011951 8.6624e-005 0.0011661 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4207 0.49699 0.15179 0.018223 12.358 0.11332 0.00014568 0.77683 0.0086812 0.0096327 0.0014034 0.98672 0.99156 3.0287e-006 1.2115e-005 0.15927 0.87467 0.89023 0.0014062 0.97143 0.46265 0.0018941 0.4236 1.9324 1.9312 16.014 144.9369 0.00020451 -85.5777 0.53995
6.644 0.98811 5.4796e-005 3.8183 0.011951 8.6637e-005 0.0011661 0.23349 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.4208 0.49704 0.15181 0.018224 12.3605 0.11333 0.0001457 0.77682 0.0086817 0.0096332 0.0014033 0.98672 0.99156 3.0284e-006 1.2113e-005 0.15928 0.87501 0.89039 0.0014061 0.9716 0.46284 0.001894 0.42362 1.9332 1.932 16.014 144.9369 0.00020427 -85.5783 0.54095
6.645 0.98811 5.4796e-005 3.8183 0.011951 8.665e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4209 0.49708 0.15182 0.018226 12.363 0.11333 0.00014571 0.77681 0.0086821 0.0096337 0.0014032 0.98672 0.99156 3.028e-006 1.2112e-005 0.15928 0.87535 0.89054 0.001406 0.97176 0.46303 0.0018939 0.42363 1.934 1.9328 16.014 144.937 0.00020404 -85.5789 0.54195
6.646 0.98811 5.4796e-005 3.8183 0.011951 8.6663e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.421 0.49713 0.15184 0.018227 12.3654 0.11334 0.00014572 0.77681 0.0086826 0.0096342 0.0014031 0.98673 0.99156 3.0277e-006 1.2111e-005 0.15929 0.87569 0.89069 0.0014059 0.97193 0.46321 0.0018938 0.42365 1.9348 1.9336 16.0139 144.937 0.0002038 -85.5795 0.54295
6.647 0.98811 5.4796e-005 3.8183 0.011951 8.6676e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4211 0.49717 0.15185 0.018228 12.3679 0.11335 0.00014573 0.7768 0.0086831 0.0096347 0.001403 0.98673 0.99156 3.0274e-006 1.211e-005 0.15929 0.87602 0.89084 0.0014059 0.97209 0.4634 0.0018937 0.42366 1.9356 1.9344 16.0139 144.937 0.00020357 -85.5801 0.54395
6.648 0.98811 5.4796e-005 3.8183 0.011951 8.6689e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4212 0.49722 0.15186 0.01823 12.3704 0.11336 0.00014574 0.77679 0.0086836 0.0096353 0.0014029 0.98673 0.99157 3.0271e-006 1.2108e-005 0.15929 0.87636 0.89099 0.0014058 0.97225 0.46359 0.0018936 0.42368 1.9364 1.9352 16.0139 144.937 0.00020334 -85.5807 0.54495
6.649 0.98811 5.4796e-005 3.8183 0.011951 8.6701e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4213 0.49727 0.15188 0.018231 12.3729 0.11336 0.00014575 0.77678 0.0086841 0.0096358 0.0014028 0.98673 0.99157 3.0268e-006 1.2107e-005 0.1593 0.8767 0.89114 0.0014058 0.97241 0.46377 0.0018935 0.42369 1.9372 1.936 16.0139 144.937 0.00020311 -85.5813 0.54595
6.65 0.98811 5.4796e-005 3.8183 0.011951 8.6714e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4214 0.49731 0.15189 0.018232 12.3754 0.11337 0.00014576 0.77677 0.0086846 0.0096363 0.0014027 0.98673 0.99157 3.0265e-006 1.2106e-005 0.1593 0.87703 0.89129 0.0014057 0.97257 0.46396 0.0018935 0.4237 1.9379 1.9368 16.0139 144.9371 0.00020287 -85.5819 0.54695
6.651 0.98811 5.4796e-005 3.8183 0.011951 8.6727e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4215 0.49736 0.15191 0.018233 12.3779 0.11338 0.00014578 0.77677 0.0086851 0.0096368 0.0014025 0.98674 0.99157 3.0261e-006 1.2105e-005 0.1593 0.87736 0.89144 0.0014056 0.97273 0.46415 0.0018934 0.42372 1.9387 1.9376 16.0139 144.9371 0.00020264 -85.5825 0.54795
6.652 0.98811 5.4796e-005 3.8183 0.011951 8.674e-005 0.0011661 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4215 0.4974 0.15192 0.018235 12.3803 0.11339 0.00014579 0.77676 0.0086855 0.0096374 0.0014024 0.98674 0.99157 3.0258e-006 1.2103e-005 0.15931 0.87769 0.89159 0.0014056 0.97289 0.46433 0.0018933 0.42373 1.9395 1.9383 16.0139 144.9371 0.00020242 -85.583 0.54895
6.653 0.98811 5.4796e-005 3.8183 0.011951 8.6753e-005 0.0011662 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4216 0.49745 0.15194 0.018236 12.3828 0.1134 0.0001458 0.77675 0.008686 0.0096379 0.0014023 0.98674 0.99157 3.0255e-006 1.2102e-005 0.15931 0.87802 0.89173 0.0014055 0.97305 0.46452 0.0018932 0.42375 1.9403 1.9391 16.0138 144.9371 0.00020219 -85.5836 0.54995
6.654 0.98811 5.4796e-005 3.8183 0.011951 8.6766e-005 0.0011662 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.4217 0.49749 0.15195 0.018237 12.3853 0.1134 0.00014581 0.77674 0.0086865 0.0096384 0.0014022 0.98674 0.99157 3.0252e-006 1.2101e-005 0.15932 0.87835 0.89188 0.0014054 0.9732 0.46471 0.0018931 0.42376 1.9411 1.9399 16.0138 144.9371 0.00020196 -85.5842 0.55095
6.655 0.98811 5.4796e-005 3.8183 0.011951 8.6779e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.4218 0.49754 0.15197 0.018239 12.3878 0.11341 0.00014582 0.77674 0.008687 0.0096389 0.001402 0.98674 0.99157 3.0249e-006 1.21e-005 0.15932 0.87868 0.89203 0.0014054 0.97336 0.46489 0.001893 0.42378 1.9419 1.9407 16.0138 144.9372 0.00020173 -85.5847 0.55195
6.656 0.98811 5.4796e-005 3.8183 0.011951 8.6792e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.4219 0.49759 0.15198 0.01824 12.3903 0.11342 0.00014583 0.77673 0.0086875 0.0096394 0.0014019 0.98674 0.99157 3.0246e-006 1.2098e-005 0.15932 0.87901 0.89217 0.0014053 0.97351 0.46508 0.0018929 0.42379 1.9426 1.9415 16.0138 144.9372 0.00020151 -85.5853 0.55295
6.657 0.98811 5.4795e-005 3.8183 0.011951 8.6805e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.422 0.49763 0.15199 0.018241 12.3928 0.11343 0.00014584 0.77672 0.008688 0.00964 0.0014017 0.98675 0.99158 3.0243e-006 1.2097e-005 0.15933 0.87934 0.89232 0.0014052 0.97367 0.46526 0.0018928 0.4238 1.9434 1.9423 16.0138 144.9372 0.00020128 -85.5859 0.55395
6.658 0.98811 5.4795e-005 3.8183 0.011951 8.6817e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4221 0.49768 0.15201 0.018242 12.3952 0.11343 0.00014586 0.77671 0.0086885 0.0096405 0.0014016 0.98675 0.99158 3.024e-006 1.2096e-005 0.15933 0.87966 0.89246 0.0014051 0.97382 0.46545 0.0018927 0.42382 1.9442 1.943 16.0138 144.9372 0.00020106 -85.5864 0.55495
6.659 0.98811 5.4795e-005 3.8183 0.011951 8.683e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4222 0.49772 0.15202 0.018244 12.3977 0.11344 0.00014587 0.7767 0.0086889 0.009641 0.0014014 0.98675 0.99158 3.0237e-006 1.2095e-005 0.15934 0.87999 0.89261 0.0014051 0.97397 0.46564 0.0018926 0.42383 1.9449 1.9438 16.0137 144.9372 0.00020084 -85.587 0.55595
6.66 0.98811 5.4795e-005 3.8183 0.011951 8.6843e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4223 0.49777 0.15204 0.018245 12.4002 0.11345 0.00014588 0.7767 0.0086894 0.0096415 0.0014013 0.98675 0.99158 3.0234e-006 1.2094e-005 0.15934 0.88031 0.89275 0.001405 0.97412 0.46582 0.0018925 0.42385 1.9457 1.9446 16.0137 144.9373 0.00020061 -85.5875 0.55695
6.661 0.98811 5.4795e-005 3.8183 0.011951 8.6856e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4224 0.49782 0.15205 0.018246 12.4027 0.11346 0.00014589 0.77669 0.0086899 0.009642 0.0014011 0.98675 0.99158 3.0231e-006 1.2092e-005 0.15934 0.88063 0.8929 0.0014049 0.97427 0.46601 0.0018925 0.42386 1.9465 1.9453 16.0137 144.9373 0.00020039 -85.5881 0.55795
6.662 0.98811 5.4795e-005 3.8183 0.011951 8.6869e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4225 0.49786 0.15207 0.018248 12.4052 0.11346 0.0001459 0.77668 0.0086904 0.0096426 0.001401 0.98675 0.99158 3.0229e-006 1.2091e-005 0.15935 0.88095 0.89304 0.0014048 0.97442 0.46619 0.0018924 0.42387 1.9472 1.9461 16.0137 144.9373 0.00020017 -85.5886 0.55895
6.663 0.98811 5.4795e-005 3.8183 0.011951 8.6882e-005 0.0011662 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4225 0.49791 0.15208 0.018249 12.4077 0.11347 0.00014591 0.77667 0.0086909 0.0096431 0.0014008 0.98676 0.99158 3.0226e-006 1.209e-005 0.15935 0.88127 0.89318 0.0014048 0.97456 0.46638 0.0018923 0.42389 1.948 1.9469 16.0137 144.9373 0.00019995 -85.5891 0.55995
6.664 0.98811 5.4795e-005 3.8183 0.011951 8.6895e-005 0.0011662 0.2335 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.4226 0.49795 0.1521 0.01825 12.4102 0.11348 0.00014592 0.77667 0.0086914 0.0096436 0.0014007 0.98676 0.99158 3.0223e-006 1.2089e-005 0.15935 0.88159 0.89332 0.0014047 0.97471 0.46656 0.0018922 0.4239 1.9488 1.9476 16.0137 144.9373 0.00019973 -85.5897 0.56095
6.665 0.98811 5.4795e-005 3.8183 0.011951 8.6908e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4227 0.498 0.15211 0.018251 12.4126 0.11349 0.00014594 0.77666 0.0086919 0.0096441 0.0014005 0.98676 0.99158 3.022e-006 1.2088e-005 0.15936 0.88191 0.89346 0.0014046 0.97486 0.46675 0.0018921 0.42392 1.9495 1.9484 16.0136 144.9374 0.00019952 -85.5902 0.56195
6.666 0.98811 5.4795e-005 3.8183 0.011951 8.6921e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4228 0.49804 0.15213 0.018253 12.4151 0.1135 0.00014595 0.77665 0.0086923 0.0096446 0.0014004 0.98676 0.99159 3.0217e-006 1.2087e-005 0.15936 0.88223 0.8936 0.0014046 0.975 0.46693 0.001892 0.42393 1.9503 1.9492 16.0136 144.9374 0.0001993 -85.5907 0.56295
6.667 0.98811 5.4795e-005 3.8183 0.011951 8.6933e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4229 0.49809 0.15214 0.018254 12.4176 0.1135 0.00014596 0.77664 0.0086928 0.0096452 0.0014003 0.98676 0.99159 3.0214e-006 1.2086e-005 0.15937 0.88254 0.89374 0.0014045 0.97514 0.46712 0.0018919 0.42395 1.951 1.9499 16.0136 144.9374 0.00019908 -85.5912 0.56395
6.668 0.98811 5.4795e-005 3.8183 0.011951 8.6946e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.423 0.49814 0.15215 0.018255 12.4201 0.11351 0.00014597 0.77663 0.0086933 0.0096457 0.0014002 0.98676 0.99159 3.0212e-006 1.2085e-005 0.15937 0.88286 0.89388 0.0014044 0.97529 0.46731 0.0018919 0.42396 1.9518 1.9507 16.0136 144.9374 0.00019887 -85.5918 0.56495
6.669 0.98811 5.4795e-005 3.8183 0.011951 8.6959e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4231 0.49818 0.15217 0.018257 12.4226 0.11352 0.00014598 0.77663 0.0086938 0.0096462 0.0014001 0.98676 0.99159 3.0209e-006 1.2083e-005 0.15937 0.88317 0.89402 0.0014044 0.97543 0.46749 0.0018918 0.42397 1.9525 1.9514 16.0136 144.9374 0.00019865 -85.5923 0.56595
6.67 0.98811 5.4794e-005 3.8183 0.011951 8.6972e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4232 0.49823 0.15218 0.018258 12.4251 0.11353 0.00014599 0.77662 0.0086943 0.0096467 0.0014 0.98677 0.99159 3.0206e-006 1.2082e-005 0.15938 0.88349 0.89416 0.0014043 0.97557 0.46768 0.0018917 0.42399 1.9533 1.9522 16.0136 144.9375 0.00019844 -85.5928 0.56695
6.671 0.98811 5.4794e-005 3.8183 0.011951 8.6985e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4233 0.49827 0.1522 0.018259 12.4276 0.11353 0.000146 0.77661 0.0086948 0.0096472 0.0013999 0.98677 0.99159 3.0203e-006 1.2081e-005 0.15938 0.8838 0.8943 0.0014042 0.97571 0.46786 0.0018916 0.424 1.954 1.9529 16.0135 144.9375 0.00019823 -85.5933 0.56795
6.672 0.98811 5.4794e-005 3.8183 0.011951 8.6998e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4234 0.49832 0.15221 0.01826 12.4301 0.11354 0.00014602 0.7766 0.0086953 0.0096478 0.0013998 0.98677 0.99159 3.0201e-006 1.208e-005 0.15938 0.88411 0.89443 0.0014042 0.97585 0.46805 0.0018915 0.42402 1.9548 1.9537 16.0135 144.9375 0.00019802 -85.5938 0.56895
6.673 0.98811 5.4794e-005 3.8183 0.011951 8.7011e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4235 0.49837 0.15223 0.018262 12.4326 0.11355 0.00014603 0.7766 0.0086957 0.0096483 0.0013997 0.98677 0.99159 3.0198e-006 1.2079e-005 0.15939 0.88442 0.89457 0.0014041 0.97598 0.46823 0.0018915 0.42403 1.9555 1.9544 16.0135 144.9375 0.0001978 -85.5943 0.56995
6.674 0.98811 5.4794e-005 3.8183 0.011951 8.7024e-005 0.0011662 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.4235 0.49841 0.15224 0.018263 12.4351 0.11356 0.00014604 0.77659 0.0086962 0.0096488 0.0013996 0.98677 0.99159 3.0195e-006 1.2078e-005 0.15939 0.88473 0.89471 0.0014041 0.97612 0.46842 0.0018914 0.42405 1.9563 1.9552 16.0135 144.9375 0.00019759 -85.5948 0.57095
6.675 0.98811 5.4794e-005 3.8183 0.011951 8.7037e-005 0.0011662 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4236 0.49846 0.15226 0.018264 12.4375 0.11357 0.00014605 0.77658 0.0086967 0.0096493 0.0013995 0.98677 0.99159 3.0193e-006 1.2077e-005 0.1594 0.88504 0.89484 0.001404 0.97626 0.4686 0.0018913 0.42406 1.957 1.9559 16.0135 144.9376 0.00019738 -85.5953 0.57195
6.676 0.98811 5.4794e-005 3.8183 0.011951 8.7049e-005 0.0011662 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4237 0.4985 0.15227 0.018265 12.44 0.11357 0.00014606 0.77657 0.0086972 0.0096498 0.0013994 0.98678 0.9916 3.019e-006 1.2076e-005 0.1594 0.88535 0.89498 0.001404 0.97639 0.46879 0.0018912 0.42407 1.9577 1.9567 16.0135 144.9376 0.00019718 -85.5958 0.57295
6.677 0.98811 5.4794e-005 3.8183 0.011951 8.7062e-005 0.0011662 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4238 0.49855 0.15229 0.018267 12.4425 0.11358 0.00014607 0.77656 0.0086977 0.0096504 0.0013993 0.98678 0.9916 3.0188e-006 1.2075e-005 0.1594 0.88565 0.89511 0.0014039 0.97653 0.46897 0.0018911 0.42409 1.9585 1.9574 16.0134 144.9376 0.00019697 -85.5963 0.57395
6.678 0.98811 5.4794e-005 3.8183 0.011951 8.7075e-005 0.0011663 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4239 0.49859 0.1523 0.018268 12.445 0.11359 0.00014608 0.77656 0.0086982 0.0096509 0.0013992 0.98678 0.9916 3.0185e-006 1.2074e-005 0.15941 0.88596 0.89525 0.0014039 0.97666 0.46916 0.0018911 0.4241 1.9592 1.9581 16.0134 144.9376 0.00019676 -85.5967 0.57495
6.679 0.98811 5.4794e-005 3.8183 0.011951 8.7088e-005 0.0011663 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.424 0.49864 0.15231 0.018269 12.4475 0.1136 0.0001461 0.77655 0.0086986 0.0096514 0.0013991 0.98678 0.9916 3.0182e-006 1.2073e-005 0.15941 0.88626 0.89538 0.0014038 0.97679 0.46934 0.001891 0.42412 1.9599 1.9589 16.0134 144.9377 0.00019655 -85.5972 0.57595
6.68 0.98811 5.4794e-005 3.8183 0.011951 8.7101e-005 0.0011663 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4241 0.49869 0.15233 0.018271 12.45 0.1136 0.00014611 0.77654 0.0086991 0.0096519 0.0013989 0.98678 0.9916 3.018e-006 1.2072e-005 0.15941 0.88657 0.89551 0.0014037 0.97693 0.46952 0.0018909 0.42413 1.9607 1.9596 16.0134 144.9377 0.00019635 -85.5977 0.57695
6.681 0.98811 5.4794e-005 3.8183 0.011951 8.7114e-005 0.0011663 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4242 0.49873 0.15234 0.018272 12.4525 0.11361 0.00014612 0.77653 0.0086996 0.0096524 0.0013988 0.98678 0.9916 3.0177e-006 1.2071e-005 0.15942 0.88687 0.89564 0.0014037 0.97706 0.46971 0.0018908 0.42414 1.9614 1.9603 16.0134 144.9377 0.00019614 -85.5982 0.57795
6.682 0.98811 5.4793e-005 3.8183 0.011951 8.7127e-005 0.0011663 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4243 0.49878 0.15236 0.018273 12.455 0.11362 0.00014613 0.77653 0.0087001 0.009653 0.0013987 0.98678 0.9916 3.0175e-006 1.207e-005 0.15942 0.88717 0.89578 0.0014036 0.97719 0.46989 0.0018908 0.42416 1.9621 1.9611 16.0134 144.9377 0.00019594 -85.5986 0.57895
6.683 0.98811 5.4793e-005 3.8183 0.011951 8.714e-005 0.0011663 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4244 0.49882 0.15237 0.018274 12.4575 0.11363 0.00014614 0.77652 0.0087006 0.0096535 0.0013986 0.98679 0.9916 3.0172e-006 1.2069e-005 0.15943 0.88747 0.89591 0.0014036 0.97732 0.47008 0.0018907 0.42417 1.9629 1.9618 16.0133 144.9377 0.00019574 -85.5991 0.57995
6.684 0.98811 5.4793e-005 3.8183 0.011951 8.7152e-005 0.0011663 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4245 0.49887 0.15239 0.018276 12.46 0.11364 0.00014615 0.77651 0.0087011 0.009654 0.0013985 0.98679 0.9916 3.017e-006 1.2068e-005 0.15943 0.88777 0.89604 0.0014035 0.97745 0.47026 0.0018906 0.42419 1.9636 1.9625 16.0133 144.9378 0.00019553 -85.5996 0.58095
6.685 0.98811 5.4793e-005 3.8183 0.011951 8.7165e-005 0.0011663 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4245 0.49892 0.1524 0.018277 12.4625 0.11364 0.00014616 0.7765 0.0087015 0.0096545 0.0013983 0.98679 0.9916 3.0167e-006 1.2067e-005 0.15943 0.88807 0.89617 0.0014035 0.97757 0.47045 0.0018905 0.4242 1.9643 1.9632 16.0133 144.9378 0.00019533 -85.6 0.58195
6.686 0.98811 5.4793e-005 3.8183 0.011951 8.7178e-005 0.0011663 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.4246 0.49896 0.15242 0.018278 12.465 0.11365 0.00014618 0.7765 0.008702 0.009655 0.0013982 0.98679 0.9916 3.0165e-006 1.2066e-005 0.15944 0.88837 0.8963 0.0014034 0.9777 0.47063 0.0018905 0.42422 1.965 1.964 16.0133 144.9378 0.00019513 -85.6005 0.58295
6.687 0.98811 5.4793e-005 3.8183 0.011951 8.7191e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4247 0.49901 0.15243 0.01828 12.4675 0.11366 0.00014619 0.77649 0.0087025 0.0096556 0.0013981 0.98679 0.99161 3.0163e-006 1.2065e-005 0.15944 0.88867 0.89643 0.0014033 0.97783 0.47082 0.0018904 0.42423 1.9657 1.9647 16.0133 144.9378 0.00019493 -85.6009 0.58395
6.688 0.98811 5.4793e-005 3.8183 0.011951 8.7204e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4248 0.49905 0.15244 0.018281 12.47 0.11367 0.0001462 0.77648 0.008703 0.0096561 0.001398 0.98679 0.99161 3.016e-006 1.2064e-005 0.15944 0.88897 0.89656 0.0014033 0.97795 0.471 0.0018903 0.42424 1.9665 1.9654 16.0132 144.9378 0.00019473 -85.6014 0.58495
6.689 0.98811 5.4793e-005 3.8183 0.01195 8.7217e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4249 0.4991 0.15246 0.018282 12.4724 0.11367 0.00014621 0.77647 0.0087035 0.0096566 0.0013979 0.98679 0.99161 3.0158e-006 1.2063e-005 0.15945 0.88926 0.89669 0.0014032 0.97808 0.47118 0.0018902 0.42426 1.9672 1.9661 16.0132 144.9379 0.00019453 -85.6018 0.58595
6.69 0.98811 5.4793e-005 3.8183 0.01195 8.723e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.425 0.49914 0.15247 0.018283 12.4749 0.11368 0.00014622 0.77646 0.008704 0.0096571 0.0013978 0.98679 0.99161 3.0155e-006 1.2062e-005 0.15945 0.88955 0.89681 0.0014032 0.9782 0.47137 0.0018902 0.42427 1.9679 1.9668 16.0132 144.9379 0.00019434 -85.6023 0.58695
6.691 0.98811 5.4793e-005 3.8183 0.01195 8.7243e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4251 0.49919 0.15249 0.018285 12.4774 0.11369 0.00014623 0.77646 0.0087044 0.0096576 0.0013977 0.9868 0.99161 3.0153e-006 1.2061e-005 0.15946 0.88985 0.89694 0.0014031 0.97832 0.47155 0.0018901 0.42429 1.9686 1.9675 16.0132 144.9379 0.00019414 -85.6027 0.58795
6.692 0.98811 5.4793e-005 3.8183 0.01195 8.7256e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4252 0.49924 0.1525 0.018286 12.4799 0.1137 0.00014624 0.77645 0.0087049 0.0096581 0.0013976 0.9868 0.99161 3.0151e-006 1.206e-005 0.15946 0.89014 0.89707 0.001403 0.97845 0.47174 0.00189 0.4243 1.9693 1.9683 16.0132 144.9379 0.00019394 -85.6032 0.58895
6.693 0.98811 5.4793e-005 3.8183 0.01195 8.7268e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4253 0.49928 0.15252 0.018287 12.4824 0.1137 0.00014626 0.77644 0.0087054 0.0096587 0.0013975 0.9868 0.99161 3.0148e-006 1.2059e-005 0.15946 0.89043 0.89719 0.001403 0.97857 0.47192 0.00189 0.42432 1.97 1.969 16.0132 144.9379 0.00019375 -85.6036 0.58995
6.694 0.98811 5.4793e-005 3.8183 0.01195 8.7281e-005 0.0011663 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.4254 0.49933 0.15253 0.018288 12.4849 0.11371 0.00014627 0.77643 0.0087059 0.0096592 0.0013974 0.9868 0.99161 3.0146e-006 1.2058e-005 0.15947 0.89072 0.89732 0.0014029 0.97869 0.4721 0.0018899 0.42433 1.9707 1.9697 16.0131 144.938 0.00019355 -85.604 0.59095
6.695 0.98811 5.4792e-005 3.8183 0.01195 8.7294e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.4255 0.49937 0.15255 0.01829 12.4874 0.11372 0.00014628 0.77643 0.0087064 0.0096597 0.0013973 0.9868 0.99161 3.0144e-006 1.2057e-005 0.15947 0.89101 0.89745 0.0014029 0.97881 0.47229 0.0018898 0.42434 1.9714 1.9704 16.0131 144.938 0.00019336 -85.6045 0.59195
6.696 0.98811 5.4792e-005 3.8183 0.01195 8.7307e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.4255 0.49942 0.15256 0.018291 12.4899 0.11373 0.00014629 0.77642 0.0087069 0.0096602 0.0013972 0.9868 0.99161 3.0142e-006 1.2057e-005 0.15947 0.8913 0.89757 0.0014028 0.97893 0.47247 0.0018898 0.42436 1.9721 1.9711 16.0131 144.938 0.00019316 -85.6049 0.59295
6.697 0.98811 5.4792e-005 3.8183 0.01195 8.732e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.4256 0.49947 0.15258 0.018292 12.4924 0.11374 0.0001463 0.77641 0.0087073 0.0096607 0.0013971 0.9868 0.99161 3.0139e-006 1.2056e-005 0.15948 0.89159 0.8977 0.0014028 0.97904 0.47265 0.0018897 0.42437 1.9728 1.9718 16.0131 144.938 0.00019297 -85.6053 0.59395
6.698 0.98811 5.4792e-005 3.8183 0.01195 8.7333e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.4257 0.49951 0.15259 0.018294 12.4949 0.11374 0.00014631 0.7764 0.0087078 0.0096613 0.001397 0.98681 0.99161 3.0137e-006 1.2055e-005 0.15948 0.89188 0.89782 0.0014027 0.97916 0.47284 0.0018896 0.42439 1.9735 1.9725 16.0131 144.938 0.00019278 -85.6057 0.59495
6.699 0.98811 5.4792e-005 3.8183 0.01195 8.7346e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4258 0.49956 0.1526 0.018295 12.4974 0.11375 0.00014632 0.7764 0.0087083 0.0096618 0.0013969 0.98681 0.99162 3.0135e-006 1.2054e-005 0.15949 0.89216 0.89794 0.0014027 0.97928 0.47302 0.0018896 0.4244 1.9742 1.9732 16.013 144.9381 0.00019259 -85.6061 0.59595
6.7 0.98811 5.4792e-005 3.8183 0.01195 8.7359e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4259 0.4996 0.15262 0.018296 12.4999 0.11376 0.00014633 0.77639 0.0087088 0.0096623 0.0013968 0.98681 0.99162 3.0133e-006 1.2053e-005 0.15949 0.89245 0.89807 0.0014026 0.97939 0.4732 0.0018895 0.42441 1.9749 1.9739 16.013 144.9381 0.0001924 -85.6066 0.59695
6.701 0.98811 5.4792e-005 3.8183 0.01195 8.7372e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.426 0.49965 0.15263 0.018297 12.5024 0.11377 0.00014635 0.77638 0.0087093 0.0096628 0.0013967 0.98681 0.99162 3.013e-006 1.2052e-005 0.15949 0.89273 0.89819 0.0014026 0.97951 0.47339 0.0018894 0.42443 1.9756 1.9746 16.013 144.9381 0.00019221 -85.607 0.59795
6.702 0.98811 5.4792e-005 3.8183 0.01195 8.7384e-005 0.0011663 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4261 0.49969 0.15265 0.018299 12.5049 0.11377 0.00014636 0.77637 0.0087098 0.0096633 0.0013966 0.98681 0.99162 3.0128e-006 1.2051e-005 0.1595 0.89302 0.89831 0.0014025 0.97962 0.47357 0.0018894 0.42444 1.9763 1.9753 16.013 144.9381 0.00019202 -85.6074 0.59895
6.703 0.98811 5.4792e-005 3.8183 0.01195 8.7397e-005 0.0011664 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4262 0.49974 0.15266 0.0183 12.5074 0.11378 0.00014637 0.77636 0.0087102 0.0096638 0.0013966 0.98681 0.99162 3.0126e-006 1.205e-005 0.1595 0.8933 0.89843 0.0014025 0.97974 0.47375 0.0018893 0.42446 1.977 1.976 16.013 144.9381 0.00019183 -85.6078 0.59995
6.704 0.98811 5.4792e-005 3.8183 0.01195 8.741e-005 0.0011664 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4263 0.49979 0.15268 0.018301 12.5099 0.11379 0.00014638 0.77636 0.0087107 0.0096644 0.0013965 0.98681 0.99162 3.0124e-006 1.205e-005 0.1595 0.89358 0.89856 0.0014024 0.97985 0.47394 0.0018892 0.42447 1.9777 1.9767 16.0129 144.9382 0.00019164 -85.6082 0.60095
6.705 0.98811 5.4792e-005 3.8183 0.01195 8.7423e-005 0.0011664 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4264 0.49983 0.15269 0.018302 12.5124 0.1138 0.00014639 0.77635 0.0087112 0.0096649 0.0013964 0.98681 0.99162 3.0122e-006 1.2049e-005 0.15951 0.89386 0.89868 0.0014024 0.97996 0.47412 0.0018892 0.42449 1.9783 1.9773 16.0129 144.9382 0.00019146 -85.6086 0.60195
6.706 0.98811 5.4792e-005 3.8183 0.01195 8.7436e-005 0.0011664 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4264 0.49988 0.15271 0.018304 12.5149 0.11381 0.0001464 0.77634 0.0087117 0.0096654 0.0013963 0.98682 0.99162 3.012e-006 1.2048e-005 0.15951 0.89414 0.8988 0.0014024 0.98007 0.4743 0.0018891 0.4245 1.979 1.978 16.0129 144.9382 0.00019127 -85.609 0.60295
6.707 0.98811 5.4792e-005 3.8183 0.01195 8.7449e-005 0.0011664 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4265 0.49992 0.15272 0.018305 12.5174 0.11381 0.00014641 0.77633 0.0087122 0.0096659 0.0013962 0.98682 0.99162 3.0118e-006 1.2047e-005 0.15952 0.89442 0.89892 0.0014023 0.98019 0.47449 0.001889 0.42451 1.9797 1.9787 16.0129 144.9382 0.00019108 -85.6094 0.60395
6.708 0.98811 5.4791e-005 3.8183 0.01195 8.7462e-005 0.0011664 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.4266 0.49997 0.15273 0.018306 12.5199 0.11382 0.00014643 0.77633 0.0087126 0.0096664 0.0013961 0.98682 0.99162 3.0116e-006 1.2046e-005 0.15952 0.8947 0.89904 0.0014023 0.9803 0.47467 0.001889 0.42453 1.9804 1.9794 16.0129 144.9382 0.0001909 -85.6098 0.60495
6.709 0.98811 5.4791e-005 3.8183 0.01195 8.7475e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.4267 0.50001 0.15275 0.018308 12.5224 0.11383 0.00014644 0.77632 0.0087131 0.0096669 0.001396 0.98682 0.99162 3.0113e-006 1.2045e-005 0.15952 0.89498 0.89916 0.0014022 0.98041 0.47485 0.0018889 0.42454 1.9811 1.9801 16.0129 144.9383 0.00019072 -85.6102 0.60595
6.71 0.98811 5.4791e-005 3.8183 0.01195 8.7488e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.4268 0.50006 0.15276 0.018309 12.5249 0.11384 0.00014645 0.77631 0.0087136 0.0096675 0.0013959 0.98682 0.99162 3.0111e-006 1.2044e-005 0.15953 0.89526 0.89927 0.0014022 0.98051 0.47503 0.0018888 0.42456 1.9818 1.9808 16.0128 144.9383 0.00019053 -85.6105 0.60695
6.711 0.98811 5.4791e-005 3.8183 0.01195 8.75e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.4269 0.50011 0.15278 0.01831 12.5274 0.11384 0.00014646 0.7763 0.0087141 0.009668 0.0013958 0.98682 0.99162 3.0109e-006 1.2044e-005 0.15953 0.89553 0.89939 0.0014021 0.98062 0.47522 0.0018888 0.42457 1.9824 1.9814 16.0128 144.9383 0.00019035 -85.6109 0.60795
6.712 0.98811 5.4791e-005 3.8183 0.01195 8.7513e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.427 0.50015 0.15279 0.018311 12.5299 0.11385 0.00014647 0.77629 0.0087146 0.0096685 0.0013957 0.98682 0.99163 3.0107e-006 1.2043e-005 0.15953 0.89581 0.89951 0.0014021 0.98073 0.4754 0.0018887 0.42458 1.9831 1.9821 16.0128 144.9383 0.00019017 -85.6113 0.60895
6.713 0.98811 5.4791e-005 3.8183 0.01195 8.7526e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.4271 0.5002 0.15281 0.018313 12.5324 0.11386 0.00014648 0.77629 0.0087151 0.009669 0.0013956 0.98682 0.99163 3.0105e-006 1.2042e-005 0.15954 0.89608 0.89963 0.001402 0.98084 0.47558 0.0018887 0.4246 1.9838 1.9828 16.0128 144.9383 0.00018999 -85.6117 0.60995
6.714 0.98811 5.4791e-005 3.8183 0.01195 8.7539e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.4272 0.50024 0.15282 0.018314 12.535 0.11387 0.00014649 0.77628 0.0087155 0.0096695 0.0013955 0.98682 0.99163 3.0103e-006 1.2041e-005 0.15954 0.89635 0.89974 0.001402 0.98094 0.47576 0.0018886 0.42461 1.9844 1.9835 16.0128 144.9384 0.0001898 -85.6121 0.61095
6.715 0.98811 5.4791e-005 3.8183 0.01195 8.7552e-005 0.0011664 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.4273 0.50029 0.15284 0.018315 12.5375 0.11387 0.00014651 0.77627 0.008716 0.00967 0.0013954 0.98683 0.99163 3.0101e-006 1.204e-005 0.15955 0.89663 0.89986 0.0014019 0.98105 0.47595 0.0018885 0.42463 1.9851 1.9841 16.0127 144.9384 0.00018962 -85.6124 0.61195
6.716 0.98811 5.4791e-005 3.8183 0.01195 8.7565e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4274 0.50034 0.15285 0.018317 12.54 0.11388 0.00014652 0.77626 0.0087165 0.0096706 0.0013953 0.98683 0.99163 3.0099e-006 1.204e-005 0.15955 0.8969 0.89998 0.0014019 0.98115 0.47613 0.0018885 0.42464 1.9858 1.9848 16.0127 144.9384 0.00018945 -85.6128 0.61295
6.717 0.98811 5.4791e-005 3.8183 0.01195 8.7578e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4274 0.50038 0.15287 0.018318 12.5425 0.11389 0.00014653 0.77626 0.008717 0.0096711 0.0013952 0.98683 0.99163 3.0097e-006 1.2039e-005 0.15955 0.89717 0.90009 0.0014018 0.98126 0.47631 0.0018884 0.42466 1.9865 1.9855 16.0127 144.9384 0.00018927 -85.6132 0.61395
6.718 0.98811 5.4791e-005 3.8183 0.01195 8.7591e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4275 0.50043 0.15288 0.018319 12.545 0.1139 0.00014654 0.77625 0.0087175 0.0096716 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.15956 0.89744 0.90021 0.0014018 0.98136 0.47649 0.0018884 0.42467 1.9871 1.9861 16.0127 144.9384 0.00018909 -85.6135 0.61495
6.719 0.98811 5.4791e-005 3.8183 0.01195 8.7603e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4276 0.50047 0.15289 0.01832 12.5475 0.11391 0.00014655 0.77624 0.0087179 0.0096721 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.15956 0.89771 0.90032 0.0014017 0.98146 0.47668 0.0018883 0.42468 1.9878 1.9868 16.0127 144.9385 0.00018891 -85.6139 0.61595
6.72 0.98811 5.4791e-005 3.8183 0.01195 8.7616e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4277 0.50052 0.15291 0.018322 12.55 0.11391 0.00014656 0.77623 0.0087184 0.0096726 0.001395 0.98683 0.99163 3.0092e-006 1.2037e-005 0.15956 0.89797 0.90044 0.0014017 0.98156 0.47686 0.0018882 0.4247 1.9884 1.9875 16.0126 144.9385 0.00018873 -85.6143 0.61695
6.721 0.98811 5.479e-005 3.8183 0.01195 8.7629e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4278 0.50056 0.15292 0.018323 12.5525 0.11392 0.00014657 0.77623 0.0087189 0.0096731 0.0013949 0.98683 0.99163 3.009e-006 1.2036e-005 0.15957 0.89824 0.90055 0.0014016 0.98166 0.47704 0.0018882 0.42471 1.9891 1.9881 16.0126 144.9385 0.00018856 -85.6146 0.61795
6.722 0.98811 5.479e-005 3.8183 0.01195 8.7642e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4279 0.50061 0.15294 0.018324 12.555 0.11393 0.00014659 0.77622 0.0087194 0.0096737 0.0013948 0.98683 0.99163 3.0088e-006 1.2035e-005 0.15957 0.89851 0.90066 0.0014016 0.98177 0.47722 0.0018881 0.42473 1.9898 1.9888 16.0126 144.9385 0.00018838 -85.615 0.61895
6.723 0.98811 5.479e-005 3.8183 0.01195 8.7655e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.428 0.50066 0.15295 0.018325 12.5575 0.11394 0.0001466 0.77621 0.0087199 0.0096742 0.0013948 0.98683 0.99163 3.0086e-006 1.2034e-005 0.15958 0.89877 0.90078 0.0014016 0.98186 0.4774 0.0018881 0.42474 1.9904 1.9895 16.0126 144.9385 0.00018821 -85.6153 0.61995
6.724 0.98811 5.479e-005 3.8183 0.01195 8.7668e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4281 0.5007 0.15297 0.018327 12.56 0.11394 0.00014661 0.7762 0.0087203 0.0096747 0.0013947 0.98684 0.99163 3.0084e-006 1.2034e-005 0.15958 0.89904 0.90089 0.0014015 0.98196 0.47759 0.001888 0.42475 1.9911 1.9901 16.0125 144.9386 0.00018803 -85.6157 0.62095
6.725 0.98811 5.479e-005 3.8183 0.01195 8.7681e-005 0.0011664 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4282 0.50075 0.15298 0.018328 12.5625 0.11395 0.00014662 0.77619 0.0087208 0.0096752 0.0013946 0.98684 0.99163 3.0082e-006 1.2033e-005 0.15958 0.8993 0.901 0.0014015 0.98206 0.47777 0.001888 0.42477 1.9917 1.9908 16.0125 144.9386 0.00018786 -85.616 0.62195
6.726 0.98811 5.479e-005 3.8183 0.01195 8.7694e-005 0.0011664 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4283 0.50079 0.153 0.018329 12.565 0.11396 0.00014663 0.77619 0.0087213 0.0096757 0.0013945 0.98684 0.99164 3.008e-006 1.2032e-005 0.15959 0.89957 0.90111 0.0014014 0.98216 0.47795 0.0018879 0.42478 1.9924 1.9914 16.0125 144.9386 0.00018769 -85.6164 0.62295
6.727 0.98811 5.479e-005 3.8183 0.01195 8.7707e-005 0.0011664 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4284 0.50084 0.15301 0.018331 12.5675 0.11397 0.00014664 0.77618 0.0087218 0.0096762 0.0013945 0.98684 0.99164 3.0079e-006 1.2031e-005 0.15959 0.89983 0.90122 0.0014014 0.98226 0.47813 0.0018879 0.4248 1.993 1.9921 16.0125 144.9386 0.00018752 -85.6167 0.62395
6.728 0.98811 5.479e-005 3.8183 0.01195 8.7719e-005 0.0011665 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4284 0.50089 0.15302 0.018332 12.57 0.11397 0.00014665 0.77617 0.0087223 0.0096767 0.0013944 0.98684 0.99164 3.0077e-006 1.2031e-005 0.15959 0.90009 0.90133 0.0014013 0.98236 0.47831 0.0018878 0.42481 1.9937 1.9927 16.0125 144.9386 0.00018734 -85.6171 0.62495
6.729 0.98811 5.479e-005 3.8183 0.01195 8.7732e-005 0.0011665 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4285 0.50093 0.15304 0.018333 12.5726 0.11398 0.00014666 0.77616 0.0087228 0.0096773 0.0013943 0.98684 0.99164 3.0075e-006 1.203e-005 0.1596 0.90035 0.90145 0.0014013 0.98245 0.47849 0.0018877 0.42482 1.9943 1.9934 16.0124 144.9387 0.00018717 -85.6174 0.62595
6.73 0.98811 5.479e-005 3.8183 0.01195 8.7745e-005 0.0011665 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.4286 0.50098 0.15305 0.018334 12.5751 0.11399 0.00014668 0.77616 0.0087232 0.0096778 0.0013942 0.98684 0.99164 3.0073e-006 1.2029e-005 0.1596 0.90061 0.90156 0.0014013 0.98255 0.47868 0.0018877 0.42484 1.995 1.994 16.0124 144.9387 0.000187 -85.6177 0.62695
6.731 0.98811 5.479e-005 3.8183 0.01195 8.7758e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.4287 0.50102 0.15307 0.018336 12.5776 0.114 0.00014669 0.77615 0.0087237 0.0096783 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.15961 0.90087 0.90166 0.0014012 0.98264 0.47886 0.0018876 0.42485 1.9956 1.9947 16.0124 144.9387 0.00018683 -85.6181 0.62795
6.732 0.98811 5.479e-005 3.8183 0.01195 8.7771e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.4288 0.50107 0.15308 0.018337 12.5801 0.11401 0.0001467 0.77614 0.0087242 0.0096788 0.0013941 0.98684 0.99164 3.007e-006 1.2028e-005 0.15961 0.90113 0.90177 0.0014012 0.98274 0.47904 0.0018876 0.42487 1.9963 1.9953 16.0124 144.9387 0.00018666 -85.6184 0.62895
6.733 0.98811 5.4789e-005 3.8183 0.01195 8.7784e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.4289 0.50111 0.1531 0.018338 12.5826 0.11401 0.00014671 0.77613 0.0087247 0.0096793 0.001394 0.98684 0.99164 3.0068e-006 1.2027e-005 0.15961 0.90138 0.90188 0.0014012 0.98283 0.47922 0.0018875 0.42488 1.9969 1.996 16.0124 144.9387 0.0001865 -85.6187 0.62995
6.734 0.98811 5.4789e-005 3.8183 0.01195 8.7797e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.429 0.50116 0.15311 0.018339 12.5851 0.11402 0.00014672 0.77613 0.0087252 0.0096798 0.0013939 0.98685 0.99164 3.0066e-006 1.2026e-005 0.15962 0.90164 0.90199 0.0014011 0.98292 0.4794 0.0018875 0.42489 1.9975 1.9966 16.0123 144.9388 0.00018633 -85.6191 0.63095
6.735 0.98811 5.4789e-005 3.8183 0.01195 8.781e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.4291 0.50121 0.15313 0.018341 12.5876 0.11403 0.00014673 0.77612 0.0087256 0.0096803 0.0013938 0.98685 0.99164 3.0064e-006 1.2026e-005 0.15962 0.9019 0.9021 0.0014011 0.98302 0.47958 0.0018874 0.42491 1.9982 1.9972 16.0123 144.9388 0.00018616 -85.6194 0.63195
6.736 0.98811 5.4789e-005 3.8183 0.01195 8.7823e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.4292 0.50125 0.15314 0.018342 12.5901 0.11404 0.00014674 0.77611 0.0087261 0.0096809 0.0013938 0.98685 0.99164 3.0063e-006 1.2025e-005 0.15962 0.90215 0.90221 0.001401 0.98311 0.47976 0.0018874 0.42492 1.9988 1.9979 16.0123 144.9388 0.000186 -85.6197 0.63295
6.737 0.98811 5.4789e-005 3.8183 0.01195 8.7835e-005 0.0011665 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.4293 0.5013 0.15315 0.018343 12.5926 0.11404 0.00014676 0.7761 0.0087266 0.0096814 0.0013937 0.98685 0.99164 3.0061e-006 1.2024e-005 0.15963 0.90241 0.90231 0.001401 0.9832 0.47995 0.0018873 0.42494 1.9994 1.9985 16.0123 144.9388 0.00018583 -85.62 0.63395
6.738 0.98811 5.4789e-005 3.8183 0.01195 8.7848e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.4294 0.50134 0.15317 0.018345 12.5952 0.11405 0.00014677 0.77609 0.0087271 0.0096819 0.0013936 0.98685 0.99164 3.0059e-006 1.2024e-005 0.15963 0.90266 0.90242 0.001401 0.98329 0.48013 0.0018873 0.42495 2.0001 1.9992 16.0123 144.9388 0.00018566 -85.6203 0.63495
6.739 0.98811 5.4789e-005 3.8183 0.01195 8.7861e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.4294 0.50139 0.15318 0.018346 12.5977 0.11406 0.00014678 0.77609 0.0087275 0.0096824 0.0013935 0.98685 0.99164 3.0058e-006 1.2023e-005 0.15964 0.90291 0.90253 0.0014009 0.98338 0.48031 0.0018872 0.42497 2.0007 1.9998 16.0122 144.9389 0.0001855 -85.6207 0.63595
6.74 0.98811 5.4789e-005 3.8183 0.01195 8.7874e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.4295 0.50143 0.1532 0.018347 12.6002 0.11407 0.00014679 0.77608 0.008728 0.0096829 0.0013934 0.98685 0.99164 3.0056e-006 1.2022e-005 0.15964 0.90316 0.90263 0.0014009 0.98347 0.48049 0.0018872 0.42498 2.0013 2.0004 16.0122 144.9389 0.00018534 -85.621 0.63695
6.741 0.98811 5.4789e-005 3.8183 0.01195 8.7887e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.4296 0.50148 0.15321 0.018348 12.6027 0.11407 0.0001468 0.77607 0.0087285 0.0096834 0.0013934 0.98685 0.99164 3.0054e-006 1.2022e-005 0.15964 0.90342 0.90274 0.0014008 0.98356 0.48067 0.0018871 0.42499 2.002 2.0011 16.0122 144.9389 0.00018517 -85.6213 0.63795
6.742 0.98811 5.4789e-005 3.8183 0.01195 8.79e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4297 0.50153 0.15323 0.01835 12.6052 0.11408 0.00014681 0.77606 0.008729 0.0096839 0.0013933 0.98685 0.99165 3.0053e-006 1.2021e-005 0.15965 0.90367 0.90284 0.0014008 0.98365 0.48085 0.0018871 0.42501 2.0026 2.0017 16.0122 144.9389 0.00018501 -85.6216 0.63895
6.743 0.98811 5.4789e-005 3.8183 0.01195 8.7913e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4298 0.50157 0.15324 0.018351 12.6077 0.11409 0.00014682 0.77606 0.0087295 0.0096845 0.0013932 0.98685 0.99165 3.0051e-006 1.202e-005 0.15965 0.90392 0.90295 0.0014008 0.98373 0.48103 0.001887 0.42502 2.0032 2.0023 16.0121 144.9389 0.00018485 -85.6219 0.63995
6.744 0.98811 5.4789e-005 3.8183 0.01195 8.7926e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4299 0.50162 0.15326 0.018352 12.6102 0.1141 0.00014683 0.77605 0.0087299 0.009685 0.0013932 0.98685 0.99165 3.0049e-006 1.202e-005 0.15965 0.90416 0.90305 0.0014007 0.98382 0.48121 0.001887 0.42504 2.0038 2.0029 16.0121 144.939 0.00018469 -85.6222 0.64095
6.745 0.98811 5.4789e-005 3.8183 0.01195 8.7938e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.43 0.50166 0.15327 0.018353 12.6128 0.11411 0.00014685 0.77604 0.0087304 0.0096855 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.15966 0.90441 0.90316 0.0014007 0.98391 0.48139 0.0018869 0.42505 2.0045 2.0036 16.0121 144.939 0.00018452 -85.6225 0.64195
6.746 0.98811 5.4788e-005 3.8183 0.01195 8.7951e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4301 0.50171 0.15328 0.018355 12.6153 0.11411 0.00014686 0.77603 0.0087309 0.009686 0.0013931 0.98686 0.99165 3.0046e-006 1.2018e-005 0.15966 0.90466 0.90326 0.0014006 0.98399 0.48157 0.0018869 0.42506 2.0051 2.0042 16.0121 144.939 0.00018436 -85.6228 0.64295
6.747 0.98811 5.4788e-005 3.8183 0.01195 8.7964e-005 0.0011665 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4302 0.50176 0.1533 0.018356 12.6178 0.11412 0.00014687 0.77603 0.0087314 0.0096865 0.001393 0.98686 0.99165 3.0044e-006 1.2018e-005 0.15967 0.90491 0.90336 0.0014006 0.98408 0.48175 0.0018868 0.42508 2.0057 2.0048 16.0121 144.939 0.0001842 -85.6231 0.64395
6.748 0.98811 5.4788e-005 3.8183 0.011949 8.7977e-005 0.0011665 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4303 0.5018 0.15331 0.018357 12.6203 0.11413 0.00014688 0.77602 0.0087319 0.009687 0.0013929 0.98686 0.99165 3.0043e-006 1.2017e-005 0.15967 0.90515 0.90347 0.0014006 0.98416 0.48193 0.0018868 0.42509 2.0063 2.0054 16.012 144.939 0.00018405 -85.6234 0.64495
6.749 0.98811 5.4788e-005 3.8183 0.011949 8.799e-005 0.0011665 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4303 0.50185 0.15333 0.018358 12.6228 0.11414 0.00014689 0.77601 0.0087323 0.0096875 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.15967 0.9054 0.90357 0.0014005 0.98425 0.48211 0.0018867 0.42511 2.0069 2.0061 16.012 144.9391 0.00018389 -85.6237 0.64595
6.75 0.98811 5.4788e-005 3.8183 0.011949 8.8003e-005 0.0011665 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4304 0.50189 0.15334 0.01836 12.6253 0.11414 0.0001469 0.776 0.0087328 0.0096881 0.0013928 0.98686 0.99165 3.004e-006 1.2016e-005 0.15968 0.90564 0.90367 0.0014005 0.98433 0.48229 0.0018867 0.42512 2.0076 2.0067 16.012 144.9391 0.00018373 -85.624 0.64695
6.751 0.98811 5.4788e-005 3.8183 0.011949 8.8016e-005 0.0011665 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4305 0.50194 0.15336 0.018361 12.6279 0.11415 0.00014691 0.776 0.0087333 0.0096886 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.15968 0.90588 0.90377 0.0014005 0.98442 0.48247 0.0018866 0.42513 2.0082 2.0073 16.012 144.9391 0.00018357 -85.6243 0.64795
6.752 0.98811 5.4788e-005 3.8183 0.011949 8.8029e-005 0.0011665 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4306 0.50198 0.15337 0.018362 12.6304 0.11416 0.00014693 0.77599 0.0087338 0.0096891 0.0013926 0.98686 0.99165 3.0037e-006 1.2015e-005 0.15968 0.90613 0.90388 0.0014004 0.9845 0.48265 0.0018866 0.42515 2.0088 2.0079 16.0119 144.9391 0.00018341 -85.6246 0.64895
6.753 0.98811 5.4788e-005 3.8183 0.011949 8.8042e-005 0.0011666 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4307 0.50203 0.15339 0.018364 12.6329 0.11417 0.00014694 0.77598 0.0087343 0.0096896 0.0013926 0.98686 0.99165 3.0035e-006 1.2014e-005 0.15969 0.90637 0.90398 0.0014004 0.98458 0.48283 0.0018866 0.42516 2.0094 2.0085 16.0119 144.9391 0.00018326 -85.6249 0.64995
6.754 0.98811 5.4788e-005 3.8183 0.011949 8.8054e-005 0.0011666 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.4308 0.50208 0.1534 0.018365 12.6354 0.11417 0.00014695 0.77597 0.0087347 0.0096901 0.0013925 0.98686 0.99165 3.0034e-006 1.2013e-005 0.15969 0.90661 0.90408 0.0014004 0.98466 0.48301 0.0018865 0.42518 2.01 2.0091 16.0119 144.9392 0.0001831 -85.6251 0.65095
6.755 0.98811 5.4788e-005 3.8183 0.011949 8.8067e-005 0.0011666 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.4309 0.50212 0.15342 0.018366 12.6379 0.11418 0.00014696 0.77596 0.0087352 0.0096906 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.1597 0.90685 0.90418 0.0014003 0.98474 0.48319 0.0018865 0.42519 2.0106 2.0097 16.0119 144.9392 0.00018295 -85.6254 0.65195
6.756 0.98811 5.4788e-005 3.8183 0.011949 8.808e-005 0.0011666 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.431 0.50217 0.15343 0.018367 12.6404 0.11419 0.00014697 0.77596 0.0087357 0.0096911 0.0013924 0.98687 0.99165 3.0031e-006 1.2012e-005 0.1597 0.90709 0.90428 0.0014003 0.98482 0.48337 0.0018864 0.4252 2.0112 2.0103 16.0119 144.9392 0.00018279 -85.6257 0.65295
6.757 0.98811 5.4788e-005 3.8183 0.011949 8.8093e-005 0.0011666 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.4311 0.50221 0.15344 0.018369 12.643 0.1142 0.00014698 0.77595 0.0087362 0.0096916 0.0013923 0.98687 0.99165 3.0029e-006 1.2012e-005 0.1597 0.90733 0.90438 0.0014003 0.98491 0.48355 0.0018864 0.42522 2.0118 2.011 16.0118 144.9392 0.00018264 -85.626 0.65395
6.758 0.98811 5.4788e-005 3.8183 0.011949 8.8106e-005 0.0011666 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.4312 0.50226 0.15346 0.01837 12.6455 0.11421 0.00014699 0.77594 0.0087366 0.0096922 0.0013922 0.98687 0.99165 3.0028e-006 1.2011e-005 0.15971 0.90757 0.90448 0.0014002 0.98498 0.48373 0.0018863 0.42523 2.0124 2.0116 16.0118 144.9392 0.00018248 -85.6263 0.65495
6.759 0.98811 5.4787e-005 3.8183 0.011949 8.8119e-005 0.0011666 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.4313 0.5023 0.15347 0.018371 12.648 0.11421 0.000147 0.77593 0.0087371 0.0096927 0.0013922 0.98687 0.99166 3.0026e-006 1.201e-005 0.15971 0.9078 0.90457 0.0014002 0.98506 0.48391 0.0018863 0.42525 2.013 2.0122 16.0118 144.9393 0.00018233 -85.6265 0.65595
6.76 0.98811 5.4787e-005 3.8183 0.011949 8.8132e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4313 0.50235 0.15349 0.018372 12.6505 0.11422 0.00014702 0.77593 0.0087376 0.0096932 0.0013921 0.98687 0.99166 3.0025e-006 1.201e-005 0.15971 0.90804 0.90467 0.0014002 0.98514 0.48409 0.0018862 0.42526 2.0136 2.0128 16.0118 144.9393 0.00018218 -85.6268 0.65695
6.761 0.98811 5.4787e-005 3.8183 0.011949 8.8145e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4314 0.5024 0.1535 0.018374 12.653 0.11423 0.00014703 0.77592 0.0087381 0.0096937 0.001392 0.98687 0.99166 3.0023e-006 1.2009e-005 0.15972 0.90828 0.90477 0.0014001 0.98522 0.48427 0.0018862 0.42527 2.0142 2.0134 16.0117 144.9393 0.00018203 -85.6271 0.65795
6.762 0.98811 5.4787e-005 3.8183 0.011949 8.8157e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4315 0.50244 0.15352 0.018375 12.6556 0.11424 0.00014704 0.77591 0.0087386 0.0096942 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.15972 0.90851 0.90487 0.0014001 0.9853 0.48445 0.0018862 0.42529 2.0148 2.014 16.0117 144.9393 0.00018188 -85.6273 0.65895
6.763 0.98811 5.4787e-005 3.8183 0.011949 8.817e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4316 0.50249 0.15353 0.018376 12.6581 0.11424 0.00014705 0.7759 0.008739 0.0096947 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.15973 0.90875 0.90497 0.0014001 0.98538 0.48463 0.0018861 0.4253 2.0154 2.0146 16.0117 144.9393 0.00018173 -85.6276 0.65995
6.764 0.98811 5.4787e-005 3.8183 0.011949 8.8183e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4317 0.50253 0.15355 0.018378 12.6606 0.11425 0.00014706 0.7759 0.0087395 0.0096952 0.0013918 0.98687 0.99166 3.0019e-006 1.2008e-005 0.15973 0.90898 0.90506 0.0014 0.98545 0.48481 0.0018861 0.42532 2.016 2.0152 16.0117 144.9394 0.00018158 -85.6279 0.66095
6.765 0.98811 5.4787e-005 3.8183 0.011949 8.8196e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4318 0.50258 0.15356 0.018379 12.6631 0.11426 0.00014707 0.77589 0.00874 0.0096957 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.15973 0.90921 0.90516 0.0014 0.98553 0.48499 0.001886 0.42533 2.0166 2.0158 16.0116 144.9394 0.00018143 -85.6281 0.66195
6.766 0.98811 5.4787e-005 3.8183 0.011949 8.8209e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4319 0.50263 0.15357 0.01838 12.6656 0.11427 0.00014708 0.77588 0.0087405 0.0096963 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.15974 0.90944 0.90526 0.0014 0.9856 0.48517 0.001886 0.42534 2.0172 2.0164 16.0116 144.9394 0.00018128 -85.6284 0.66295
6.767 0.98811 5.4787e-005 3.8183 0.011949 8.8222e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.432 0.50267 0.15359 0.018381 12.6682 0.11427 0.0001471 0.77587 0.0087409 0.0096968 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.15974 0.90968 0.90535 0.0013999 0.98568 0.48535 0.0018859 0.42536 2.0178 2.017 16.0116 144.9394 0.00018113 -85.6287 0.66395
6.768 0.98811 5.4787e-005 3.8183 0.011949 8.8235e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4321 0.50272 0.1536 0.018383 12.6707 0.11428 0.00014711 0.77586 0.0087414 0.0096973 0.0013916 0.98688 0.99166 3.0014e-006 1.2005e-005 0.15974 0.90991 0.90545 0.0013999 0.98575 0.48553 0.0018859 0.42537 2.0184 2.0175 16.0116 144.9395 0.00018098 -85.6289 0.66495
6.769 0.98811 5.4787e-005 3.8183 0.011949 8.8248e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4322 0.50276 0.15362 0.018384 12.6732 0.11429 0.00014712 0.77586 0.0087419 0.0096978 0.0013916 0.98688 0.99166 3.0012e-006 1.2005e-005 0.15975 0.91014 0.90554 0.0013999 0.98583 0.48571 0.0018859 0.42539 2.019 2.0181 16.0116 144.9395 0.00018083 -85.6292 0.66595
6.77 0.98811 5.4787e-005 3.8183 0.011949 8.8261e-005 0.0011666 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4322 0.50281 0.15363 0.018385 12.6757 0.1143 0.00014713 0.77585 0.0087424 0.0096983 0.0013915 0.98688 0.99166 3.0011e-006 1.2004e-005 0.15975 0.91037 0.90564 0.0013998 0.9859 0.48589 0.0018858 0.4254 2.0196 2.0187 16.0115 144.9395 0.00018069 -85.6294 0.66695
6.771 0.98811 5.4786e-005 3.8183 0.011949 8.8273e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4323 0.50285 0.15365 0.018386 12.6783 0.11431 0.00014714 0.77584 0.0087429 0.0096988 0.0013914 0.98688 0.99166 3.001e-006 1.2004e-005 0.15975 0.91059 0.90573 0.0013998 0.98597 0.48607 0.0018858 0.42541 2.0202 2.0193 16.0115 144.9395 0.00018054 -85.6297 0.66795
6.772 0.98811 5.4786e-005 3.8183 0.011949 8.8286e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4324 0.5029 0.15366 0.018388 12.6808 0.11431 0.00014715 0.77583 0.0087433 0.0096993 0.0013914 0.98688 0.99166 3.0008e-006 1.2003e-005 0.15976 0.91082 0.90583 0.0013998 0.98605 0.48625 0.0018857 0.42543 2.0207 2.0199 16.0115 144.9395 0.00018039 -85.6299 0.66895
6.773 0.98811 5.4786e-005 3.8183 0.011949 8.8299e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4325 0.50295 0.15368 0.018389 12.6833 0.11432 0.00014716 0.77583 0.0087438 0.0096998 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.15976 0.91105 0.90592 0.0013997 0.98612 0.48642 0.0018857 0.42544 2.0213 2.0205 16.0115 144.9396 0.00018025 -85.6302 0.66995
6.774 0.98811 5.4786e-005 3.8183 0.011949 8.8312e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4326 0.50299 0.15369 0.01839 12.6858 0.11433 0.00014717 0.77582 0.0087443 0.0097003 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.15977 0.91128 0.90601 0.0013997 0.98619 0.4866 0.0018857 0.42546 2.0219 2.0211 16.0114 144.9396 0.0001801 -85.6304 0.67095
6.775 0.98811 5.4786e-005 3.8183 0.011949 8.8325e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4327 0.50304 0.1537 0.018391 12.6884 0.11434 0.00014719 0.77581 0.0087448 0.0097009 0.0013912 0.98688 0.99166 3.0004e-006 1.2002e-005 0.15977 0.9115 0.90611 0.0013997 0.98626 0.48678 0.0018856 0.42547 2.0225 2.0216 16.0114 144.9396 0.00017996 -85.6307 0.67195
6.776 0.98811 5.4786e-005 3.8183 0.011949 8.8338e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4328 0.50308 0.15372 0.018393 12.6909 0.11434 0.0001472 0.7758 0.0087452 0.0097014 0.0013912 0.98688 0.99166 3.0003e-006 1.2001e-005 0.15977 0.91173 0.9062 0.0013996 0.98633 0.48696 0.0018856 0.42548 2.0231 2.0222 16.0114 144.9396 0.00017982 -85.6309 0.67295
6.777 0.98811 5.4786e-005 3.8183 0.011949 8.8351e-005 0.0011666 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.4329 0.50313 0.15373 0.018394 12.6934 0.11435 0.00014721 0.7758 0.0087457 0.0097019 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.15978 0.91195 0.90629 0.0013996 0.9864 0.48714 0.0018855 0.4255 2.0236 2.0228 16.0114 144.9396 0.00017967 -85.6312 0.67395
6.778 0.98811 5.4786e-005 3.8183 0.011949 8.8364e-005 0.0011667 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.433 0.50317 0.15375 0.018395 12.6959 0.11436 0.00014722 0.77579 0.0087462 0.0097024 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.15978 0.91217 0.90638 0.0013996 0.98647 0.48732 0.0018855 0.42551 2.0242 2.0234 16.0113 144.9397 0.00017953 -85.6314 0.67495
6.779 0.98811 5.4786e-005 3.8183 0.011949 8.8377e-005 0.0011667 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.4331 0.50322 0.15376 0.018396 12.6985 0.11437 0.00014723 0.77578 0.0087467 0.0097029 0.001391 0.98688 0.99167 2.9999e-006 1.2e-005 0.15978 0.9124 0.90648 0.0013996 0.98654 0.4875 0.0018855 0.42553 2.0248 2.024 16.0113 144.9397 0.00017939 -85.6316 0.67595
6.78 0.98811 5.4786e-005 3.8183 0.011949 8.8389e-005 0.0011667 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.4332 0.50327 0.15378 0.018398 12.701 0.11437 0.00014724 0.77577 0.0087471 0.0097034 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.15979 0.91262 0.90657 0.0013995 0.98661 0.48767 0.0018854 0.42554 2.0254 2.0245 16.0113 144.9397 0.00017925 -85.6319 0.67695
6.781 0.98811 5.4786e-005 3.8183 0.011949 8.8402e-005 0.0011667 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.4332 0.50331 0.15379 0.018399 12.7035 0.11438 0.00014725 0.77577 0.0087476 0.0097039 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.15979 0.91284 0.90666 0.0013995 0.98668 0.48785 0.0018854 0.42555 2.0259 2.0251 16.0113 144.9397 0.00017911 -85.6321 0.67795
6.782 0.98811 5.4786e-005 3.8183 0.011949 8.8415e-005 0.0011667 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.4333 0.50336 0.15381 0.0184 12.706 0.11439 0.00014727 0.77576 0.0087481 0.0097044 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.1598 0.91306 0.90675 0.0013995 0.98675 0.48803 0.0018853 0.42557 2.0265 2.0257 16.0112 144.9397 0.00017896 -85.6323 0.67895
6.783 0.98811 5.4786e-005 3.8183 0.011949 8.8428e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.4334 0.5034 0.15382 0.018402 12.7086 0.1144 0.00014728 0.77575 0.0087486 0.0097049 0.0013908 0.98689 0.99167 2.9994e-006 1.1998e-005 0.1598 0.91328 0.90684 0.0013995 0.98682 0.48821 0.0018853 0.42558 2.0271 2.0263 16.0112 144.9398 0.00017882 -85.6326 0.67995
6.784 0.98811 5.4785e-005 3.8183 0.011949 8.8441e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.4335 0.50345 0.15383 0.018403 12.7111 0.1144 0.00014729 0.77574 0.008749 0.0097055 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.1598 0.9135 0.90693 0.0013994 0.98688 0.48839 0.0018853 0.42559 2.0276 2.0268 16.0112 144.9398 0.00017869 -85.6328 0.68095
6.785 0.98811 5.4785e-005 3.8183 0.011949 8.8454e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.4336 0.50349 0.15385 0.018404 12.7136 0.11441 0.0001473 0.77573 0.0087495 0.009706 0.0013906 0.98689 0.99167 2.9992e-006 1.1997e-005 0.15981 0.91372 0.90702 0.0013994 0.98695 0.48857 0.0018852 0.42561 2.0282 2.0274 16.0112 144.9398 0.00017855 -85.633 0.68195
6.786 0.98811 5.4785e-005 3.8183 0.011949 8.8467e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.4337 0.50354 0.15386 0.018405 12.7162 0.11442 0.00014731 0.77573 0.00875 0.0097065 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.15981 0.91394 0.90711 0.0013994 0.98702 0.48874 0.0018852 0.42562 2.0288 2.028 16.0112 144.9398 0.00017841 -85.6333 0.68295
6.787 0.98811 5.4785e-005 3.8183 0.011949 8.848e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.4338 0.50359 0.15388 0.018407 12.7187 0.11443 0.00014732 0.77572 0.0087505 0.009707 0.0013905 0.98689 0.99167 2.9989e-006 1.1996e-005 0.15981 0.91416 0.9072 0.0013994 0.98708 0.48892 0.0018852 0.42564 2.0293 2.0285 16.0111 144.9398 0.00017827 -85.6335 0.68395
6.788 0.98811 5.4785e-005 3.8183 0.011949 8.8492e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4339 0.50363 0.15389 0.018408 12.7212 0.11444 0.00014733 0.77571 0.008751 0.0097075 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.15982 0.91437 0.90729 0.0013993 0.98715 0.4891 0.0018851 0.42565 2.0299 2.0291 16.0111 144.9399 0.00017813 -85.6337 0.68495
6.789 0.98811 5.4785e-005 3.8183 0.011949 8.8505e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.434 0.50368 0.15391 0.018409 12.7238 0.11444 0.00014734 0.7757 0.0087514 0.009708 0.0013904 0.98689 0.99167 2.9987e-006 1.1995e-005 0.15982 0.91459 0.90738 0.0013993 0.98721 0.48928 0.0018851 0.42566 2.0305 2.0297 16.0111 144.9399 0.00017799 -85.6339 0.68595
6.79 0.98811 5.4785e-005 3.8183 0.011949 8.8518e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4341 0.50372 0.15392 0.01841 12.7263 0.11445 0.00014736 0.7757 0.0087519 0.0097085 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.15983 0.9148 0.90746 0.0013993 0.98728 0.48946 0.0018851 0.42568 2.031 2.0302 16.0111 144.9399 0.00017786 -85.6342 0.68695
6.791 0.98811 5.4785e-005 3.8183 0.011949 8.8531e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4341 0.50377 0.15394 0.018412 12.7288 0.11446 0.00014737 0.77569 0.0087524 0.009709 0.0013903 0.98689 0.99167 2.9985e-006 1.1994e-005 0.15983 0.91502 0.90755 0.0013992 0.98734 0.48963 0.001885 0.42569 2.0316 2.0308 16.011 144.9399 0.00017772 -85.6344 0.68795
6.792 0.98811 5.4785e-005 3.8183 0.011949 8.8544e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4342 0.50381 0.15395 0.018413 12.7313 0.11447 0.00014738 0.77568 0.0087529 0.0097095 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.15983 0.91523 0.90764 0.0013992 0.98741 0.48981 0.001885 0.42571 2.0321 2.0314 16.011 144.9399 0.00017759 -85.6346 0.68895
6.793 0.98811 5.4785e-005 3.8183 0.011949 8.8557e-005 0.0011667 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4343 0.50386 0.15396 0.018414 12.7339 0.11447 0.00014739 0.77567 0.0087533 0.00971 0.0013902 0.98689 0.99167 2.9982e-006 1.1993e-005 0.15984 0.91545 0.90773 0.0013992 0.98747 0.48999 0.001885 0.42572 2.0327 2.0319 16.011 144.94 0.00017745 -85.6348 0.68995
6.794 0.98811 5.4785e-005 3.8183 0.011949 8.857e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4344 0.50391 0.15398 0.018415 12.7364 0.11448 0.0001474 0.77567 0.0087538 0.0097106 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.15984 0.91566 0.90781 0.0013991 0.98753 0.49017 0.0018849 0.42573 2.0333 2.0325 16.011 144.94 0.00017732 -85.635 0.69095
6.795 0.98811 5.4785e-005 3.8183 0.011949 8.8583e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4345 0.50395 0.15399 0.018417 12.7389 0.11449 0.00014741 0.77566 0.0087543 0.0097111 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.15984 0.91587 0.9079 0.0013991 0.9876 0.49034 0.0018849 0.42575 2.0338 2.033 16.0109 144.94 0.00017718 -85.6352 0.69195
6.796 0.98811 5.4785e-005 3.8183 0.011949 8.8595e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4346 0.504 0.15401 0.018418 12.7415 0.1145 0.00014742 0.77565 0.0087548 0.0097116 0.0013901 0.98689 0.99167 2.9979e-006 1.1991e-005 0.15985 0.91608 0.90799 0.0013991 0.98766 0.49052 0.0018849 0.42576 2.0344 2.0336 16.0109 144.94 0.00017705 -85.6355 0.69295
6.797 0.98811 5.4784e-005 3.8183 0.011949 8.8608e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4347 0.50404 0.15402 0.018419 12.744 0.1145 0.00014743 0.77564 0.0087552 0.0097121 0.0013901 0.9869 0.99167 2.9978e-006 1.1991e-005 0.15985 0.91629 0.90807 0.0013991 0.98772 0.4907 0.0018848 0.42578 2.0349 2.0341 16.0109 144.94 0.00017692 -85.6357 0.69395
6.798 0.98811 5.4784e-005 3.8183 0.011949 8.8621e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4348 0.50409 0.15404 0.018421 12.7465 0.11451 0.00014745 0.77564 0.0087557 0.0097126 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.15986 0.9165 0.90816 0.001399 0.98778 0.49088 0.0018848 0.42579 2.0355 2.0347 16.0109 144.9401 0.00017678 -85.6359 0.69495
6.799 0.98811 5.4784e-005 3.8183 0.011949 8.8634e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4349 0.50414 0.15405 0.018422 12.7491 0.11452 0.00014746 0.77563 0.0087562 0.0097131 0.00139 0.9869 0.99167 2.9976e-006 1.199e-005 0.15986 0.91671 0.90824 0.001399 0.98784 0.49105 0.0018848 0.4258 2.036 2.0352 16.0108 144.9401 0.00017665 -85.6361 0.69595
6.8 0.98811 5.4784e-005 3.8183 0.011949 8.8647e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.435 0.50418 0.15407 0.018423 12.7516 0.11453 0.00014747 0.77562 0.0087567 0.0097136 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.15986 0.91692 0.90833 0.001399 0.9879 0.49123 0.0018847 0.42582 2.0366 2.0358 16.0108 144.9401 0.00017652 -85.6363 0.69695
6.801 0.98811 5.4784e-005 3.8183 0.011949 8.866e-005 0.0011667 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4351 0.50423 0.15408 0.018424 12.7541 0.11453 0.00014748 0.77561 0.0087571 0.0097141 0.0013899 0.9869 0.99167 2.9973e-006 1.1989e-005 0.15987 0.91713 0.90841 0.0013989 0.98796 0.49141 0.0018847 0.42583 2.0371 2.0363 16.0108 144.9401 0.00017639 -85.6365 0.69795
6.802 0.98811 5.4784e-005 3.8183 0.011949 8.8673e-005 0.0011668 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4351 0.50427 0.15409 0.018426 12.7567 0.11454 0.00014749 0.77561 0.0087576 0.0097146 0.0013898 0.9869 0.99167 2.9972e-006 1.1989e-005 0.15987 0.91734 0.9085 0.0013989 0.98802 0.49159 0.0018847 0.42584 2.0377 2.0369 16.0108 144.9401 0.00017626 -85.6367 0.69895
6.803 0.98811 5.4784e-005 3.8183 0.011949 8.8686e-005 0.0011668 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.4352 0.50432 0.15411 0.018427 12.7592 0.11455 0.0001475 0.7756 0.0087581 0.0097151 0.0013898 0.9869 0.99168 2.9971e-006 1.1988e-005 0.15987 0.91755 0.90858 0.0013989 0.98808 0.49176 0.0018846 0.42586 2.0382 2.0374 16.0107 144.9402 0.00017613 -85.6369 0.69995
6.804 0.98811 5.4784e-005 3.8183 0.011949 8.8699e-005 0.0011668 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.4353 0.50436 0.15412 0.018428 12.7617 0.11456 0.00014751 0.77559 0.0087586 0.0097156 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.15988 0.91775 0.90867 0.0013989 0.98814 0.49194 0.0018846 0.42587 2.0387 2.038 16.0107 144.9402 0.000176 -85.6371 0.70095
6.805 0.98811 5.4784e-005 3.8183 0.011949 8.8711e-005 0.0011668 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.4354 0.50441 0.15414 0.018429 12.7643 0.11457 0.00014752 0.77558 0.008759 0.0097162 0.0013897 0.9869 0.99168 2.9969e-006 1.1988e-005 0.15988 0.91796 0.90875 0.0013989 0.9882 0.49212 0.0018846 0.42589 2.0393 2.0385 16.0107 144.9402 0.00017587 -85.6373 0.70195
6.806 0.98811 5.4784e-005 3.8183 0.011949 8.8724e-005 0.0011668 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.4355 0.50446 0.15415 0.018431 12.7668 0.11457 0.00014754 0.77557 0.0087595 0.0097167 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.15988 0.91816 0.90883 0.0013988 0.98826 0.49229 0.0018845 0.4259 2.0398 2.0391 16.0107 144.9402 0.00017574 -85.6375 0.70295
6.807 0.98811 5.4784e-005 3.8183 0.011948 8.8737e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4356 0.5045 0.15417 0.018432 12.7694 0.11458 0.00014755 0.77557 0.00876 0.0097172 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.15989 0.91837 0.90892 0.0013988 0.98832 0.49247 0.0018845 0.42591 2.0404 2.0396 16.0106 144.9402 0.00017561 -85.6377 0.70395
6.808 0.98811 5.4784e-005 3.8183 0.011948 8.875e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4357 0.50455 0.15418 0.018433 12.7719 0.11459 0.00014756 0.77556 0.0087604 0.0097177 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.15989 0.91857 0.909 0.0013988 0.98837 0.49265 0.0018845 0.42593 2.0409 2.0401 16.0106 144.9403 0.00017548 -85.6379 0.70495
6.809 0.98811 5.4783e-005 3.8183 0.011948 8.8763e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4358 0.50459 0.15419 0.018434 12.7744 0.1146 0.00014757 0.77555 0.0087609 0.0097182 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.1599 0.91877 0.90908 0.0013988 0.98843 0.49282 0.0018844 0.42594 2.0414 2.0407 16.0106 144.9403 0.00017535 -85.6381 0.70595
6.81 0.98811 5.4783e-005 3.8183 0.011948 8.8776e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4359 0.50464 0.15421 0.018436 12.777 0.1146 0.00014758 0.77554 0.0087614 0.0097187 0.0013894 0.9869 0.99168 2.9964e-006 1.1985e-005 0.1599 0.91898 0.90916 0.0013988 0.98849 0.493 0.0018844 0.42596 2.042 2.0412 16.0106 144.9403 0.00017523 -85.6383 0.70695
6.811 0.98811 5.4783e-005 3.8183 0.011948 8.8789e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.436 0.50468 0.15422 0.018437 12.7795 0.11461 0.00014759 0.77554 0.0087619 0.0097192 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.1599 0.91918 0.90925 0.0013987 0.98855 0.49318 0.0018844 0.42597 2.0425 2.0418 16.0105 144.9403 0.0001751 -85.6385 0.70795
6.812 0.98811 5.4783e-005 3.8183 0.011948 8.8802e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.436 0.50473 0.15424 0.018438 12.782 0.11462 0.0001476 0.77553 0.0087623 0.0097197 0.0013893 0.9869 0.99168 2.9962e-006 1.1985e-005 0.15991 0.91938 0.90933 0.0013987 0.9886 0.49335 0.0018843 0.42598 2.0431 2.0423 16.0105 144.9403 0.00017497 -85.6387 0.70895
6.813 0.98811 5.4783e-005 3.8183 0.011948 8.8814e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4361 0.50478 0.15425 0.018439 12.7846 0.11463 0.00014761 0.77552 0.0087628 0.0097202 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.15991 0.91958 0.90941 0.0013987 0.98866 0.49353 0.0018843 0.426 2.0436 2.0428 16.0105 144.9404 0.00017485 -85.6388 0.70995
6.814 0.98811 5.4783e-005 3.8183 0.011948 8.8827e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4362 0.50482 0.15427 0.018441 12.7871 0.11463 0.00014763 0.77551 0.0087633 0.0097207 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.15991 0.91978 0.90949 0.0013987 0.98871 0.49371 0.0018843 0.42601 2.0441 2.0434 16.0105 144.9404 0.00017472 -85.639 0.71095
6.815 0.98811 5.4783e-005 3.8183 0.011948 8.884e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4363 0.50487 0.15428 0.018442 12.7897 0.11464 0.00014764 0.77551 0.0087638 0.0097212 0.0013892 0.98691 0.99168 2.9959e-006 1.1983e-005 0.15992 0.91998 0.90957 0.0013987 0.98877 0.49388 0.0018842 0.42602 2.0446 2.0439 16.0104 144.9404 0.0001746 -85.6392 0.71195
6.816 0.98811 5.4783e-005 3.8183 0.011948 8.8853e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4364 0.50491 0.1543 0.018443 12.7922 0.11465 0.00014765 0.7755 0.0087642 0.0097217 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.15992 0.92018 0.90965 0.0013986 0.98882 0.49406 0.0018842 0.42604 2.0452 2.0444 16.0104 144.9404 0.00017447 -85.6394 0.71295
6.817 0.98811 5.4783e-005 3.8183 0.011948 8.8866e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4365 0.50496 0.15431 0.018444 12.7947 0.11466 0.00014766 0.77549 0.0087647 0.0097223 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.15993 0.92037 0.90973 0.0013986 0.98888 0.49424 0.0018842 0.42605 2.0457 2.045 16.0104 144.9405 0.00017435 -85.6396 0.71395
6.818 0.98811 5.4783e-005 3.8183 0.011948 8.8879e-005 0.0011668 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4366 0.505 0.15432 0.018446 12.7973 0.11466 0.00014767 0.77548 0.0087652 0.0097228 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.15993 0.92057 0.90981 0.0013986 0.98893 0.49441 0.0018842 0.42607 2.0462 2.0455 16.0103 144.9405 0.00017423 -85.6398 0.71495
6.819 0.98811 5.4783e-005 3.8183 0.011948 8.8892e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4367 0.50505 0.15434 0.018447 12.7998 0.11467 0.00014768 0.77548 0.0087657 0.0097233 0.0013891 0.98691 0.99168 2.9955e-006 1.1982e-005 0.15993 0.92077 0.90989 0.0013985 0.98898 0.49459 0.0018841 0.42608 2.0468 2.046 16.0103 144.9405 0.0001741 -85.64 0.71595
6.82 0.98811 5.4783e-005 3.8183 0.011948 8.8905e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4368 0.5051 0.15435 0.018448 12.8024 0.11468 0.00014769 0.77547 0.0087661 0.0097238 0.001389 0.98691 0.99168 2.9954e-006 1.1982e-005 0.15994 0.92096 0.90997 0.0013985 0.98904 0.49476 0.0018841 0.42609 2.0473 2.0465 16.0103 144.9405 0.00017398 -85.6401 0.71695
6.821 0.98811 5.4783e-005 3.8183 0.011948 8.8918e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4369 0.50514 0.15437 0.01845 12.8049 0.11469 0.00014771 0.77546 0.0087666 0.0097243 0.001389 0.98691 0.99168 2.9953e-006 1.1981e-005 0.15994 0.92116 0.91005 0.0013985 0.98909 0.49494 0.0018841 0.42611 2.0478 2.0471 16.0103 144.9405 0.00017386 -85.6403 0.71795
6.822 0.98811 5.4782e-005 3.8183 0.011948 8.893e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4369 0.50519 0.15438 0.018451 12.8074 0.11469 0.00014772 0.77545 0.0087671 0.0097248 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.15994 0.92135 0.91013 0.0013985 0.98914 0.49512 0.001884 0.42612 2.0483 2.0476 16.0102 144.9406 0.00017374 -85.6405 0.71895
6.823 0.98811 5.4782e-005 3.8183 0.011948 8.8943e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.437 0.50523 0.1544 0.018452 12.81 0.1147 0.00014773 0.77545 0.0087676 0.0097253 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.15995 0.92155 0.9102 0.0013984 0.98919 0.49529 0.001884 0.42613 2.0488 2.0481 16.0102 144.9406 0.00017362 -85.6407 0.71995
6.824 0.98811 5.4782e-005 3.8183 0.011948 8.8956e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4371 0.50528 0.15441 0.018453 12.8125 0.11471 0.00014774 0.77544 0.008768 0.0097258 0.0013889 0.98691 0.99168 2.995e-006 1.198e-005 0.15995 0.92174 0.91028 0.0013984 0.98925 0.49547 0.001884 0.42615 2.0494 2.0486 16.0102 144.9406 0.00017349 -85.6408 0.72095
6.825 0.98811 5.4782e-005 3.8183 0.011948 8.8969e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4372 0.50532 0.15443 0.018455 12.8151 0.11472 0.00014775 0.77543 0.0087685 0.0097263 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.15995 0.92194 0.91036 0.0013984 0.9893 0.49564 0.001884 0.42616 2.0499 2.0492 16.0102 144.9406 0.00017337 -85.641 0.72195
6.826 0.98811 5.4782e-005 3.8183 0.011948 8.8982e-005 0.0011668 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4373 0.50537 0.15444 0.018456 12.8176 0.11473 0.00014776 0.77542 0.008769 0.0097268 0.0013888 0.98691 0.99168 2.9949e-006 1.1979e-005 0.15996 0.92213 0.91044 0.0013984 0.98935 0.49582 0.0018839 0.42618 2.0504 2.0497 16.0101 144.9406 0.00017325 -85.6412 0.72295
6.827 0.98811 5.4782e-005 3.8183 0.011948 8.8995e-005 0.0011669 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4374 0.50542 0.15445 0.018457 12.8201 0.11473 0.00014777 0.77541 0.0087694 0.0097273 0.0013887 0.98691 0.99168 2.9948e-006 1.1979e-005 0.15996 0.92232 0.91051 0.0013984 0.9894 0.49599 0.0018839 0.42619 2.0509 2.0502 16.0101 144.9407 0.00017313 -85.6414 0.72395
6.828 0.98811 5.4782e-005 3.8183 0.011948 8.9008e-005 0.0011669 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.4375 0.50546 0.15447 0.018458 12.8227 0.11474 0.00014778 0.77541 0.0087699 0.0097278 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.15997 0.92251 0.91059 0.0013983 0.98945 0.49617 0.0018839 0.4262 2.0514 2.0507 16.0101 144.9407 0.00017302 -85.6415 0.72495
6.829 0.98811 5.4782e-005 3.8183 0.011948 8.9021e-005 0.0011669 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.4376 0.50551 0.15448 0.01846 12.8252 0.11475 0.0001478 0.7754 0.0087704 0.0097283 0.0013886 0.98691 0.99168 2.9946e-006 1.1978e-005 0.15997 0.9227 0.91067 0.0013983 0.9895 0.49634 0.0018839 0.42622 2.052 2.0512 16.0101 144.9407 0.0001729 -85.6417 0.72595
6.83 0.98811 5.4782e-005 3.8183 0.011948 8.9033e-005 0.0011669 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.4377 0.50555 0.1545 0.018461 12.8278 0.11476 0.00014781 0.77539 0.0087709 0.0097288 0.0013886 0.98691 0.99168 2.9945e-006 1.1978e-005 0.15997 0.92289 0.91074 0.0013983 0.98955 0.49652 0.0018838 0.42623 2.0525 2.0517 16.01 144.9407 0.00017278 -85.6419 0.72695
6.831 0.98811 5.4782e-005 3.8183 0.011948 8.9046e-005 0.0011669 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.4378 0.5056 0.15451 0.018462 12.8303 0.11476 0.00014782 0.77538 0.0087713 0.0097294 0.0013886 0.98691 0.99169 2.9944e-006 1.1978e-005 0.15998 0.92308 0.91082 0.0013983 0.9896 0.4967 0.0018838 0.42624 2.053 2.0523 16.01 144.9407 0.00017266 -85.642 0.72795
6.832 0.98811 5.4782e-005 3.8183 0.011948 8.9059e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.4379 0.50564 0.15453 0.018463 12.8329 0.11477 0.00014783 0.77538 0.0087718 0.0097299 0.0013885 0.98691 0.99169 2.9943e-006 1.1977e-005 0.15998 0.92327 0.9109 0.0013983 0.98965 0.49687 0.0018838 0.42626 2.0535 2.0528 16.01 144.9408 0.00017254 -85.6422 0.72895
6.833 0.98811 5.4782e-005 3.8183 0.011948 8.9072e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.4379 0.50569 0.15454 0.018465 12.8354 0.11478 0.00014784 0.77537 0.0087723 0.0097304 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.15998 0.92346 0.91097 0.0013983 0.9897 0.49705 0.0018837 0.42627 2.054 2.0533 16.01 144.9408 0.00017243 -85.6424 0.72995
6.834 0.98811 5.4782e-005 3.8183 0.011948 8.9085e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.438 0.50574 0.15456 0.018466 12.838 0.11479 0.00014785 0.77536 0.0087728 0.0097309 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.15999 0.92365 0.91105 0.0013983 0.98975 0.49722 0.0018837 0.42629 2.0545 2.0538 16.0099 144.9408 0.00017231 -85.6425 0.73095
6.835 0.98811 5.4781e-005 3.8183 0.011948 8.9098e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.4381 0.50578 0.15457 0.018467 12.8405 0.11479 0.00014786 0.77535 0.0087732 0.0097314 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.15999 0.92383 0.91112 0.0013983 0.9898 0.4974 0.0018837 0.4263 2.055 2.0543 16.0099 144.9408 0.00017219 -85.6427 0.73195
6.836 0.98811 5.4781e-005 3.8183 0.011948 8.9111e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.4382 0.50583 0.15458 0.018468 12.8431 0.1148 0.00014787 0.77535 0.0087737 0.0097319 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.16 0.92402 0.9112 0.0013983 0.98984 0.49757 0.0018837 0.42631 2.0555 2.0548 16.0099 144.9408 0.00017208 -85.6428 0.73295
6.837 0.98811 5.4781e-005 3.8183 0.011948 8.9124e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4383 0.50587 0.1546 0.01847 12.8456 0.11481 0.00014789 0.77534 0.0087742 0.0097324 0.0013883 0.98692 0.99169 2.9939e-006 1.1975e-005 0.16 0.92421 0.91127 0.0013982 0.98989 0.49775 0.0018836 0.42633 2.056 2.0553 16.0098 144.9409 0.00017196 -85.643 0.73395
6.838 0.98811 5.4781e-005 3.8183 0.011948 8.9136e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4384 0.50592 0.15461 0.018471 12.8481 0.11482 0.0001479 0.77533 0.0087746 0.0097329 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.16 0.92439 0.91135 0.0013982 0.98994 0.49792 0.0018836 0.42634 2.0565 2.0558 16.0098 144.9409 0.00017185 -85.6432 0.73495
6.839 0.98811 5.4781e-005 3.8183 0.011948 8.9149e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4385 0.50596 0.15463 0.018472 12.8507 0.11482 0.00014791 0.77532 0.0087751 0.0097334 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.16001 0.92458 0.91142 0.0013982 0.98999 0.4981 0.0018836 0.42635 2.057 2.0563 16.0098 144.9409 0.00017173 -85.6433 0.73595
6.84 0.98811 5.4781e-005 3.8183 0.011948 8.9162e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4386 0.50601 0.15464 0.018473 12.8532 0.11483 0.00014792 0.77532 0.0087756 0.0097339 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16001 0.92476 0.91149 0.0013981 0.99003 0.49827 0.0018836 0.42637 2.0575 2.0568 16.0098 144.9409 0.00017162 -85.6435 0.73695
6.841 0.98811 5.4781e-005 3.8183 0.011948 8.9175e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4387 0.50606 0.15466 0.018475 12.8558 0.11484 0.00014793 0.77531 0.0087761 0.0097344 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16001 0.92494 0.91157 0.0013981 0.99008 0.49845 0.0018835 0.42638 2.058 2.0573 16.0097 144.9409 0.0001715 -85.6436 0.73795
6.842 0.98811 5.4781e-005 3.8183 0.011948 8.9188e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4388 0.5061 0.15467 0.018476 12.8583 0.11485 0.00014794 0.7753 0.0087765 0.0097349 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.16002 0.92513 0.91164 0.0013981 0.99012 0.49862 0.0018835 0.42639 2.0585 2.0578 16.0097 144.941 0.00017139 -85.6438 0.73895
6.843 0.98811 5.4781e-005 3.8183 0.011948 8.9201e-005 0.0011669 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4388 0.50615 0.15468 0.018477 12.8609 0.11485 0.00014795 0.77529 0.008777 0.0097354 0.0013881 0.98692 0.99169 2.9934e-006 1.1973e-005 0.16002 0.92531 0.91171 0.0013981 0.99017 0.4988 0.0018835 0.42641 2.059 2.0583 16.0097 144.941 0.00017128 -85.6439 0.73995
6.844 0.98811 5.4781e-005 3.8183 0.011948 8.9214e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4389 0.50619 0.1547 0.018478 12.8634 0.11486 0.00014796 0.77529 0.0087775 0.0097359 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.16002 0.92549 0.91179 0.001398 0.99022 0.49897 0.0018835 0.42642 2.0595 2.0588 16.0097 144.941 0.00017116 -85.6441 0.74095
6.845 0.98811 5.4781e-005 3.8183 0.011948 8.9227e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.439 0.50624 0.15471 0.01848 12.866 0.11487 0.00014797 0.77528 0.0087779 0.0097364 0.0013881 0.98692 0.99169 2.9932e-006 1.1973e-005 0.16003 0.92567 0.91186 0.001398 0.99026 0.49914 0.0018834 0.42644 2.06 2.0593 16.0096 144.941 0.00017105 -85.6442 0.74195
6.846 0.98811 5.4781e-005 3.8183 0.011948 8.924e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4391 0.50629 0.15473 0.018481 12.8685 0.11488 0.00014799 0.77527 0.0087784 0.0097369 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.16003 0.92585 0.91193 0.001398 0.99031 0.49932 0.0018834 0.42645 2.0605 2.0598 16.0096 144.941 0.00017094 -85.6444 0.74295
6.847 0.98811 5.478e-005 3.8183 0.011948 8.9252e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4392 0.50633 0.15474 0.018482 12.8711 0.11488 0.000148 0.77526 0.0087789 0.0097374 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.16004 0.92603 0.912 0.0013979 0.99035 0.49949 0.0018834 0.42646 2.061 2.0603 16.0096 144.9411 0.00017083 -85.6445 0.74395
6.848 0.98811 5.478e-005 3.8183 0.011948 8.9265e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4393 0.50638 0.15476 0.018484 12.8736 0.11489 0.00014801 0.77526 0.0087794 0.0097379 0.001388 0.98692 0.99169 2.993e-006 1.1972e-005 0.16004 0.92621 0.91207 0.0013979 0.9904 0.49967 0.0018834 0.42648 2.0615 2.0608 16.0096 144.9411 0.00017072 -85.6447 0.74495
6.849 0.98811 5.478e-005 3.8183 0.011948 8.9278e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4394 0.50642 0.15477 0.018485 12.8762 0.1149 0.00014802 0.77525 0.0087798 0.0097385 0.0013879 0.98692 0.99169 2.9929e-006 1.1972e-005 0.16004 0.92639 0.91214 0.0013979 0.99044 0.49984 0.0018834 0.42649 2.062 2.0613 16.0095 144.9411 0.00017061 -85.6448 0.74595
6.85 0.98811 5.478e-005 3.8183 0.011948 8.9291e-005 0.0011669 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4395 0.50647 0.15479 0.018486 12.8787 0.11491 0.00014803 0.77524 0.0087803 0.009739 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.16005 0.92657 0.91222 0.0013979 0.99048 0.50002 0.0018833 0.4265 2.0625 2.0618 16.0095 144.9411 0.0001705 -85.645 0.74695
6.851 0.98811 5.478e-005 3.8183 0.011948 8.9304e-005 0.001167 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4396 0.50651 0.1548 0.018487 12.8813 0.11492 0.00014804 0.77523 0.0087808 0.0097395 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.16005 0.92675 0.91229 0.0013979 0.99053 0.50019 0.0018833 0.42652 2.063 2.0623 16.0095 144.9411 0.00017039 -85.6451 0.74795
6.852 0.98811 5.478e-005 3.8183 0.011948 8.9317e-005 0.001167 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4397 0.50656 0.15481 0.018489 12.8838 0.11492 0.00014805 0.77523 0.0087812 0.00974 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.16005 0.92693 0.91236 0.0013979 0.99057 0.50036 0.0018833 0.42653 2.0635 2.0628 16.0094 144.9412 0.00017028 -85.6452 0.74895
6.853 0.98811 5.478e-005 3.8183 0.011948 8.933e-005 0.001167 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4397 0.50661 0.15483 0.01849 12.8864 0.11493 0.00014806 0.77522 0.0087817 0.0097405 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.16006 0.9271 0.91243 0.0013978 0.99061 0.50054 0.0018833 0.42654 2.064 2.0633 16.0094 144.9412 0.00017017 -85.6454 0.74995
6.854 0.98811 5.478e-005 3.8183 0.011948 8.9343e-005 0.001167 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4398 0.50665 0.15484 0.018491 12.8889 0.11494 0.00014808 0.77521 0.0087822 0.009741 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.16006 0.92728 0.9125 0.0013978 0.99066 0.50071 0.0018832 0.42656 2.0645 2.0638 16.0094 144.9412 0.00017006 -85.6455 0.75095
6.855 0.98811 5.478e-005 3.8183 0.011948 8.9355e-005 0.001167 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.4399 0.5067 0.15486 0.018492 12.8915 0.11495 0.00014809 0.7752 0.0087827 0.0097415 0.0013877 0.98693 0.99169 2.9925e-006 1.197e-005 0.16006 0.92746 0.91257 0.0013978 0.9907 0.50089 0.0018832 0.42657 2.0649 2.0643 16.0094 144.9412 0.00016995 -85.6457 0.75195
6.856 0.98811 5.478e-005 3.8183 0.011948 8.9368e-005 0.001167 0.23358 0.00065931 0.23423 0.21615 0 0.032265 0.0389 0 1.44 0.50674 0.15487 0.018494 12.894 0.11495 0.0001481 0.77519 0.0087831 0.009742 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.16007 0.92763 0.91264 0.0013978 0.99074 0.50106 0.0018832 0.42659 2.0654 2.0647 16.0093 144.9412 0.00016984 -85.6458 0.75295
6.857 0.98811 5.478e-005 3.8183 0.011948 8.9381e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4401 0.50679 0.15489 0.018495 12.8966 0.11496 0.00014811 0.77519 0.0087836 0.0097425 0.0013877 0.98693 0.99169 2.9923e-006 1.1969e-005 0.16007 0.92781 0.91271 0.0013978 0.99078 0.50123 0.0018832 0.4266 2.0659 2.0652 16.0093 144.9413 0.00016974 -85.6459 0.75395
6.858 0.98811 5.478e-005 3.8183 0.011948 8.9394e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4402 0.50683 0.1549 0.018496 12.8992 0.11497 0.00014812 0.77518 0.0087841 0.009743 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.16008 0.92798 0.91278 0.0013978 0.99082 0.50141 0.0018832 0.42661 2.0664 2.0657 16.0093 144.9413 0.00016963 -85.6461 0.75495
6.859 0.98811 5.478e-005 3.8183 0.011948 8.9407e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4403 0.50688 0.15492 0.018497 12.9017 0.11498 0.00014813 0.77517 0.0087845 0.0097435 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.16008 0.92815 0.91285 0.0013978 0.99086 0.50158 0.0018831 0.42663 2.0669 2.0662 16.0093 144.9413 0.00016952 -85.6462 0.75595
6.86 0.98811 5.4779e-005 3.8183 0.011948 8.942e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4404 0.50693 0.15493 0.018499 12.9043 0.11498 0.00014814 0.77516 0.008785 0.009744 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.16008 0.92833 0.91291 0.0013978 0.99091 0.50176 0.0018831 0.42664 2.0674 2.0667 16.0092 144.9413 0.00016942 -85.6464 0.75695
6.861 0.98811 5.4779e-005 3.8183 0.011948 8.9433e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4405 0.50697 0.15494 0.0185 12.9068 0.11499 0.00014815 0.77516 0.0087855 0.0097445 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16009 0.9285 0.91298 0.0013978 0.99095 0.50193 0.0018831 0.42665 2.0678 2.0672 16.0092 144.9414 0.00016931 -85.6465 0.75795
6.862 0.98811 5.4779e-005 3.8183 0.011948 8.9446e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4406 0.50702 0.15496 0.018501 12.9094 0.115 0.00014817 0.77515 0.0087859 0.009745 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16009 0.92867 0.91305 0.0013978 0.99099 0.5021 0.0018831 0.42667 2.0683 2.0676 16.0092 144.9414 0.0001692 -85.6466 0.75895
6.863 0.98811 5.4779e-005 3.8183 0.011948 8.9458e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4407 0.50706 0.15497 0.018502 12.9119 0.11501 0.00014818 0.77514 0.0087864 0.0097455 0.0013875 0.98693 0.99169 2.9919e-006 1.1967e-005 0.16009 0.92884 0.91312 0.0013978 0.99103 0.50228 0.001883 0.42668 2.0688 2.0681 16.0091 144.9414 0.0001691 -85.6468 0.75995
6.864 0.98811 5.4779e-005 3.8183 0.011948 8.9471e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4407 0.50711 0.15499 0.018504 12.9145 0.11501 0.00014819 0.77513 0.0087869 0.009746 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.1601 0.92901 0.91319 0.0013977 0.99107 0.50245 0.001883 0.42669 2.0693 2.0686 16.0091 144.9414 0.00016899 -85.6469 0.76095
6.865 0.98811 5.4779e-005 3.8183 0.011948 8.9484e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4408 0.50715 0.155 0.018505 12.917 0.11502 0.0001482 0.77513 0.0087874 0.0097465 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.1601 0.92918 0.91325 0.0013977 0.99111 0.50262 0.001883 0.42671 2.0697 2.0691 16.0091 144.9414 0.00016889 -85.647 0.76195
6.866 0.98811 5.4779e-005 3.8183 0.011947 8.9497e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4409 0.5072 0.15502 0.018506 12.9196 0.11503 0.00014821 0.77512 0.0087878 0.009747 0.0013874 0.98693 0.9917 2.9917e-006 1.1967e-005 0.1601 0.92935 0.91332 0.0013977 0.99115 0.5028 0.001883 0.42672 2.0702 2.0696 16.0091 144.9415 0.00016878 -85.6471 0.76295
6.867 0.98811 5.4779e-005 3.8183 0.011947 8.951e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.441 0.50725 0.15503 0.018507 12.9222 0.11504 0.00014822 0.77511 0.0087883 0.0097475 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.16011 0.92952 0.91339 0.0013977 0.99119 0.50297 0.001883 0.42673 2.0707 2.07 16.009 144.9415 0.00016868 -85.6473 0.76395
6.868 0.98811 5.4779e-005 3.8183 0.011947 8.9523e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4411 0.50729 0.15504 0.018509 12.9247 0.11504 0.00014823 0.7751 0.0087888 0.009748 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.16011 0.92969 0.91345 0.0013976 0.99122 0.50314 0.0018829 0.42675 2.0712 2.0705 16.009 144.9415 0.00016858 -85.6474 0.76495
6.869 0.98811 5.4779e-005 3.8183 0.011947 8.9536e-005 0.001167 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4412 0.50734 0.15506 0.01851 12.9273 0.11505 0.00014824 0.7751 0.0087892 0.0097485 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.16012 0.92986 0.91352 0.0013976 0.99126 0.50332 0.0018829 0.42676 2.0716 2.071 16.009 144.9415 0.00016847 -85.6475 0.76595
6.87 0.98811 5.4779e-005 3.8183 0.011947 8.9549e-005 0.001167 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4413 0.50738 0.15507 0.018511 12.9298 0.11506 0.00014826 0.77509 0.0087897 0.009749 0.0013873 0.98693 0.9917 2.9914e-006 1.1966e-005 0.16012 0.93003 0.91359 0.0013976 0.9913 0.50349 0.0018829 0.42677 2.0721 2.0715 16.0089 144.9415 0.00016837 -85.6477 0.76695
6.871 0.98811 5.4779e-005 3.8183 0.011947 8.9561e-005 0.001167 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4414 0.50743 0.15509 0.018512 12.9324 0.11507 0.00014827 0.77508 0.0087902 0.0097495 0.0013872 0.98693 0.9917 2.9914e-006 1.1965e-005 0.16012 0.9302 0.91365 0.0013976 0.99134 0.50366 0.0018829 0.42679 2.0726 2.0719 16.0089 144.9416 0.00016827 -85.6478 0.76795
6.872 0.98811 5.4779e-005 3.8183 0.011947 8.9574e-005 0.001167 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4415 0.50747 0.1551 0.018514 12.9349 0.11507 0.00014828 0.77507 0.0087906 0.00975 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16013 0.93036 0.91372 0.0013975 0.99138 0.50383 0.0018829 0.4268 2.0731 2.0724 16.0089 144.9416 0.00016817 -85.6479 0.76895
6.873 0.98811 5.4778e-005 3.8183 0.011947 8.9587e-005 0.001167 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4416 0.50752 0.15512 0.018515 12.9375 0.11508 0.00014829 0.77507 0.0087911 0.0097505 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.16013 0.93053 0.91378 0.0013975 0.99142 0.50401 0.0018828 0.42682 2.0735 2.0729 16.0089 144.9416 0.00016806 -85.648 0.76995
6.874 0.98811 5.4778e-005 3.8183 0.011947 8.96e-005 0.001167 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4416 0.50757 0.15513 0.018516 12.9401 0.11509 0.0001483 0.77506 0.0087916 0.009751 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.16013 0.93069 0.91385 0.0013975 0.99145 0.50418 0.0018828 0.42683 2.074 2.0733 16.0088 144.9416 0.00016796 -85.6481 0.77095
6.875 0.98811 5.4778e-005 3.8183 0.011947 8.9613e-005 0.001167 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4417 0.50761 0.15515 0.018517 12.9426 0.1151 0.00014831 0.77505 0.0087921 0.0097516 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.16014 0.93086 0.91391 0.0013975 0.99149 0.50435 0.0018828 0.42684 2.0745 2.0738 16.0088 144.9416 0.00016786 -85.6483 0.77195
6.876 0.98811 5.4778e-005 3.8183 0.011947 8.9626e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4418 0.50766 0.15516 0.018519 12.9452 0.1151 0.00014832 0.77504 0.0087925 0.0097521 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16014 0.93102 0.91398 0.0013975 0.99153 0.50453 0.0018828 0.42686 2.0749 2.0743 16.0088 144.9417 0.00016776 -85.6484 0.77295
6.877 0.98811 5.4778e-005 3.8183 0.011947 8.9639e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4419 0.5077 0.15517 0.01852 12.9477 0.11511 0.00014833 0.77504 0.008793 0.0097526 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16015 0.93119 0.91404 0.0013975 0.99156 0.5047 0.0018828 0.42687 2.0754 2.0747 16.0087 144.9417 0.00016766 -85.6485 0.77395
6.878 0.98811 5.4778e-005 3.8183 0.011947 8.9652e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.442 0.50775 0.15519 0.018521 12.9503 0.11512 0.00014835 0.77503 0.0087935 0.0097531 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.16015 0.93135 0.91411 0.0013974 0.9916 0.50487 0.0018827 0.42688 2.0759 2.0752 16.0087 144.9417 0.00016756 -85.6486 0.77495
6.879 0.98811 5.4778e-005 3.8183 0.011947 8.9664e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4421 0.50779 0.1552 0.018522 12.9529 0.11513 0.00014836 0.77502 0.0087939 0.0097536 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.16015 0.93151 0.91417 0.0013974 0.99164 0.50504 0.0018827 0.4269 2.0763 2.0757 16.0087 144.9417 0.00016746 -85.6487 0.77595
6.88 0.98811 5.4778e-005 3.8183 0.011947 8.9677e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4422 0.50784 0.15522 0.018524 12.9554 0.11514 0.00014837 0.77501 0.0087944 0.0097541 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.16016 0.93168 0.91424 0.0013974 0.99167 0.50522 0.0018827 0.42691 2.0768 2.0761 16.0087 144.9417 0.00016736 -85.6489 0.77695
6.881 0.98811 5.4778e-005 3.8183 0.011947 8.969e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4423 0.50789 0.15523 0.018525 12.958 0.11514 0.00014838 0.77501 0.0087949 0.0097546 0.001387 0.98693 0.9917 2.9907e-006 1.1963e-005 0.16016 0.93184 0.9143 0.0013974 0.99171 0.50539 0.0018827 0.42692 2.0772 2.0766 16.0086 144.9418 0.00016726 -85.649 0.77795
6.882 0.98811 5.4778e-005 3.8183 0.011947 8.9703e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4424 0.50793 0.15525 0.018526 12.9605 0.11515 0.00014839 0.775 0.0087953 0.0097551 0.0013869 0.98694 0.9917 2.9907e-006 1.1963e-005 0.16016 0.932 0.91436 0.0013974 0.99174 0.50556 0.0018827 0.42694 2.0777 2.0771 16.0086 144.9418 0.00016716 -85.6491 0.77895
6.883 0.98811 5.4778e-005 3.8183 0.011947 8.9716e-005 0.0011671 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.4425 0.50798 0.15526 0.018527 12.9631 0.11516 0.0001484 0.77499 0.0087958 0.0097556 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16017 0.93216 0.91443 0.0013974 0.99178 0.50573 0.0018827 0.42695 2.0782 2.0775 16.0086 144.9418 0.00016707 -85.6492 0.77995
6.884 0.98811 5.4778e-005 3.8183 0.011947 8.9729e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.4425 0.50802 0.15527 0.018529 12.9657 0.11517 0.00014841 0.77498 0.0087963 0.0097561 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16017 0.93232 0.91449 0.0013974 0.99181 0.5059 0.0018826 0.42696 2.0786 2.078 16.0085 144.9418 0.00016697 -85.6493 0.78095
6.885 0.98811 5.4777e-005 3.8183 0.011947 8.9742e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.4426 0.50807 0.15529 0.01853 12.9682 0.11517 0.00014842 0.77498 0.0087967 0.0097566 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16017 0.93248 0.91455 0.0013974 0.99185 0.50608 0.0018826 0.42698 2.0791 2.0784 16.0085 144.9418 0.00016687 -85.6494 0.78195
6.886 0.98811 5.4777e-005 3.8183 0.011947 8.9755e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.4427 0.50811 0.1553 0.018531 12.9708 0.11518 0.00014843 0.77497 0.0087972 0.0097571 0.0013868 0.98694 0.9917 2.9904e-006 1.1962e-005 0.16018 0.93264 0.91462 0.0013974 0.99188 0.50625 0.0018826 0.42699 2.0795 2.0789 16.0085 144.9419 0.00016677 -85.6495 0.78295
6.887 0.98811 5.4777e-005 3.8183 0.011947 8.9768e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.4428 0.50816 0.15532 0.018532 12.9734 0.11519 0.00014845 0.77496 0.0087977 0.0097576 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.16018 0.9328 0.91468 0.0013974 0.99192 0.50642 0.0018826 0.427 2.08 2.0793 16.0085 144.9419 0.00016668 -85.6497 0.78395
6.888 0.98811 5.4777e-005 3.8183 0.011947 8.978e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.4429 0.5082 0.15533 0.018534 12.9759 0.1152 0.00014846 0.77495 0.0087981 0.0097581 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16019 0.93296 0.91474 0.0013974 0.99195 0.50659 0.0018826 0.42702 2.0804 2.0798 16.0084 144.9419 0.00016658 -85.6498 0.78495
6.889 0.98811 5.4777e-005 3.8183 0.011947 8.9793e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.443 0.50825 0.15535 0.018535 12.9785 0.1152 0.00014847 0.77495 0.0087986 0.0097586 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16019 0.93312 0.9148 0.0013974 0.99199 0.50676 0.0018825 0.42703 2.0809 2.0803 16.0084 144.9419 0.00016648 -85.6499 0.78595
6.89 0.98811 5.4777e-005 3.8183 0.011947 8.9806e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4431 0.5083 0.15536 0.018536 12.9811 0.11521 0.00014848 0.77494 0.0087991 0.0097591 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16019 0.93328 0.91486 0.0013974 0.99202 0.50694 0.0018825 0.42704 2.0813 2.0807 16.0084 144.9419 0.00016639 -85.65 0.78695
6.891 0.98811 5.4777e-005 3.8183 0.011947 8.9819e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4432 0.50834 0.15538 0.018537 12.9836 0.11522 0.00014849 0.77493 0.0087996 0.0097596 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.1602 0.93343 0.91493 0.0013973 0.99205 0.50711 0.0018825 0.42706 2.0818 2.0812 16.0083 144.942 0.00016629 -85.6501 0.78795
6.892 0.98811 5.4777e-005 3.8183 0.011947 8.9832e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4433 0.50839 0.15539 0.018539 12.9862 0.11523 0.0001485 0.77492 0.0088 0.0097601 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.1602 0.93359 0.91499 0.0013973 0.99209 0.50728 0.0018825 0.42707 2.0822 2.0816 16.0083 144.942 0.0001662 -85.6502 0.78895
6.893 0.98811 5.4777e-005 3.8183 0.011947 8.9845e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4434 0.50843 0.1554 0.01854 12.9888 0.11523 0.00014851 0.77492 0.0088005 0.0097606 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.1602 0.93375 0.91505 0.0013973 0.99212 0.50745 0.0018825 0.42708 2.0827 2.0821 16.0083 144.942 0.0001661 -85.6503 0.78995
6.894 0.98811 5.4777e-005 3.8183 0.011947 8.9858e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4434 0.50848 0.15542 0.018541 12.9913 0.11524 0.00014852 0.77491 0.008801 0.0097611 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.16021 0.9339 0.91511 0.0013973 0.99215 0.50762 0.0018825 0.4271 2.0831 2.0825 16.0083 144.942 0.00016601 -85.6504 0.79095
6.895 0.98811 5.4777e-005 3.8183 0.011947 8.9871e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4435 0.50852 0.15543 0.018542 12.9939 0.11525 0.00014854 0.7749 0.0088014 0.0097616 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.16021 0.93406 0.91517 0.0013973 0.99219 0.50779 0.0018824 0.42711 2.0836 2.083 16.0082 144.942 0.00016591 -85.6505 0.79195
6.896 0.98811 5.4777e-005 3.8183 0.011947 8.9883e-005 0.0011671 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4436 0.50857 0.15545 0.018544 12.9965 0.11526 0.00014855 0.77489 0.0088019 0.0097621 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.16021 0.93421 0.91523 0.0013972 0.99222 0.50797 0.0018824 0.42712 2.084 2.0834 16.0082 144.9421 0.00016582 -85.6506 0.79295
6.897 0.98811 5.4777e-005 3.8183 0.011947 8.9896e-005 0.0011671 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4437 0.50862 0.15546 0.018545 12.999 0.11526 0.00014856 0.77488 0.0088024 0.0097626 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.16022 0.93436 0.91529 0.0013972 0.99225 0.50814 0.0018824 0.42714 2.0845 2.0839 16.0082 144.9421 0.00016573 -85.6507 0.79395
6.898 0.98811 5.4776e-005 3.8183 0.011947 8.9909e-005 0.0011671 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4438 0.50866 0.15548 0.018546 13.0016 0.11527 0.00014857 0.77488 0.0088028 0.0097631 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.16022 0.93452 0.91535 0.0013972 0.99228 0.50831 0.0018824 0.42715 2.0849 2.0843 16.0081 144.9421 0.00016563 -85.6508 0.79495
6.899 0.98811 5.4776e-005 3.8183 0.011947 8.9922e-005 0.0011671 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4439 0.50871 0.15549 0.018547 13.0042 0.11528 0.00014858 0.77487 0.0088033 0.0097636 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.16023 0.93467 0.91541 0.0013972 0.99231 0.50848 0.0018824 0.42716 2.0854 2.0848 16.0081 144.9421 0.00016554 -85.6509 0.79595
6.9 0.98811 5.4776e-005 3.8183 0.011947 8.9935e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.444 0.50875 0.1555 0.018549 13.0067 0.11529 0.00014859 0.77486 0.0088038 0.0097641 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16023 0.93482 0.91547 0.0013972 0.99235 0.50865 0.0018824 0.42718 2.0858 2.0852 16.0081 144.9422 0.00016545 -85.651 0.79695
6.901 0.98811 5.4776e-005 3.8183 0.011947 8.9948e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4441 0.5088 0.15552 0.01855 13.0093 0.11529 0.0001486 0.77485 0.0088042 0.0097646 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16023 0.93498 0.91553 0.0013972 0.99238 0.50882 0.0018823 0.42719 2.0863 2.0856 16.0081 144.9422 0.00016535 -85.6511 0.79795
6.902 0.98811 5.4776e-005 3.8183 0.011947 8.9961e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4442 0.50884 0.15553 0.018551 13.0119 0.1153 0.00014861 0.77485 0.0088047 0.0097651 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16024 0.93513 0.91559 0.0013971 0.99241 0.50899 0.0018823 0.4272 2.0867 2.0861 16.008 144.9422 0.00016526 -85.6512 0.79895
6.903 0.98811 5.4776e-005 3.8183 0.011947 8.9974e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4443 0.50889 0.15555 0.018552 13.0144 0.11531 0.00014862 0.77484 0.0088052 0.0097656 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16024 0.93528 0.91565 0.0013971 0.99244 0.50916 0.0018823 0.42722 2.0871 2.0865 16.008 144.9422 0.00016517 -85.6513 0.79995
6.904 0.98811 5.4776e-005 3.8183 0.011947 8.9986e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4443 0.50894 0.15556 0.018554 13.017 0.11532 0.00014864 0.77483 0.0088056 0.0097661 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.16024 0.93543 0.91571 0.0013971 0.99247 0.50934 0.0018823 0.42723 2.0876 2.087 16.008 144.9422 0.00016508 -85.6514 0.80095
6.905 0.98811 5.4776e-005 3.8183 0.011947 8.9999e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4444 0.50898 0.15558 0.018555 13.0196 0.11532 0.00014865 0.77482 0.0088061 0.0097666 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.16025 0.93558 0.91577 0.0013971 0.9925 0.50951 0.0018823 0.42724 2.088 2.0874 16.0079 144.9423 0.00016499 -85.6515 0.80195
6.906 0.98811 5.4776e-005 3.8183 0.011947 9.0012e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4445 0.50903 0.15559 0.018556 13.0221 0.11533 0.00014866 0.77482 0.0088066 0.0097671 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16025 0.93573 0.91582 0.0013971 0.99253 0.50968 0.0018823 0.42726 2.0885 2.0878 16.0079 144.9423 0.0001649 -85.6516 0.80295
6.907 0.98811 5.4776e-005 3.8183 0.011947 9.0025e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4446 0.50907 0.1556 0.018557 13.0247 0.11534 0.00014867 0.77481 0.008807 0.0097676 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16025 0.93588 0.91588 0.0013971 0.99256 0.50985 0.0018822 0.42727 2.0889 2.0883 16.0079 144.9423 0.00016481 -85.6517 0.80395
6.908 0.98811 5.4776e-005 3.8183 0.011947 9.0038e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4447 0.50912 0.15562 0.018559 13.0273 0.11535 0.00014868 0.7748 0.0088075 0.0097681 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16026 0.93603 0.91594 0.0013971 0.99259 0.51002 0.0018822 0.42728 2.0893 2.0887 16.0079 144.9423 0.00016472 -85.6518 0.80495
6.909 0.98811 5.4776e-005 3.8183 0.011947 9.0051e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4448 0.50916 0.15563 0.01856 13.0299 0.11535 0.00014869 0.77479 0.008808 0.0097686 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16026 0.93618 0.916 0.0013971 0.99262 0.51019 0.0018822 0.4273 2.0898 2.0892 16.0078 144.9423 0.00016463 -85.6519 0.80595
6.91 0.98811 5.4776e-005 3.8183 0.011947 9.0064e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.4449 0.50921 0.15565 0.018561 13.0324 0.11536 0.0001487 0.77479 0.0088084 0.0097691 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.16027 0.93633 0.91606 0.0013971 0.99265 0.51036 0.0018822 0.42731 2.0902 2.0896 16.0078 144.9424 0.00016454 -85.652 0.80695
6.911 0.98811 5.4775e-005 3.8183 0.011947 9.0077e-005 0.0011672 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.445 0.50926 0.15566 0.018562 13.035 0.11537 0.00014871 0.77478 0.0088089 0.0097696 0.0013862 0.98694 0.9917 2.9891e-006 1.1956e-005 0.16027 0.93647 0.91611 0.0013971 0.99268 0.51053 0.0018822 0.42732 2.0906 2.09 16.0078 144.9424 0.00016445 -85.6521 0.80795
6.912 0.98811 5.4775e-005 3.8183 0.011947 9.0089e-005 0.0011672 0.2336 0.00065931 0.23426 0.21616 0 0.032264 0.0389 0 1.4451 0.5093 0.15568 0.018564 13.0376 0.11538 0.00014873 0.77477 0.0088094 0.0097701 0.0013862 0.98694 0.9917 2.989e-006 1.1956e-005 0.16027 0.93662 0.91617 0.0013971 0.99271 0.5107 0.0018822 0.42734 2.0911 2.0905 16.0077 144.9424 0.00016436 -85.6522 0.80895
6.913 0.98811 5.4775e-005 3.8183 0.011947 9.0102e-005 0.0011672 0.2336 0.00065931 0.23426 0.21616 0 0.032264 0.0389 0 1.4452 0.50935 0.15569 0.018565 13.0401 0.11538 0.00014874 0.77476 0.0088098 0.0097706 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16028 0.93677 0.91623 0.0013971 0.99274 0.51087 0.0018822 0.42735 2.0915 2.0909 16.0077 144.9424 0.00016427 -85.6523 0.80995
6.914 0.98811 5.4775e-005 3.8183 0.011947 9.0115e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4452 0.50939 0.15571 0.018566 13.0427 0.11539 0.00014875 0.77476 0.0088103 0.0097711 0.0013862 0.98695 0.99171 2.9889e-006 1.1956e-005 0.16028 0.93691 0.91628 0.0013971 0.99277 0.51104 0.0018821 0.42736 2.0919 2.0913 16.0077 144.9424 0.00016418 -85.6524 0.81095
6.915 0.98811 5.4775e-005 3.8183 0.011947 9.0128e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4453 0.50944 0.15572 0.018567 13.0453 0.1154 0.00014876 0.77475 0.0088108 0.0097716 0.0013861 0.98695 0.99171 2.9889e-006 1.1955e-005 0.16028 0.93706 0.91634 0.0013971 0.9928 0.51121 0.0018821 0.42738 2.0924 2.0918 16.0076 144.9425 0.0001641 -85.6525 0.81195
6.916 0.98811 5.4775e-005 3.8183 0.011947 9.0141e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4454 0.50948 0.15573 0.018569 13.0479 0.11541 0.00014877 0.77474 0.0088112 0.0097721 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16029 0.9372 0.9164 0.001397 0.99282 0.51138 0.0018821 0.42739 2.0928 2.0922 16.0076 144.9425 0.00016401 -85.6526 0.81295
6.917 0.98811 5.4775e-005 3.8183 0.011947 9.0154e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4455 0.50953 0.15575 0.01857 13.0504 0.11541 0.00014878 0.77473 0.0088117 0.0097726 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16029 0.93735 0.91645 0.001397 0.99285 0.51155 0.0018821 0.4274 2.0932 2.0926 16.0076 144.9425 0.00016392 -85.6526 0.81395
6.918 0.98811 5.4775e-005 3.8183 0.011947 9.0167e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4456 0.50958 0.15576 0.018571 13.053 0.11542 0.00014879 0.77473 0.0088122 0.0097731 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16029 0.93749 0.91651 0.001397 0.99288 0.51172 0.0018821 0.42742 2.0937 2.0931 16.0076 144.9425 0.00016383 -85.6527 0.81495
6.919 0.98811 5.4775e-005 3.8183 0.011947 9.018e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4457 0.50962 0.15578 0.018572 13.0556 0.11543 0.0001488 0.77472 0.0088126 0.0097736 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.1603 0.93764 0.91657 0.001397 0.99291 0.51189 0.0018821 0.42743 2.0941 2.0935 16.0075 144.9425 0.00016375 -85.6528 0.81595
6.92 0.98811 5.4775e-005 3.8183 0.011947 9.0192e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4458 0.50967 0.15579 0.018574 13.0582 0.11544 0.00014881 0.77471 0.0088131 0.0097741 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.1603 0.93778 0.91662 0.001397 0.99294 0.51206 0.0018821 0.42744 2.0945 2.0939 16.0075 144.9426 0.00016366 -85.6529 0.81695
6.921 0.98811 5.4775e-005 3.8183 0.011947 9.0205e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4459 0.50971 0.15581 0.018575 13.0607 0.11544 0.00014883 0.7747 0.0088136 0.0097746 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.1603 0.93792 0.91668 0.001397 0.99296 0.51223 0.001882 0.42746 2.0949 2.0943 16.0075 144.9426 0.00016357 -85.653 0.81795
6.922 0.98811 5.4775e-005 3.8183 0.011947 9.0218e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.446 0.50976 0.15582 0.018576 13.0633 0.11545 0.00014884 0.7747 0.008814 0.0097751 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16031 0.93807 0.91673 0.0013969 0.99299 0.5124 0.001882 0.42747 2.0954 2.0948 16.0074 144.9426 0.00016349 -85.6531 0.81895
6.923 0.98811 5.4774e-005 3.8183 0.011947 9.0231e-005 0.0011672 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4461 0.5098 0.15583 0.018577 13.0659 0.11546 0.00014885 0.77469 0.0088145 0.0097756 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16031 0.93821 0.91679 0.0013969 0.99302 0.51257 0.001882 0.42748 2.0958 2.0952 16.0074 144.9426 0.0001634 -85.6532 0.81995
6.924 0.98811 5.4774e-005 3.8183 0.011947 9.0244e-005 0.0011673 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4461 0.50985 0.15585 0.018579 13.0685 0.11547 0.00014886 0.77468 0.008815 0.0097761 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16032 0.93835 0.91684 0.0013969 0.99305 0.51274 0.001882 0.4275 2.0962 2.0956 16.0074 144.9426 0.00016332 -85.6532 0.82095
6.925 0.98811 5.4774e-005 3.8183 0.011946 9.0257e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4462 0.5099 0.15586 0.01858 13.071 0.11547 0.00014887 0.77467 0.0088154 0.0097766 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.16032 0.93849 0.9169 0.0013969 0.99307 0.51291 0.001882 0.42751 2.0966 2.096 16.0073 144.9427 0.00016323 -85.6533 0.82195
6.926 0.98811 5.4774e-005 3.8183 0.011946 9.027e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4463 0.50994 0.15588 0.018581 13.0736 0.11548 0.00014888 0.77467 0.0088159 0.0097771 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.16032 0.93863 0.91695 0.0013969 0.9931 0.51308 0.001882 0.42752 2.097 2.0965 16.0073 144.9427 0.00016315 -85.6534 0.82295
6.927 0.98811 5.4774e-005 3.8183 0.011946 9.0283e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4464 0.50999 0.15589 0.018582 13.0762 0.11549 0.00014889 0.77466 0.0088164 0.0097776 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16033 0.93877 0.91701 0.0013969 0.99313 0.51325 0.001882 0.42754 2.0975 2.0969 16.0073 144.9427 0.00016306 -85.6535 0.82395
6.928 0.98811 5.4774e-005 3.8183 0.011946 9.0295e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4465 0.51003 0.15591 0.018584 13.0788 0.1155 0.0001489 0.77465 0.0088168 0.0097781 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16033 0.93891 0.91706 0.0013969 0.99315 0.51342 0.001882 0.42755 2.0979 2.0973 16.0073 144.9427 0.00016298 -85.6536 0.82495
6.929 0.98811 5.4774e-005 3.8183 0.011946 9.0308e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4466 0.51008 0.15592 0.018585 13.0814 0.1155 0.00014891 0.77464 0.0088173 0.0097786 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16033 0.93905 0.91711 0.0013968 0.99318 0.51359 0.0018819 0.42756 2.0983 2.0977 16.0072 144.9427 0.0001629 -85.6537 0.82595
6.93 0.98811 5.4774e-005 3.8183 0.011946 9.0321e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4467 0.51012 0.15593 0.018586 13.0839 0.11551 0.00014893 0.77464 0.0088177 0.0097791 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16034 0.93919 0.91717 0.0013968 0.9932 0.51376 0.0018819 0.42758 2.0987 2.0981 16.0072 144.9428 0.00016281 -85.6537 0.82695
6.931 0.98811 5.4774e-005 3.8183 0.011946 9.0334e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4468 0.51017 0.15595 0.018587 13.0865 0.11552 0.00014894 0.77463 0.0088182 0.0097796 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16034 0.93933 0.91722 0.0013968 0.99323 0.51393 0.0018819 0.42759 2.0991 2.0986 16.0072 144.9428 0.00016273 -85.6538 0.82795
6.932 0.98811 5.4774e-005 3.8183 0.011946 9.0347e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4469 0.51022 0.15596 0.018589 13.0891 0.11553 0.00014895 0.77462 0.0088187 0.0097801 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16034 0.93947 0.91727 0.0013968 0.99326 0.5141 0.0018819 0.4276 2.0996 2.099 16.0071 144.9428 0.00016265 -85.6539 0.82895
6.933 0.98811 5.4774e-005 3.8183 0.011946 9.036e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.447 0.51026 0.15598 0.01859 13.0917 0.11554 0.00014896 0.77461 0.0088191 0.0097806 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16035 0.93961 0.91733 0.0013968 0.99328 0.51427 0.0018819 0.42762 2.1 2.0994 16.0071 144.9428 0.00016256 -85.654 0.82995
6.934 0.98811 5.4774e-005 3.8183 0.011946 9.0373e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.447 0.51031 0.15599 0.018591 13.0942 0.11554 0.00014897 0.77461 0.0088196 0.0097811 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16035 0.93974 0.91738 0.0013968 0.99331 0.51444 0.0018819 0.42763 2.1004 2.0998 16.0071 144.9428 0.00016248 -85.6541 0.83095
6.935 0.98811 5.4774e-005 3.8183 0.011946 9.0386e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4471 0.51035 0.15601 0.018592 13.0968 0.11555 0.00014898 0.7746 0.0088201 0.0097816 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16036 0.93988 0.91743 0.0013968 0.99333 0.51461 0.0018819 0.42764 2.1008 2.1002 16.007 144.9429 0.0001624 -85.6541 0.83195
6.936 0.98811 5.4773e-005 3.8183 0.011946 9.0398e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4472 0.5104 0.15602 0.018594 13.0994 0.11556 0.00014899 0.77459 0.0088205 0.0097821 0.0013857 0.98695 0.99171 2.988e-006 1.1952e-005 0.16036 0.94002 0.91749 0.0013968 0.99336 0.51478 0.0018818 0.42766 2.1012 2.1006 16.007 144.9429 0.00016232 -85.6542 0.83295
6.937 0.98811 5.4773e-005 3.8183 0.011946 9.0411e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4473 0.51044 0.15604 0.018595 13.102 0.11557 0.000149 0.77458 0.008821 0.0097826 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.16036 0.94015 0.91754 0.0013968 0.99338 0.51495 0.0018818 0.42767 2.1016 2.1011 16.007 144.9429 0.00016223 -85.6543 0.83395
6.938 0.98811 5.4773e-005 3.8183 0.011946 9.0424e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4474 0.51049 0.15605 0.018596 13.1046 0.11557 0.00014902 0.77458 0.0088215 0.0097831 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.16037 0.94029 0.91759 0.0013968 0.99341 0.51511 0.0018818 0.42768 2.102 2.1015 16.007 144.9429 0.00016215 -85.6544 0.83495
6.939 0.98811 5.4773e-005 3.8183 0.011946 9.0437e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4475 0.51053 0.15606 0.018597 13.1072 0.11558 0.00014903 0.77457 0.0088219 0.0097836 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16037 0.94042 0.91764 0.0013968 0.99343 0.51528 0.0018818 0.4277 2.1025 2.1019 16.0069 144.943 0.00016207 -85.6544 0.83595
6.94 0.98811 5.4773e-005 3.8183 0.011946 9.045e-005 0.0011673 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.4476 0.51058 0.15608 0.018599 13.1097 0.11559 0.00014904 0.77456 0.0088224 0.0097841 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16037 0.94056 0.9177 0.0013968 0.99346 0.51545 0.0018818 0.42771 2.1029 2.1023 16.0069 144.943 0.00016199 -85.6545 0.83695
6.941 0.98811 5.4773e-005 3.8183 0.011946 9.0463e-005 0.0011673 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.4477 0.51063 0.15609 0.0186 13.1123 0.1156 0.00014905 0.77455 0.0088229 0.0097846 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16038 0.94069 0.91775 0.0013968 0.99348 0.51562 0.0018818 0.42772 2.1033 2.1027 16.0069 144.943 0.00016191 -85.6546 0.83795
6.942 0.98811 5.4773e-005 3.8183 0.011946 9.0476e-005 0.0011673 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.4478 0.51067 0.15611 0.018601 13.1149 0.1156 0.00014906 0.77455 0.0088233 0.0097851 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16038 0.94083 0.9178 0.0013968 0.9935 0.51579 0.0018818 0.42773 2.1037 2.1031 16.0068 144.943 0.00016183 -85.6547 0.83895
6.943 0.98811 5.4773e-005 3.8183 0.011946 9.0489e-005 0.0011673 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.4479 0.51072 0.15612 0.018602 13.1175 0.11561 0.00014907 0.77454 0.0088238 0.0097855 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16038 0.94096 0.91785 0.0013968 0.99353 0.51596 0.0018818 0.42775 2.1041 2.1035 16.0068 144.943 0.00016175 -85.6547 0.83995
6.944 0.98811 5.4773e-005 3.8183 0.011946 9.0501e-005 0.0011673 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.4479 0.51076 0.15614 0.018604 13.1201 0.11562 0.00014908 0.77453 0.0088243 0.009786 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16039 0.94109 0.9179 0.0013968 0.99355 0.51613 0.0018818 0.42776 2.1045 2.1039 16.0068 144.9431 0.00016167 -85.6548 0.84095
6.945 0.98811 5.4773e-005 3.8183 0.011946 9.0514e-005 0.0011673 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.448 0.51081 0.15615 0.018605 13.1227 0.11563 0.00014909 0.77452 0.0088247 0.0097865 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16039 0.94122 0.91795 0.0013967 0.99357 0.5163 0.0018817 0.42777 2.1049 2.1043 16.0067 144.9431 0.00016159 -85.6549 0.84195
6.946 0.98811 5.4773e-005 3.8183 0.011946 9.0527e-005 0.0011673 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.4481 0.51085 0.15616 0.018606 13.1252 0.11563 0.0001491 0.77452 0.0088252 0.009787 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.1604 0.94136 0.918 0.0013967 0.9936 0.51646 0.0018817 0.42779 2.1053 2.1047 16.0067 144.9431 0.00016151 -85.655 0.84295
6.947 0.98811 5.4773e-005 3.8183 0.011946 9.054e-005 0.0011673 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.4482 0.5109 0.15618 0.018607 13.1278 0.11564 0.00014912 0.77451 0.0088256 0.0097875 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.1604 0.94149 0.91805 0.0013967 0.99362 0.51663 0.0018817 0.4278 2.1057 2.1052 16.0067 144.9431 0.00016143 -85.655 0.84395
6.948 0.98812 5.4773e-005 3.8183 0.011946 9.0553e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4483 0.51095 0.15619 0.018608 13.1304 0.11565 0.00014913 0.7745 0.0088261 0.009788 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.1604 0.94162 0.9181 0.0013967 0.99364 0.5168 0.0018817 0.42781 2.1061 2.1056 16.0066 144.9431 0.00016136 -85.6551 0.84495
6.949 0.98812 5.4772e-005 3.8183 0.011946 9.0566e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4484 0.51099 0.15621 0.01861 13.133 0.11566 0.00014914 0.77449 0.0088266 0.0097885 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.16041 0.94175 0.91815 0.0013967 0.99367 0.51697 0.0018817 0.42783 2.1065 2.106 16.0066 144.9432 0.00016128 -85.6552 0.84595
6.95 0.98812 5.4772e-005 3.8183 0.011946 9.0579e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4485 0.51104 0.15622 0.018611 13.1356 0.11566 0.00014915 0.77449 0.008827 0.009789 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.16041 0.94188 0.9182 0.0013967 0.99369 0.51714 0.0018817 0.42784 2.1069 2.1064 16.0066 144.9432 0.0001612 -85.6552 0.84695
6.951 0.98812 5.4772e-005 3.8183 0.011946 9.0592e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4486 0.51108 0.15624 0.018612 13.1382 0.11567 0.00014916 0.77448 0.0088275 0.0097895 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.16041 0.94201 0.91825 0.0013967 0.99371 0.51731 0.0018817 0.42785 2.1073 2.1068 16.0066 144.9432 0.00016112 -85.6553 0.84795
6.952 0.98812 5.4772e-005 3.8183 0.011946 9.0604e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4487 0.51113 0.15625 0.018613 13.1407 0.11568 0.00014917 0.77447 0.008828 0.00979 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16042 0.94214 0.9183 0.0013966 0.99374 0.51747 0.0018817 0.42787 2.1077 2.1072 16.0065 144.9432 0.00016104 -85.6554 0.84895
6.953 0.98812 5.4772e-005 3.8183 0.011946 9.0617e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4488 0.51117 0.15626 0.018615 13.1433 0.11569 0.00014918 0.77446 0.0088284 0.0097905 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16042 0.94227 0.91835 0.0013966 0.99376 0.51764 0.0018817 0.42788 2.1081 2.1076 16.0065 144.9432 0.00016097 -85.6555 0.84995
6.954 0.98812 5.4772e-005 3.8183 0.011946 9.063e-005 0.0011674 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4488 0.51122 0.15628 0.018616 13.1459 0.11569 0.00014919 0.77446 0.0088289 0.009791 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16042 0.9424 0.9184 0.0013966 0.99378 0.51781 0.0018816 0.42789 2.1085 2.108 16.0065 144.9433 0.00016089 -85.6555 0.85095
6.955 0.98812 5.4772e-005 3.8183 0.011946 9.0643e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4489 0.51127 0.15629 0.018617 13.1485 0.1157 0.0001492 0.77445 0.0088294 0.0097915 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16043 0.94253 0.91845 0.0013966 0.9938 0.51798 0.0018816 0.42791 2.1089 2.1084 16.0064 144.9433 0.00016081 -85.6556 0.85195
6.956 0.98812 5.4772e-005 3.8183 0.011946 9.0656e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.449 0.51131 0.15631 0.018618 13.1511 0.11571 0.00014922 0.77444 0.0088298 0.009792 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16043 0.94266 0.9185 0.0013966 0.99382 0.51815 0.0018816 0.42792 2.1093 2.1088 16.0064 144.9433 0.00016074 -85.6557 0.85295
6.957 0.98812 5.4772e-005 3.8183 0.011946 9.0669e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4491 0.51136 0.15632 0.01862 13.1537 0.11572 0.00014923 0.77443 0.0088303 0.0097925 0.0013854 0.98696 0.99171 2.9872e-006 1.1949e-005 0.16043 0.94278 0.91855 0.0013966 0.99385 0.51831 0.0018816 0.42793 2.1097 2.1092 16.0064 144.9433 0.00016066 -85.6557 0.85395
6.958 0.98812 5.4772e-005 3.8183 0.011946 9.0682e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4492 0.5114 0.15634 0.018621 13.1563 0.11572 0.00014924 0.77443 0.0088307 0.009793 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16044 0.94291 0.9186 0.0013966 0.99387 0.51848 0.0018816 0.42794 2.1101 2.1096 16.0063 144.9433 0.00016058 -85.6558 0.85495
6.959 0.98812 5.4772e-005 3.8183 0.011946 9.0695e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4493 0.51145 0.15635 0.018622 13.1589 0.11573 0.00014925 0.77442 0.0088312 0.0097935 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16044 0.94304 0.91865 0.0013966 0.99389 0.51865 0.0018816 0.42796 2.1105 2.11 16.0063 144.9434 0.00016051 -85.6558 0.85595
6.96 0.98812 5.4772e-005 3.8183 0.011946 9.0707e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4494 0.51149 0.15636 0.018623 13.1614 0.11574 0.00014926 0.77441 0.0088317 0.009794 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16045 0.94317 0.9187 0.0013966 0.99391 0.51882 0.0018816 0.42797 2.1109 2.1104 16.0063 144.9434 0.00016043 -85.6559 0.85695
6.961 0.98812 5.4771e-005 3.8183 0.011946 9.072e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4495 0.51154 0.15638 0.018625 13.164 0.11575 0.00014927 0.7744 0.0088321 0.0097945 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16045 0.94329 0.91875 0.0013966 0.99393 0.51898 0.0018816 0.42798 2.1113 2.1108 16.0062 144.9434 0.00016036 -85.656 0.85795
6.962 0.98812 5.4771e-005 3.8183 0.011946 9.0733e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4496 0.51158 0.15639 0.018626 13.1666 0.11575 0.00014928 0.7744 0.0088326 0.009795 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16045 0.94342 0.91879 0.0013966 0.99395 0.51915 0.0018816 0.428 2.1117 2.1112 16.0062 144.9434 0.00016028 -85.656 0.85895
6.963 0.98812 5.4771e-005 3.8183 0.011946 9.0746e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4497 0.51163 0.15641 0.018627 13.1692 0.11576 0.00014929 0.77439 0.0088331 0.0097955 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16046 0.94354 0.91884 0.0013966 0.99397 0.51932 0.0018815 0.42801 2.1121 2.1115 16.0062 144.9434 0.00016021 -85.6561 0.85995
6.964 0.98812 5.4771e-005 3.8183 0.011946 9.0759e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4497 0.51168 0.15642 0.018628 13.1718 0.11577 0.0001493 0.77438 0.0088335 0.009796 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16046 0.94367 0.91889 0.0013966 0.99399 0.51949 0.0018815 0.42802 2.1125 2.1119 16.0062 144.9435 0.00016013 -85.6562 0.86095
6.965 0.98812 5.4771e-005 3.8183 0.011946 9.0772e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4498 0.51172 0.15644 0.01863 13.1744 0.11578 0.00014932 0.77437 0.008834 0.0097965 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16046 0.94379 0.91894 0.0013966 0.99402 0.51965 0.0018815 0.42804 2.1129 2.1123 16.0061 144.9435 0.00016006 -85.6562 0.86195
6.966 0.98812 5.4771e-005 3.8183 0.011946 9.0785e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4499 0.51177 0.15645 0.018631 13.177 0.11578 0.00014933 0.77437 0.0088344 0.009797 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16047 0.94392 0.91898 0.0013966 0.99404 0.51982 0.0018815 0.42805 2.1133 2.1127 16.0061 144.9435 0.00015999 -85.6563 0.86295
6.967 0.98812 5.4771e-005 3.8183 0.011946 9.0798e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.45 0.51181 0.15646 0.018632 13.1796 0.11579 0.00014934 0.77436 0.0088349 0.0097975 0.0013853 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16047 0.94404 0.91903 0.0013966 0.99406 0.51999 0.0018815 0.42806 2.1137 2.1131 16.0061 144.9435 0.00015991 -85.6564 0.86395
6.968 0.98812 5.4771e-005 3.8183 0.011946 9.081e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4501 0.51186 0.15648 0.018633 13.1822 0.1158 0.00014935 0.77435 0.0088354 0.009798 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16047 0.94416 0.91908 0.0013966 0.99408 0.52016 0.0018815 0.42807 2.114 2.1135 16.006 144.9435 0.00015984 -85.6564 0.86495
6.969 0.98812 5.4771e-005 3.8183 0.011946 9.0823e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4502 0.5119 0.15649 0.018635 13.1848 0.11581 0.00014936 0.77434 0.0088358 0.0097984 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16048 0.94429 0.91913 0.0013966 0.9941 0.52032 0.0018815 0.42809 2.1144 2.1139 16.006 144.9436 0.00015977 -85.6565 0.86595
6.97 0.98812 5.4771e-005 3.8183 0.011946 9.0836e-005 0.0011674 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.4503 0.51195 0.15651 0.018636 13.1874 0.11581 0.00014937 0.77434 0.0088363 0.0097989 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16048 0.94441 0.91917 0.0013965 0.99412 0.52049 0.0018815 0.4281 2.1148 2.1143 16.006 144.9436 0.00015969 -85.6565 0.86695
6.971 0.98812 5.4771e-005 3.8183 0.011946 9.0849e-005 0.0011674 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.4504 0.512 0.15652 0.018637 13.1899 0.11582 0.00014938 0.77433 0.0088368 0.0097994 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16049 0.94453 0.91922 0.0013965 0.99414 0.52066 0.0018815 0.42811 2.1152 2.1147 16.0059 144.9436 0.00015962 -85.6566 0.86795
6.972 0.98812 5.4771e-005 3.8183 0.011946 9.0862e-005 0.0011675 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.4505 0.51204 0.15654 0.018638 13.1925 0.11583 0.00014939 0.77432 0.0088372 0.0097999 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16049 0.94465 0.91927 0.0013965 0.99416 0.52082 0.0018815 0.42813 2.1156 2.1151 16.0059 144.9436 0.00015955 -85.6567 0.86895
6.973 0.98812 5.4771e-005 3.8183 0.011946 9.0875e-005 0.0011675 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.4506 0.51209 0.15655 0.01864 13.1951 0.11584 0.0001494 0.77431 0.0088377 0.0098004 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16049 0.94478 0.91931 0.0013965 0.99418 0.52099 0.0018815 0.42814 2.116 2.1155 16.0059 144.9437 0.00015948 -85.6567 0.86995
6.974 0.98812 5.477e-005 3.8183 0.011946 9.0888e-005 0.0011675 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.4506 0.51213 0.15657 0.018641 13.1977 0.11584 0.00014942 0.77431 0.0088381 0.0098009 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.1605 0.9449 0.91936 0.0013965 0.9942 0.52116 0.0018814 0.42815 2.1164 2.1158 16.0058 144.9437 0.0001594 -85.6568 0.87095
6.975 0.98812 5.477e-005 3.8183 0.011946 9.0901e-005 0.0011675 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.4507 0.51218 0.15658 0.018642 13.2003 0.11585 0.00014943 0.7743 0.0088386 0.0098014 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.1605 0.94502 0.91941 0.0013965 0.99421 0.52133 0.0018814 0.42817 2.1168 2.1162 16.0058 144.9437 0.00015933 -85.6568 0.87195
6.976 0.98812 5.477e-005 3.8183 0.011946 9.0913e-005 0.0011675 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.4508 0.51222 0.15659 0.018643 13.2029 0.11586 0.00014944 0.77429 0.0088391 0.0098019 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.1605 0.94514 0.91945 0.0013965 0.99423 0.52149 0.0018814 0.42818 2.1171 2.1166 16.0058 144.9437 0.00015926 -85.6569 0.87295
6.977 0.98812 5.477e-005 3.8183 0.011946 9.0926e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4509 0.51227 0.15661 0.018645 13.2055 0.11587 0.00014945 0.77428 0.0088395 0.0098024 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16051 0.94526 0.9195 0.0013965 0.99425 0.52166 0.0018814 0.42819 2.1175 2.117 16.0057 144.9437 0.00015919 -85.6569 0.87395
6.978 0.98812 5.477e-005 3.8183 0.011946 9.0939e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.451 0.51232 0.15662 0.018646 13.2081 0.11587 0.00014946 0.77428 0.00884 0.0098029 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16051 0.94538 0.91954 0.0013965 0.99427 0.52183 0.0018814 0.4282 2.1179 2.1174 16.0057 144.9438 0.00015912 -85.657 0.87495
6.979 0.98812 5.477e-005 3.8183 0.011946 9.0952e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4511 0.51236 0.15664 0.018647 13.2107 0.11588 0.00014947 0.77427 0.0088405 0.0098034 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16051 0.9455 0.91959 0.0013964 0.99429 0.52199 0.0018814 0.42822 2.1183 2.1178 16.0057 144.9438 0.00015905 -85.657 0.87595
6.98 0.98812 5.477e-005 3.8183 0.011946 9.0965e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4512 0.51241 0.15665 0.018648 13.2133 0.11589 0.00014948 0.77426 0.0088409 0.0098039 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.16052 0.94562 0.91963 0.0013964 0.99431 0.52216 0.0018814 0.42823 2.1187 2.1181 16.0057 144.9438 0.00015898 -85.6571 0.87695
6.981 0.98812 5.477e-005 3.8183 0.011946 9.0978e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4513 0.51245 0.15667 0.018649 13.2159 0.1159 0.00014949 0.77425 0.0088414 0.0098044 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.16052 0.94573 0.91968 0.0013964 0.99433 0.52233 0.0018814 0.42824 2.119 2.1185 16.0056 144.9438 0.00015891 -85.6572 0.87795
6.982 0.98812 5.477e-005 3.8183 0.011946 9.0991e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4514 0.5125 0.15668 0.018651 13.2185 0.1159 0.0001495 0.77425 0.0088418 0.0098049 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.16052 0.94585 0.91972 0.0013964 0.99435 0.52249 0.0018814 0.42826 2.1194 2.1189 16.0056 144.9438 0.00015884 -85.6572 0.87895
6.983 0.98812 5.477e-005 3.8183 0.011946 9.1003e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4514 0.51254 0.15669 0.018652 13.2211 0.11591 0.00014952 0.77424 0.0088423 0.0098054 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.16053 0.94597 0.91977 0.0013964 0.99437 0.52266 0.0018814 0.42827 2.1198 2.1193 16.0056 144.9439 0.00015877 -85.6573 0.87995
6.984 0.98812 5.477e-005 3.8183 0.011945 9.1016e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4515 0.51259 0.15671 0.018653 13.2237 0.11592 0.00014953 0.77423 0.0088428 0.0098059 0.001385 0.98696 0.99171 2.9863e-006 1.1945e-005 0.16053 0.94609 0.91981 0.0013964 0.99438 0.52282 0.0018814 0.42828 2.1202 2.1197 16.0055 144.9439 0.0001587 -85.6573 0.88095
6.985 0.98812 5.477e-005 3.8183 0.011945 9.1029e-005 0.0011675 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4516 0.51263 0.15672 0.018654 13.2263 0.11593 0.00014954 0.77422 0.0088432 0.0098064 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16054 0.9462 0.91986 0.0013964 0.9944 0.52299 0.0018813 0.42829 2.1206 2.12 16.0055 144.9439 0.00015863 -85.6574 0.88195
6.986 0.98812 5.4769e-005 3.8183 0.011945 9.1042e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4517 0.51268 0.15674 0.018656 13.2289 0.11593 0.00014955 0.77422 0.0088437 0.0098068 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16054 0.94632 0.9199 0.0013964 0.99442 0.52316 0.0018813 0.42831 2.1209 2.1204 16.0055 144.9439 0.00015856 -85.6574 0.88295
6.987 0.98812 5.4769e-005 3.8183 0.011945 9.1055e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4518 0.51273 0.15675 0.018657 13.2315 0.11594 0.00014956 0.77421 0.0088441 0.0098073 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16054 0.94644 0.91995 0.0013964 0.99444 0.52332 0.0018813 0.42832 2.1213 2.1208 16.0054 144.9439 0.00015849 -85.6575 0.88395
6.988 0.98812 5.4769e-005 3.8183 0.011945 9.1068e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4519 0.51277 0.15677 0.018658 13.2341 0.11595 0.00014957 0.7742 0.0088446 0.0098078 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16055 0.94655 0.91999 0.0013964 0.99446 0.52349 0.0018813 0.42833 2.1217 2.1212 16.0054 144.944 0.00015842 -85.6575 0.88495
6.989 0.98812 5.4769e-005 3.8183 0.011945 9.1081e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.452 0.51282 0.15678 0.018659 13.2367 0.11595 0.00014958 0.77419 0.0088451 0.0098083 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16055 0.94667 0.92003 0.0013964 0.99447 0.52365 0.0018813 0.42835 2.1221 2.1216 16.0054 144.944 0.00015835 -85.6576 0.88595
6.99 0.98812 5.4769e-005 3.8183 0.011945 9.1094e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4521 0.51286 0.15679 0.018661 13.2393 0.11596 0.00014959 0.77419 0.0088455 0.0098088 0.001385 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16055 0.94678 0.92008 0.0013964 0.99449 0.52382 0.0018813 0.42836 2.1224 2.1219 16.0053 144.944 0.00015829 -85.6576 0.88695
6.991 0.98812 5.4769e-005 3.8183 0.011945 9.1106e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4522 0.51291 0.15681 0.018662 13.2419 0.11597 0.0001496 0.77418 0.008846 0.0098093 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16056 0.9469 0.92012 0.0013964 0.99451 0.52399 0.0018813 0.42837 2.1228 2.1223 16.0053 144.944 0.00015822 -85.6577 0.88795
6.992 0.98812 5.4769e-005 3.8183 0.011945 9.1119e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4523 0.51295 0.15682 0.018663 13.2445 0.11598 0.00014961 0.77417 0.0088464 0.0098098 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16056 0.94701 0.92017 0.0013964 0.99453 0.52415 0.0018813 0.42838 2.1232 2.1227 16.0053 144.944 0.00015815 -85.6577 0.88895
6.993 0.98812 5.4769e-005 3.8183 0.011945 9.1132e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4523 0.513 0.15684 0.018664 13.2471 0.11598 0.00014963 0.77416 0.0088469 0.0098103 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16056 0.94713 0.92021 0.0013964 0.99454 0.52432 0.0018813 0.4284 2.1236 2.1231 16.0052 144.9441 0.00015808 -85.6578 0.88995
6.994 0.98812 5.4769e-005 3.8183 0.011945 9.1145e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4524 0.51305 0.15685 0.018666 13.2497 0.11599 0.00014964 0.77416 0.0088474 0.0098108 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16057 0.94724 0.92025 0.0013964 0.99456 0.52448 0.0018813 0.42841 2.1239 2.1234 16.0052 144.9441 0.00015802 -85.6578 0.89095
6.995 0.98812 5.4769e-005 3.8183 0.011945 9.1158e-005 0.0011675 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4525 0.51309 0.15687 0.018667 13.2523 0.116 0.00014965 0.77415 0.0088478 0.0098113 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16057 0.94735 0.92029 0.0013964 0.99458 0.52465 0.0018813 0.42842 2.1243 2.1238 16.0052 144.9441 0.00015795 -85.6579 0.89195
6.996 0.98812 5.4769e-005 3.8183 0.011945 9.1171e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4526 0.51314 0.15688 0.018668 13.2549 0.11601 0.00014966 0.77414 0.0088483 0.0098118 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16057 0.94747 0.92034 0.0013964 0.99459 0.52482 0.0018813 0.42844 2.1247 2.1242 16.0051 144.9441 0.00015788 -85.6579 0.89295
6.997 0.98812 5.4769e-005 3.8183 0.011945 9.1184e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4527 0.51318 0.15689 0.018669 13.2575 0.11601 0.00014967 0.77413 0.0088487 0.0098123 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16058 0.94758 0.92038 0.0013964 0.99461 0.52498 0.0018812 0.42845 2.125 2.1245 16.0051 144.9441 0.00015782 -85.658 0.89395
6.998 0.98812 5.4769e-005 3.8183 0.011945 9.1197e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4528 0.51323 0.15691 0.018671 13.2601 0.11602 0.00014968 0.77413 0.0088492 0.0098128 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16058 0.94769 0.92042 0.0013964 0.99463 0.52515 0.0018812 0.42846 2.1254 2.1249 16.0051 144.9442 0.00015775 -85.658 0.89495
6.999 0.98812 5.4768e-005 3.8183 0.011945 9.1209e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4529 0.51327 0.15692 0.018672 13.2627 0.11603 0.00014969 0.77412 0.0088497 0.0098133 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16059 0.94781 0.92047 0.0013963 0.99464 0.52531 0.0018812 0.42847 2.1258 2.1253 16.005 144.9442 0.00015768 -85.6581 0.89595
7 0.98812 5.4768e-005 3.8183 0.011945 9.1222e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.453 0.51332 0.15694 0.018673 13.2653 0.11604 0.0001497 0.77411 0.0088501 0.0098138 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16059 0.94792 0.92051 0.0013963 0.99466 0.52548 0.0018812 0.42849 2.1262 2.1256 16.005 144.9442 0.00015762 -85.6581 0.89695
7.001 0.98812 5.4768e-005 3.8183 0.011945 9.1235e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4531 0.51336 0.15695 0.018674 13.2679 0.11604 0.00014971 0.77411 0.0088506 0.0098142 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16059 0.94803 0.92055 0.0013963 0.99468 0.52564 0.0018812 0.4285 2.1265 2.126 16.005 144.9442 0.00015755 -85.6582 0.89795
7.002 0.98812 5.4768e-005 3.8183 0.011945 9.1248e-005 0.0011676 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.4532 0.51341 0.15697 0.018675 13.2705 0.11605 0.00014973 0.7741 0.008851 0.0098147 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.1606 0.94814 0.92059 0.0013963 0.99469 0.52581 0.0018812 0.42851 2.1269 2.1264 16.005 144.9442 0.00015749 -85.6582 0.89895
7.003 0.98812 5.4768e-005 3.8183 0.011945 9.1261e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4532 0.51346 0.15698 0.018677 13.2731 0.11606 0.00014974 0.77409 0.0088515 0.0098152 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.1606 0.94825 0.92063 0.0013963 0.99471 0.52597 0.0018812 0.42853 2.1273 2.1268 16.0049 144.9443 0.00015742 -85.6583 0.89995
7.004 0.98812 5.4768e-005 3.8183 0.011945 9.1274e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4533 0.5135 0.15699 0.018678 13.2757 0.11607 0.00014975 0.77408 0.008852 0.0098157 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.1606 0.94836 0.92068 0.0013963 0.99472 0.52614 0.0018812 0.42854 2.1276 2.1271 16.0049 144.9443 0.00015736 -85.6583 0.90095
7.005 0.98812 5.4768e-005 3.8183 0.011945 9.1287e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4534 0.51355 0.15701 0.018679 13.2783 0.11607 0.00014976 0.77408 0.0088524 0.0098162 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16061 0.94847 0.92072 0.0013963 0.99474 0.5263 0.0018812 0.42855 2.128 2.1275 16.0049 144.9443 0.00015729 -85.6584 0.90195
7.006 0.98812 5.4768e-005 3.8183 0.011945 9.13e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4535 0.51359 0.15702 0.01868 13.2809 0.11608 0.00014977 0.77407 0.0088529 0.0098167 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16061 0.94858 0.92076 0.0013963 0.99476 0.52647 0.0018812 0.42856 2.1283 2.1278 16.0048 144.9443 0.00015723 -85.6584 0.90295
7.007 0.98812 5.4768e-005 3.8183 0.011945 9.1312e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4536 0.51364 0.15704 0.018682 13.2835 0.11609 0.00014978 0.77406 0.0088533 0.0098172 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16061 0.94869 0.9208 0.0013963 0.99477 0.52663 0.0018812 0.42858 2.1287 2.1282 16.0048 144.9443 0.00015716 -85.6584 0.90395
7.008 0.98812 5.4768e-005 3.8183 0.011945 9.1325e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4537 0.51368 0.15705 0.018683 13.2861 0.1161 0.00014979 0.77405 0.0088538 0.0098177 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16062 0.9488 0.92084 0.0013963 0.99479 0.5268 0.0018812 0.42859 2.1291 2.1286 16.0048 144.9444 0.0001571 -85.6585 0.90495
7.009 0.98812 5.4768e-005 3.8183 0.011945 9.1338e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4538 0.51373 0.15707 0.018684 13.2887 0.1161 0.0001498 0.77405 0.0088543 0.0098182 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16062 0.94891 0.92088 0.0013963 0.9948 0.52696 0.0018812 0.4286 2.1294 2.1289 16.0047 144.9444 0.00015703 -85.6585 0.90595
7.01 0.98812 5.4768e-005 3.8183 0.011945 9.1351e-005 0.0011676 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.4539 0.51378 0.15708 0.018685 13.2913 0.11611 0.00014981 0.77404 0.0088547 0.0098187 0.0013847 0.98696 0.99172 2.9857e-006 1.1942e-005 0.16062 0.94901 0.92092 0.0013962 0.99482 0.52713 0.0018812 0.42862 2.1298 2.1293 16.0047 144.9444 0.00015697 -85.6586 0.90695
7.011 0.98812 5.4768e-005 3.8183 0.011945 9.1364e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032263 0.0389 0 1.454 0.51382 0.15709 0.018687 13.2939 0.11612 0.00014983 0.77403 0.0088552 0.0098192 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16063 0.94912 0.92096 0.0013962 0.99483 0.52729 0.0018811 0.42863 2.1302 2.1297 16.0047 144.9444 0.00015691 -85.6586 0.90795
7.012 0.98812 5.4767e-005 3.8183 0.011945 9.1377e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4541 0.51387 0.15711 0.018688 13.2965 0.11613 0.00014984 0.77402 0.0088556 0.0098197 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16063 0.94923 0.921 0.0013962 0.99485 0.52746 0.0018811 0.42864 2.1305 2.13 16.0046 144.9445 0.00015684 -85.6587 0.90895
7.013 0.98812 5.4767e-005 3.8183 0.011945 9.139e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4541 0.51391 0.15712 0.018689 13.2991 0.11613 0.00014985 0.77402 0.0088561 0.0098201 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16064 0.94934 0.92105 0.0013962 0.99486 0.52762 0.0018811 0.42865 2.1309 2.1304 16.0046 144.9445 0.00015678 -85.6587 0.90995
7.014 0.98812 5.4767e-005 3.8183 0.011945 9.1403e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4542 0.51396 0.15714 0.01869 13.3018 0.11614 0.00014986 0.77401 0.0088566 0.0098206 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16064 0.94944 0.92109 0.0013962 0.99488 0.52779 0.0018811 0.42867 2.1312 2.1307 16.0046 144.9445 0.00015672 -85.6587 0.91095
7.015 0.98812 5.4767e-005 3.8183 0.011945 9.1415e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4543 0.514 0.15715 0.018692 13.3044 0.11615 0.00014987 0.774 0.008857 0.0098211 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16064 0.94955 0.92113 0.0013962 0.99489 0.52795 0.0018811 0.42868 2.1316 2.1311 16.0045 144.9445 0.00015665 -85.6588 0.91195
7.016 0.98812 5.4767e-005 3.8183 0.011945 9.1428e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4544 0.51405 0.15717 0.018693 13.307 0.11616 0.00014988 0.77399 0.0088575 0.0098216 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16065 0.94966 0.92117 0.0013962 0.99491 0.52812 0.0018811 0.42869 2.132 2.1315 16.0045 144.9445 0.00015659 -85.6588 0.91295
7.017 0.98812 5.4767e-005 3.8183 0.011945 9.1441e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4545 0.51409 0.15718 0.018694 13.3096 0.11616 0.00014989 0.77399 0.0088579 0.0098221 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16065 0.94976 0.92121 0.0013962 0.99492 0.52828 0.0018811 0.4287 2.1323 2.1318 16.0045 144.9446 0.00015653 -85.6589 0.91395
7.018 0.98812 5.4767e-005 3.8183 0.011945 9.1454e-005 0.0011676 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4546 0.51414 0.15719 0.018695 13.3122 0.11617 0.0001499 0.77398 0.0088584 0.0098226 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16065 0.94987 0.92125 0.0013962 0.99494 0.52844 0.0018811 0.42872 2.1327 2.1322 16.0044 144.9446 0.00015647 -85.6589 0.91495
7.019 0.98812 5.4767e-005 3.8183 0.011945 9.1467e-005 0.0011676 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4547 0.51419 0.15721 0.018696 13.3148 0.11618 0.00014991 0.77397 0.0088589 0.0098231 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16066 0.94997 0.92129 0.0013962 0.99495 0.52861 0.0018811 0.42873 2.133 2.1325 16.0044 144.9446 0.00015641 -85.6589 0.91595
7.02 0.98812 5.4767e-005 3.8183 0.011945 9.148e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4548 0.51423 0.15722 0.018698 13.3174 0.11619 0.00014992 0.77396 0.0088593 0.0098236 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.16066 0.95008 0.92132 0.0013962 0.99497 0.52877 0.0018811 0.42874 2.1334 2.1329 16.0044 144.9446 0.00015634 -85.659 0.91695
7.021 0.98812 5.4767e-005 3.8183 0.011945 9.1493e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4549 0.51428 0.15724 0.018699 13.32 0.11619 0.00014994 0.77396 0.0088598 0.0098241 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.16066 0.95018 0.92136 0.0013962 0.99498 0.52894 0.0018811 0.42876 2.1337 2.1333 16.0043 144.9446 0.00015628 -85.659 0.91795
7.022 0.98812 5.4767e-005 3.8183 0.011945 9.1505e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4549 0.51432 0.15725 0.0187 13.3226 0.1162 0.00014995 0.77395 0.0088602 0.0098246 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16067 0.95029 0.9214 0.0013962 0.995 0.5291 0.0018811 0.42877 2.1341 2.1336 16.0043 144.9447 0.00015622 -85.6591 0.91895
7.023 0.98812 5.4767e-005 3.8183 0.011945 9.1518e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.455 0.51437 0.15727 0.018701 13.3252 0.11621 0.00014996 0.77394 0.0088607 0.0098251 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16067 0.95039 0.92144 0.0013962 0.99501 0.52927 0.0018811 0.42878 2.1344 2.134 16.0043 144.9447 0.00015616 -85.6591 0.91995
7.024 0.98812 5.4766e-005 3.8183 0.011945 9.1531e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4551 0.51441 0.15728 0.018703 13.3278 0.11622 0.00014997 0.77393 0.0088611 0.0098255 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16067 0.95049 0.92148 0.0013962 0.99502 0.52943 0.0018811 0.42879 2.1348 2.1343 16.0042 144.9447 0.0001561 -85.6591 0.92095
7.025 0.98812 5.4766e-005 3.8183 0.011945 9.1544e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4552 0.51446 0.15729 0.018704 13.3305 0.11622 0.00014998 0.77393 0.0088616 0.009826 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16068 0.9506 0.92152 0.0013962 0.99504 0.52959 0.0018811 0.42881 2.1352 2.1347 16.0042 144.9447 0.00015604 -85.6592 0.92195
7.026 0.98812 5.4766e-005 3.8183 0.011945 9.1557e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4553 0.51451 0.15731 0.018705 13.3331 0.11623 0.00014999 0.77392 0.0088621 0.0098265 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16068 0.9507 0.92156 0.0013962 0.99505 0.52976 0.001881 0.42882 2.1355 2.135 16.0042 144.9447 0.00015598 -85.6592 0.92295
7.027 0.98812 5.4766e-005 3.8183 0.011945 9.157e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4554 0.51455 0.15732 0.018706 13.3357 0.11624 0.00015 0.77391 0.0088625 0.009827 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16069 0.9508 0.9216 0.0013962 0.99507 0.52992 0.001881 0.42883 2.1359 2.1354 16.0041 144.9448 0.00015592 -85.6593 0.92395
7.028 0.98812 5.4766e-005 3.8183 0.011945 9.1583e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4555 0.5146 0.15734 0.018708 13.3383 0.11625 0.00015001 0.7739 0.008863 0.0098275 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16069 0.95091 0.92164 0.0013962 0.99508 0.53008 0.001881 0.42884 2.1362 2.1357 16.0041 144.9448 0.00015586 -85.6593 0.92495
7.029 0.98812 5.4766e-005 3.8183 0.011945 9.1596e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4556 0.51464 0.15735 0.018709 13.3409 0.11625 0.00015002 0.7739 0.0088634 0.009828 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16069 0.95101 0.92168 0.0013962 0.99509 0.53025 0.001881 0.42886 2.1366 2.1361 16.0041 144.9448 0.0001558 -85.6593 0.92595
7.03 0.98812 5.4766e-005 3.8183 0.011945 9.1608e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4557 0.51469 0.15737 0.01871 13.3435 0.11626 0.00015004 0.77389 0.0088639 0.0098285 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1607 0.95111 0.92171 0.0013962 0.99511 0.53041 0.001881 0.42887 2.1369 2.1364 16.004 144.9448 0.00015574 -85.6594 0.92695
7.031 0.98812 5.4766e-005 3.8183 0.011945 9.1621e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4558 0.51473 0.15738 0.018711 13.3461 0.11627 0.00015005 0.77388 0.0088644 0.009829 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1607 0.95121 0.92175 0.0013962 0.99512 0.53058 0.001881 0.42888 2.1373 2.1368 16.004 144.9448 0.00015568 -85.6594 0.92795
7.032 0.98812 5.4766e-005 3.8183 0.011945 9.1634e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4558 0.51478 0.15739 0.018712 13.3487 0.11628 0.00015006 0.77387 0.0088648 0.0098295 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1607 0.95131 0.92179 0.0013961 0.99513 0.53074 0.001881 0.4289 2.1376 2.1371 16.004 144.9449 0.00015562 -85.6594 0.92895
7.033 0.98812 5.4766e-005 3.8183 0.011945 9.1647e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4559 0.51482 0.15741 0.018714 13.3514 0.11628 0.00015007 0.77387 0.0088653 0.00983 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16071 0.95141 0.92183 0.0013961 0.99515 0.5309 0.001881 0.42891 2.138 2.1375 16.0039 144.9449 0.00015556 -85.6595 0.92995
7.034 0.98812 5.4766e-005 3.8183 0.011945 9.166e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.456 0.51487 0.15742 0.018715 13.354 0.11629 0.00015008 0.77386 0.0088657 0.0098304 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16071 0.95151 0.92187 0.0013961 0.99516 0.53107 0.001881 0.42892 2.1383 2.1378 16.0039 144.9449 0.0001555 -85.6595 0.93095
7.035 0.98812 5.4766e-005 3.8183 0.011945 9.1673e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4561 0.51492 0.15744 0.018716 13.3566 0.1163 0.00015009 0.77385 0.0088662 0.0098309 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16071 0.95161 0.9219 0.0013961 0.99517 0.53123 0.001881 0.42893 2.1386 2.1382 16.0039 144.9449 0.00015544 -85.6596 0.93195
7.036 0.98812 5.4766e-005 3.8183 0.011945 9.1686e-005 0.0011677 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.4562 0.51496 0.15745 0.018717 13.3592 0.11631 0.0001501 0.77384 0.0088666 0.0098314 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16072 0.95171 0.92194 0.0013961 0.99519 0.53139 0.001881 0.42895 2.139 2.1385 16.0038 144.9449 0.00015539 -85.6596 0.93295
7.037 0.98812 5.4765e-005 3.8183 0.011945 9.1699e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4563 0.51501 0.15747 0.018719 13.3618 0.11631 0.00015011 0.77384 0.0088671 0.0098319 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16072 0.95181 0.92198 0.0013961 0.9952 0.53156 0.001881 0.42896 2.1393 2.1389 16.0038 144.945 0.00015533 -85.6596 0.93395
7.038 0.98812 5.4765e-005 3.8183 0.011945 9.1711e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4564 0.51505 0.15748 0.01872 13.3644 0.11632 0.00015012 0.77383 0.0088676 0.0098324 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16072 0.95191 0.92201 0.0013961 0.99521 0.53172 0.001881 0.42897 2.1397 2.1392 16.0038 144.945 0.00015527 -85.6597 0.93495
7.039 0.98812 5.4765e-005 3.8183 0.011945 9.1724e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4565 0.5151 0.15749 0.018721 13.367 0.11633 0.00015013 0.77382 0.008868 0.0098329 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16073 0.95201 0.92205 0.0013961 0.99522 0.53188 0.001881 0.42898 2.14 2.1396 16.0037 144.945 0.00015521 -85.6597 0.93595
7.04 0.98812 5.4765e-005 3.8183 0.011945 9.1737e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4566 0.51514 0.15751 0.018722 13.3697 0.11634 0.00015015 0.77382 0.0088685 0.0098334 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16073 0.95211 0.92209 0.0013961 0.99524 0.53205 0.001881 0.429 2.1404 2.1399 16.0037 144.945 0.00015515 -85.6597 0.93695
7.041 0.98812 5.4765e-005 3.8183 0.011945 9.175e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4567 0.51519 0.15752 0.018724 13.3723 0.11634 0.00015016 0.77381 0.0088689 0.0098339 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16074 0.95221 0.92213 0.0013961 0.99525 0.53221 0.001881 0.42901 2.1407 2.1402 16.0037 144.945 0.0001551 -85.6598 0.93795
7.042 0.98812 5.4765e-005 3.8183 0.011944 9.1763e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4567 0.51524 0.15754 0.018725 13.3749 0.11635 0.00015017 0.7738 0.0088694 0.0098344 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16074 0.9523 0.92216 0.0013961 0.99526 0.53237 0.001881 0.42902 2.1411 2.1406 16.0036 144.9451 0.00015504 -85.6598 0.93895
7.043 0.98812 5.4765e-005 3.8183 0.011944 9.1776e-005 0.0011677 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4568 0.51528 0.15755 0.018726 13.3775 0.11636 0.00015018 0.77379 0.0088698 0.0098349 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.16074 0.9524 0.9222 0.0013961 0.99527 0.53253 0.001881 0.42903 2.1414 2.1409 16.0036 144.9451 0.00015498 -85.6598 0.93995
7.044 0.98812 5.4765e-005 3.8183 0.011944 9.1789e-005 0.0011678 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4569 0.51533 0.15756 0.018727 13.3801 0.11636 0.00015019 0.77379 0.0088703 0.0098353 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.16075 0.9525 0.92224 0.0013961 0.99529 0.5327 0.0018809 0.42905 2.1417 2.1413 16.0036 144.9451 0.00015493 -85.6599 0.94095
7.045 0.98812 5.4765e-005 3.8183 0.011944 9.1802e-005 0.0011678 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.457 0.51537 0.15758 0.018729 13.3828 0.11637 0.0001502 0.77378 0.0088708 0.0098358 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.16075 0.9526 0.92227 0.0013961 0.9953 0.53286 0.0018809 0.42906 2.1421 2.1416 16.0035 144.9451 0.00015487 -85.6599 0.94195
7.046 0.98812 5.4765e-005 3.8183 0.011944 9.1814e-005 0.0011678 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.4571 0.51542 0.15759 0.01873 13.3854 0.11638 0.00015021 0.77377 0.0088712 0.0098363 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16075 0.95269 0.92231 0.0013961 0.99531 0.53302 0.0018809 0.42907 2.1424 2.142 16.0035 144.9452 0.00015481 -85.6599 0.94295
7.047 0.98812 5.4765e-005 3.8183 0.011944 9.1827e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4572 0.51546 0.15761 0.018731 13.388 0.11639 0.00015022 0.77376 0.0088717 0.0098368 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16076 0.95279 0.92234 0.0013961 0.99532 0.53319 0.0018809 0.42908 2.1428 2.1423 16.0035 144.9452 0.00015476 -85.66 0.94395
7.048 0.98812 5.4765e-005 3.8183 0.011944 9.184e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4573 0.51551 0.15762 0.018732 13.3906 0.11639 0.00015023 0.77376 0.0088721 0.0098373 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16076 0.95289 0.92238 0.0013961 0.99534 0.53335 0.0018809 0.4291 2.1431 2.1426 16.0034 144.9452 0.0001547 -85.66 0.94495
7.049 0.98812 5.4764e-005 3.8183 0.011944 9.1853e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4574 0.51555 0.15764 0.018733 13.3932 0.1164 0.00015024 0.77375 0.0088726 0.0098378 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16076 0.95298 0.92242 0.0013961 0.99535 0.53351 0.0018809 0.42911 2.1434 2.143 16.0034 144.9452 0.00015464 -85.66 0.94595
7.05 0.98812 5.4764e-005 3.8183 0.011944 9.1866e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4575 0.5156 0.15765 0.018735 13.3958 0.11641 0.00015026 0.77374 0.008873 0.0098383 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16077 0.95308 0.92245 0.0013961 0.99536 0.53367 0.0018809 0.42912 2.1438 2.1433 16.0034 144.9452 0.00015459 -85.66 0.94695
7.051 0.98812 5.4764e-005 3.8183 0.011944 9.1879e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4575 0.51565 0.15766 0.018736 13.3985 0.11642 0.00015027 0.77373 0.0088735 0.0098388 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16077 0.95317 0.92249 0.0013961 0.99537 0.53384 0.0018809 0.42913 2.1441 2.1437 16.0033 144.9453 0.00015453 -85.6601 0.94795
7.052 0.98812 5.4764e-005 3.8183 0.011944 9.1892e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4576 0.51569 0.15768 0.018737 13.4011 0.11642 0.00015028 0.77373 0.0088739 0.0098392 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16077 0.95327 0.92252 0.0013961 0.99538 0.534 0.0018809 0.42915 2.1445 2.144 16.0033 144.9453 0.00015448 -85.6601 0.94895
7.053 0.98812 5.4764e-005 3.8183 0.011944 9.1904e-005 0.0011678 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4577 0.51574 0.15769 0.018738 13.4037 0.11643 0.00015029 0.77372 0.0088744 0.0098397 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16078 0.95336 0.92256 0.0013961 0.99539 0.53416 0.0018809 0.42916 2.1448 2.1443 16.0033 144.9453 0.00015442 -85.6601 0.94995
7.054 0.98812 5.4764e-005 3.8183 0.011944 9.1917e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4578 0.51578 0.15771 0.01874 13.4063 0.11644 0.0001503 0.77371 0.0088749 0.0098402 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16078 0.95346 0.92259 0.0013961 0.99541 0.53432 0.0018809 0.42917 2.1451 2.1447 16.0032 144.9453 0.00015437 -85.6602 0.95095
7.055 0.98812 5.4764e-005 3.8183 0.011944 9.193e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4579 0.51583 0.15772 0.018741 13.4089 0.11645 0.00015031 0.7737 0.0088753 0.0098407 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16078 0.95355 0.92263 0.0013961 0.99542 0.53448 0.0018809 0.42918 2.1455 2.145 16.0032 144.9453 0.00015431 -85.6602 0.95195
7.056 0.98812 5.4764e-005 3.8183 0.011944 9.1943e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.458 0.51587 0.15774 0.018742 13.4116 0.11645 0.00015032 0.7737 0.0088758 0.0098412 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16079 0.95364 0.92266 0.0013961 0.99543 0.53465 0.0018809 0.4292 2.1458 2.1453 16.0032 144.9454 0.00015426 -85.6602 0.95295
7.057 0.98812 5.4764e-005 3.8183 0.011944 9.1956e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4581 0.51592 0.15775 0.018743 13.4142 0.11646 0.00015033 0.77369 0.0088762 0.0098417 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16079 0.95374 0.9227 0.0013961 0.99544 0.53481 0.0018809 0.42921 2.1461 2.1457 16.0031 144.9454 0.0001542 -85.6603 0.95395
7.058 0.98812 5.4764e-005 3.8183 0.011944 9.1969e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4582 0.51596 0.15776 0.018745 13.4168 0.11647 0.00015034 0.77368 0.0088767 0.0098422 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.1608 0.95383 0.92273 0.0013961 0.99545 0.53497 0.0018809 0.42922 2.1465 2.146 16.0031 144.9454 0.00015415 -85.6603 0.95495
7.059 0.98812 5.4764e-005 3.8183 0.011944 9.1982e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4583 0.51601 0.15778 0.018746 13.4194 0.11648 0.00015036 0.77367 0.0088771 0.0098427 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.1608 0.95392 0.92277 0.0013961 0.99546 0.53513 0.0018809 0.42923 2.1468 2.1463 16.0031 144.9454 0.0001541 -85.6603 0.95595
7.06 0.98812 5.4764e-005 3.8183 0.011944 9.1995e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4584 0.51606 0.15779 0.018747 13.4221 0.11648 0.00015037 0.77367 0.0088776 0.0098432 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.1608 0.95402 0.9228 0.001396 0.99547 0.5353 0.0018809 0.42925 2.1471 2.1467 16.003 144.9454 0.00015404 -85.6603 0.95695
7.061 0.98812 5.4764e-005 3.8183 0.011944 9.2007e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4584 0.5161 0.15781 0.018748 13.4247 0.11649 0.00015038 0.77366 0.008878 0.0098436 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16081 0.95411 0.92284 0.001396 0.99549 0.53546 0.0018809 0.42926 2.1475 2.147 16.003 144.9455 0.00015399 -85.6604 0.95795
7.062 0.98812 5.4763e-005 3.8183 0.011944 9.202e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4585 0.51615 0.15782 0.018749 13.4273 0.1165 0.00015039 0.77365 0.0088785 0.0098441 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16081 0.9542 0.92287 0.001396 0.9955 0.53562 0.0018809 0.42927 2.1478 2.1473 16.003 144.9455 0.00015393 -85.6604 0.95895
7.063 0.98812 5.4763e-005 3.8183 0.011944 9.2033e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4586 0.51619 0.15784 0.018751 13.4299 0.11651 0.0001504 0.77364 0.008879 0.0098446 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16081 0.95429 0.92291 0.001396 0.99551 0.53578 0.0018809 0.42928 2.1481 2.1477 16.0029 144.9455 0.00015388 -85.6604 0.95995
7.064 0.98812 5.4763e-005 3.8183 0.011944 9.2046e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4587 0.51624 0.15785 0.018752 13.4326 0.11651 0.00015041 0.77364 0.0088794 0.0098451 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16082 0.95438 0.92294 0.001396 0.99552 0.53594 0.0018809 0.4293 2.1485 2.148 16.0029 144.9455 0.00015383 -85.6604 0.96095
7.065 0.98812 5.4763e-005 3.8183 0.011944 9.2059e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4588 0.51628 0.15786 0.018753 13.4352 0.11652 0.00015042 0.77363 0.0088799 0.0098456 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16082 0.95447 0.92297 0.001396 0.99553 0.5361 0.0018808 0.42931 2.1488 2.1483 16.0029 144.9455 0.00015377 -85.6605 0.96195
7.066 0.98812 5.4763e-005 3.8183 0.011944 9.2072e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4589 0.51633 0.15788 0.018754 13.4378 0.11653 0.00015043 0.77362 0.0088803 0.0098461 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16082 0.95457 0.92301 0.001396 0.99554 0.53627 0.0018808 0.42932 2.1491 2.1487 16.0028 144.9456 0.00015372 -85.6605 0.96295
7.067 0.98812 5.4763e-005 3.8183 0.011944 9.2085e-005 0.0011678 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.459 0.51637 0.15789 0.018756 13.4404 0.11654 0.00015044 0.77361 0.0088808 0.0098466 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16083 0.95466 0.92304 0.001396 0.99555 0.53643 0.0018808 0.42933 2.1495 2.149 16.0028 144.9456 0.00015367 -85.6605 0.96395
7.068 0.98812 5.4763e-005 3.8183 0.011944 9.2097e-005 0.0011679 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4591 0.51642 0.15791 0.018757 13.4431 0.11654 0.00015045 0.77361 0.0088812 0.0098471 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16083 0.95475 0.92308 0.001396 0.99556 0.53659 0.0018808 0.42935 2.1498 2.1493 16.0028 144.9456 0.00015362 -85.6606 0.96495
7.069 0.98812 5.4763e-005 3.8183 0.011944 9.211e-005 0.0011679 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4592 0.51647 0.15792 0.018758 13.4457 0.11655 0.00015047 0.7736 0.0088817 0.0098475 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16083 0.95484 0.92311 0.001396 0.99557 0.53675 0.0018808 0.42936 2.1501 2.1497 16.0027 144.9456 0.00015356 -85.6606 0.96595
7.07 0.98812 5.4763e-005 3.8183 0.011944 9.2123e-005 0.0011679 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4592 0.51651 0.15794 0.018759 13.4483 0.11656 0.00015048 0.77359 0.0088821 0.009848 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16084 0.95493 0.92314 0.001396 0.99558 0.53691 0.0018808 0.42937 2.1504 2.15 16.0027 144.9456 0.00015351 -85.6606 0.96695
7.071 0.98812 5.4763e-005 3.8183 0.011944 9.2136e-005 0.0011679 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4593 0.51656 0.15795 0.01876 13.4509 0.11657 0.00015049 0.77359 0.0088826 0.0098485 0.0013843 0.98697 0.99172 2.9846e-006 1.1938e-005 0.16084 0.95501 0.92318 0.001396 0.99559 0.53707 0.0018808 0.42938 2.1508 2.1503 16.0027 144.9457 0.00015346 -85.6606 0.96795
7.072 0.98812 5.4763e-005 3.8183 0.011944 9.2149e-005 0.0011679 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.4594 0.5166 0.15796 0.018762 13.4536 0.11657 0.0001505 0.77358 0.0088831 0.009849 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16084 0.9551 0.92321 0.001396 0.9956 0.53723 0.0018808 0.4294 2.1511 2.1506 16.0026 144.9457 0.00015341 -85.6607 0.96895
7.073 0.98812 5.4763e-005 3.8183 0.011944 9.2162e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4595 0.51665 0.15798 0.018763 13.4562 0.11658 0.00015051 0.77357 0.0088835 0.0098495 0.0013843 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16085 0.95519 0.92324 0.001396 0.99561 0.5374 0.0018808 0.42941 2.1514 2.151 16.0026 144.9457 0.00015336 -85.6607 0.96995
7.074 0.98812 5.4763e-005 3.8183 0.011944 9.2175e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4596 0.51669 0.15799 0.018764 13.4588 0.11659 0.00015052 0.77356 0.008884 0.00985 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16085 0.95528 0.92328 0.001396 0.99562 0.53756 0.0018808 0.42942 2.1517 2.1513 16.0026 144.9457 0.00015331 -85.6607 0.97095
7.075 0.98812 5.4762e-005 3.8183 0.011944 9.2188e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4597 0.51674 0.15801 0.018765 13.4614 0.11659 0.00015053 0.77356 0.0088844 0.0098505 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16086 0.95537 0.92331 0.001396 0.99563 0.53772 0.0018808 0.42943 2.1521 2.1516 16.0025 144.9457 0.00015325 -85.6607 0.97195
7.076 0.98812 5.4762e-005 3.8183 0.011944 9.22e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4598 0.51679 0.15802 0.018767 13.4641 0.1166 0.00015054 0.77355 0.0088849 0.0098509 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16086 0.95546 0.92334 0.001396 0.99564 0.53788 0.0018808 0.42945 2.1524 2.152 16.0025 144.9458 0.0001532 -85.6608 0.97295
7.077 0.98812 5.4762e-005 3.8183 0.011944 9.2213e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4599 0.51683 0.15804 0.018768 13.4667 0.11661 0.00015055 0.77354 0.0088853 0.0098514 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16086 0.95555 0.92337 0.001396 0.99565 0.53804 0.0018808 0.42946 2.1527 2.1523 16.0025 144.9458 0.00015315 -85.6608 0.97395
7.078 0.98812 5.4762e-005 3.8183 0.011944 9.2226e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.46 0.51688 0.15805 0.018769 13.4693 0.11662 0.00015056 0.77353 0.0088858 0.0098519 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16087 0.95563 0.92341 0.001396 0.99566 0.5382 0.0018808 0.42947 2.153 2.1526 16.0024 144.9458 0.0001531 -85.6608 0.97495
7.079 0.98812 5.4762e-005 3.8183 0.011944 9.2239e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4601 0.51692 0.15806 0.01877 13.472 0.11662 0.00015058 0.77353 0.0088862 0.0098524 0.0013842 0.98697 0.99172 2.9845e-006 1.1938e-005 0.16087 0.95572 0.92344 0.001396 0.99567 0.53836 0.0018808 0.42948 2.1534 2.1529 16.0024 144.9458 0.00015305 -85.6608 0.97595
7.08 0.98812 5.4762e-005 3.8183 0.011944 9.2252e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4601 0.51697 0.15808 0.018772 13.4746 0.11663 0.00015059 0.77352 0.0088867 0.0098529 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.16087 0.95581 0.92347 0.001396 0.99568 0.53852 0.0018808 0.4295 2.1537 2.1533 16.0024 144.9459 0.000153 -85.6609 0.97695
7.081 0.98812 5.4762e-005 3.8183 0.011944 9.2265e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4602 0.51701 0.15809 0.018773 13.4772 0.11664 0.0001506 0.77351 0.0088871 0.0098534 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.16088 0.95589 0.9235 0.001396 0.99569 0.53868 0.0018808 0.42951 2.154 2.1536 16.0023 144.9459 0.00015295 -85.6609 0.97795
7.082 0.98812 5.4762e-005 3.8183 0.011944 9.2278e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.4603 0.51706 0.15811 0.018774 13.4799 0.11665 0.00015061 0.7735 0.0088876 0.0098539 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.16088 0.95598 0.92354 0.001396 0.9957 0.53884 0.0018808 0.42952 2.1543 2.1539 16.0023 144.9459 0.0001529 -85.6609 0.97895
7.083 0.98812 5.4762e-005 3.8183 0.011944 9.2291e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032261 0.0389 0 1.4604 0.5171 0.15812 0.018775 13.4825 0.11665 0.00015062 0.7735 0.0088881 0.0098543 0.0013842 0.98697 0.99172 2.9844e-006 1.1938e-005 0.16088 0.95607 0.92357 0.001396 0.99571 0.539 0.0018808 0.42953 2.1547 2.1542 16.0023 144.9459 0.00015285 -85.6609 0.97995
7.084 0.98812 5.4762e-005 3.8183 0.011944 9.2303e-005 0.0011679 0.23365 0.00065931 0.23431 0.21621 0 0.032261 0.0389 0 1.4605 0.51715 0.15813 0.018776 13.4851 0.11666 0.00015063 0.77349 0.0088885 0.0098548 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.16089 0.95615 0.9236 0.001396 0.99572 0.53916 0.0018808 0.42954 2.155 2.1545 16.0022 144.9459 0.0001528 -85.6609 0.98095
7.085 0.98812 5.4762e-005 3.8183 0.011944 9.2316e-005 0.0011679 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4606 0.5172 0.15815 0.018778 13.4878 0.11667 0.00015064 0.77348 0.008889 0.0098553 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.16089 0.95624 0.92363 0.001396 0.99573 0.53933 0.0018808 0.42956 2.1553 2.1549 16.0022 144.946 0.00015275 -85.661 0.98195
7.086 0.98812 5.4762e-005 3.8183 0.011944 9.2329e-005 0.0011679 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4607 0.51724 0.15816 0.018779 13.4904 0.11668 0.00015065 0.77347 0.0088894 0.0098558 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.16089 0.95632 0.92366 0.001396 0.99574 0.53949 0.0018808 0.42957 2.1556 2.1552 16.0022 144.946 0.0001527 -85.661 0.98295
7.087 0.98812 5.4761e-005 3.8183 0.011944 9.2342e-005 0.0011679 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4608 0.51729 0.15818 0.01878 13.493 0.11668 0.00015066 0.77347 0.0088899 0.0098563 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.1609 0.95641 0.9237 0.0013959 0.99575 0.53965 0.0018808 0.42958 2.1559 2.1555 16.0021 144.946 0.00015265 -85.661 0.98395
7.088 0.98812 5.4761e-005 3.8183 0.011944 9.2355e-005 0.0011679 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4609 0.51733 0.15819 0.018781 13.4956 0.11669 0.00015067 0.77346 0.0088903 0.0098568 0.0013842 0.98697 0.99172 2.9844e-006 1.1937e-005 0.1609 0.95649 0.92373 0.0013959 0.99576 0.53981 0.0018808 0.42959 2.1563 2.1558 16.0021 144.946 0.0001526 -85.661 0.98495
7.089 0.98812 5.4761e-005 3.8183 0.011944 9.2368e-005 0.0011679 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4609 0.51738 0.15821 0.018783 13.4983 0.1167 0.00015068 0.77345 0.0088908 0.0098573 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.1609 0.95658 0.92376 0.0013959 0.99577 0.53997 0.0018808 0.42961 2.1566 2.1561 16.0021 144.946 0.00015255 -85.6611 0.98595
7.09 0.98812 5.4761e-005 3.8183 0.011944 9.2381e-005 0.0011679 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.461 0.51742 0.15822 0.018784 13.5009 0.11671 0.0001507 0.77345 0.0088912 0.0098577 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16091 0.95666 0.92379 0.0013959 0.99578 0.54013 0.0018808 0.42962 2.1569 2.1565 16.002 144.9461 0.0001525 -85.6611 0.98695
7.091 0.98812 5.4761e-005 3.8183 0.011944 9.2393e-005 0.0011679 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4611 0.51747 0.15823 0.018785 13.5035 0.11671 0.00015071 0.77344 0.0088917 0.0098582 0.0013842 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16091 0.95675 0.92382 0.0013959 0.99578 0.54029 0.0018807 0.42963 2.1572 2.1568 16.002 144.9461 0.00015246 -85.6611 0.98795
7.092 0.98812 5.4761e-005 3.8183 0.011944 9.2406e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4612 0.51751 0.15825 0.018786 13.5062 0.11672 0.00015072 0.77343 0.0088921 0.0098587 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16092 0.95683 0.92385 0.0013959 0.99579 0.54045 0.0018807 0.42964 2.1575 2.1571 16.002 144.9461 0.00015241 -85.6611 0.98895
7.093 0.98812 5.4761e-005 3.8183 0.011944 9.2419e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4613 0.51756 0.15826 0.018787 13.5088 0.11673 0.00015073 0.77342 0.0088926 0.0098592 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16092 0.95691 0.92388 0.0013959 0.9958 0.54061 0.0018807 0.42966 2.1578 2.1574 16.0019 144.9461 0.00015236 -85.6611 0.98995
7.094 0.98812 5.4761e-005 3.8183 0.011944 9.2432e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4614 0.51761 0.15828 0.018789 13.5115 0.11674 0.00015074 0.77342 0.008893 0.0098597 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16092 0.957 0.92391 0.0013959 0.99581 0.54077 0.0018807 0.42967 2.1582 2.1577 16.0019 144.9461 0.00015231 -85.6612 0.99095
7.095 0.98812 5.4761e-005 3.8183 0.011944 9.2445e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4615 0.51765 0.15829 0.01879 13.5141 0.11674 0.00015075 0.77341 0.0088935 0.0098602 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16093 0.95708 0.92394 0.0013959 0.99582 0.54093 0.0018807 0.42968 2.1585 2.158 16.0019 144.9462 0.00015226 -85.6612 0.99195
7.096 0.98812 5.4761e-005 3.8183 0.011944 9.2458e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4616 0.5177 0.15831 0.018791 13.5167 0.11675 0.00015076 0.7734 0.0088939 0.0098607 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16093 0.95716 0.92397 0.0013959 0.99583 0.54109 0.0018807 0.42969 2.1588 2.1584 16.0018 144.9462 0.00015222 -85.6612 0.99295
7.097 0.98812 5.4761e-005 3.8183 0.011944 9.2471e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4617 0.51774 0.15832 0.018792 13.5194 0.11676 0.00015077 0.77339 0.0088944 0.0098611 0.0013841 0.98697 0.99172 2.9843e-006 1.1937e-005 0.16093 0.95724 0.92401 0.0013959 0.99584 0.54125 0.0018807 0.42971 2.1591 2.1587 16.0018 144.9462 0.00015217 -85.6612 0.99395
7.098 0.98812 5.4761e-005 3.8183 0.011944 9.2484e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4618 0.51779 0.15833 0.018794 13.522 0.11676 0.00015078 0.77339 0.0088949 0.0098616 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.16094 0.95733 0.92404 0.0013959 0.99585 0.54141 0.0018807 0.42972 2.1594 2.159 16.0018 144.9462 0.00015212 -85.6612 0.99495
7.099 0.98812 5.4761e-005 3.8183 0.011944 9.2496e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4618 0.51783 0.15835 0.018795 13.5246 0.11677 0.00015079 0.77338 0.0088953 0.0098621 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.16094 0.95741 0.92407 0.0013959 0.99586 0.54157 0.0018807 0.42973 2.1597 2.1593 16.0017 144.9462 0.00015207 -85.6613 0.99595
7.1 0.98812 5.476e-005 3.8183 0.011944 9.2509e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4619 0.51788 0.15836 0.018796 13.5273 0.11678 0.00015081 0.77337 0.0088958 0.0098626 0.0013841 0.98697 0.99172 2.9842e-006 1.1937e-005 0.16094 0.95749 0.9241 0.0013959 0.99586 0.54173 0.0018807 0.42974 2.16 2.1596 16.0017 144.9463 0.00015203 -85.659 0.99695
7.101 0.98812 5.476e-005 3.8183 0.011943 9.2522e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.462 0.51792 0.15838 0.018797 13.5299 0.11679 0.00015082 0.77336 0.0088962 0.0098631 0.0064782 0.98322 0.99099 1.453e-005 5.3377e-005 0.16095 0.95752 0.92413 0.0027742 0.99586 0.54187 0.0023961 0.4297 2.1604 2.1599 16.0016 144.9463 0.00015199 -76.1558 0.99795
7.102 0.98812 5.476e-005 3.8183 0.011943 9.2535e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4621 0.51797 0.15839 0.018798 13.5325 0.11679 0.00015083 0.77336 0.0088967 0.0098636 0.02624 0.9717 0.98766 6.6031e-005 0.00022967 0.16095 0.95733 0.92416 0.0053024 0.99581 0.54198 0.0033369 0.42958 2.1607 2.1602 16.0016 144.9462 0.00015197 -67.142 0.99895
7.103 0.98812 5.476e-005 3.8183 0.011943 9.2548e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4622 0.51802 0.15841 0.0188 13.5352 0.1168 0.00015084 0.77335 0.0088971 0.009864 0.094939 0.9472 0.97731 0.00028463 0.00091381 0.16095 0.95659 0.92419 0.0092501 0.99554 0.54209 0.0044257 0.42942 2.161 2.1606 16.0015 144.9462 0.00015198 -58.01 0.99995
7.104 0.98812 5.476e-005 3.8183 0.011943 9.2561e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4623 0.51806 0.15842 0.018801 13.5378 0.11681 0.00015085 0.77334 0.0088976 0.0098645 0.48883 0.85604 0.93867 0.0021849 0.0054876 0.16096 0.95459 0.92421 0.015759 0.99143 0.54213 0.0056248 0.42923 2.1613 2.1609 16.0022 144.9462 0.00015201 -37.1731 0.15522
7.105 0.98812 5.476e-005 3.8183 0.011943 9.2574e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4624 0.51811 0.15843 0.018802 13.5405 0.11682 0.00015086 0.77333 0.008898 0.009865 0.99963 0.0021564 0.71199 0.94299 0.99658 0.16096 0.92126 0.92115 0.33565 0.96401 0.53022 0.044504 0.42903 2.1064 0.96705 16.0061 144.9459 0.00024677 25.0917 0.001946
7.106 0.98812 5.476e-005 3.8183 0.011943 9.2586e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4625 0.51815 0.15845 0.018803 13.5431 0.11682 0.00015087 0.77333 0.0088985 0.0098655 0.99952 1.303e-006 0.52805 0.99822 0.99959 0.16096 0.88135 0.90277 0.6266 0.93686 0.51537 0.10056 0.42882 1.8972 0.61415 16.0057 144.9445 0.00036344 21.9716 0.002946
7.107 0.98812 5.476e-005 3.8183 0.011943 9.2599e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4626 0.5182 0.15846 0.018805 13.5457 0.11683 0.00015088 0.77332 0.0088989 0.009866 0.99919 9.9959e-010 0.39188 0.99661 0.99905 0.16097 0.84355 0.87894 0.75413 0.91047 0.50107 0.1444 0.42862 1.7017 0.59819 16.0054 144.9427 0.00043947 17.0368 0.003946
7.108 0.98812 5.476e-005 3.8183 0.011943 9.2612e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4626 0.51824 0.15848 0.018806 13.5484 0.11684 0.00015089 0.77331 0.0088994 0.0098665 0.99883 -9.4567e-011 0.29108 0.99378 0.99825 0.16097 0.80818 0.85219 0.81009 0.88483 0.48742 0.17904 0.42841 1.5397 0.64497 16.005 144.9408 0.00049744 13.6041 0.004946
7.109 0.98812 5.476e-005 3.8183 0.011943 9.2625e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4627 0.51829 0.15849 0.018807 13.551 0.11685 0.0001509 0.7733 0.0088998 0.0098669 0.9985 -3.1386e-011 0.2164 0.99052 0.99736 0.16098 0.77522 0.82378 0.83468 0.85991 0.47442 0.2081 0.42821 1.4115 0.71157 16.0047 144.939 0.00054263 11.3342 0.005946
7.11 0.98812 5.476e-005 3.8183 0.011943 9.2638e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4628 0.51833 0.1585 0.018808 13.5537 0.11685 0.00015092 0.7733 0.0089003 0.0098674 0.99819 -1.82e-010 0.16099 0.98706 0.99641 0.16098 0.74443 0.7946 0.84385 0.8357 0.46204 0.23344 0.428 1.3135 0.78223 16.0044 144.9372 0.00057763 9.6459 0.006946
7.111 0.98812 5.476e-005 3.8183 0.011943 9.2651e-005 0.001168 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.4629 0.51838 0.15852 0.018809 13.5563 0.11686 0.00015093 0.77329 0.0089007 0.0098679 0.99789 -4.5978e-012 0.11986 0.98336 0.99539 0.16098 0.7156 0.7653 0.84462 0.81217 0.45025 0.25596 0.4278 1.2411 0.84866 16.0041 144.9354 0.00060453 8.2345 0.007946
7.112 0.98812 5.4759e-005 3.8183 0.011943 9.2664e-005 0.001168 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.463 0.51843 0.15853 0.018811 13.5589 0.11687 0.00015094 0.77328 0.0089012 0.0098684 0.99758 -2.9407e-011 0.089291 0.97929 0.99425 0.16099 0.6886 0.73638 0.84041 0.78931 0.43903 0.27614 0.4276 1.1892 0.90635 16.0037 144.9338 0.00062523 6.9576 0.008946
7.113 0.98812 5.4759e-005 3.8183 0.011943 9.2677e-005 0.001168 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4631 0.51847 0.15855 0.018812 13.5616 0.11688 0.00015095 0.77328 0.0089016 0.0098689 0.99724 2.6419e-011 0.06657 0.9747 0.99294 0.16099 0.66331 0.70817 0.83301 0.76709 0.42839 0.2943 0.42739 1.1533 0.95353 16.0034 144.9322 0.00064135 5.7448 0.009946
7.114 0.98812 5.4759e-005 3.8183 0.011943 9.2689e-005 0.001168 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4632 0.51852 0.15856 0.018813 13.5642 0.11688 0.00015096 0.77327 0.0089021 0.0098694 0.99686 -5.9348e-011 0.049669 0.96942 0.99138 0.16099 0.63966 0.68092 0.82338 0.7455 0.41832 0.31063 0.42719 1.1292 0.99037 16.0032 144.9307 0.00065415 4.5576 0.010946
7.115 0.98812 5.4759e-005 3.8183 0.011943 9.2702e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4633 0.51856 0.15858 0.018814 13.5669 0.11689 0.00015097 0.77326 0.0089025 0.0098698 0.99642 2.9388e-011 0.037092 0.96324 0.98954 0.161 0.61756 0.65479 0.81206 0.72453 0.40883 0.32531 0.42699 1.1137 1.0182 16.0029 144.9293 0.00066459 3.3716 0.011946
7.116 0.98812 5.4759e-005 3.8183 0.011943 9.2715e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4634 0.51861 0.15859 0.018816 13.5695 0.1169 0.00015098 0.77325 0.008903 0.0098703 0.99592 1.1102e-011 0.027727 0.95594 0.98727 0.161 0.59696 0.62991 0.79931 0.70414 0.39992 0.33844 0.42678 1.1042 1.0387 16.0026 144.9279 0.00067334 2.1682 0.012946
7.117 0.98812 5.4759e-005 3.8183 0.011943 9.2728e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4634 0.51865 0.1586 0.018817 13.5721 0.1169 0.00015099 0.77325 0.0089034 0.0098708 0.99532 4.1032e-012 0.020749 0.94724 0.98453 0.161 0.57782 0.60637 0.78525 0.68434 0.39162 0.35013 0.42658 1.0988 1.0537 16.0023 144.9267 0.00068084 0.93075 0.013946
7.118 0.98812 5.4759e-005 3.8183 0.011943 9.2741e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4635 0.5187 0.15862 0.018818 13.5748 0.11691 0.000151 0.77324 0.0089039 0.0098713 0.99461 1.217e-011 0.015548 0.93678 0.98111 0.16101 0.56009 0.58425 0.76989 0.6651 0.38394 0.36046 0.42638 1.0962 1.0647 16.0021 144.9255 0.00068738 -0.35902 0.014946
7.119 0.98812 5.4759e-005 3.8183 0.011943 9.2754e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4636 0.51874 0.15863 0.018819 13.5774 0.11692 0.00015101 0.77323 0.0089043 0.0098718 0.99374 -1.2773e-011 0.011669 0.92408 0.97681 0.16101 0.54375 0.56362 0.75316 0.64641 0.37689 0.36947 0.42618 1.0955 1.0729 16.0018 144.9243 0.00069315 -1.7234 0.015946
7.12 0.98812 5.4759e-005 3.8183 0.011943 9.2767e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4637 0.51879 0.15865 0.01882 13.5801 0.11693 0.00015102 0.77322 0.0089048 0.0098723 0.99263 4.3039e-012 0.0087737 0.9085 0.97131 0.16101 0.52879 0.54456 0.73491 0.62826 0.37051 0.37721 0.42597 1.096 1.0792 16.0015 144.9233 0.00069823 -3.1914 0.016946
7.121 0.98812 5.4759e-005 3.8183 0.011943 9.2779e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4638 0.51884 0.15866 0.018822 13.5827 0.11693 0.00015104 0.77322 0.0089053 0.0098727 0.99119 -4.2501e-012 0.0066123 0.88914 0.96414 0.16102 0.5152 0.52716 0.71492 0.61064 0.36482 0.3837 0.42577 1.0973 1.0842 16.0013 144.9223 0.00070269 -4.8031 0.017946
7.122 0.98812 5.4759e-005 3.8183 0.011943 9.2792e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4639 0.51888 0.15868 0.018823 13.5854 0.11694 0.00015105 0.77321 0.0089057 0.0098732 0.98923 3.7345e-012 0.0049983 0.86469 0.95456 0.16102 0.50301 0.51154 0.6929 0.59353 0.35985 0.38896 0.42557 1.099 1.0884 16.0011 144.9214 0.00070653 -6.6149 0.018946
7.123 0.98812 5.4759e-005 3.8183 0.011943 9.2805e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.464 0.51893 0.15869 0.018824 13.588 0.11695 0.00015106 0.7732 0.0089062 0.0098737 0.98641 -2.9138e-012 0.0037934 0.8333 0.94142 0.16102 0.49225 0.49782 0.66845 0.57693 0.35565 0.39296 0.42536 1.1011 1.092 16.0008 144.9206 0.00070972 -8.7069 0.019946
7.124 0.98812 5.4759e-005 3.8183 0.011943 9.2818e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4641 0.51897 0.1587 0.018825 13.5907 0.11696 0.00015107 0.77319 0.0089066 0.0098742 0.98208 3.6575e-012 0.0028951 0.79219 0.92285 0.16103 0.48298 0.48616 0.64111 0.56084 0.35223 0.39568 0.42516 1.1034 1.0953 16.0006 144.9199 0.00071221 -11.1923 0.020946
7.125 0.98812 5.4758e-005 3.8183 0.011943 9.2831e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4642 0.51902 0.15872 0.018827 13.5933 0.11696 0.00015108 0.77319 0.0089071 0.0098747 0.97488 -5.1259e-012 0.0022277 0.73734 0.89578 0.16103 0.47526 0.47672 0.61045 0.54529 0.34961 0.39711 0.42496 1.1058 1.0983 16.0004 144.9192 0.00071391 -14.2226 0.021946
7.126 0.98812 5.4758e-005 3.8183 0.011943 9.2844e-005 0.0011681 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.4643 0.51906 0.15873 0.018828 13.5959 0.11697 0.00015109 0.77318 0.0089075 0.0098752 0.96183 1.9632e-012 0.0017362 0.66318 0.85522 0.16103 0.46911 0.46962 0.57619 0.53033 0.34774 0.39726 0.42476 1.1084 1.1012 16.0002 144.9186 0.0007147 -17.9733 0.022946
7.127 0.98812 5.4758e-005 3.8183 0.011943 9.2857e-005 0.0011681 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4643 0.51911 0.15875 0.018829 13.5986 0.11698 0.0001511 0.77317 0.008908 0.0098756 0.93636 1.0261e-012 0.0013805 0.56323 0.79357 0.16104 0.46447 0.46485 0.53839 0.51613 0.34654 0.3962 0.42456 1.1109 1.104 16.0001 144.9181 0.00071449 -22.5637 0.023946
7.128 0.98812 5.4758e-005 3.8183 0.011943 9.287e-005 0.0011681 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4644 0.51915 0.15876 0.01883 13.6012 0.11699 0.00015111 0.77317 0.0089084 0.0098761 0.88577 -6.248e-012 0.0011313 0.43425 0.70133 0.16104 0.4611 0.46207 0.49724 0.50308 0.34585 0.39406 0.42436 1.1135 1.1068 15.9999 144.9177 0.00071333 -27.8697 0.024946
7.129 0.98812 5.4758e-005 3.8183 0.011943 9.2882e-005 0.0011681 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4645 0.5192 0.15877 0.018831 13.6039 0.11699 0.00015112 0.77316 0.0089089 0.0098766 0.79518 3.5006e-012 0.00096385 0.28675 0.57294 0.16105 0.45867 0.46065 0.45204 0.49208 0.3455 0.39093 0.42416 1.1161 1.1095 15.9998 144.9174 0.0007115 -33.3557 0.025946
7.13 0.98812 5.4758e-005 3.8183 0.011943 9.2895e-005 0.0011681 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4646 0.51925 0.15879 0.018833 13.6065 0.117 0.00015113 0.77315 0.0089093 0.0098771 0.6666 3.8278e-012 0.00085387 0.15215 0.41838 0.16105 0.45688 0.45996 0.40088 0.48446 0.34536 0.38662 0.42396 1.1188 1.1122 15.9997 144.9171 0.00070936 -38.3527 0.026946
7.131 0.98812 5.4758e-005 3.8183 0.011943 9.2908e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4647 0.51929 0.1588 0.018834 13.6092 0.11701 0.00015115 0.77314 0.0089098 0.0098776 0.52661 0.00027128 0.00086823 0.062152 0.26591 0.16105 0.45554 0.45994 0.34268 0.48094 0.34535 0.38077 0.42376 1.1214 1.1149 15.9996 144.9169 0.00070711 -42.5772 0.027946
7.132 0.98812 5.4758e-005 3.8183 0.011943 9.2921e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4648 0.51934 0.15882 0.018835 13.6118 0.11702 0.00015116 0.77314 0.0089102 0.0098781 0.40294 0.00090707 0.0011255 0.019761 0.14498 0.16106 0.45456 0.4609 0.27923 0.48063 0.34542 0.37301 0.42357 1.124 1.1176 15.9996 144.9167 0.00070482 -46.0677 0.028946
7.133 0.98812 5.4758e-005 3.8183 0.011943 9.2934e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4649 0.51938 0.15883 0.018836 13.6145 0.11702 0.00015117 0.77313 0.0089107 0.0098785 0.30764 0.0019177 0.0016429 0.0056418 0.068047 0.16106 0.45391 0.46296 0.21532 0.48197 0.34553 0.3631 0.42337 1.1267 1.1202 15.9995 144.9166 0.00070248 -48.9284 0.029946
7.134 0.98812 5.4758e-005 3.8183 0.011943 9.2947e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.465 0.51943 0.15885 0.018838 13.6171 0.11703 0.00015118 0.77312 0.0089111 0.009879 0.23914 0.0033978 0.0024429 0.0020392 0.028428 0.16106 0.45352 0.46583 0.15696 0.4839 0.34566 0.35097 0.42318 1.1293 1.1229 15.9995 144.9165 0.00070012 -51.2699 0.030946
7.135 0.98812 5.4758e-005 3.8183 0.011943 9.296e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4651 0.51947 0.15886 0.018839 13.6198 0.11704 0.00015119 0.77311 0.0089116 0.0098795 0.19067 0.0054176 0.0035353 0.0011234 0.011513 0.16107 0.45337 0.46913 0.10886 0.48594 0.34581 0.33675 0.423 1.1319 1.1255 15.9995 144.9164 0.00069774 -53.2054 0.031946
7.136 0.98812 5.4758e-005 3.8183 0.011943 9.2972e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4651 0.51952 0.15887 0.01884 13.6224 0.11704 0.0001512 0.77311 0.008912 0.00988 0.15571 0.0080304 0.0049226 0.00077922 0.005225 0.16107 0.45342 0.47258 0.072888 0.48792 0.34596 0.32069 0.42281 1.1345 1.1282 15.9995 144.9163 0.00069534 -54.8424 0.032946
7.137 0.98812 5.4757e-005 3.8183 0.011943 9.2985e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4652 0.51956 0.15889 0.018841 13.6251 0.11705 0.00015121 0.7731 0.0089125 0.0098805 0.12954 0.011284 0.0066069 0.0005875 0.0029769 0.16107 0.45364 0.47606 0.048254 0.48981 0.34612 0.30308 0.42263 1.1372 1.1308 15.9995 144.9163 0.00069292 -56.2717 0.033946
7.138 0.98812 5.4757e-005 3.8183 0.011943 9.2998e-005 0.0011681 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4653 0.51961 0.1589 0.018842 13.6277 0.11706 0.00015122 0.77309 0.0089129 0.0098809 0.10915 0.015236 0.0085941 0.00045977 0.0020651 0.16108 0.454 0.47952 0.032591 0.49159 0.34628 0.28421 0.42246 1.1398 1.1335 15.9995 144.9163 0.00069051 -57.5622 0.034946
7.139 0.98812 5.4757e-005 3.8183 0.011943 9.3011e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4654 0.51966 0.15892 0.018844 13.6304 0.11707 0.00015123 0.77308 0.0089134 0.0098814 0.092731 0.019955 0.010896 0.00036819 0.0015831 0.16108 0.4545 0.48296 0.023182 0.49326 0.34644 0.26437 0.42228 1.1424 1.1361 15.9995 144.9162 0.00068808 -58.7612 0.035946
7.14 0.98812 5.4757e-005 3.8183 0.011943 9.3024e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4655 0.5197 0.15893 0.018845 13.633 0.11707 0.00015124 0.77308 0.0089138 0.0098819 0.079189 0.02553 0.013532 0.00029901 0.0012635 0.16108 0.4551 0.48636 0.017693 0.49485 0.3466 0.24382 0.42211 1.145 1.1387 15.9996 144.9162 0.00068565 -59.8983 0.036946
7.141 0.98812 5.4757e-005 3.8183 0.011943 9.3037e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4656 0.51975 0.15894 0.018846 13.6357 0.11708 0.00015125 0.77307 0.0089143 0.0098824 0.067859 0.032065 0.016524 0.00024467 0.0010264 0.16109 0.45581 0.48973 0.014451 0.49636 0.34677 0.22283 0.42194 1.1477 1.1414 15.9996 144.9162 0.00068322 -60.9906 0.037946
7.142 0.98812 5.4757e-005 3.8183 0.011943 9.305e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4657 0.51979 0.15896 0.018847 13.6383 0.11709 0.00015127 0.77306 0.0089147 0.0098829 0.058304 0.03968 0.019899 0.00020218 0.00084229 0.16109 0.45661 0.49306 0.012411 0.4978 0.34693 0.20168 0.42177 1.1503 1.144 15.9996 144.9162 0.00068078 -62.0474 0.038946
7.143 0.98812 5.4757e-005 3.8183 0.011943 9.3063e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4658 0.51984 0.15897 0.018849 13.641 0.1171 0.00015128 0.77306 0.0089152 0.0098833 0.05021 0.048502 0.023686 0.00016787 0.00069632 0.16109 0.4575 0.49635 0.010989 0.49918 0.3471 0.18064 0.42161 1.1529 1.1467 15.9997 144.9161 0.00067834 -63.0737 0.039946
7.144 0.98812 5.4757e-005 3.8183 0.011943 9.3075e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4659 0.51988 0.15899 0.01885 13.6436 0.1171 0.00015129 0.77305 0.0089156 0.0098838 0.043338 0.058669 0.027918 0.00014023 0.00057927 0.1611 0.45846 0.49961 0.0098932 0.50051 0.34726 0.16002 0.42145 1.1555 1.1493 15.9997 144.9161 0.0006759 -64.0722 0.040946
7.145 0.98812 5.4757e-005 3.8183 0.011943 9.3088e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4659 0.51993 0.159 0.018851 13.6463 0.11711 0.0001513 0.77304 0.0089161 0.0098843 0.037492 0.070322 0.032628 0.00011771 0.00048463 0.1611 0.4595 0.50284 0.0089863 0.5018 0.34743 0.1401 0.4213 1.1581 1.1519 15.9998 144.9161 0.00067346 -65.0443 0.041946
7.146 0.98812 5.4757e-005 3.8183 0.011943 9.3101e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.466 0.51997 0.15902 0.018852 13.6489 0.11712 0.00015131 0.77303 0.0089165 0.0098848 0.032514 0.083604 0.037853 9.9292e-005 0.0004076 0.1611 0.46059 0.50603 0.0082061 0.50306 0.34759 0.12116 0.42115 1.1607 1.1545 15.9998 144.916 0.00067101 -65.9911 0.042946
7.147 0.98812 5.4757e-005 3.8183 0.011943 9.3114e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4661 0.52002 0.15903 0.018853 13.6516 0.11713 0.00015132 0.77303 0.008917 0.0098853 0.028267 0.098654 0.043633 8.4155e-005 0.00034455 0.16111 0.46174 0.50918 0.0075222 0.5043 0.34776 0.10344 0.421 1.1633 1.1572 15.9999 144.916 0.00066857 -66.913 0.043946
7.148 0.98812 5.4757e-005 3.8183 0.011943 9.3127e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4662 0.52007 0.15904 0.018855 13.6542 0.11713 0.00015133 0.77302 0.0089174 0.0098858 0.024641 0.1156 0.050012 7.1694e-005 0.0002927 0.16111 0.46294 0.5123 0.0069176 0.50552 0.34792 0.087144 0.42086 1.166 1.1598 15.9999 144.916 0.00066613 -67.8104 0.044946
7.149 0.98812 5.4757e-005 3.8183 0.011943 9.314e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4663 0.52011 0.15906 0.018856 13.6569 0.11714 0.00015134 0.77301 0.0089179 0.0098862 0.02154 0.13457 0.057036 6.128e-005 0.00024984 0.16111 0.46418 0.51539 0.00638 0.50673 0.34809 0.072432 0.42073 1.1686 1.1624 16 144.916 0.00066369 -68.6832 0.045946
7.15 0.98812 5.4756e-005 3.8183 0.011943 9.3153e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4664 0.52016 0.15907 0.018857 13.6595 0.11715 0.00015135 0.773 0.0089183 0.0098867 0.018886 0.15565 0.064757 5.2631e-005 0.00021428 0.16112 0.46545 0.51844 0.0059006 0.50793 0.34825 0.0594 0.42059 1.1712 1.165 16.0001 144.9159 0.00066125 -69.5314 0.046946
7.151 0.98812 5.4756e-005 3.8183 0.011943 9.3165e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4665 0.5202 0.15909 0.018858 13.6622 0.11715 0.00015136 0.773 0.0089188 0.0098872 0.016611 0.17892 0.07323 4.5451e-005 0.00018466 0.16112 0.46677 0.52145 0.005472 0.50914 0.34842 0.048085 0.42047 1.1738 1.1676 16.0001 144.9159 0.00065881 -70.3544 0.047946
7.152 0.98812 5.4756e-005 3.8183 0.011943 9.3178e-005 0.0011682 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.4666 0.52025 0.1591 0.01886 13.6649 0.11716 0.00015137 0.77299 0.0089192 0.0098877 0.014659 0.20441 0.082515 3.942e-005 0.00015992 0.16113 0.46811 0.52444 0.0050882 0.51035 0.34859 0.038463 0.42035 1.1764 1.1703 16.0002 144.9159 0.00065637 -71.1516 0.048946
7.153 0.98812 5.4756e-005 3.8183 0.011943 9.3191e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4667 0.52029 0.15912 0.018861 13.6675 0.11717 0.00015139 0.77298 0.0089197 0.0098882 0.012982 0.23211 0.092673 3.4349e-005 0.00013917 0.16113 0.46947 0.52739 0.0047439 0.51158 0.34876 0.030452 0.42023 1.1789 1.1729 16.0003 144.9158 0.00065394 -71.9223 0.049946
7.154 0.98812 5.4756e-005 3.8183 0.011943 9.3204e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4668 0.52034 0.15913 0.018862 13.6702 0.11718 0.0001514 0.77297 0.0089201 0.0098886 0.011541 0.26195 0.10377 3.0085e-005 0.00012174 0.16113 0.47086 0.53031 0.0044349 0.51282 0.34893 0.023927 0.42012 1.1815 1.1755 16.0004 144.9158 0.00065151 -72.6656 0.050946
7.155 0.98812 5.4756e-005 3.8183 0.011943 9.3217e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4668 0.52038 0.15914 0.018863 13.6728 0.11718 0.00015141 0.77297 0.0089206 0.0098891 0.010302 0.29383 0.11585 2.648e-005 0.00010705 0.16114 0.47227 0.5332 0.0041574 0.51408 0.3491 0.018728 0.42001 1.1841 1.1781 16.0005 144.9158 0.00064909 -73.3806 0.051946
7.156 0.98812 5.4756e-005 3.8183 0.011943 9.323e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4669 0.52043 0.15916 0.018864 13.6755 0.11719 0.00015142 0.77296 0.008921 0.0098896 0.0092344 0.32756 0.12898 2.3433e-005 9.4632e-005 0.16114 0.47369 0.53605 0.0039081 0.51537 0.34927 0.014675 0.41991 1.1867 1.1807 16.0006 144.9158 0.00064666 -74.0663 0.052946
7.157 0.98812 5.4756e-005 3.8183 0.011943 9.3243e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.467 0.52047 0.15917 0.018866 13.6781 0.1172 0.00015143 0.77295 0.0089214 0.0098901 0.0083147 0.3629 0.1432 2.0849e-005 8.412e-005 0.16114 0.47512 0.53888 0.0036843 0.51669 0.34945 0.01158 0.41981 1.1893 1.1833 16.0006 144.9157 0.00064425 -74.7218 0.053946
7.158 0.98812 5.4756e-005 3.8183 0.011943 9.3255e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4671 0.52052 0.15919 0.018867 13.6808 0.11721 0.00015144 0.77295 0.0089219 0.0098906 0.0075213 0.39955 0.15853 1.8652e-005 7.5198e-005 0.16115 0.47657 0.54167 0.0034833 0.51804 0.34962 0.0092629 0.41972 1.1919 1.1859 16.0007 144.9157 0.00064184 -75.3464 0.054946
7.159 0.98812 5.4756e-005 3.8183 0.011942 9.3268e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4672 0.52057 0.1592 0.018868 13.6834 0.11721 0.00015145 0.77294 0.0089223 0.009891 0.0068363 0.43716 0.17496 1.6783e-005 6.7607e-005 0.16115 0.47803 0.54443 0.0033028 0.51943 0.3498 0.0075573 0.41964 1.1945 1.1885 16.0008 144.9157 0.00063943 -75.9395 0.055946
7.16 0.98812 5.4756e-005 3.8183 0.011942 9.3281e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4673 0.52061 0.15921 0.018869 13.6861 0.11722 0.00015146 0.77293 0.0089228 0.0098915 0.0062442 0.47533 0.19249 1.5186e-005 6.1134e-005 0.16115 0.47949 0.54717 0.0031409 0.52085 0.34998 0.0063187 0.41956 1.197 1.1911 16.0009 144.9157 0.00063703 -76.5006 0.056946
7.161 0.98812 5.4756e-005 3.8183 0.011942 9.3294e-005 0.0011682 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4674 0.52066 0.15923 0.01887 13.6888 0.11723 0.00015147 0.77292 0.0089232 0.009892 0.0057316 0.51366 0.21106 1.382e-005 5.5602e-005 0.16116 0.48097 0.54987 0.0029957 0.52231 0.35016 0.0054265 0.41948 1.1996 1.1937 16.001 144.9156 0.00063464 -77.0298 0.057946
7.162 0.98812 5.4755e-005 3.8183 0.011942 9.3307e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4675 0.5207 0.15924 0.018872 13.6914 0.11724 0.00015148 0.77292 0.0089237 0.0098925 0.0052876 0.55171 0.23059 1.2651e-005 5.0863e-005 0.16116 0.48244 0.55255 0.0028655 0.52381 0.35034 0.004785 0.41941 1.2022 1.1963 16.0011 144.9156 0.00063226 -77.527 0.058946
7.163 0.98812 5.4755e-005 3.8183 0.011942 9.332e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4676 0.52075 0.15926 0.018873 13.6941 0.11724 0.00015149 0.77291 0.0089241 0.009893 0.0049022 0.58906 0.25101 1.1644e-005 4.6792e-005 0.16116 0.48392 0.55519 0.0027489 0.52535 0.35052 0.0043209 0.41934 1.2047 1.1988 16.0013 144.9156 0.00062988 -77.9926 0.059946
7.164 0.98812 5.4755e-005 3.8183 0.011942 9.3333e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.4676 0.52079 0.15927 0.018874 13.6967 0.11725 0.00015151 0.7729 0.0089246 0.0098934 0.0045672 0.62533 0.27218 1.0776e-005 4.3288e-005 0.16117 0.48541 0.55781 0.0026443 0.52693 0.35071 0.0039803 0.41928 1.2073 1.2014 16.0014 144.9156 0.00062751 -78.4274 0.060946
7.165 0.98812 5.4755e-005 3.8183 0.011942 9.3346e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.4677 0.52084 0.15929 0.018875 13.6994 0.11726 0.00015152 0.77289 0.008925 0.0098939 0.0042755 0.66016 0.29398 1.0028e-005 4.0263e-005 0.16117 0.48689 0.56041 0.0025507 0.52856 0.35089 0.0037247 0.41922 1.2099 1.204 16.0015 144.9155 0.00062515 -78.8321 0.061946
7.166 0.98812 5.4755e-005 3.8183 0.011942 9.3358e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.4678 0.52088 0.1593 0.018877 13.7021 0.11726 0.00015153 0.77289 0.0089255 0.0098944 0.0040211 0.69324 0.31629 9.3793e-006 3.7646e-005 0.16117 0.48838 0.56297 0.0024667 0.53022 0.35108 0.0035274 0.41917 1.2124 1.2066 16.0016 144.9155 0.0006228 -79.2077 0.062946
7.167 0.98812 5.4755e-005 3.8183 0.011942 9.3371e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.4679 0.52093 0.15931 0.018878 13.7047 0.11727 0.00015154 0.77288 0.0089259 0.0098949 0.0037987 0.72435 0.33895 8.8165e-006 3.5375e-005 0.16118 0.48987 0.56551 0.0023916 0.53192 0.35127 0.0033707 0.41912 1.215 1.2092 16.0017 144.9155 0.00062046 -79.5555 0.063946
7.168 0.98812 5.4755e-005 3.8183 0.011942 9.3384e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.468 0.52098 0.15933 0.018879 13.7074 0.11728 0.00015155 0.77287 0.0089264 0.0098953 0.0036041 0.7533 0.36183 8.3271e-006 3.34e-005 0.16118 0.49136 0.56802 0.0023242 0.53366 0.35146 0.0032427 0.41907 1.2175 1.2117 16.0018 144.9155 0.00061813 -79.8767 0.064946
7.169 0.98812 5.4755e-005 3.8183 0.011942 9.3397e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.4681 0.52102 0.15934 0.01888 13.71 0.11729 0.00015156 0.77286 0.0089268 0.0098958 0.0034333 0.77998 0.38481 7.8999e-006 3.1678e-005 0.16118 0.49284 0.5705 0.0022638 0.53543 0.35165 0.0031355 0.41903 1.2201 1.2143 16.0019 144.9155 0.0006158 -80.1728 0.065946
7.17 0.98812 5.4755e-005 3.8183 0.011942 9.341e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.4682 0.52107 0.15936 0.018881 13.7127 0.11729 0.00015157 0.77286 0.0089273 0.0098963 0.0032831 0.80436 0.40775 7.5262e-006 3.0172e-005 0.16119 0.49433 0.57296 0.0022097 0.53724 0.35185 0.0030439 0.41899 1.2226 1.2169 16.002 144.9155 0.00061349 -80.4453 0.066946
7.171 0.98812 5.4755e-005 3.8183 0.011942 9.3423e-005 0.0011683 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.4683 0.52111 0.15937 0.018883 13.7154 0.1173 0.00015158 0.77285 0.0089277 0.0098968 0.0031509 0.82644 0.43055 7.1987e-006 2.8853e-005 0.16119 0.49581 0.5754 0.0021612 0.53908 0.35204 0.0029644 0.41895 1.2252 1.2194 16.0022 144.9155 0.00061119 -80.6955 0.067946
7.172 0.98812 5.4755e-005 3.8183 0.011942 9.3436e-005 0.0011683 0.23367 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4684 0.52116 0.15938 0.018884 13.718 0.11731 0.00015159 0.77284 0.0089282 0.0098973 0.0030342 0.84627 0.4531 6.9109e-006 2.7693e-005 0.16119 0.4973 0.57781 0.0021176 0.54094 0.35224 0.0028949 0.41891 1.2277 1.222 16.0023 144.9154 0.0006089 -80.9251 0.068946
7.173 0.98812 5.4755e-005 3.8183 0.011942 9.3448e-005 0.0011683 0.23367 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4684 0.5212 0.1594 0.018885 13.7207 0.11732 0.0001516 0.77284 0.0089286 0.0098977 0.002931 0.86394 0.47532 6.6573e-006 2.6672e-005 0.1612 0.49878 0.58019 0.0020784 0.54284 0.35243 0.0028335 0.41888 1.2303 1.2245 16.0024 144.9154 0.00060662 -81.1354 0.069946
7.174 0.98812 5.4755e-005 3.8183 0.011942 9.3461e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4685 0.52125 0.15941 0.018886 13.7233 0.11732 0.00015161 0.77283 0.0089291 0.0098982 0.0028395 0.87959 0.49712 6.4331e-006 2.577e-005 0.1612 0.50026 0.58255 0.0020432 0.54476 0.35263 0.0027791 0.41885 1.2328 1.2271 16.0025 144.9154 0.00060435 -81.328 0.070946
7.175 0.98812 5.4754e-005 3.8183 0.011942 9.3474e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4686 0.52129 0.15943 0.018887 13.726 0.11733 0.00015163 0.77282 0.0089295 0.0098987 0.0027582 0.89336 0.51844 6.2346e-006 2.4972e-005 0.16121 0.50173 0.58489 0.0020116 0.5467 0.35283 0.0027308 0.41882 1.2353 1.2297 16.0026 144.9154 0.0006021 -81.5042 0.071946
7.176 0.98812 5.4754e-005 3.8183 0.011942 9.3487e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4687 0.52134 0.15944 0.018889 13.7287 0.11734 0.00015164 0.77281 0.00893 0.0098992 0.0026859 0.9054 0.53924 6.0587e-006 2.4264e-005 0.16121 0.5032 0.5872 0.001983 0.54867 0.35303 0.0026876 0.41879 1.2379 1.2322 16.0027 144.9154 0.00059985 -81.6654 0.072946
7.177 0.98812 5.4754e-005 3.8183 0.011942 9.35e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4688 0.52139 0.15946 0.01889 13.7313 0.11735 0.00015165 0.77281 0.0089304 0.0098997 0.0026214 0.91587 0.55945 5.9022e-006 2.3634e-005 0.16121 0.50467 0.58949 0.0019573 0.55065 0.35323 0.0026489 0.41876 1.2404 1.2347 16.0028 144.9154 0.00059762 -81.8128 0.073946
7.178 0.98812 5.4754e-005 3.8183 0.011942 9.3513e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4689 0.52143 0.15947 0.018891 13.734 0.11735 0.00015166 0.7728 0.0089309 0.0099001 0.0025638 0.92493 0.57907 5.7625e-006 2.3072e-005 0.16122 0.50614 0.59175 0.0019341 0.55265 0.35343 0.0026141 0.41874 1.2429 1.2373 16.003 144.9154 0.0005954 -81.9476 0.074946
7.179 0.98812 5.4754e-005 3.8183 0.011942 9.3526e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.469 0.52148 0.15948 0.018892 13.7367 0.11736 0.00015167 0.77279 0.0089313 0.0099006 0.002512 0.93274 0.59805 5.6374e-006 2.257e-005 0.16122 0.5076 0.594 0.0019131 0.55466 0.35363 0.0025829 0.41871 1.2454 1.2398 16.0031 144.9154 0.00059319 -82.0709 0.075946
7.18 0.98812 5.4754e-005 3.8183 0.011942 9.3538e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4691 0.52152 0.1595 0.018894 13.7393 0.11737 0.00015168 0.77278 0.0089317 0.0099011 0.0024656 0.93945 0.61638 5.5255e-006 2.212e-005 0.16122 0.50907 0.59622 0.0018941 0.55669 0.35383 0.0025548 0.41869 1.248 1.2424 16.0032 144.9154 0.00059099 -82.1838 0.076946
7.181 0.98812 5.4754e-005 3.8183 0.011942 9.3551e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4692 0.52157 0.15951 0.018895 13.742 0.11737 0.00015169 0.77278 0.0089322 0.0099016 0.0024239 0.94519 0.63406 5.4252e-006 2.1716e-005 0.16123 0.51052 0.59841 0.0018769 0.55872 0.35403 0.0025295 0.41867 1.2505 1.2449 16.0033 144.9154 0.0005888 -82.2871 0.077946
7.182 0.98812 5.4754e-005 3.8183 0.011942 9.3564e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4692 0.52161 0.15953 0.018896 13.7447 0.11738 0.0001517 0.77277 0.0089326 0.009902 0.0023863 0.95009 0.65107 5.3348e-006 2.1352e-005 0.16123 0.51198 0.60059 0.0018612 0.56077 0.35424 0.0025066 0.41865 1.253 1.2474 16.0034 144.9154 0.00058663 -82.3819 0.078946
7.183 0.98812 5.4754e-005 3.8183 0.011942 9.3577e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4693 0.52166 0.15954 0.018897 13.7473 0.11739 0.00015171 0.77276 0.0089331 0.0099025 0.002352 0.95427 0.66741 5.2526e-006 2.1023e-005 0.16123 0.51343 0.60275 0.0018469 0.56282 0.35444 0.0024858 0.41863 1.2555 1.2499 16.0035 144.9154 0.00058446 -82.4689 0.079946
7.184 0.98812 5.4754e-005 3.8183 0.011942 9.359e-005 0.0011683 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4694 0.5217 0.15955 0.018898 13.75 0.1174 0.00015172 0.77276 0.0089335 0.009903 0.0023212 0.95782 0.6831 5.1786e-006 2.0726e-005 0.16124 0.51487 0.60488 0.0018339 0.56488 0.35464 0.002467 0.41862 1.258 1.2525 16.0037 144.9154 0.00058231 -82.5488 0.080946
7.185 0.98812 5.4754e-005 3.8183 0.011942 9.3603e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4695 0.52175 0.15957 0.0189 13.7526 0.1174 0.00015173 0.77275 0.008934 0.0099035 0.0022933 0.96083 0.69814 5.1116e-006 2.0456e-005 0.16124 0.51631 0.60699 0.0018221 0.56694 0.35485 0.0024498 0.4186 1.2605 1.255 16.0038 144.9154 0.00058018 -82.6224 0.081946
7.186 0.98812 5.4754e-005 3.8183 0.011942 9.3616e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4696 0.52179 0.15958 0.018901 13.7553 0.11741 0.00015175 0.77274 0.0089344 0.009904 0.0022676 0.96338 0.71255 5.0503e-006 2.021e-005 0.16124 0.51775 0.60909 0.0018112 0.56901 0.35505 0.0024342 0.41858 1.263 1.2575 16.0039 144.9154 0.00057805 -82.6902 0.082946
7.187 0.98812 5.4753e-005 3.8183 0.011942 9.3629e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4697 0.52184 0.1596 0.018902 13.758 0.11742 0.00015176 0.77273 0.0089349 0.0099044 0.0022443 0.96555 0.72632 4.9945e-006 1.9986e-005 0.16125 0.51919 0.61116 0.0018012 0.57108 0.35526 0.0024199 0.41857 1.2655 1.26 16.004 144.9154 0.00057593 -82.7529 0.083946
7.188 0.98812 5.4753e-005 3.8183 0.011942 9.3641e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4698 0.52189 0.15961 0.018903 13.7606 0.11743 0.00015177 0.77273 0.0089353 0.0099049 0.0022229 0.96739 0.73949 4.9434e-006 1.9781e-005 0.16125 0.52062 0.61321 0.001792 0.57316 0.35546 0.0024067 0.41855 1.268 1.2625 16.0041 144.9154 0.00057383 -82.8108 0.084946
7.189 0.98812 5.4753e-005 3.8183 0.011942 9.3654e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4699 0.52193 0.15963 0.018904 13.7633 0.11743 0.00015178 0.77272 0.0089358 0.0099054 0.0022031 0.96895 0.75206 4.8964e-006 1.9592e-005 0.16125 0.52204 0.61524 0.0017835 0.57523 0.35567 0.0023947 0.41854 1.2705 1.265 16.0042 144.9154 0.00057174 -82.8646 0.085946
7.19 0.98812 5.4753e-005 3.8183 0.011942 9.3667e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.47 0.52198 0.15964 0.018906 13.766 0.11744 0.00015179 0.77271 0.0089362 0.0099059 0.002185 0.97028 0.76406 4.8531e-006 1.9419e-005 0.16126 0.52346 0.61726 0.0017757 0.57731 0.35587 0.0023836 0.41852 1.273 1.2675 16.0043 144.9154 0.00056966 -82.9146 0.086946
7.191 0.98812 5.4753e-005 3.8183 0.011942 9.368e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.47 0.52202 0.15965 0.018907 13.7686 0.11745 0.0001518 0.7727 0.0089367 0.0099063 0.0021682 0.97141 0.7755 4.8132e-006 1.9258e-005 0.16126 0.52488 0.61925 0.0017684 0.57938 0.35608 0.0023733 0.41851 1.2754 1.27 16.0044 144.9154 0.00056759 -82.9612 0.087946
7.192 0.98812 5.4753e-005 3.8183 0.011942 9.3693e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4701 0.52207 0.15967 0.018908 13.7713 0.11746 0.00015181 0.7727 0.0089371 0.0099068 0.0021525 0.97237 0.78641 4.7761e-006 1.911e-005 0.16126 0.5263 0.62123 0.0017616 0.58145 0.35629 0.0023638 0.4185 1.2779 1.2725 16.0046 144.9154 0.00056554 -83.0047 0.088946
7.193 0.98812 5.4753e-005 3.8183 0.011942 9.3706e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4702 0.52211 0.15968 0.018909 13.774 0.11746 0.00015182 0.77269 0.0089376 0.0099073 0.0021381 0.97319 0.7968 4.7417e-006 1.8972e-005 0.16127 0.52771 0.62318 0.0017553 0.58352 0.35649 0.002355 0.41849 1.2804 1.275 16.0047 144.9154 0.00056349 -83.0455 0.089946
7.194 0.98812 5.4753e-005 3.8183 0.011942 9.3719e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4703 0.52216 0.1597 0.018911 13.7767 0.11747 0.00015183 0.77268 0.008938 0.0099078 0.0021247 0.9739 0.80669 4.7096e-006 1.8843e-005 0.16127 0.52911 0.62512 0.0017494 0.58559 0.3567 0.0023468 0.41847 1.2829 1.2775 16.0048 144.9154 0.00056146 -83.0838 0.090946
7.195 0.98812 5.4753e-005 3.8183 0.011942 9.3731e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4704 0.5222 0.15971 0.018912 13.7793 0.11748 0.00015184 0.77267 0.0089384 0.0099082 0.0021119 0.97451 0.8161 4.6796e-006 1.8723e-005 0.16127 0.53052 0.62704 0.0017439 0.58765 0.35691 0.0023391 0.41846 1.2853 1.28 16.0049 144.9154 0.00055944 -83.1198 0.091946
7.196 0.98812 5.4753e-005 3.8183 0.011942 9.3744e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4705 0.52225 0.15972 0.018913 13.782 0.11748 0.00015185 0.77267 0.0089389 0.0099087 0.0021 0.97503 0.82505 4.6514e-006 1.861e-005 0.16128 0.53191 0.62894 0.0017386 0.58972 0.35711 0.0023318 0.41845 1.2878 1.2825 16.005 144.9154 0.00055743 -83.1539 0.092946
7.197 0.98812 5.4753e-005 3.8183 0.011942 9.3757e-005 0.0011684 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.4706 0.5223 0.15974 0.018914 13.7847 0.11749 0.00015186 0.77266 0.0089393 0.0099092 0.0020889 0.97549 0.83356 4.6249e-006 1.8504e-005 0.16128 0.53331 0.63082 0.0017337 0.59177 0.35732 0.0023251 0.41844 1.2903 1.285 16.0051 144.9154 0.00055543 -83.1861 0.093946
7.198 0.98812 5.4753e-005 3.8183 0.011942 9.377e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4707 0.52234 0.15975 0.018915 13.7873 0.1175 0.00015188 0.77265 0.0089398 0.0099097 0.0020783 0.97589 0.84165 4.5999e-006 1.8403e-005 0.16129 0.5347 0.63269 0.0017291 0.59383 0.35753 0.0023186 0.41843 1.2927 1.2874 16.0052 144.9154 0.00055344 -83.2167 0.094946
7.199 0.98812 5.4753e-005 3.8183 0.011942 9.3783e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4708 0.52239 0.15977 0.018917 13.79 0.11751 0.00015189 0.77265 0.0089402 0.0099102 0.0020683 0.97624 0.84934 4.5762e-006 1.8308e-005 0.16129 0.53608 0.63453 0.0017246 0.59588 0.35773 0.0023126 0.41842 1.2952 1.2899 16.0053 144.9154 0.00055147 -83.2459 0.095946
7.2 0.98812 5.4752e-005 3.8183 0.011942 9.3796e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4709 0.52243 0.15978 0.018918 13.7927 0.11751 0.0001519 0.77264 0.0089407 0.0099106 0.0020588 0.97655 0.85664 4.5537e-006 1.8218e-005 0.16129 0.53747 0.63636 0.0017204 0.59792 0.35794 0.0023068 0.41841 1.2976 1.2924 16.0054 144.9154 0.0005495 -83.2737 0.096946
7.201 0.98812 5.4752e-005 3.8183 0.011942 9.3809e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4709 0.52248 0.1598 0.018919 13.7953 0.11752 0.00015191 0.77263 0.0089411 0.0099111 0.0020497 0.97683 0.86358 4.5323e-006 1.8132e-005 0.1613 0.53884 0.63818 0.0017164 0.59996 0.35815 0.0023014 0.4184 1.3001 1.2948 16.0055 144.9154 0.00054755 -83.3003 0.097946
7.202 0.98812 5.4752e-005 3.8183 0.011942 9.3821e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.471 0.52252 0.15981 0.01892 13.798 0.11753 0.00015192 0.77262 0.0089416 0.0099116 0.0020411 0.97707 0.87016 4.5118e-006 1.805e-005 0.1613 0.54022 0.63997 0.0017126 0.60199 0.35836 0.0022962 0.41839 1.3025 1.2973 16.0056 144.9154 0.00054561 -83.3258 0.098946
7.203 0.98812 5.4752e-005 3.8183 0.011942 9.3834e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4711 0.52257 0.15982 0.018921 13.8007 0.11754 0.00015193 0.77262 0.008942 0.0099121 0.0020328 0.9773 0.87641 4.4923e-006 1.7972e-005 0.1613 0.54159 0.64176 0.0017089 0.60402 0.35856 0.0022912 0.41839 1.305 1.2997 16.0057 144.9154 0.00054368 -83.3504 0.099946
7.204 0.98812 5.4752e-005 3.8183 0.011942 9.3847e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4712 0.52261 0.15984 0.018923 13.8034 0.11754 0.00015194 0.77261 0.0089425 0.0099125 0.0020248 0.9775 0.88234 4.4735e-006 1.7896e-005 0.16131 0.54295 0.64352 0.0017053 0.60605 0.35877 0.0022864 0.41838 1.3074 1.3022 16.0058 144.9154 0.00054176 -83.374 0.10095
7.205 0.98812 5.4752e-005 3.8183 0.011942 9.386e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4713 0.52266 0.15985 0.018924 13.806 0.11755 0.00015195 0.7726 0.0089429 0.009913 0.0020172 0.97768 0.88797 4.4554e-006 1.7824e-005 0.16131 0.54431 0.64527 0.0017019 0.60806 0.35898 0.0022818 0.41837 1.3098 1.3047 16.0059 144.9154 0.00053985 -83.3969 0.10195
7.206 0.98812 5.4752e-005 3.8183 0.011942 9.3873e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4714 0.5227 0.15987 0.018925 13.8087 0.11756 0.00015196 0.77259 0.0089433 0.0099135 0.0020098 0.97785 0.8933 4.438e-006 1.7754e-005 0.16131 0.54567 0.647 0.0016986 0.61007 0.35919 0.0022774 0.41836 1.3123 1.3071 16.0061 144.9154 0.00053795 -83.419 0.10295
7.207 0.98812 5.4752e-005 3.8183 0.011942 9.3886e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4715 0.52275 0.15988 0.018926 13.8114 0.11756 0.00015197 0.77259 0.0089438 0.009914 0.0020027 0.978 0.89837 4.4212e-006 1.7687e-005 0.16132 0.54702 0.64872 0.0016954 0.61208 0.35939 0.0022731 0.41835 1.3147 1.3095 16.0062 144.9154 0.00053606 -83.4404 0.10395
7.208 0.98812 5.4752e-005 3.8183 0.011942 9.3899e-005 0.0011684 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4716 0.5228 0.15989 0.018927 13.8141 0.11757 0.00015198 0.77258 0.0089442 0.0099144 0.0019957 0.97815 0.90317 4.4049e-006 1.7622e-005 0.16132 0.54837 0.65042 0.0016923 0.61408 0.3596 0.002269 0.41835 1.3171 1.312 16.0063 144.9154 0.00053418 -83.4612 0.10495
7.209 0.98812 5.4752e-005 3.8183 0.011942 9.3912e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4717 0.52284 0.15991 0.018929 13.8167 0.11758 0.000152 0.77257 0.0089447 0.0099149 0.001989 0.97828 0.90772 4.3891e-006 1.7558e-005 0.16132 0.54972 0.6521 0.0016893 0.61607 0.35981 0.0022649 0.41834 1.3195 1.3144 16.0064 144.9154 0.00053232 -83.4815 0.10595
7.21 0.98812 5.4752e-005 3.8183 0.011942 9.3924e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4717 0.52289 0.15992 0.01893 13.8194 0.11759 0.00015201 0.77257 0.0089451 0.0099154 0.0019825 0.97841 0.91203 4.3737e-006 1.7497e-005 0.16133 0.55106 0.65377 0.0016864 0.61806 0.36002 0.002261 0.41833 1.3219 1.3168 16.0065 144.9154 0.00053046 -83.5013 0.10695
7.211 0.98812 5.4752e-005 3.8183 0.011942 9.3937e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4718 0.52293 0.15994 0.018931 13.8221 0.11759 0.00015202 0.77256 0.0089456 0.0099159 0.0019762 0.97853 0.91612 4.3588e-006 1.7437e-005 0.16133 0.5524 0.65543 0.0016836 0.62004 0.36023 0.0022573 0.41833 1.3244 1.3193 16.0066 144.9155 0.00052862 -83.5206 0.10795
7.212 0.98812 5.4752e-005 3.8183 0.011942 9.395e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4719 0.52298 0.15995 0.018932 13.8248 0.1176 0.00015203 0.77255 0.008946 0.0099163 0.00197 0.97865 0.92 4.3443e-006 1.7379e-005 0.16133 0.55373 0.65707 0.0016808 0.62201 0.36044 0.0022536 0.41832 1.3268 1.3217 16.0067 144.9155 0.00052678 -83.5395 0.10895
7.213 0.98812 5.4751e-005 3.8183 0.011942 9.3963e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.472 0.52302 0.15997 0.018934 13.8274 0.11761 0.00015204 0.77254 0.0089465 0.0099168 0.001964 0.97875 0.92367 4.3301e-006 1.7322e-005 0.16134 0.55506 0.6587 0.001678 0.62398 0.36064 0.00225 0.41831 1.3292 1.3241 16.0068 144.9155 0.00052496 -83.558 0.10995
7.214 0.98812 5.4751e-005 3.8183 0.011942 9.3976e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4721 0.52307 0.15998 0.018935 13.8301 0.11762 0.00015205 0.77254 0.0089469 0.0099173 0.0019581 0.97886 0.92716 4.3162e-006 1.7267e-005 0.16134 0.55638 0.66031 0.0016754 0.62593 0.36085 0.0022464 0.41831 1.3316 1.3265 16.0069 144.9155 0.00052314 -83.5761 0.11095
7.215 0.98812 5.4751e-005 3.8183 0.011942 9.3989e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4722 0.52311 0.15999 0.018936 13.8328 0.11762 0.00015206 0.77253 0.0089474 0.0099178 0.0019524 0.97896 0.93045 4.3026e-006 1.7212e-005 0.16134 0.5577 0.66191 0.0016728 0.62789 0.36106 0.002243 0.4183 1.334 1.329 16.007 144.9155 0.00052134 -83.5939 0.11195
7.216 0.98812 5.4751e-005 3.8183 0.011942 9.4002e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4723 0.52316 0.16001 0.018937 13.8355 0.11763 0.00015207 0.77252 0.0089478 0.0099182 0.0019467 0.97905 0.93358 4.2894e-006 1.7159e-005 0.16135 0.55902 0.66349 0.0016702 0.62983 0.36127 0.0022396 0.4183 1.3364 1.3314 16.007 144.9155 0.00051954 -83.6113 0.11295
7.217 0.98812 5.4751e-005 3.8183 0.011941 9.4014e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4724 0.52321 0.16002 0.018938 13.8381 0.11764 0.00015208 0.77251 0.0089482 0.0099187 0.0019412 0.97914 0.93654 4.2764e-006 1.7107e-005 0.16135 0.56033 0.66506 0.0016677 0.63177 0.36148 0.0022363 0.41829 1.3387 1.3338 16.0071 144.9155 0.00051776 -83.6285 0.11395
7.218 0.98812 5.4751e-005 3.8183 0.011941 9.4027e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4725 0.52325 0.16004 0.01894 13.8408 0.11764 0.00015209 0.77251 0.0089487 0.0099192 0.0019358 0.97923 0.93934 4.2636e-006 1.7056e-005 0.16135 0.56164 0.66662 0.0016653 0.6337 0.36169 0.0022331 0.41829 1.3411 1.3362 16.0072 144.9155 0.00051598 -83.6453 0.11495
7.219 0.98812 5.4751e-005 3.8183 0.011941 9.404e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4725 0.5233 0.16005 0.018941 13.8435 0.11765 0.0001521 0.7725 0.0089491 0.0099197 0.0019304 0.97932 0.94199 4.2511e-006 1.7006e-005 0.16136 0.56295 0.66816 0.0016628 0.63563 0.36189 0.0022299 0.41828 1.3435 1.3386 16.0073 144.9155 0.00051422 -83.662 0.11595
7.22 0.98812 5.4751e-005 3.8183 0.011941 9.4053e-005 0.0011685 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4726 0.52334 0.16006 0.018942 13.8462 0.11766 0.00015211 0.77249 0.0089496 0.0099201 0.0019252 0.9794 0.94451 4.2388e-006 1.6957e-005 0.16136 0.56425 0.66969 0.0016605 0.63755 0.3621 0.0022267 0.41828 1.3459 1.341 16.0074 144.9155 0.00051247 -83.6783 0.11695
7.221 0.98812 5.4751e-005 3.8183 0.011941 9.4066e-005 0.0011685 0.23369 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.4727 0.52339 0.16008 0.018943 13.8488 0.11767 0.00015213 0.77249 0.00895 0.0099206 0.00192 0.97948 0.94689 4.2267e-006 1.6908e-005 0.16136 0.56555 0.6712 0.0016581 0.63946 0.36231 0.0022237 0.41827 1.3483 1.3434 16.0075 144.9155 0.00051072 -83.6945 0.11795
7.222 0.98812 5.4751e-005 3.8183 0.011941 9.4079e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4728 0.52343 0.16009 0.018944 13.8515 0.11767 0.00015214 0.77248 0.0089505 0.0099211 0.001915 0.97956 0.94914 4.2148e-006 1.6861e-005 0.16137 0.56684 0.67271 0.0016558 0.64136 0.36252 0.0022206 0.41827 1.3506 1.3457 16.0076 144.9155 0.00050899 -83.7104 0.11895
7.223 0.98812 5.4751e-005 3.8183 0.011941 9.4092e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4729 0.52348 0.16011 0.018946 13.8542 0.11768 0.00015215 0.77247 0.0089509 0.0099216 0.00191 0.97964 0.95128 4.2031e-006 1.6814e-005 0.16137 0.56813 0.6742 0.0016535 0.64326 0.36273 0.0022176 0.41826 1.353 1.3481 16.0077 144.9155 0.00050726 -83.7261 0.11995
7.224 0.98812 5.4751e-005 3.8183 0.011941 9.4104e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.473 0.52352 0.16012 0.018947 13.8569 0.11769 0.00015216 0.77246 0.0089513 0.009922 0.0019051 0.97972 0.9533 4.1915e-006 1.6768e-005 0.16137 0.56942 0.67567 0.0016513 0.64515 0.36294 0.0022147 0.41826 1.3554 1.3505 16.0078 144.9155 0.00050554 -83.7416 0.12095
7.225 0.98812 5.475e-005 3.8183 0.011941 9.4117e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4731 0.52357 0.16013 0.018948 13.8596 0.1177 0.00015217 0.77246 0.0089518 0.0099225 0.0019002 0.97979 0.95521 4.1801e-006 1.6722e-005 0.16138 0.5707 0.67714 0.0016491 0.64703 0.36315 0.0022118 0.41825 1.3577 1.3529 16.0079 144.9155 0.00050384 -83.757 0.12195
7.226 0.98812 5.475e-005 3.8183 0.011941 9.413e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4732 0.52361 0.16015 0.018949 13.8622 0.1177 0.00015218 0.77245 0.0089522 0.009923 0.0018955 0.97987 0.95702 4.1689e-006 1.6677e-005 0.16138 0.57197 0.67859 0.0016469 0.6489 0.36335 0.0022089 0.41825 1.3601 1.3552 16.008 144.9155 0.00050214 -83.7721 0.12295
7.227 0.98812 5.475e-005 3.8183 0.011941 9.4143e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4733 0.52366 0.16016 0.01895 13.8649 0.11771 0.00015219 0.77244 0.0089527 0.0099235 0.0018908 0.97994 0.95874 4.1579e-006 1.6633e-005 0.16139 0.57325 0.68003 0.0016447 0.65077 0.36356 0.0022061 0.41825 1.3624 1.3576 16.0081 144.9155 0.00050045 -83.7871 0.12395
7.228 0.98812 5.475e-005 3.8183 0.011941 9.4156e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4733 0.52371 0.16018 0.018952 13.8676 0.11772 0.0001522 0.77243 0.0089531 0.0099239 0.0018861 0.98001 0.96036 4.147e-006 1.6589e-005 0.16139 0.57452 0.68146 0.0016426 0.65263 0.36377 0.0022033 0.41824 1.3648 1.36 16.0082 144.9156 0.00049878 -83.802 0.12495
7.229 0.98812 5.475e-005 3.8183 0.011941 9.4169e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4734 0.52375 0.16019 0.018953 13.8703 0.11772 0.00015221 0.77243 0.0089536 0.0099244 0.0018815 0.98008 0.9619 4.1363e-006 1.6546e-005 0.16139 0.57578 0.68288 0.0016405 0.65448 0.36398 0.0022005 0.41824 1.3671 1.3623 16.0083 144.9156 0.00049711 -83.8166 0.12595
7.23 0.98812 5.475e-005 3.8183 0.011941 9.4182e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4735 0.5238 0.16021 0.018954 13.873 0.11773 0.00015222 0.77242 0.008954 0.0099249 0.001877 0.98015 0.96335 4.1257e-006 1.6504e-005 0.1614 0.57705 0.68428 0.0016384 0.65633 0.36419 0.0021978 0.41824 1.3695 1.3647 16.0083 144.9156 0.00049545 -83.8311 0.12695
7.231 0.98812 5.475e-005 3.8183 0.011941 9.4194e-005 0.0011685 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4736 0.52384 0.16022 0.018955 13.8756 0.11774 0.00015223 0.77241 0.0089545 0.0099254 0.0018725 0.98021 0.96473 4.1152e-006 1.6462e-005 0.1614 0.5783 0.68567 0.0016363 0.65817 0.3644 0.0021951 0.41823 1.3718 1.367 16.0084 144.9156 0.0004938 -83.8455 0.12795
7.232 0.98812 5.475e-005 3.8183 0.011941 9.4207e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4737 0.52389 0.16023 0.018957 13.8783 0.11775 0.00015224 0.77241 0.0089549 0.0099258 0.0018681 0.98028 0.96603 4.1048e-006 1.6421e-005 0.1614 0.57956 0.68705 0.0016343 0.66 0.36461 0.0021924 0.41823 1.3741 1.3694 16.0085 144.9156 0.00049216 -83.8597 0.12895
7.233 0.98812 5.475e-005 3.8183 0.011941 9.422e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4738 0.52393 0.16025 0.018958 13.881 0.11775 0.00015226 0.7724 0.0089553 0.0099263 0.0018638 0.98035 0.96726 4.0946e-006 1.638e-005 0.16141 0.58081 0.68842 0.0016323 0.66182 0.36482 0.0021898 0.41823 1.3765 1.3717 16.0086 144.9156 0.00049052 -83.8738 0.12995
7.234 0.98812 5.475e-005 3.8183 0.011941 9.4233e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4739 0.52398 0.16026 0.018959 13.8837 0.11776 0.00015227 0.77239 0.0089558 0.0099268 0.0018594 0.98041 0.96843 4.0845e-006 1.6339e-005 0.16141 0.58206 0.68978 0.0016303 0.66364 0.36503 0.0021872 0.41823 1.3788 1.3741 16.0087 144.9156 0.0004889 -83.8878 0.13095
7.235 0.98812 5.475e-005 3.8183 0.011941 9.4246e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.474 0.52402 0.16028 0.01896 13.8864 0.11777 0.00015228 0.77238 0.0089562 0.0099273 0.0018552 0.98047 0.96953 4.0746e-006 1.63e-005 0.16141 0.5833 0.69113 0.0016283 0.66545 0.36523 0.0021846 0.41822 1.3811 1.3764 16.0088 144.9156 0.00048728 -83.9016 0.13195
7.236 0.98812 5.475e-005 3.8183 0.011941 9.4259e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4741 0.52407 0.16029 0.018961 13.8891 0.11778 0.00015229 0.77238 0.0089567 0.0099277 0.001851 0.98054 0.97058 4.0647e-006 1.626e-005 0.16142 0.58454 0.69246 0.0016264 0.66725 0.36544 0.002182 0.41822 1.3834 1.3787 16.0089 144.9156 0.00048568 -83.9152 0.13295
7.237 0.98812 5.475e-005 3.8183 0.011941 9.4272e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4741 0.52411 0.1603 0.018963 13.8917 0.11778 0.0001523 0.77237 0.0089571 0.0099282 0.0018468 0.9806 0.97157 4.055e-006 1.6221e-005 0.16142 0.58578 0.69379 0.0016244 0.66904 0.36565 0.0021795 0.41822 1.3857 1.3811 16.009 144.9156 0.00048408 -83.9288 0.13395
7.238 0.98812 5.4749e-005 3.8183 0.011941 9.4284e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4742 0.52416 0.16032 0.018964 13.8944 0.11779 0.00015231 0.77236 0.0089576 0.0099287 0.0018427 0.98066 0.97251 4.0453e-006 1.6183e-005 0.16142 0.58701 0.6951 0.0016225 0.67083 0.36586 0.002177 0.41822 1.388 1.3834 16.009 144.9156 0.00048249 -83.9422 0.13495
7.239 0.98812 5.4749e-005 3.8183 0.011941 9.4297e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4743 0.52421 0.16033 0.018965 13.8971 0.1178 0.00015232 0.77235 0.008958 0.0099292 0.0018386 0.98072 0.97339 4.0358e-006 1.6145e-005 0.16143 0.58824 0.69641 0.0016206 0.67261 0.36607 0.0021746 0.41822 1.3903 1.3857 16.0091 144.9156 0.00048091 -83.9555 0.13595
7.24 0.98812 5.4749e-005 3.8183 0.011941 9.431e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4744 0.52425 0.16035 0.018966 13.8998 0.1178 0.00015233 0.77235 0.0089584 0.0099296 0.0018346 0.98078 0.97423 4.0264e-006 1.6107e-005 0.16143 0.58946 0.6977 0.0016188 0.67438 0.36628 0.0021721 0.41821 1.3926 1.388 16.0092 144.9156 0.00047934 -83.9687 0.13695
7.241 0.98812 5.4749e-005 3.8183 0.011941 9.4323e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4745 0.5243 0.16036 0.018967 13.9025 0.11781 0.00015234 0.77234 0.0089589 0.0099301 0.0018306 0.98083 0.97502 4.0171e-006 1.607e-005 0.16143 0.59068 0.69898 0.0016169 0.67615 0.36649 0.0021697 0.41821 1.3949 1.3903 16.0093 144.9156 0.00047778 -83.9818 0.13795
7.242 0.98812 5.4749e-005 3.8183 0.011941 9.4336e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4746 0.52434 0.16037 0.018969 13.9052 0.11782 0.00015235 0.77233 0.0089593 0.0099306 0.0018267 0.98089 0.97577 4.0079e-006 1.6033e-005 0.16144 0.5919 0.70026 0.0016151 0.67791 0.3667 0.0021673 0.41821 1.3972 1.3926 16.0094 144.9157 0.00047623 -83.9947 0.13895
7.243 0.98812 5.4749e-005 3.8183 0.011941 9.4349e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4747 0.52439 0.16039 0.01897 13.9079 0.11783 0.00015236 0.77233 0.0089598 0.009931 0.0018228 0.98095 0.97648 3.9988e-006 1.5996e-005 0.16144 0.59311 0.70152 0.0016133 0.67966 0.36691 0.0021649 0.41821 1.3995 1.3949 16.0095 144.9157 0.00047468 -84.0076 0.13995
7.244 0.98812 5.4749e-005 3.8183 0.011941 9.4362e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4748 0.52443 0.1604 0.018971 13.9105 0.11783 0.00015237 0.77232 0.0089602 0.0099315 0.001819 0.98101 0.97716 3.9898e-006 1.596e-005 0.16144 0.59432 0.70277 0.0016115 0.6814 0.36712 0.0021626 0.41821 1.4018 1.3972 16.0095 144.9157 0.00047314 -84.0203 0.14095
7.245 0.98812 5.4749e-005 3.8183 0.011941 9.4375e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4749 0.52448 0.16042 0.018972 13.9132 0.11784 0.00015239 0.77231 0.0089607 0.009932 0.0018152 0.98106 0.97779 3.9809e-006 1.5925e-005 0.16145 0.59553 0.70401 0.0016097 0.68314 0.36732 0.0021602 0.41821 1.4041 1.3995 16.0096 144.9157 0.00047161 -84.0329 0.14195
7.246 0.98812 5.4749e-005 3.8183 0.011941 9.4387e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.4749 0.52452 0.16043 0.018973 13.9159 0.11785 0.0001524 0.7723 0.0089611 0.0099325 0.0018114 0.98112 0.9784 3.9721e-006 1.589e-005 0.16145 0.59673 0.70524 0.0016079 0.68486 0.36753 0.0021579 0.41821 1.4064 1.4018 16.0097 144.9157 0.00047009 -84.0454 0.14295
7.247 0.98812 5.4749e-005 3.8183 0.011941 9.44e-005 0.0011686 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.475 0.52457 0.16045 0.018975 13.9186 0.11786 0.00015241 0.7723 0.0089615 0.0099329 0.0018077 0.98117 0.97897 3.9634e-006 1.5855e-005 0.16145 0.59793 0.70647 0.0016062 0.68658 0.36774 0.0021557 0.41821 1.4086 1.4041 16.0098 144.9157 0.00046858 -84.0578 0.14395
7.248 0.98812 5.4749e-005 3.8183 0.011941 9.4413e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4751 0.52462 0.16046 0.018976 13.9213 0.11786 0.00015242 0.77229 0.008962 0.0099334 0.001804 0.98122 0.97951 3.9548e-006 1.582e-005 0.16146 0.59912 0.70768 0.0016045 0.6883 0.36795 0.0021534 0.41821 1.4109 1.4064 16.0099 144.9157 0.00046708 -84.0701 0.14495
7.249 0.98812 5.4749e-005 3.8183 0.011941 9.4426e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4752 0.52466 0.16047 0.018977 13.924 0.11787 0.00015243 0.77228 0.0089624 0.0099339 0.0018003 0.98128 0.98002 3.9463e-006 1.5786e-005 0.16146 0.60031 0.70888 0.0016028 0.69 0.36816 0.0021512 0.41821 1.4132 1.4087 16.0099 144.9157 0.00046558 -84.0823 0.14595
7.25 0.98812 5.4748e-005 3.8183 0.011941 9.4439e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4753 0.52471 0.16049 0.018978 13.9267 0.11788 0.00015244 0.77227 0.0089629 0.0099344 0.0017967 0.98133 0.9805 3.9378e-006 1.5752e-005 0.16146 0.6015 0.71008 0.0016011 0.6917 0.36837 0.0021489 0.41821 1.4154 1.4109 16.01 144.9157 0.00046409 -84.0944 0.14695
7.251 0.98812 5.4748e-005 3.8183 0.011941 9.4452e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4754 0.52475 0.1605 0.018979 13.9294 0.11788 0.00015245 0.77227 0.0089633 0.0099348 0.0017931 0.98138 0.98096 3.9295e-006 1.5719e-005 0.16147 0.60268 0.71126 0.0015994 0.6934 0.36858 0.0021468 0.41821 1.4177 1.4132 16.0101 144.9157 0.00046261 -84.1064 0.14795
7.252 0.98812 5.4748e-005 3.8183 0.011941 9.4465e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4755 0.5248 0.16052 0.018981 13.932 0.11789 0.00015246 0.77226 0.0089638 0.0099353 0.0017896 0.98143 0.9814 3.9212e-006 1.5686e-005 0.16147 0.60386 0.71244 0.0015977 0.69508 0.36879 0.0021446 0.41821 1.4199 1.4155 16.0102 144.9157 0.00046114 -84.1183 0.14895
7.253 0.98812 5.4748e-005 3.8183 0.011941 9.4477e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4756 0.52484 0.16053 0.018982 13.9347 0.1179 0.00015247 0.77225 0.0089642 0.0099358 0.0017861 0.98148 0.98181 3.913e-006 1.5653e-005 0.16147 0.60504 0.71361 0.0015961 0.69676 0.369 0.0021424 0.41821 1.4222 1.4177 16.0102 144.9158 0.00045968 -84.1301 0.14995
7.254 0.98812 5.4748e-005 3.8183 0.011941 9.449e-005 0.0011686 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4757 0.52489 0.16054 0.018983 13.9374 0.11791 0.00015248 0.77225 0.0089646 0.0099362 0.0017826 0.98153 0.9822 3.9049e-006 1.5621e-005 0.16148 0.60621 0.71476 0.0015944 0.69843 0.36921 0.0021403 0.41821 1.4244 1.42 16.0103 144.9158 0.00045822 -84.1418 0.15095
7.255 0.98812 5.4748e-005 3.8183 0.011941 9.4503e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4757 0.52493 0.16056 0.018984 13.9401 0.11791 0.00015249 0.77224 0.0089651 0.0099367 0.0017792 0.98158 0.98257 3.8969e-006 1.5589e-005 0.16148 0.60738 0.71591 0.0015928 0.70009 0.36942 0.0021382 0.41821 1.4267 1.4223 16.0104 144.9158 0.00045677 -84.1534 0.15195
7.256 0.98812 5.4748e-005 3.8183 0.011941 9.4516e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4758 0.52498 0.16057 0.018985 13.9428 0.11792 0.0001525 0.77223 0.0089655 0.0099372 0.0017758 0.98163 0.98292 3.889e-006 1.5557e-005 0.16148 0.60855 0.71705 0.0015912 0.70174 0.36963 0.0021361 0.41821 1.4289 1.4245 16.0105 144.9158 0.00045533 -84.1649 0.15295
7.257 0.98812 5.4748e-005 3.8183 0.011941 9.4529e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4759 0.52502 0.16059 0.018987 13.9455 0.11793 0.00015251 0.77222 0.008966 0.0099377 0.0017724 0.98168 0.98325 3.8811e-006 1.5526e-005 0.16149 0.60971 0.71818 0.0015896 0.70339 0.36984 0.002134 0.41821 1.4311 1.4267 16.0105 144.9158 0.0004539 -84.1763 0.15395
7.258 0.98812 5.4748e-005 3.8183 0.011941 9.4542e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.476 0.52507 0.1606 0.018988 13.9482 0.11794 0.00015253 0.77222 0.0089664 0.0099381 0.0017691 0.98173 0.98357 3.8734e-006 1.5494e-005 0.16149 0.61087 0.71931 0.0015881 0.70503 0.37004 0.0021319 0.41821 1.4333 1.429 16.0106 144.9158 0.00045247 -84.1876 0.15495
7.259 0.98812 5.4748e-005 3.8183 0.011941 9.4555e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4761 0.52512 0.16061 0.018989 13.9509 0.11794 0.00015254 0.77221 0.0089668 0.0099386 0.0017658 0.98178 0.98386 3.8657e-006 1.5464e-005 0.16149 0.61203 0.72042 0.0015865 0.70667 0.37025 0.0021299 0.41821 1.4356 1.4312 16.0107 144.9158 0.00045105 -84.1989 0.15595
7.26 0.98812 5.4748e-005 3.8183 0.011941 9.4567e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4762 0.52516 0.16063 0.01899 13.9536 0.11795 0.00015255 0.7722 0.0089673 0.0099391 0.0017625 0.98182 0.98415 3.8581e-006 1.5433e-005 0.1615 0.61318 0.72153 0.001585 0.70829 0.37046 0.0021279 0.41821 1.4378 1.4335 16.0108 144.9158 0.00044964 -84.21 0.15695
7.261 0.98812 5.4748e-005 3.8183 0.011941 9.458e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4763 0.52521 0.16064 0.018991 13.9563 0.11796 0.00015256 0.7722 0.0089677 0.0099396 0.0017593 0.98187 0.98441 3.8506e-006 1.5403e-005 0.1615 0.61433 0.72262 0.0015834 0.70991 0.37067 0.0021259 0.41821 1.44 1.4357 16.0108 144.9158 0.00044824 -84.221 0.15795
7.262 0.98812 5.4748e-005 3.8183 0.011941 9.4593e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.4764 0.52525 0.16066 0.018993 13.9589 0.11796 0.00015257 0.77219 0.0089682 0.00994 0.0017561 0.98191 0.98467 3.8431e-006 1.5373e-005 0.16151 0.61547 0.72371 0.0015819 0.71152 0.37088 0.0021239 0.41822 1.4422 1.4379 16.0109 144.9158 0.00044684 -84.232 0.15895
7.263 0.98812 5.4747e-005 3.8183 0.011941 9.4606e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4765 0.5253 0.16067 0.018994 13.9616 0.11797 0.00015258 0.77218 0.0089686 0.0099405 0.0017529 0.98196 0.98491 3.8357e-006 1.5344e-005 0.16151 0.61661 0.72479 0.0015804 0.71312 0.37109 0.0021219 0.41822 1.4444 1.4401 16.011 144.9158 0.00044545 -84.2429 0.15995
7.264 0.98812 5.4747e-005 3.8183 0.011941 9.4619e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4765 0.52534 0.16069 0.018995 13.9643 0.11798 0.00015259 0.77217 0.008969 0.009941 0.0017498 0.982 0.98514 3.8284e-006 1.5314e-005 0.16151 0.61775 0.72587 0.0015789 0.71472 0.3713 0.00212 0.41822 1.4466 1.4423 16.0111 144.9159 0.00044407 -84.2536 0.16095
7.265 0.98812 5.4747e-005 3.8183 0.011941 9.4632e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4766 0.52539 0.1607 0.018996 13.967 0.11799 0.0001526 0.77217 0.0089695 0.0099414 0.0017467 0.98205 0.98536 3.8212e-006 1.5286e-005 0.16152 0.61889 0.72693 0.0015774 0.71631 0.37151 0.0021181 0.41822 1.4488 1.4445 16.0111 144.9159 0.0004427 -84.2643 0.16195
7.266 0.98812 5.4747e-005 3.8183 0.011941 9.4645e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4767 0.52543 0.16071 0.018997 13.9697 0.11799 0.00015261 0.77216 0.0089699 0.0099419 0.0017436 0.98209 0.98556 3.814e-006 1.5257e-005 0.16152 0.62002 0.72799 0.001576 0.71789 0.37172 0.0021161 0.41822 1.451 1.4468 16.0112 144.9159 0.00044133 -84.2749 0.16295
7.267 0.98812 5.4747e-005 3.8183 0.011941 9.4657e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4768 0.52548 0.16073 0.018999 13.9724 0.118 0.00015262 0.77215 0.0089704 0.0099424 0.0017406 0.98214 0.98576 3.8069e-006 1.5228e-005 0.16152 0.62114 0.72904 0.0015745 0.71947 0.37193 0.0021142 0.41822 1.4532 1.449 16.0113 144.9159 0.00043998 -84.2855 0.16395
7.268 0.98812 5.4747e-005 3.8183 0.011941 9.467e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4769 0.52552 0.16074 0.019 13.9751 0.11801 0.00015263 0.77214 0.0089708 0.0099428 0.0017376 0.98218 0.98594 3.7999e-006 1.52e-005 0.16153 0.62227 0.73008 0.0015731 0.72104 0.37214 0.0021124 0.41823 1.4554 1.4512 16.0113 144.9159 0.00043862 -84.2959 0.16495
7.269 0.98812 5.4747e-005 3.8183 0.011941 9.4683e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.477 0.52557 0.16076 0.019001 13.9778 0.11802 0.00015264 0.77214 0.0089713 0.0099433 0.0017346 0.98222 0.98612 3.7929e-006 1.5173e-005 0.16153 0.62339 0.73111 0.0015717 0.7226 0.37235 0.0021105 0.41823 1.4575 1.4533 16.0114 144.9159 0.00043728 -84.3062 0.16595
7.27 0.98812 5.4747e-005 3.8183 0.011941 9.4696e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4771 0.52562 0.16077 0.019002 13.9805 0.11802 0.00015266 0.77213 0.0089717 0.0099438 0.0017316 0.98226 0.98629 3.7861e-006 1.5145e-005 0.16153 0.6245 0.73214 0.0015703 0.72415 0.37256 0.0021087 0.41823 1.4597 1.4555 16.0115 144.9159 0.00043594 -84.3165 0.16695
7.271 0.98812 5.4747e-005 3.8183 0.011941 9.4709e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4772 0.52566 0.16078 0.019004 13.9832 0.11803 0.00015267 0.77212 0.0089721 0.0099443 0.0017287 0.9823 0.98645 3.7793e-006 1.5118e-005 0.16154 0.62562 0.73316 0.0015689 0.7257 0.37277 0.0021068 0.41823 1.4619 1.4577 16.0115 144.9159 0.00043461 -84.3267 0.16795
7.272 0.98812 5.4747e-005 3.8183 0.011941 9.4722e-005 0.0011687 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4773 0.52571 0.1608 0.019005 13.9859 0.11804 0.00015268 0.77212 0.0089726 0.0099447 0.0017258 0.98235 0.9866 3.7725e-006 1.5091e-005 0.16154 0.62673 0.73417 0.0015675 0.72724 0.37297 0.002105 0.41824 1.4641 1.4599 16.0116 144.9159 0.00043329 -84.3368 0.16895
7.273 0.98812 5.4747e-005 3.8183 0.011941 9.4735e-005 0.0011687 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4773 0.52575 0.16081 0.019006 13.9886 0.11804 0.00015269 0.77211 0.008973 0.0099452 0.0017229 0.98239 0.98674 3.7658e-006 1.5064e-005 0.16154 0.62784 0.73518 0.0015661 0.72877 0.37318 0.0021032 0.41824 1.4662 1.4621 16.0117 144.9159 0.00043197 -84.3468 0.16995
7.274 0.98812 5.4747e-005 3.8183 0.011941 9.4747e-005 0.0011687 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4774 0.5258 0.16083 0.019007 13.9913 0.11805 0.0001527 0.7721 0.0089735 0.0099457 0.0017201 0.98243 0.98688 3.7592e-006 1.5038e-005 0.16155 0.62894 0.73617 0.0015647 0.73029 0.37339 0.0021014 0.41824 1.4684 1.4642 16.0117 144.916 0.00043066 -84.3567 0.17095
7.275 0.98812 5.4746e-005 3.8183 0.011941 9.476e-005 0.0011687 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4775 0.52584 0.16084 0.019008 13.994 0.11806 0.00015271 0.77209 0.0089739 0.0099461 0.0017172 0.98247 0.98701 3.7526e-006 1.5011e-005 0.16155 0.63004 0.73716 0.0015634 0.73181 0.3736 0.0020997 0.41825 1.4705 1.4664 16.0118 144.916 0.00042936 -84.3666 0.17195
7.276 0.98812 5.4746e-005 3.8183 0.01194 9.4773e-005 0.0011687 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.4776 0.52589 0.16085 0.01901 13.9967 0.11807 0.00015272 0.77209 0.0089743 0.0099466 0.0017144 0.98251 0.98714 3.7461e-006 1.4985e-005 0.16155 0.63114 0.73815 0.001562 0.73332 0.37381 0.0020979 0.41825 1.4727 1.4686 16.0119 144.916 0.00042806 -84.3764 0.17295
7.277 0.98812 5.4746e-005 3.8183 0.01194 9.4786e-005 0.0011687 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4777 0.52593 0.16087 0.019011 13.9994 0.11807 0.00015273 0.77208 0.0089748 0.0099471 0.0017117 0.98255 0.98726 3.7397e-006 1.4959e-005 0.16156 0.63223 0.73912 0.0015607 0.73483 0.37402 0.0020962 0.41825 1.4748 1.4707 16.0119 144.916 0.00042677 -84.3861 0.17395
7.278 0.98812 5.4746e-005 3.8183 0.01194 9.4799e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4778 0.52598 0.16088 0.019012 14.0021 0.11808 0.00015274 0.77207 0.0089752 0.0099476 0.0017089 0.98258 0.98737 3.7333e-006 1.4934e-005 0.16156 0.63332 0.74009 0.0015594 0.73632 0.37423 0.0020945 0.41825 1.477 1.4729 16.012 144.916 0.00042549 -84.3957 0.17495
7.279 0.98812 5.4746e-005 3.8183 0.01194 9.4812e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4779 0.52602 0.1609 0.019013 14.0048 0.11809 0.00015275 0.77207 0.0089757 0.009948 0.0017062 0.98262 0.98748 3.727e-006 1.4909e-005 0.16156 0.63441 0.74105 0.0015581 0.73781 0.37444 0.0020928 0.41826 1.4791 1.475 16.0121 144.916 0.00042421 -84.4053 0.17595
7.28 0.98812 5.4746e-005 3.8183 0.01194 9.4825e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.478 0.52607 0.16091 0.019014 14.0075 0.11809 0.00015276 0.77206 0.0089761 0.0099485 0.0017036 0.98266 0.98758 3.7208e-006 1.4884e-005 0.16157 0.63549 0.74201 0.0015568 0.73929 0.37465 0.0020911 0.41826 1.4812 1.4772 16.0121 144.916 0.00042295 -84.4147 0.17695
7.281 0.98812 5.4746e-005 3.8183 0.01194 9.4837e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4781 0.52612 0.16093 0.019016 14.0102 0.1181 0.00015277 0.77205 0.0089765 0.009949 0.0017009 0.9827 0.98768 3.7147e-006 1.4859e-005 0.16157 0.63657 0.74296 0.0015555 0.74077 0.37486 0.0020894 0.41827 1.4834 1.4793 16.0122 144.916 0.00042168 -84.4241 0.17795
7.282 0.98812 5.4746e-005 3.8183 0.01194 9.485e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4781 0.52616 0.16094 0.019017 14.0129 0.11811 0.00015278 0.77204 0.008977 0.0099494 0.0016983 0.98274 0.98777 3.7086e-006 1.4835e-005 0.16157 0.63765 0.7439 0.0015543 0.74224 0.37507 0.0020878 0.41827 1.4855 1.4815 16.0123 144.916 0.00042043 -84.4335 0.17895
7.283 0.98812 5.4746e-005 3.8183 0.01194 9.4863e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4782 0.52621 0.16095 0.019018 14.0156 0.11812 0.0001528 0.77204 0.0089774 0.0099499 0.0016957 0.98277 0.98786 3.7025e-006 1.4811e-005 0.16158 0.63872 0.74483 0.001553 0.7437 0.37528 0.0020861 0.41827 1.4876 1.4836 16.0123 144.9161 0.00041918 -84.4427 0.17995
7.284 0.98812 5.4746e-005 3.8183 0.01194 9.4876e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4783 0.52625 0.16097 0.019019 14.0183 0.11812 0.00015281 0.77203 0.0089779 0.0099504 0.0016931 0.98281 0.98795 3.6964e-006 1.4786e-005 0.16158 0.63979 0.74576 0.0015518 0.74515 0.37549 0.0020845 0.41828 1.4897 1.4857 16.0124 144.9161 0.00041793 -84.4519 0.18095
7.285 0.98812 5.4746e-005 3.8183 0.01194 9.4889e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4784 0.5263 0.16098 0.01902 14.021 0.11813 0.00015282 0.77202 0.0089783 0.0099508 0.0016904 0.98284 0.98803 3.6904e-006 1.4762e-005 0.16158 0.64086 0.74668 0.0015505 0.7466 0.3757 0.0020829 0.41828 1.4918 1.4878 16.0125 144.9161 0.0004167 -84.461 0.18195
7.286 0.98812 5.4746e-005 3.8183 0.01194 9.4902e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4785 0.52634 0.161 0.019022 14.0237 0.11814 0.00015283 0.77201 0.0089787 0.0099513 0.0016879 0.98288 0.9881 3.6844e-006 1.4738e-005 0.16159 0.64192 0.7476 0.0015493 0.74804 0.3759 0.0020813 0.41828 1.4939 1.49 16.0125 144.9161 0.00041547 -84.47 0.18295
7.287 0.98812 5.4746e-005 3.8183 0.01194 9.4915e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4786 0.52639 0.16101 0.019023 14.0264 0.11815 0.00015284 0.77201 0.0089792 0.0099518 0.0016853 0.98292 0.98818 3.6786e-006 1.4715e-005 0.16159 0.64298 0.74851 0.0015481 0.74947 0.37611 0.0020797 0.41829 1.496 1.4921 16.0126 144.9161 0.00041424 -84.479 0.18395
7.288 0.98812 5.4745e-005 3.8183 0.01194 9.4927e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4787 0.52643 0.16102 0.019024 14.0291 0.11815 0.00015285 0.772 0.0089796 0.0099523 0.0016829 0.98295 0.98825 3.6728e-006 1.4692e-005 0.16159 0.64404 0.74941 0.0015469 0.7509 0.37632 0.0020781 0.41829 1.4981 1.4942 16.0126 144.9161 0.00041303 -84.4879 0.18495
7.289 0.98812 5.4745e-005 3.8183 0.01194 9.494e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4788 0.52648 0.16104 0.019025 14.0318 0.11816 0.00015286 0.77199 0.0089801 0.0099527 0.0016805 0.98299 0.98832 3.6672e-006 1.4669e-005 0.1616 0.64509 0.75031 0.0015457 0.75232 0.37653 0.0020765 0.4183 1.5002 1.4963 16.0127 144.9161 0.00041181 -84.4967 0.18595
7.29 0.98812 5.4745e-005 3.8183 0.01194 9.4953e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4789 0.52652 0.16105 0.019026 14.0345 0.11817 0.00015287 0.77199 0.0089805 0.0099532 0.0016782 0.98302 0.98839 3.6617e-006 1.4647e-005 0.1616 0.64614 0.7512 0.0015445 0.75373 0.37674 0.002075 0.4183 1.5023 1.4984 16.0128 144.9161 0.00041061 -84.5054 0.18695
7.291 0.98812 5.4745e-005 3.8183 0.01194 9.4966e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4789 0.52657 0.16107 0.019028 14.0372 0.11817 0.00015288 0.77198 0.0089809 0.0099537 0.0016759 0.98305 0.98845 3.6562e-006 1.4625e-005 0.1616 0.64719 0.75209 0.0015434 0.75514 0.37695 0.0020735 0.41831 1.5044 1.5005 16.0128 144.9161 0.00040941 -84.5141 0.18795
7.292 0.98812 5.4745e-005 3.8183 0.01194 9.4979e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.479 0.52661 0.16108 0.019029 14.0399 0.11818 0.00015289 0.77197 0.0089814 0.0099541 0.0016735 0.98309 0.98851 3.6507e-006 1.4603e-005 0.16161 0.64823 0.75296 0.0015422 0.75654 0.37716 0.002072 0.41831 1.5065 1.5026 16.0129 144.9162 0.00040822 -84.5227 0.18895
7.293 0.98812 5.4745e-005 3.8183 0.01194 9.4992e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4791 0.52666 0.16109 0.01903 14.0426 0.11819 0.0001529 0.77196 0.0089818 0.0099546 0.0016711 0.98312 0.98857 3.6452e-006 1.4581e-005 0.16161 0.64927 0.75384 0.0015411 0.75793 0.37737 0.0020704 0.41832 1.5085 1.5047 16.0129 144.9162 0.00040703 -84.5313 0.18995
7.294 0.98812 5.4745e-005 3.8183 0.01194 9.5005e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4792 0.52671 0.16111 0.019031 14.0453 0.1182 0.00015291 0.77196 0.0089823 0.0099551 0.0016687 0.98315 0.98862 3.6396e-006 1.4559e-005 0.16161 0.65031 0.7547 0.0015399 0.75931 0.37758 0.002069 0.41832 1.5106 1.5068 16.013 144.9162 0.00040585 -84.5398 0.19095
7.295 0.98812 5.4745e-005 3.8183 0.01194 9.5017e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4793 0.52675 0.16112 0.019032 14.048 0.1182 0.00015292 0.77195 0.0089827 0.0099555 0.0016663 0.98319 0.98868 3.6341e-006 1.4537e-005 0.16162 0.65135 0.75556 0.0015388 0.76069 0.37779 0.0020675 0.41833 1.5127 1.5088 16.0131 144.9162 0.00040468 -84.5482 0.19195
7.296 0.98812 5.4745e-005 3.8183 0.01194 9.503e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4794 0.5268 0.16114 0.019034 14.0507 0.11821 0.00015294 0.77194 0.0089831 0.009956 0.0016639 0.98322 0.98873 3.6286e-006 1.4515e-005 0.16162 0.65238 0.75642 0.0015376 0.76206 0.378 0.002066 0.41833 1.5147 1.5109 16.0131 144.9162 0.00040351 -84.5565 0.19295
7.297 0.98812 5.4745e-005 3.8183 0.01194 9.5043e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4795 0.52684 0.16115 0.019035 14.0534 0.11822 0.00015295 0.77194 0.0089836 0.0099565 0.0016616 0.98325 0.98878 3.6233e-006 1.4494e-005 0.16162 0.65341 0.75727 0.0015365 0.76343 0.37821 0.0020645 0.41834 1.5168 1.513 16.0132 144.9162 0.00040235 -84.5648 0.19395
7.298 0.98812 5.4745e-005 3.8183 0.01194 9.5056e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4796 0.52689 0.16116 0.019036 14.0561 0.11822 0.00015296 0.77193 0.008984 0.0099569 0.0016593 0.98328 0.98882 3.618e-006 1.4473e-005 0.16163 0.65443 0.75811 0.0015354 0.76479 0.37841 0.0020631 0.41834 1.5189 1.515 16.0132 144.9162 0.00040119 -84.573 0.19495
7.299 0.98812 5.4745e-005 3.8183 0.01194 9.5069e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4797 0.52693 0.16118 0.019037 14.0588 0.11823 0.00015297 0.77192 0.0089844 0.0099574 0.001657 0.98331 0.98887 3.6127e-006 1.4452e-005 0.16163 0.65545 0.75895 0.0015343 0.76614 0.37862 0.0020617 0.41835 1.5209 1.5171 16.0133 144.9162 0.00040004 -84.5812 0.19595
7.3 0.98812 5.4744e-005 3.8183 0.01194 9.5082e-005 0.0011688 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4797 0.52698 0.16119 0.019038 14.0615 0.11824 0.00015298 0.77191 0.0089849 0.0099579 0.0016548 0.98334 0.98891 3.6076e-006 1.4431e-005 0.16163 0.65647 0.75978 0.0015332 0.76748 0.37883 0.0020602 0.41835 1.5229 1.5192 16.0133 144.9163 0.0003989 -84.5892 0.19695
7.301 0.98812 5.4744e-005 3.8183 0.01194 9.5095e-005 0.0011689 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4798 0.52702 0.16121 0.01904 14.0642 0.11825 0.00015299 0.77191 0.0089853 0.0099584 0.0016525 0.98337 0.98896 3.6025e-006 1.441e-005 0.16164 0.65749 0.76061 0.0015321 0.76882 0.37904 0.0020588 0.41836 1.525 1.5212 16.0134 144.9163 0.00039776 -84.5973 0.19795
7.302 0.98812 5.4744e-005 3.8183 0.01194 9.5107e-005 0.0011689 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.4799 0.52707 0.16122 0.019041 14.0669 0.11825 0.000153 0.7719 0.0089858 0.0099588 0.0016503 0.9834 0.989 3.5974e-006 1.439e-005 0.16164 0.6585 0.76143 0.0015311 0.77015 0.37925 0.0020574 0.41836 1.527 1.5233 16.0134 144.9163 0.00039663 -84.6052 0.19895
7.303 0.98812 5.4744e-005 3.8183 0.01194 9.512e-005 0.0011689 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.48 0.52711 0.16124 0.019042 14.0696 0.11826 0.00015301 0.77189 0.0089862 0.0099593 0.0016482 0.98344 0.98904 3.5924e-006 1.437e-005 0.16164 0.65951 0.76225 0.00153 0.77148 0.37946 0.0020561 0.41837 1.529 1.5253 16.0135 144.9163 0.0003955 -84.6131 0.19995
7.304 0.98812 5.4744e-005 3.8183 0.01194 9.5133e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4801 0.52716 0.16125 0.019043 14.0723 0.11827 0.00015302 0.77188 0.0089866 0.0099598 0.0016461 0.98346 0.98908 3.5874e-006 1.435e-005 0.16165 0.66052 0.76306 0.001529 0.77279 0.37967 0.0020547 0.41837 1.5311 1.5273 16.0136 144.9163 0.00039438 -84.621 0.20095
7.305 0.98812 5.4744e-005 3.8183 0.01194 9.5146e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4802 0.52721 0.16126 0.019044 14.075 0.11828 0.00015303 0.77188 0.0089871 0.0099602 0.001644 0.98349 0.98911 3.5825e-006 1.4331e-005 0.16165 0.66152 0.76387 0.0015279 0.7741 0.37988 0.0020533 0.41838 1.5331 1.5294 16.0136 144.9163 0.00039326 -84.6287 0.20195
7.306 0.98812 5.4744e-005 3.8183 0.01194 9.5159e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4803 0.52725 0.16128 0.019046 14.0777 0.11828 0.00015304 0.77187 0.0089875 0.0099607 0.0016419 0.98352 0.98915 3.5777e-006 1.4311e-005 0.16166 0.66252 0.76467 0.0015269 0.77541 0.38009 0.002052 0.41839 1.5351 1.5314 16.0137 144.9163 0.00039215 -84.6365 0.20295
7.307 0.98812 5.4744e-005 3.8183 0.01194 9.5172e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4804 0.5273 0.16129 0.019047 14.0804 0.11829 0.00015305 0.77186 0.008988 0.0099612 0.0016398 0.98355 0.98919 3.5728e-006 1.4292e-005 0.16166 0.66352 0.76546 0.0015259 0.77671 0.3803 0.0020507 0.41839 1.5371 1.5334 16.0137 144.9163 0.00039105 -84.6441 0.20395
7.308 0.98812 5.4744e-005 3.8183 0.01194 9.5185e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4804 0.52734 0.16131 0.019048 14.0832 0.1183 0.00015306 0.77186 0.0089884 0.0099616 0.0016378 0.98358 0.98922 3.568e-006 1.4273e-005 0.16166 0.66451 0.76625 0.0015249 0.778 0.3805 0.0020493 0.4184 1.5391 1.5354 16.0138 144.9164 0.00038995 -84.6517 0.20495
7.309 0.98812 5.4744e-005 3.8183 0.01194 9.5197e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4805 0.52739 0.16132 0.019049 14.0859 0.1183 0.00015308 0.77185 0.0089888 0.0099621 0.0016357 0.98361 0.98925 3.5633e-006 1.4254e-005 0.16167 0.6655 0.76704 0.0015239 0.77928 0.38071 0.002048 0.4184 1.5411 1.5375 16.0138 144.9164 0.00038886 -84.6592 0.20595
7.31 0.98812 5.4744e-005 3.8183 0.01194 9.521e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4806 0.52743 0.16133 0.01905 14.0886 0.11831 0.00015309 0.77184 0.0089893 0.0099626 0.0016337 0.98364 0.98928 3.5585e-006 1.4235e-005 0.16167 0.66649 0.76782 0.0015229 0.78056 0.38092 0.0020467 0.41841 1.5431 1.5395 16.0139 144.9164 0.00038777 -84.6667 0.20695
7.311 0.98812 5.4744e-005 3.8183 0.01194 9.5223e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4807 0.52748 0.16135 0.019052 14.0913 0.11832 0.0001531 0.77183 0.0089897 0.009963 0.0016316 0.98367 0.98931 3.5539e-006 1.4216e-005 0.16167 0.66748 0.76859 0.0015219 0.78183 0.38113 0.0020454 0.41842 1.5451 1.5415 16.0139 144.9164 0.00038669 -84.6741 0.20795
7.312 0.98812 5.4744e-005 3.8183 0.01194 9.5236e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4808 0.52752 0.16136 0.019053 14.094 0.11833 0.00015311 0.77183 0.0089901 0.0099635 0.0016296 0.98369 0.98934 3.5492e-006 1.4197e-005 0.16168 0.66846 0.76936 0.0015209 0.7831 0.38134 0.0020441 0.41842 1.5471 1.5435 16.014 144.9164 0.00038561 -84.6815 0.20895
7.313 0.98812 5.4743e-005 3.8183 0.01194 9.5249e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4809 0.52757 0.16138 0.019054 14.0967 0.11833 0.00015312 0.77182 0.0089906 0.009964 0.0016277 0.98372 0.98937 3.5446e-006 1.4179e-005 0.16168 0.66944 0.77012 0.0015199 0.78436 0.38155 0.0020429 0.41843 1.5491 1.5455 16.014 144.9164 0.00038454 -84.6888 0.20995
7.314 0.98812 5.4743e-005 3.8183 0.01194 9.5262e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.481 0.52761 0.16139 0.019055 14.0994 0.11834 0.00015313 0.77181 0.008991 0.0099644 0.0016257 0.98375 0.9894 3.5401e-006 1.4161e-005 0.16168 0.67041 0.77088 0.001519 0.78561 0.38176 0.0020416 0.41844 1.5511 1.5475 16.0141 144.9164 0.00038347 -84.696 0.21095
7.315 0.98812 5.4743e-005 3.8183 0.01194 9.5275e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4811 0.52766 0.1614 0.019056 14.1021 0.11835 0.00015314 0.77181 0.0089915 0.0099649 0.0016237 0.98377 0.98943 3.5356e-006 1.4143e-005 0.16169 0.67138 0.77164 0.001518 0.78686 0.38197 0.0020404 0.41844 1.5531 1.5495 16.0141 144.9164 0.00038241 -84.7032 0.21195
7.316 0.98812 5.4743e-005 3.8183 0.01194 9.5287e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4812 0.52771 0.16142 0.019057 14.1048 0.11835 0.00015315 0.7718 0.0089919 0.0099654 0.0016218 0.9838 0.98946 3.5311e-006 1.4125e-005 0.16169 0.67235 0.77239 0.0015171 0.78809 0.38217 0.0020391 0.41845 1.555 1.5515 16.0142 144.9165 0.00038136 -84.7104 0.21295
7.317 0.98812 5.4743e-005 3.8183 0.01194 9.53e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4812 0.52775 0.16143 0.019059 14.1075 0.11836 0.00015316 0.77179 0.0089923 0.0099658 0.0016199 0.98383 0.98948 3.5267e-006 1.4107e-005 0.16169 0.67332 0.77314 0.0015161 0.78933 0.38238 0.0020379 0.41846 1.557 1.5534 16.0142 144.9165 0.00038031 -84.7174 0.21395
7.318 0.98812 5.4743e-005 3.8183 0.01194 9.5313e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4813 0.5278 0.16145 0.01906 14.1103 0.11837 0.00015317 0.77178 0.0089928 0.0099663 0.001618 0.98385 0.98951 3.5223e-006 1.409e-005 0.1617 0.67429 0.77388 0.0015152 0.79055 0.38259 0.0020367 0.41846 1.559 1.5554 16.0143 144.9165 0.00037926 -84.7245 0.21495
7.319 0.98812 5.4743e-005 3.8183 0.01194 9.5326e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4814 0.52784 0.16146 0.019061 14.113 0.11838 0.00015318 0.77178 0.0089932 0.0099668 0.0016161 0.98388 0.98953 3.518e-006 1.4072e-005 0.1617 0.67525 0.77461 0.0015143 0.79177 0.3828 0.0020355 0.41847 1.5609 1.5574 16.0143 144.9165 0.00037822 -84.7314 0.21595
7.32 0.98812 5.4743e-005 3.8183 0.01194 9.5339e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4815 0.52789 0.16147 0.019062 14.1157 0.11838 0.00015319 0.77177 0.0089936 0.0099672 0.0016143 0.98391 0.98956 3.5137e-006 1.4055e-005 0.1617 0.6762 0.77534 0.0015133 0.79299 0.38301 0.0020343 0.41848 1.5629 1.5593 16.0144 144.9165 0.00037719 -84.7384 0.21695
7.321 0.98812 5.4743e-005 3.8183 0.01194 9.5352e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4816 0.52793 0.16149 0.019063 14.1184 0.11839 0.0001532 0.77176 0.0089941 0.0099677 0.0016124 0.98393 0.98958 3.5094e-006 1.4038e-005 0.16171 0.67716 0.77607 0.0015124 0.7942 0.38322 0.0020331 0.41849 1.5648 1.5613 16.0144 144.9165 0.00037616 -84.7452 0.21795
7.322 0.98812 5.4743e-005 3.8183 0.01194 9.5365e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4817 0.52798 0.1615 0.019065 14.1211 0.1184 0.00015322 0.77176 0.0089945 0.0099682 0.0016106 0.98396 0.98961 3.5052e-006 1.4021e-005 0.16171 0.67811 0.77679 0.0015115 0.7954 0.38343 0.0020319 0.41849 1.5668 1.5633 16.0145 144.9165 0.00037514 -84.752 0.21895
7.323 0.98812 5.4743e-005 3.8183 0.01194 9.5377e-005 0.0011689 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4818 0.52802 0.16152 0.019066 14.1238 0.11841 0.00015323 0.77175 0.008995 0.0099686 0.0016088 0.98398 0.98963 3.501e-006 1.4004e-005 0.16171 0.67906 0.77751 0.0015106 0.79659 0.38364 0.0020307 0.4185 1.5687 1.5652 16.0145 144.9166 0.00037412 -84.7588 0.21995
7.324 0.98812 5.4743e-005 3.8183 0.01194 9.539e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4819 0.52807 0.16153 0.019067 14.1265 0.11841 0.00015324 0.77174 0.0089954 0.0099691 0.001607 0.98401 0.98965 3.4969e-006 1.3988e-005 0.16172 0.68001 0.77823 0.0015098 0.79778 0.38384 0.0020296 0.41851 1.5707 1.5672 16.0146 144.9166 0.00037311 -84.7655 0.22095
7.325 0.98812 5.4742e-005 3.8183 0.01194 9.5403e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.482 0.52811 0.16154 0.019068 14.1292 0.11842 0.00015325 0.77173 0.0089958 0.0099696 0.0016052 0.98403 0.98967 3.4927e-006 1.3971e-005 0.16172 0.68095 0.77893 0.0015089 0.79896 0.38405 0.0020284 0.41851 1.5726 1.5691 16.0146 144.9166 0.0003721 -84.7721 0.22195
7.326 0.98812 5.4742e-005 3.8183 0.01194 9.5416e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.482 0.52816 0.16156 0.019069 14.132 0.11843 0.00015326 0.77173 0.0089963 0.00997 0.0016035 0.98405 0.98969 3.4887e-006 1.3955e-005 0.16172 0.68189 0.77964 0.001508 0.80014 0.38426 0.0020273 0.41852 1.5745 1.5711 16.0147 144.9166 0.0003711 -84.7787 0.22295
7.327 0.98812 5.4742e-005 3.8183 0.01194 9.5429e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4821 0.5282 0.16157 0.019071 14.1347 0.11843 0.00015327 0.77172 0.0089967 0.0099705 0.0016017 0.98408 0.98971 3.4846e-006 1.3939e-005 0.16173 0.68283 0.78034 0.0015071 0.80131 0.38447 0.0020262 0.41853 1.5764 1.573 16.0147 144.9166 0.0003701 -84.7853 0.22395
7.328 0.98812 5.4742e-005 3.8183 0.01194 9.5442e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4822 0.52825 0.16159 0.019072 14.1374 0.11844 0.00015328 0.77171 0.0089971 0.009971 0.0016 0.9841 0.98974 3.4806e-006 1.3923e-005 0.16173 0.68376 0.78104 0.0015063 0.80248 0.38468 0.002025 0.41854 1.5784 1.5749 16.0147 144.9166 0.0003691 -84.7918 0.22495
7.329 0.98812 5.4742e-005 3.8183 0.01194 9.5455e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4823 0.5283 0.1616 0.019073 14.1401 0.11845 0.00015329 0.7717 0.0089976 0.0099714 0.0015983 0.98413 0.98976 3.4767e-006 1.3907e-005 0.16173 0.68469 0.78173 0.0015054 0.80363 0.38489 0.0020239 0.41854 1.5803 1.5768 16.0148 144.9166 0.00036812 -84.7982 0.22595
7.33 0.98812 5.4742e-005 3.8183 0.01194 9.5467e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4824 0.52834 0.16162 0.019074 14.1428 0.11846 0.0001533 0.7717 0.008998 0.0099719 0.0015966 0.98415 0.98978 3.4727e-006 1.3891e-005 0.16174 0.68562 0.78242 0.0015046 0.80479 0.38509 0.0020228 0.41855 1.5822 1.5788 16.0148 144.9167 0.00036713 -84.8046 0.22695
7.331 0.98812 5.4742e-005 3.8183 0.01194 9.548e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4825 0.52839 0.16163 0.019075 14.1455 0.11846 0.00015331 0.77169 0.0089984 0.0099724 0.0015949 0.98417 0.98979 3.4688e-006 1.3876e-005 0.16174 0.68655 0.7831 0.0015038 0.80593 0.3853 0.0020217 0.41856 1.5841 1.5807 16.0149 144.9167 0.00036615 -84.811 0.22795
7.332 0.98812 5.4742e-005 3.8183 0.01194 9.5493e-005 0.001169 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4826 0.52843 0.16164 0.019077 14.1482 0.11847 0.00015332 0.77168 0.0089989 0.0099728 0.0015932 0.98419 0.98981 3.465e-006 1.386e-005 0.16174 0.68747 0.78378 0.0015029 0.80707 0.38551 0.0020206 0.41857 1.586 1.5826 16.0149 144.9167 0.00036518 -84.8173 0.22895
7.333 0.98812 5.4742e-005 3.8183 0.01194 9.5506e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4827 0.52848 0.16166 0.019078 14.151 0.11848 0.00015333 0.77168 0.0089993 0.0099733 0.0015915 0.98422 0.98983 3.4611e-006 1.3845e-005 0.16175 0.68839 0.78445 0.0015021 0.8082 0.38572 0.0020196 0.41858 1.5879 1.5845 16.015 144.9167 0.00036421 -84.8235 0.22995
7.334 0.98812 5.4742e-005 3.8183 0.011939 9.5519e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4828 0.52852 0.16167 0.019079 14.1537 0.11848 0.00015334 0.77167 0.0089998 0.0099738 0.0015899 0.98424 0.98985 3.4573e-006 1.383e-005 0.16175 0.68931 0.78513 0.0015013 0.80933 0.38593 0.0020185 0.41858 1.5898 1.5864 16.015 144.9167 0.00036325 -84.8298 0.23095
7.335 0.98812 5.4742e-005 3.8183 0.011939 9.5532e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4828 0.52857 0.16169 0.01908 14.1564 0.11849 0.00015335 0.77166 0.0090002 0.0099742 0.0015883 0.98426 0.98987 3.4535e-006 1.3815e-005 0.16175 0.69023 0.78579 0.0015005 0.81045 0.38614 0.0020174 0.41859 1.5917 1.5883 16.0151 144.9167 0.00036229 -84.8359 0.23195
7.336 0.98812 5.4742e-005 3.8183 0.011939 9.5545e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4829 0.52861 0.1617 0.019081 14.1591 0.1185 0.00015337 0.77165 0.0090006 0.0099747 0.0015867 0.98428 0.98989 3.4498e-006 1.38e-005 0.16176 0.69114 0.78646 0.0014997 0.81157 0.38634 0.0020164 0.4186 1.5935 1.5902 16.0151 144.9167 0.00036133 -84.842 0.23295
7.337 0.98812 5.4741e-005 3.8183 0.011939 9.5557e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.483 0.52866 0.16171 0.019083 14.1618 0.11851 0.00015338 0.77165 0.0090011 0.0099752 0.0015851 0.98431 0.9899 3.4461e-006 1.3785e-005 0.16176 0.69205 0.78712 0.0014989 0.81268 0.38655 0.0020154 0.41861 1.5954 1.5921 16.0151 144.9168 0.00036038 -84.8481 0.23395
7.338 0.98812 5.4741e-005 3.8183 0.011939 9.557e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4831 0.5287 0.16173 0.019084 14.1646 0.11851 0.00015339 0.77164 0.0090015 0.0099756 0.0015835 0.98433 0.98992 3.4424e-006 1.377e-005 0.16176 0.69295 0.78777 0.0014981 0.81378 0.38676 0.0020143 0.41862 1.5973 1.594 16.0152 144.9168 0.00035944 -84.8541 0.23495
7.339 0.98812 5.4741e-005 3.8183 0.011939 9.5583e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4832 0.52875 0.16174 0.019085 14.1673 0.11852 0.0001534 0.77163 0.0090019 0.0099761 0.0015819 0.98435 0.98994 3.4388e-006 1.3756e-005 0.16177 0.69386 0.78842 0.0014973 0.81488 0.38697 0.0020133 0.41863 1.5992 1.5959 16.0152 144.9168 0.0003585 -84.8601 0.23595
7.34 0.98812 5.4741e-005 3.8183 0.011939 9.5596e-005 0.001169 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.4833 0.5288 0.16176 0.019086 14.17 0.11853 0.00015341 0.77163 0.0090024 0.0099766 0.0015803 0.98437 0.98995 3.4352e-006 1.3741e-005 0.16177 0.69476 0.78907 0.0014965 0.81597 0.38718 0.0020123 0.41863 1.601 1.5977 16.0153 144.9168 0.00035756 -84.866 0.23695
7.341 0.98812 5.4741e-005 3.8183 0.011939 9.5609e-005 0.001169 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4834 0.52884 0.16177 0.019087 14.1727 0.11853 0.00015342 0.77162 0.0090028 0.009977 0.0015788 0.98439 0.98997 3.4316e-006 1.3727e-005 0.16177 0.69565 0.78971 0.0014958 0.81706 0.38739 0.0020113 0.41864 1.6029 1.5996 16.0153 144.9168 0.00035663 -84.8719 0.23795
7.342 0.98812 5.4741e-005 3.8183 0.011939 9.5622e-005 0.001169 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4835 0.52889 0.16178 0.019089 14.1754 0.11854 0.00015343 0.77161 0.0090032 0.0099775 0.0015772 0.98441 0.98999 3.4281e-006 1.3713e-005 0.16178 0.69655 0.79035 0.001495 0.81814 0.38759 0.0020103 0.41865 1.6048 1.6015 16.0153 144.9168 0.00035571 -84.8777 0.23895
7.343 0.98812 5.4741e-005 3.8183 0.011939 9.5635e-005 0.001169 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4836 0.52893 0.1618 0.01909 14.1781 0.11855 0.00015344 0.7716 0.0090037 0.009978 0.0015757 0.98443 0.99 3.4246e-006 1.3699e-005 0.16178 0.69744 0.79099 0.0014942 0.81921 0.3878 0.0020093 0.41866 1.6066 1.6033 16.0154 144.9168 0.00035478 -84.8835 0.23995
7.344 0.98812 5.4741e-005 3.8183 0.011939 9.5647e-005 0.001169 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4836 0.52898 0.16181 0.019091 14.1809 0.11856 0.00015345 0.7716 0.0090041 0.0099784 0.0015742 0.98445 0.99002 3.4211e-006 1.3685e-005 0.16178 0.69833 0.79162 0.0014935 0.82028 0.38801 0.0020083 0.41867 1.6085 1.6052 16.0154 144.9169 0.00035387 -84.8892 0.24095
7.345 0.98812 5.4741e-005 3.8183 0.011939 9.566e-005 0.001169 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4837 0.52902 0.16183 0.019092 14.1836 0.11856 0.00015346 0.77159 0.0090046 0.0099789 0.0015727 0.98447 0.99003 3.4176e-006 1.3671e-005 0.16179 0.69922 0.79225 0.0014928 0.82134 0.38822 0.0020073 0.41868 1.6103 1.6071 16.0155 144.9169 0.00035295 -84.8949 0.24195
7.346 0.98812 5.4741e-005 3.8183 0.011939 9.5673e-005 0.001169 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4838 0.52907 0.16184 0.019093 14.1863 0.11857 0.00015347 0.77158 0.009005 0.0099794 0.0015713 0.98449 0.99005 3.4142e-006 1.3657e-005 0.16179 0.7001 0.79288 0.001492 0.8224 0.38843 0.0020064 0.41869 1.6121 1.6089 16.0155 144.9169 0.00035205 -84.9006 0.24295
7.347 0.98812 5.4741e-005 3.8183 0.011939 9.5686e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4839 0.52911 0.16185 0.019095 14.189 0.11858 0.00015348 0.77158 0.0090054 0.0099798 0.0015698 0.98451 0.99006 3.4108e-006 1.3644e-005 0.16179 0.70098 0.7935 0.0014913 0.82345 0.38863 0.0020054 0.41869 1.614 1.6107 16.0155 144.9169 0.00035114 -84.9062 0.24395
7.348 0.98812 5.4741e-005 3.8183 0.011939 9.5699e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.484 0.52916 0.16187 0.019096 14.1918 0.11858 0.00015349 0.77157 0.0090059 0.0099803 0.0015684 0.98453 0.99008 3.4075e-006 1.363e-005 0.1618 0.70186 0.79411 0.0014906 0.8245 0.38884 0.0020045 0.4187 1.6158 1.6126 16.0156 144.9169 0.00035024 -84.9118 0.24495
7.349 0.98812 5.4741e-005 3.8183 0.011939 9.5712e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4841 0.5292 0.16188 0.019097 14.1945 0.11859 0.00015351 0.77156 0.0090063 0.0099808 0.0015669 0.98455 0.99009 3.4041e-006 1.3617e-005 0.1618 0.70274 0.79473 0.0014899 0.82554 0.38905 0.0020035 0.41871 1.6176 1.6144 16.0156 144.9169 0.00034935 -84.9173 0.24595
7.35 0.98812 5.474e-005 3.8183 0.011939 9.5725e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4842 0.52925 0.1619 0.019098 14.1972 0.1186 0.00015352 0.77155 0.0090067 0.0099812 0.0015655 0.98457 0.99011 3.4008e-006 1.3604e-005 0.1618 0.70361 0.79534 0.0014891 0.82657 0.38926 0.0020026 0.41872 1.6194 1.6163 16.0157 144.9169 0.00034846 -84.9228 0.24695
7.351 0.98812 5.474e-005 3.8183 0.011939 9.5737e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4843 0.52929 0.16191 0.019099 14.1999 0.11861 0.00015353 0.77155 0.0090072 0.0099817 0.001564 0.98459 0.99012 3.3976e-006 1.3591e-005 0.16181 0.70448 0.79595 0.0014884 0.8276 0.38946 0.0020017 0.41873 1.6213 1.6181 16.0157 144.917 0.00034757 -84.9283 0.24795
7.352 0.98812 5.474e-005 3.8183 0.011939 9.575e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4843 0.52934 0.16192 0.019101 14.2026 0.11861 0.00015354 0.77154 0.0090076 0.0099822 0.0015626 0.98461 0.99014 3.3943e-006 1.3578e-005 0.16181 0.70535 0.79655 0.0014877 0.82862 0.38967 0.0020007 0.41874 1.6231 1.6199 16.0157 144.917 0.00034669 -84.9337 0.24895
7.353 0.98812 5.474e-005 3.8183 0.011939 9.5763e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4844 0.52939 0.16194 0.019102 14.2054 0.11862 0.00015355 0.77153 0.009008 0.0099826 0.0015612 0.98463 0.99015 3.3911e-006 1.3565e-005 0.16181 0.70622 0.79715 0.001487 0.82964 0.38988 0.0019998 0.41875 1.6249 1.6217 16.0158 144.917 0.00034581 -84.939 0.24995
7.354 0.98812 5.474e-005 3.8183 0.011939 9.5776e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4845 0.52943 0.16195 0.019103 14.2081 0.11863 0.00015356 0.77153 0.0090085 0.0099831 0.0015598 0.98465 0.99016 3.3879e-006 1.3552e-005 0.16182 0.70708 0.79775 0.0014863 0.83065 0.39009 0.0019989 0.41876 1.6267 1.6235 16.0158 144.917 0.00034494 -84.9443 0.25095
7.355 0.98812 5.474e-005 3.8183 0.011939 9.5789e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4846 0.52948 0.16197 0.019104 14.2108 0.11864 0.00015357 0.77152 0.0090089 0.0099835 0.0015585 0.98467 0.99018 3.3847e-006 1.3539e-005 0.16182 0.70794 0.79834 0.0014856 0.83166 0.3903 0.001998 0.41877 1.6285 1.6253 16.0158 144.917 0.00034407 -84.9496 0.25195
7.356 0.98812 5.474e-005 3.8183 0.011939 9.5802e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4847 0.52952 0.16198 0.019105 14.2135 0.11864 0.00015358 0.77151 0.0090093 0.009984 0.0015571 0.98469 0.99019 3.3816e-006 1.3527e-005 0.16182 0.7088 0.79893 0.0014849 0.83266 0.3905 0.0019971 0.41878 1.6303 1.6272 16.0159 144.917 0.0003432 -84.9549 0.25295
7.357 0.98812 5.474e-005 3.8183 0.011939 9.5815e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4848 0.52957 0.16199 0.019106 14.2163 0.11865 0.00015359 0.7715 0.0090098 0.0099845 0.0015558 0.9847 0.9902 3.3785e-006 1.3514e-005 0.16183 0.70965 0.79952 0.0014843 0.83366 0.39071 0.0019962 0.41879 1.6321 1.629 16.0159 144.917 0.00034234 -84.9601 0.25395
7.358 0.98812 5.474e-005 3.8183 0.011939 9.5827e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4849 0.52961 0.16201 0.019108 14.219 0.11866 0.0001536 0.7715 0.0090102 0.0099849 0.0015544 0.98472 0.99022 3.3754e-006 1.3502e-005 0.16183 0.7105 0.8001 0.0014836 0.83465 0.39092 0.0019954 0.4188 1.6339 1.6308 16.016 144.9171 0.00034149 -84.9652 0.25495
7.359 0.98812 5.474e-005 3.8183 0.011939 9.584e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.485 0.52966 0.16202 0.019109 14.2217 0.11866 0.00015361 0.77149 0.0090106 0.0099854 0.0015531 0.98474 0.99023 3.3724e-006 1.349e-005 0.16183 0.71135 0.80068 0.0014829 0.83563 0.39113 0.0019945 0.41881 1.6356 1.6325 16.016 144.9171 0.00034063 -84.9704 0.25595
7.36 0.98812 5.474e-005 3.8183 0.011939 9.5853e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4851 0.5297 0.16204 0.01911 14.2244 0.11867 0.00015362 0.77148 0.0090111 0.0099859 0.0015518 0.98476 0.99024 3.3693e-006 1.3478e-005 0.16184 0.7122 0.80126 0.0014823 0.83661 0.39133 0.0019936 0.41882 1.6374 1.6343 16.016 144.9171 0.00033979 -84.9754 0.25695
7.361 0.98812 5.474e-005 3.8183 0.011939 9.5866e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4851 0.52975 0.16205 0.019111 14.2272 0.11868 0.00015363 0.77148 0.0090115 0.0099863 0.0015505 0.98478 0.99025 3.3663e-006 1.3465e-005 0.16184 0.71304 0.80183 0.0014816 0.83758 0.39154 0.0019928 0.41882 1.6392 1.6361 16.0161 144.9171 0.00033894 -84.9805 0.25795
7.362 0.98812 5.4739e-005 3.8183 0.011939 9.5879e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4852 0.52979 0.16206 0.019112 14.2299 0.11869 0.00015364 0.77147 0.0090119 0.0099868 0.0015492 0.98479 0.99027 3.3633e-006 1.3454e-005 0.16184 0.71388 0.8024 0.001481 0.83855 0.39175 0.0019919 0.41883 1.6409 1.6379 16.0161 144.9171 0.0003381 -84.9855 0.25895
7.363 0.98812 5.4739e-005 3.8183 0.011939 9.5892e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4853 0.52984 0.16208 0.019114 14.2326 0.11869 0.00015365 0.77146 0.0090124 0.0099873 0.0015479 0.98481 0.99028 3.3604e-006 1.3442e-005 0.16185 0.71472 0.80297 0.0014803 0.83951 0.39196 0.0019911 0.41884 1.6427 1.6397 16.0161 144.9171 0.00033727 -84.9905 0.25995
7.364 0.98812 5.4739e-005 3.8183 0.011939 9.5905e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4854 0.52988 0.16209 0.019115 14.2353 0.1187 0.00015367 0.77145 0.0090128 0.0099877 0.0015466 0.98483 0.99029 3.3574e-006 1.343e-005 0.16185 0.71556 0.80353 0.0014797 0.84047 0.39216 0.0019903 0.41885 1.6445 1.6414 16.0162 144.9172 0.00033643 -84.9954 0.26095
7.365 0.98812 5.4739e-005 3.8183 0.011939 9.5917e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4855 0.52993 0.16211 0.019116 14.2381 0.11871 0.00015368 0.77145 0.0090132 0.0099882 0.0015454 0.98484 0.9903 3.3545e-006 1.3418e-005 0.16185 0.71639 0.80409 0.001479 0.84142 0.39237 0.0019894 0.41886 1.6462 1.6432 16.0162 144.9172 0.00033561 -85.0003 0.26195
7.366 0.98812 5.4739e-005 3.8183 0.011939 9.593e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4856 0.52998 0.16212 0.019117 14.2408 0.11871 0.00015369 0.77144 0.0090137 0.0099886 0.0015441 0.98486 0.99031 3.3517e-006 1.3407e-005 0.16186 0.71722 0.80465 0.0014784 0.84237 0.39258 0.0019886 0.41887 1.648 1.645 16.0162 144.9172 0.00033478 -85.0051 0.26295
7.367 0.98812 5.4739e-005 3.8183 0.011939 9.5943e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4857 0.53002 0.16214 0.019118 14.2435 0.11872 0.0001537 0.77143 0.0090141 0.0099891 0.0015429 0.98488 0.99033 3.3488e-006 1.3395e-005 0.16186 0.71805 0.8052 0.0014778 0.84331 0.39278 0.0019878 0.41888 1.6497 1.6467 16.0163 144.9172 0.00033396 -85.01 0.26395
7.368 0.98812 5.4739e-005 3.8183 0.011939 9.5956e-005 0.0011691 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.4858 0.53007 0.16215 0.01912 14.2463 0.11873 0.00015371 0.77143 0.0090145 0.0099896 0.0015416 0.98489 0.99034 3.346e-006 1.3384e-005 0.16186 0.71888 0.80575 0.0014772 0.84425 0.39299 0.001987 0.41889 1.6515 1.6485 16.0163 144.9172 0.00033315 -85.0148 0.26495
7.369 0.98812 5.4739e-005 3.8183 0.011939 9.5969e-005 0.0011691 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4859 0.53011 0.16216 0.019121 14.249 0.11874 0.00015372 0.77142 0.009015 0.00999 0.0015404 0.98491 0.99035 3.3431e-006 1.3373e-005 0.16187 0.7197 0.8063 0.0014765 0.84518 0.3932 0.0019862 0.4189 1.6532 1.6502 16.0163 144.9172 0.00033233 -85.0195 0.26595
7.37 0.98812 5.4739e-005 3.8183 0.011939 9.5982e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4859 0.53016 0.16218 0.019122 14.2517 0.11874 0.00015373 0.77141 0.0090154 0.0099905 0.0015392 0.98493 0.99036 3.3404e-006 1.3362e-005 0.16187 0.72052 0.80685 0.0014759 0.8461 0.39341 0.0019854 0.41891 1.6549 1.652 16.0164 144.9172 0.00033153 -85.0242 0.26695
7.371 0.98812 5.4739e-005 3.8183 0.011939 9.5995e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.486 0.5302 0.16219 0.019123 14.2544 0.11875 0.00015374 0.7714 0.0090159 0.009991 0.001538 0.98494 0.99037 3.3376e-006 1.3351e-005 0.16187 0.72134 0.80739 0.0014753 0.84702 0.39361 0.0019846 0.41892 1.6567 1.6537 16.0164 144.9173 0.00033072 -85.0289 0.26795
7.372 0.98812 5.4739e-005 3.8183 0.011939 9.6007e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4861 0.53025 0.16221 0.019124 14.2572 0.11876 0.00015375 0.7714 0.0090163 0.0099914 0.0015368 0.98496 0.99038 3.3349e-006 1.334e-005 0.16188 0.72216 0.80793 0.0014748 0.84794 0.39382 0.0019838 0.41893 1.6584 1.6554 16.0164 144.9173 0.00032992 -85.0335 0.26895
7.373 0.98812 5.4739e-005 3.8183 0.011939 9.602e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4862 0.53029 0.16222 0.019126 14.2599 0.11876 0.00015376 0.77139 0.0090167 0.0099919 0.0015357 0.98498 0.99039 3.3321e-006 1.3329e-005 0.16188 0.72297 0.80847 0.0014742 0.84885 0.39403 0.001983 0.41894 1.6601 1.6572 16.0165 144.9173 0.00032912 -85.0381 0.26995
7.374 0.98812 5.4739e-005 3.8183 0.011939 9.6033e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4863 0.53034 0.16223 0.019127 14.2626 0.11877 0.00015377 0.77138 0.0090172 0.0099924 0.0015345 0.98499 0.99041 3.3294e-006 1.3318e-005 0.16188 0.72378 0.809 0.0014736 0.84975 0.39423 0.0019823 0.41896 1.6618 1.6589 16.0165 144.9173 0.00032833 -85.0427 0.27095
7.375 0.98812 5.4738e-005 3.8183 0.011939 9.6046e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4864 0.53038 0.16225 0.019128 14.2654 0.11878 0.00015378 0.77138 0.0090176 0.0099928 0.0015333 0.98501 0.99042 3.3268e-006 1.3307e-005 0.16189 0.72459 0.80953 0.001473 0.85065 0.39444 0.0019815 0.41897 1.6635 1.6606 16.0165 144.9173 0.00032754 -85.0472 0.27195
7.376 0.98812 5.4738e-005 3.8183 0.011939 9.6059e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4865 0.53043 0.16226 0.019129 14.2681 0.11879 0.00015379 0.77137 0.009018 0.0099933 0.0015322 0.98502 0.99043 3.3241e-006 1.3297e-005 0.16189 0.7254 0.81006 0.0014724 0.85155 0.39465 0.0019807 0.41898 1.6652 1.6623 16.0165 144.9173 0.00032676 -85.0517 0.27295
7.377 0.98812 5.4738e-005 3.8183 0.011939 9.6072e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4866 0.53047 0.16228 0.01913 14.2708 0.11879 0.0001538 0.77136 0.0090185 0.0099937 0.0015311 0.98504 0.99044 3.3215e-006 1.3286e-005 0.16189 0.7262 0.81058 0.0014718 0.85244 0.39485 0.00198 0.41899 1.6669 1.664 16.0166 144.9174 0.00032598 -85.0562 0.27395
7.378 0.98812 5.4738e-005 3.8183 0.011939 9.6085e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4866 0.53052 0.16229 0.019131 14.2736 0.1188 0.00015382 0.77135 0.0090189 0.0099942 0.0015299 0.98505 0.99045 3.3189e-006 1.3276e-005 0.1619 0.727 0.8111 0.0014713 0.85332 0.39506 0.0019792 0.419 1.6686 1.6658 16.0166 144.9174 0.0003252 -85.0606 0.27495
7.379 0.98812 5.4738e-005 3.8183 0.011939 9.6097e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4867 0.53057 0.1623 0.019133 14.2763 0.11881 0.00015383 0.77135 0.0090193 0.0099947 0.0015288 0.98507 0.99046 3.3163e-006 1.3265e-005 0.1619 0.7278 0.81162 0.0014707 0.8542 0.39527 0.0019785 0.41901 1.6703 1.6675 16.0166 144.9174 0.00032443 -85.065 0.27595
7.38 0.98812 5.4738e-005 3.8183 0.011939 9.611e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4868 0.53061 0.16232 0.019134 14.279 0.11881 0.00015384 0.77134 0.0090198 0.0099951 0.0015277 0.98508 0.99047 3.3137e-006 1.3255e-005 0.1619 0.72859 0.81214 0.0014701 0.85508 0.39547 0.0019778 0.41902 1.672 1.6692 16.0167 144.9174 0.00032366 -85.0694 0.27695
7.381 0.98812 5.4738e-005 3.8183 0.011939 9.6123e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4869 0.53066 0.16233 0.019135 14.2818 0.11882 0.00015385 0.77133 0.0090202 0.0099956 0.0015266 0.9851 0.99048 3.3112e-006 1.3245e-005 0.16191 0.72939 0.81265 0.0014696 0.85595 0.39568 0.001977 0.41903 1.6737 1.6709 16.0167 144.9174 0.00032289 -85.0737 0.27795
7.382 0.98812 5.4738e-005 3.8183 0.011939 9.6136e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.487 0.5307 0.16235 0.019136 14.2845 0.11883 0.00015386 0.77133 0.0090206 0.0099961 0.0015255 0.98511 0.99049 3.3087e-006 1.3235e-005 0.16191 0.73018 0.81316 0.001469 0.85681 0.39589 0.0019763 0.41904 1.6754 1.6725 16.0167 144.9174 0.00032213 -85.0781 0.27895
7.383 0.98812 5.4738e-005 3.8183 0.011939 9.6149e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4871 0.53075 0.16236 0.019137 14.2872 0.11884 0.00015387 0.77132 0.009021 0.0099965 0.0015244 0.98513 0.9905 3.3062e-006 1.3225e-005 0.16191 0.73097 0.81367 0.0014685 0.85767 0.39609 0.0019756 0.41905 1.6771 1.6742 16.0168 144.9175 0.00032137 -85.0823 0.27995
7.384 0.98812 5.4738e-005 3.8183 0.011939 9.6162e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4872 0.53079 0.16237 0.019139 14.29 0.11884 0.00015388 0.77131 0.0090215 0.009997 0.0015233 0.98514 0.99051 3.3037e-006 1.3215e-005 0.16192 0.73175 0.81418 0.0014679 0.85853 0.3963 0.0019749 0.41906 1.6787 1.6759 16.0168 144.9175 0.00032061 -85.0866 0.28095
7.385 0.98812 5.4738e-005 3.8183 0.011939 9.6174e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4873 0.53084 0.16239 0.01914 14.2927 0.11885 0.00015389 0.7713 0.0090219 0.0099974 0.0015223 0.98516 0.99052 3.3012e-006 1.3205e-005 0.16192 0.73254 0.81468 0.0014674 0.85938 0.39651 0.0019742 0.41907 1.6804 1.6776 16.0168 144.9175 0.00031986 -85.0908 0.28195
7.386 0.98812 5.4738e-005 3.8183 0.011939 9.6187e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4874 0.53088 0.1624 0.019141 14.2954 0.11886 0.0001539 0.7713 0.0090223 0.0099979 0.0015212 0.98517 0.99053 3.2988e-006 1.3195e-005 0.16192 0.73332 0.81518 0.0014668 0.86023 0.39671 0.0019735 0.41908 1.6821 1.6793 16.0168 144.9175 0.00031911 -85.0949 0.28295
7.387 0.98812 5.4737e-005 3.8183 0.011939 9.62e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4874 0.53093 0.16242 0.019142 14.2982 0.11886 0.00015391 0.77129 0.0090228 0.0099984 0.0015201 0.98518 0.99054 3.2964e-006 1.3186e-005 0.16193 0.7341 0.81568 0.0014663 0.86107 0.39692 0.0019728 0.41909 1.6837 1.6809 16.0169 144.9175 0.00031837 -85.0991 0.28395
7.388 0.98812 5.4737e-005 3.8183 0.011939 9.6213e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4875 0.53097 0.16243 0.019143 14.3009 0.11887 0.00015392 0.77128 0.0090232 0.0099988 0.0015191 0.9852 0.99055 3.294e-006 1.3176e-005 0.16193 0.73487 0.81617 0.0014658 0.8619 0.39713 0.0019721 0.4191 1.6854 1.6826 16.0169 144.9175 0.00031763 -85.1032 0.28495
7.389 0.98812 5.4737e-005 3.8183 0.011939 9.6226e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.4876 0.53102 0.16244 0.019145 14.3036 0.11888 0.00015393 0.77128 0.0090236 0.0099993 0.0015181 0.98521 0.99056 3.2916e-006 1.3167e-005 0.16193 0.73565 0.81667 0.0014653 0.86273 0.39733 0.0019714 0.41911 1.687 1.6843 16.0169 144.9175 0.00031689 -85.1073 0.28595
7.39 0.98812 5.4737e-005 3.8183 0.011939 9.6239e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4877 0.53106 0.16246 0.019146 14.3064 0.11889 0.00015394 0.77127 0.0090241 0.0099998 0.001517 0.98523 0.99057 3.2893e-006 1.3157e-005 0.16194 0.73642 0.81715 0.0014647 0.86356 0.39754 0.0019707 0.41913 1.6887 1.6859 16.0169 144.9176 0.00031615 -85.1113 0.28695
7.391 0.98812 5.4737e-005 3.8183 0.011939 9.6252e-005 0.0011692 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4878 0.53111 0.16247 0.019147 14.3091 0.11889 0.00015395 0.77126 0.0090245 0.01 0.001516 0.98524 0.99058 3.2869e-006 1.3148e-005 0.16194 0.73719 0.81764 0.0014642 0.86438 0.39775 0.0019701 0.41914 1.6903 1.6876 16.017 144.9176 0.00031542 -85.1153 0.28795
7.392 0.98812 5.4737e-005 3.8183 0.011938 9.6264e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4879 0.53116 0.16249 0.019148 14.3118 0.1189 0.00015396 0.77125 0.0090249 0.010001 0.001515 0.98525 0.99058 3.2846e-006 1.3139e-005 0.16194 0.73796 0.81813 0.0014637 0.8652 0.39795 0.0019694 0.41915 1.692 1.6892 16.017 144.9176 0.0003147 -85.1193 0.28895
7.393 0.98812 5.4737e-005 3.8183 0.011938 9.6277e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.488 0.5312 0.1625 0.019149 14.3146 0.11891 0.00015398 0.77125 0.0090254 0.010001 0.001514 0.98527 0.99059 3.2823e-006 1.3129e-005 0.16195 0.73872 0.81861 0.0014632 0.86601 0.39816 0.0019687 0.41916 1.6936 1.6909 16.017 144.9176 0.00031397 -85.1233 0.28995
7.394 0.98812 5.4737e-005 3.8183 0.011938 9.629e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4881 0.53125 0.16251 0.01915 14.3173 0.11891 0.00015399 0.77124 0.0090258 0.010002 0.001513 0.98528 0.9906 3.28e-006 1.312e-005 0.16195 0.73948 0.81909 0.0014627 0.86682 0.39836 0.0019681 0.41917 1.6952 1.6925 16.017 144.9176 0.00031325 -85.1272 0.29095
7.395 0.98812 5.4737e-005 3.8183 0.011938 9.6303e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4882 0.53129 0.16253 0.019152 14.32 0.11892 0.000154 0.77123 0.0090262 0.010002 0.0015121 0.98529 0.99061 3.2777e-006 1.3111e-005 0.16195 0.74024 0.81956 0.0014622 0.86762 0.39857 0.0019674 0.41918 1.6969 1.6941 16.0171 144.9176 0.00031253 -85.1311 0.29195
7.396 0.98812 5.4737e-005 3.8183 0.011938 9.6316e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4882 0.53134 0.16254 0.019153 14.3228 0.11893 0.00015401 0.77123 0.0090267 0.010003 0.0015111 0.98531 0.99062 3.2755e-006 1.3102e-005 0.16196 0.741 0.82004 0.0014617 0.86842 0.39878 0.0019668 0.41919 1.6985 1.6958 16.0171 144.9177 0.00031182 -85.135 0.29295
7.397 0.98812 5.4737e-005 3.8183 0.011938 9.6329e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4883 0.53138 0.16256 0.019154 14.3255 0.11894 0.00015402 0.77122 0.0090271 0.010003 0.0015101 0.98532 0.99063 3.2733e-006 1.3093e-005 0.16196 0.74175 0.82051 0.0014612 0.86921 0.39898 0.0019661 0.4192 1.7001 1.6974 16.0171 144.9177 0.00031111 -85.1388 0.29395
7.398 0.98812 5.4737e-005 3.8183 0.011938 9.6342e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4884 0.53143 0.16257 0.019155 14.3283 0.11894 0.00015403 0.77121 0.0090275 0.010003 0.0015092 0.98533 0.99064 3.2711e-006 1.3084e-005 0.16197 0.74251 0.82098 0.0014607 0.87 0.39919 0.0019655 0.41922 1.7017 1.699 16.0171 144.9177 0.0003104 -85.1427 0.29495
7.399 0.98812 5.4737e-005 3.8183 0.011938 9.6354e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4885 0.53147 0.16258 0.019156 14.331 0.11895 0.00015404 0.7712 0.009028 0.010004 0.0015082 0.98534 0.99065 3.2689e-006 1.3076e-005 0.16197 0.74326 0.82145 0.0014603 0.87079 0.39939 0.0019648 0.41923 1.7033 1.7006 16.0172 144.9177 0.0003097 -85.1464 0.29595
7.4 0.98812 5.4736e-005 3.8183 0.011938 9.6367e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4886 0.53152 0.1626 0.019158 14.3337 0.11896 0.00015405 0.7712 0.0090284 0.010004 0.0015073 0.98536 0.99066 3.2667e-006 1.3067e-005 0.16197 0.74401 0.82191 0.0014598 0.87157 0.3996 0.0019642 0.41924 1.7049 1.7022 16.0172 144.9177 0.000309 -85.1502 0.29695
7.401 0.98812 5.4736e-005 3.8183 0.011938 9.638e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4887 0.53156 0.16261 0.019159 14.3365 0.11896 0.00015406 0.77119 0.0090288 0.010005 0.0015063 0.98537 0.99066 3.2646e-006 1.3058e-005 0.16198 0.74475 0.82237 0.0014593 0.87234 0.39981 0.0019636 0.41925 1.7065 1.7039 16.0172 144.9177 0.0003083 -85.1539 0.29795
7.402 0.98812 5.4736e-005 3.8183 0.011938 9.6393e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4888 0.53161 0.16263 0.01916 14.3392 0.11897 0.00015407 0.77118 0.0090293 0.010005 0.0015054 0.98538 0.99067 3.2624e-006 1.305e-005 0.16198 0.7455 0.82283 0.0014588 0.87311 0.40001 0.001963 0.41926 1.7081 1.7055 16.0172 144.9178 0.00030761 -85.1576 0.29895
7.403 0.98812 5.4736e-005 3.8183 0.011938 9.6406e-005 0.0011693 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4889 0.53165 0.16264 0.019161 14.342 0.11898 0.00015408 0.77118 0.0090297 0.010006 0.0015045 0.98539 0.99068 3.2603e-006 1.3041e-005 0.16198 0.74624 0.82329 0.0014583 0.87388 0.40022 0.0019624 0.41927 1.7097 1.7071 16.0173 144.9178 0.00030692 -85.1613 0.29995
7.404 0.98812 5.4736e-005 3.8183 0.011938 9.6419e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4889 0.5317 0.16265 0.019162 14.3447 0.11899 0.00015409 0.77117 0.0090301 0.010006 0.0015036 0.98541 0.99069 3.2582e-006 1.3033e-005 0.16199 0.74698 0.82375 0.0014579 0.87464 0.40042 0.0019618 0.41928 1.7113 1.7087 16.0173 144.9178 0.00030623 -85.165 0.30095
7.405 0.98812 5.4736e-005 3.8183 0.011938 9.6432e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.489 0.53175 0.16267 0.019164 14.3474 0.11899 0.0001541 0.77116 0.0090306 0.010007 0.0015026 0.98542 0.9907 3.2561e-006 1.3025e-005 0.16199 0.74771 0.8242 0.0014574 0.8754 0.40063 0.0019612 0.4193 1.7129 1.7103 16.0173 144.9178 0.00030555 -85.1686 0.30195
7.406 0.98812 5.4736e-005 3.8183 0.011938 9.6444e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4891 0.53179 0.16268 0.019165 14.3502 0.119 0.00015411 0.77115 0.009031 0.010007 0.0015018 0.98543 0.9907 3.254e-006 1.3016e-005 0.16199 0.74845 0.82465 0.001457 0.87615 0.40083 0.0019606 0.41931 1.7145 1.7118 16.0173 144.9178 0.00030487 -85.1722 0.30295
7.407 0.98812 5.4736e-005 3.8183 0.011938 9.6457e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4892 0.53184 0.1627 0.019166 14.3529 0.11901 0.00015412 0.77115 0.0090314 0.010008 0.0015009 0.98544 0.99071 3.252e-006 1.3008e-005 0.162 0.74918 0.8251 0.0014565 0.8769 0.40104 0.00196 0.41932 1.716 1.7134 16.0174 144.9178 0.00030419 -85.1757 0.30395
7.408 0.98812 5.4736e-005 3.8183 0.011938 9.647e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4893 0.53188 0.16271 0.019167 14.3557 0.11901 0.00015414 0.77114 0.0090319 0.010008 0.0015 0.98545 0.99072 3.2499e-006 1.3e-005 0.162 0.74991 0.82554 0.0014561 0.87765 0.40125 0.0019594 0.41933 1.7176 1.715 16.0174 144.9179 0.00030352 -85.1793 0.30495
7.409 0.98812 5.4736e-005 3.8183 0.011938 9.6483e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4894 0.53193 0.16272 0.019168 14.3584 0.11902 0.00015415 0.77113 0.0090323 0.010009 0.0014991 0.98547 0.99073 3.2479e-006 1.2992e-005 0.162 0.75064 0.82599 0.0014556 0.87839 0.40145 0.0019588 0.41934 1.7192 1.7166 16.0174 144.9179 0.00030284 -85.1828 0.30595
7.41 0.98812 5.4736e-005 3.8183 0.011938 9.6496e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4895 0.53197 0.16274 0.019169 14.3612 0.11903 0.00015416 0.77113 0.0090327 0.010009 0.0014982 0.98548 0.99074 3.2459e-006 1.2984e-005 0.16201 0.75136 0.82643 0.0014552 0.87912 0.40166 0.0019582 0.41935 1.7207 1.7182 16.0174 144.9179 0.00030218 -85.1863 0.30695
7.411 0.98812 5.4736e-005 3.8183 0.011938 9.6509e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4896 0.53202 0.16275 0.019171 14.3639 0.11904 0.00015417 0.77112 0.0090331 0.010009 0.0014974 0.98549 0.99074 3.2439e-006 1.2976e-005 0.16201 0.75208 0.82687 0.0014547 0.87986 0.40186 0.0019576 0.41937 1.7223 1.7197 16.0174 144.9179 0.00030151 -85.1897 0.30795
7.412 0.98812 5.4735e-005 3.8183 0.011938 9.6522e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4897 0.53206 0.16277 0.019172 14.3666 0.11904 0.00015418 0.77111 0.0090336 0.01001 0.0014965 0.9855 0.99075 3.242e-006 1.2968e-005 0.16201 0.75281 0.8273 0.0014543 0.88058 0.40207 0.0019571 0.41938 1.7239 1.7213 16.0175 144.9179 0.00030085 -85.1932 0.30895
7.413 0.98812 5.4735e-005 3.8183 0.011938 9.6534e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4897 0.53211 0.16278 0.019173 14.3694 0.11905 0.00015419 0.7711 0.009034 0.01001 0.0014957 0.98551 0.99076 3.24e-006 1.296e-005 0.16202 0.75352 0.82774 0.0014539 0.88131 0.40227 0.0019565 0.41939 1.7254 1.7228 16.0175 144.9179 0.00030019 -85.1966 0.30995
7.414 0.98812 5.4735e-005 3.8183 0.011938 9.6547e-005 0.0011693 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4898 0.53215 0.16279 0.019174 14.3721 0.11906 0.0001542 0.7711 0.0090344 0.010011 0.0014948 0.98552 0.99077 3.2381e-006 1.2952e-005 0.16202 0.75424 0.82817 0.0014534 0.88202 0.40248 0.0019559 0.4194 1.727 1.7244 16.0175 144.918 0.00029953 -85.2 0.31095
7.415 0.98812 5.4735e-005 3.8183 0.011938 9.656e-005 0.0011694 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.4899 0.5322 0.16281 0.019175 14.3749 0.11906 0.00015421 0.77109 0.0090349 0.010011 0.001494 0.98553 0.99077 3.2361e-006 1.2945e-005 0.16202 0.75495 0.8286 0.001453 0.88274 0.40268 0.0019554 0.41941 1.7285 1.726 16.0175 144.918 0.00029888 -85.2033 0.31195
7.416 0.98812 5.4735e-005 3.8183 0.011938 9.6573e-005 0.0011694 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.49 0.53224 0.16282 0.019177 14.3776 0.11907 0.00015422 0.77108 0.0090353 0.010012 0.0014931 0.98554 0.99078 3.2342e-006 1.2937e-005 0.16203 0.75567 0.82903 0.0014526 0.88345 0.40289 0.0019548 0.41943 1.73 1.7275 16.0175 144.918 0.00029823 -85.2066 0.31295
7.417 0.98812 5.4735e-005 3.8183 0.011938 9.6586e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4901 0.53229 0.16284 0.019178 14.3804 0.11908 0.00015423 0.77108 0.0090357 0.010012 0.0014923 0.98556 0.99079 3.2323e-006 1.293e-005 0.16203 0.75638 0.82945 0.0014522 0.88416 0.40309 0.0019543 0.41944 1.7316 1.729 16.0176 144.918 0.00029759 -85.2099 0.31395
7.418 0.98812 5.4735e-005 3.8183 0.011938 9.6599e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4902 0.53233 0.16285 0.019179 14.3831 0.11909 0.00015424 0.77107 0.0090362 0.010013 0.0014915 0.98557 0.9908 3.2305e-006 1.2922e-005 0.16203 0.75708 0.82988 0.0014517 0.88486 0.4033 0.0019537 0.41945 1.7331 1.7306 16.0176 144.918 0.00029694 -85.2132 0.31495
7.419 0.98812 5.4735e-005 3.8183 0.011938 9.6611e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4903 0.53238 0.16286 0.01918 14.3859 0.11909 0.00015425 0.77106 0.0090366 0.010013 0.0014907 0.98558 0.9908 3.2286e-006 1.2915e-005 0.16204 0.75779 0.8303 0.0014513 0.88556 0.4035 0.0019532 0.41946 1.7346 1.7321 16.0176 144.918 0.0002963 -85.2165 0.31595
7.42 0.98812 5.4735e-005 3.8183 0.011938 9.6624e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4904 0.53243 0.16288 0.019181 14.3886 0.1191 0.00015426 0.77105 0.009037 0.010014 0.0014899 0.98559 0.99081 3.2268e-006 1.2907e-005 0.16204 0.75849 0.83072 0.0014509 0.88625 0.40371 0.0019526 0.41947 1.7361 1.7336 16.0176 144.9181 0.00029566 -85.2197 0.31695
7.421 0.98812 5.4735e-005 3.8183 0.011938 9.6637e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4904 0.53247 0.16289 0.019183 14.3913 0.11911 0.00015427 0.77105 0.0090374 0.010014 0.0014891 0.9856 0.99082 3.2249e-006 1.29e-005 0.16204 0.75919 0.83114 0.0014505 0.88694 0.40391 0.0019521 0.41949 1.7377 1.7352 16.0176 144.9181 0.00029503 -85.2229 0.31795
7.422 0.98812 5.4735e-005 3.8183 0.011938 9.665e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4905 0.53252 0.16291 0.019184 14.3941 0.11911 0.00015428 0.77104 0.0090379 0.010014 0.0014883 0.98561 0.99083 3.2231e-006 1.2893e-005 0.16205 0.75989 0.83155 0.0014501 0.88763 0.40412 0.0019516 0.4195 1.7392 1.7367 16.0177 144.9181 0.0002944 -85.2261 0.31895
7.423 0.98812 5.4735e-005 3.8183 0.011938 9.6663e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4906 0.53256 0.16292 0.019185 14.3968 0.11912 0.0001543 0.77103 0.0090383 0.010015 0.0014875 0.98562 0.99083 3.2213e-006 1.2885e-005 0.16205 0.76059 0.83197 0.0014497 0.88831 0.40432 0.0019511 0.41951 1.7407 1.7382 16.0177 144.9181 0.00029377 -85.2293 0.31995
7.424 0.98812 5.4735e-005 3.8183 0.011938 9.6676e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4907 0.53261 0.16293 0.019186 14.3996 0.11913 0.00015431 0.77103 0.0090387 0.010015 0.0014867 0.98563 0.99084 3.2195e-006 1.2878e-005 0.16205 0.76128 0.83238 0.0014493 0.88899 0.40453 0.0019505 0.41952 1.7422 1.7397 16.0177 144.9181 0.00029314 -85.2324 0.32095
7.425 0.98812 5.4734e-005 3.8183 0.011938 9.6689e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4908 0.53265 0.16295 0.019187 14.4023 0.11914 0.00015432 0.77102 0.0090392 0.010016 0.001486 0.98564 0.99085 3.2177e-006 1.2871e-005 0.16206 0.76198 0.83279 0.0014489 0.88966 0.40473 0.00195 0.41953 1.7437 1.7412 16.0177 144.9182 0.00029252 -85.2355 0.32195
7.426 0.98812 5.4734e-005 3.8183 0.011938 9.6701e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4909 0.5327 0.16296 0.019188 14.4051 0.11914 0.00015433 0.77101 0.0090396 0.010016 0.0014852 0.98565 0.99085 3.216e-006 1.2864e-005 0.16206 0.76267 0.83319 0.0014485 0.89033 0.40494 0.0019495 0.41955 1.7452 1.7427 16.0177 144.9182 0.0002919 -85.2386 0.32295
7.427 0.98812 5.4734e-005 3.8183 0.011938 9.6714e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.491 0.53274 0.16298 0.01919 14.4078 0.11915 0.00015434 0.771 0.00904 0.010017 0.0014844 0.98566 0.99086 3.2142e-006 1.2857e-005 0.16206 0.76335 0.8336 0.0014481 0.891 0.40514 0.001949 0.41956 1.7467 1.7443 16.0177 144.9182 0.00029128 -85.2417 0.32395
7.428 0.98812 5.4734e-005 3.8183 0.011938 9.6727e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4911 0.53279 0.16299 0.019191 14.4106 0.11916 0.00015435 0.771 0.0090405 0.010017 0.0014837 0.98567 0.99087 3.2125e-006 1.285e-005 0.16207 0.76404 0.834 0.0014477 0.89166 0.40534 0.0019485 0.41957 1.7482 1.7457 16.0178 144.9182 0.00029067 -85.2448 0.32495
7.429 0.98812 5.4734e-005 3.8183 0.011938 9.674e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4912 0.53283 0.163 0.019192 14.4133 0.11916 0.00015436 0.77099 0.0090409 0.010018 0.0014829 0.98568 0.99087 3.2108e-006 1.2843e-005 0.16207 0.76472 0.8344 0.0014474 0.89232 0.40555 0.001948 0.41958 1.7497 1.7472 16.0178 144.9182 0.00029006 -85.2478 0.32595
7.43 0.98812 5.4734e-005 3.8183 0.011938 9.6753e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4912 0.53288 0.16302 0.019193 14.4161 0.11917 0.00015437 0.77098 0.0090413 0.010018 0.0014822 0.98569 0.99088 3.2091e-006 1.2836e-005 0.16207 0.7654 0.8348 0.001447 0.89297 0.40575 0.0019475 0.4196 1.7511 1.7487 16.0178 144.9182 0.00028945 -85.2508 0.32695
7.431 0.98812 5.4734e-005 3.8183 0.011938 9.6766e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4913 0.53292 0.16303 0.019194 14.4188 0.11918 0.00015438 0.77098 0.0090417 0.010019 0.0014815 0.9857 0.99089 3.2074e-006 1.283e-005 0.16208 0.76608 0.8352 0.0014466 0.89362 0.40596 0.001947 0.41961 1.7526 1.7502 16.0178 144.9183 0.00028884 -85.2538 0.32795
7.432 0.98812 5.4734e-005 3.8183 0.011938 9.6779e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4914 0.53297 0.16305 0.019196 14.4216 0.11919 0.00015439 0.77097 0.0090422 0.010019 0.0014807 0.98571 0.99089 3.2057e-006 1.2823e-005 0.16208 0.76676 0.8356 0.0014463 0.89427 0.40616 0.0019465 0.41962 1.7541 1.7517 16.0178 144.9183 0.00028824 -85.2567 0.32895
7.433 0.98812 5.4734e-005 3.8183 0.011938 9.6791e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4915 0.53301 0.16306 0.019197 14.4243 0.11919 0.0001544 0.77096 0.0090426 0.01002 0.00148 0.98572 0.9909 3.204e-006 1.2816e-005 0.16208 0.76744 0.83599 0.0014459 0.89491 0.40637 0.001946 0.41963 1.7556 1.7532 16.0179 144.9183 0.00028764 -85.2597 0.32995
7.434 0.98812 5.4734e-005 3.8183 0.011938 9.6804e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4916 0.53306 0.16307 0.019198 14.4271 0.1192 0.00015441 0.77096 0.009043 0.01002 0.0014793 0.98573 0.99091 3.2024e-006 1.281e-005 0.16209 0.76811 0.83638 0.0014455 0.89555 0.40657 0.0019455 0.41965 1.757 1.7547 16.0179 144.9183 0.00028704 -85.2626 0.33095
7.435 0.98812 5.4734e-005 3.8183 0.011938 9.6817e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4917 0.53311 0.16309 0.019199 14.4298 0.11921 0.00015442 0.77095 0.0090435 0.01002 0.0014786 0.98574 0.99091 3.2007e-006 1.2803e-005 0.16209 0.76878 0.83677 0.0014451 0.89618 0.40678 0.0019451 0.41966 1.7585 1.7561 16.0179 144.9183 0.00028644 -85.2655 0.33195
7.436 0.98812 5.4734e-005 3.8183 0.011938 9.683e-005 0.0011694 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4918 0.53315 0.1631 0.0192 14.4326 0.11921 0.00015443 0.77094 0.0090439 0.010021 0.0014779 0.98575 0.99092 3.1991e-006 1.2797e-005 0.16209 0.76945 0.83716 0.0014448 0.89681 0.40698 0.0019446 0.41967 1.76 1.7576 16.0179 144.9183 0.00028585 -85.2683 0.33295
7.437 0.98812 5.4733e-005 3.8183 0.011938 9.6843e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4919 0.5332 0.16312 0.019201 14.4353 0.11922 0.00015444 0.77093 0.0090443 0.010021 0.0014772 0.98576 0.99092 3.1975e-006 1.279e-005 0.1621 0.77012 0.83755 0.0014444 0.89744 0.40718 0.0019441 0.41968 1.7614 1.7591 16.0179 144.9184 0.00028526 -85.2712 0.33395
7.438 0.98812 5.4733e-005 3.8183 0.011938 9.6856e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4919 0.53324 0.16313 0.019203 14.4381 0.11923 0.00015445 0.77093 0.0090448 0.010022 0.0014765 0.98577 0.99093 3.1959e-006 1.2784e-005 0.1621 0.77078 0.83793 0.0014441 0.89807 0.40739 0.0019436 0.4197 1.7629 1.7605 16.0179 144.9184 0.00028468 -85.274 0.33495
7.439 0.98812 5.4733e-005 3.8183 0.011938 9.6869e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.492 0.53329 0.16314 0.019204 14.4408 0.11923 0.00015447 0.77092 0.0090452 0.010022 0.0014758 0.98578 0.99094 3.1943e-006 1.2777e-005 0.1621 0.77145 0.83831 0.0014437 0.89869 0.40759 0.0019432 0.41971 1.7643 1.762 16.0179 144.9184 0.00028409 -85.2768 0.33595
7.44 0.98812 5.4733e-005 3.8183 0.011938 9.6881e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4921 0.53333 0.16316 0.019205 14.4436 0.11924 0.00015448 0.77091 0.0090456 0.010023 0.0014751 0.98578 0.99094 3.1927e-006 1.2771e-005 0.1621 0.77211 0.83869 0.0014433 0.8993 0.4078 0.0019427 0.41972 1.7658 1.7634 16.018 144.9184 0.00028351 -85.2796 0.33695
7.441 0.98812 5.4733e-005 3.8183 0.011938 9.6894e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4922 0.53338 0.16317 0.019206 14.4463 0.11925 0.00015449 0.77091 0.009046 0.010023 0.0014744 0.98579 0.99095 3.1912e-006 1.2765e-005 0.16211 0.77277 0.83907 0.001443 0.89991 0.408 0.0019423 0.41973 1.7672 1.7649 16.018 144.9184 0.00028293 -85.2824 0.33795
7.442 0.98812 5.4733e-005 3.8183 0.011938 9.6907e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4923 0.53342 0.16319 0.019207 14.4491 0.11926 0.0001545 0.7709 0.0090465 0.010024 0.0014737 0.9858 0.99095 3.1896e-006 1.2759e-005 0.16211 0.77342 0.83945 0.0014426 0.90052 0.4082 0.0019418 0.41975 1.7686 1.7663 16.018 144.9184 0.00028236 -85.2851 0.33895
7.443 0.98812 5.4733e-005 3.8183 0.011938 9.692e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4924 0.53347 0.1632 0.019209 14.4519 0.11926 0.00015451 0.77089 0.0090469 0.010024 0.0014731 0.98581 0.99096 3.1881e-006 1.2752e-005 0.16211 0.77408 0.83982 0.0014423 0.90113 0.40841 0.0019414 0.41976 1.7701 1.7677 16.018 144.9185 0.00028178 -85.2879 0.33995
7.444 0.98812 5.4733e-005 3.8183 0.011938 9.6933e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4925 0.53351 0.16321 0.01921 14.4546 0.11927 0.00015452 0.77088 0.0090473 0.010025 0.0014724 0.98582 0.99097 3.1866e-006 1.2746e-005 0.16212 0.77473 0.8402 0.001442 0.90173 0.40861 0.0019409 0.41977 1.7715 1.7692 16.018 144.9185 0.00028121 -85.2906 0.34095
7.445 0.98812 5.4733e-005 3.8183 0.011938 9.6946e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4926 0.53356 0.16323 0.019211 14.4574 0.11928 0.00015453 0.77088 0.0090478 0.010025 0.0014717 0.98583 0.99097 3.185e-006 1.274e-005 0.16212 0.77538 0.84057 0.0014416 0.90233 0.40881 0.0019405 0.41978 1.7729 1.7706 16.018 144.9185 0.00028064 -85.2933 0.34195
7.446 0.98812 5.4733e-005 3.8183 0.011938 9.6958e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4927 0.5336 0.16324 0.019212 14.4601 0.11928 0.00015454 0.77087 0.0090482 0.010025 0.0014711 0.98584 0.99098 3.1835e-006 1.2734e-005 0.16212 0.77603 0.84094 0.0014413 0.90292 0.40902 0.00194 0.4198 1.7743 1.772 16.018 144.9185 0.00028008 -85.2959 0.34295
7.447 0.98812 5.4733e-005 3.8183 0.011938 9.6971e-005 0.0011695 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.4927 0.53365 0.16326 0.019213 14.4629 0.11929 0.00015455 0.77086 0.0090486 0.010026 0.0014704 0.98585 0.99098 3.182e-006 1.2728e-005 0.16213 0.77668 0.84131 0.001441 0.90351 0.40922 0.0019396 0.41981 1.7757 1.7735 16.0181 144.9185 0.00027951 -85.2986 0.34395
7.448 0.98812 5.4733e-005 3.8183 0.011938 9.6984e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4928 0.53369 0.16327 0.019214 14.4656 0.1193 0.00015456 0.77086 0.009049 0.010026 0.0014698 0.98585 0.99099 3.1806e-006 1.2722e-005 0.16213 0.77732 0.84167 0.0014406 0.9041 0.40943 0.0019392 0.41982 1.7772 1.7749 16.0181 144.9186 0.00027895 -85.3012 0.34495
7.449 0.98812 5.4732e-005 3.8183 0.011937 9.6997e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4929 0.53374 0.16328 0.019216 14.4684 0.11931 0.00015457 0.77085 0.0090495 0.010027 0.0014692 0.98586 0.99099 3.1791e-006 1.2716e-005 0.16213 0.77796 0.84204 0.0014403 0.90469 0.40963 0.0019387 0.41984 1.7786 1.7763 16.0181 144.9186 0.00027839 -85.3038 0.34595
7.45 0.98812 5.4732e-005 3.8183 0.011937 9.701e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.493 0.53379 0.1633 0.019217 14.4711 0.11931 0.00015458 0.77084 0.0090499 0.010027 0.0014685 0.98587 0.991 3.1776e-006 1.2711e-005 0.16214 0.7786 0.8424 0.00144 0.90527 0.40983 0.0019383 0.41985 1.78 1.7777 16.0181 144.9186 0.00027784 -85.3064 0.34695
7.451 0.98812 5.4732e-005 3.8183 0.011937 9.7023e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4931 0.53383 0.16331 0.019218 14.4739 0.11932 0.00015459 0.77083 0.0090503 0.010028 0.0014679 0.98588 0.99101 3.1762e-006 1.2705e-005 0.16214 0.77924 0.84276 0.0014397 0.90584 0.41004 0.0019379 0.41986 1.7814 1.7791 16.0181 144.9186 0.00027729 -85.309 0.34795
7.452 0.98812 5.4732e-005 3.8183 0.011937 9.7036e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4932 0.53388 0.16333 0.019219 14.4767 0.11933 0.0001546 0.77083 0.0090508 0.010028 0.0014673 0.98589 0.99101 3.1748e-006 1.2699e-005 0.16214 0.77988 0.84312 0.0014393 0.90642 0.41024 0.0019375 0.41988 1.7828 1.7805 16.0181 144.9186 0.00027674 -85.3115 0.34895
7.453 0.98812 5.4732e-005 3.8183 0.011937 9.7048e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4933 0.53392 0.16334 0.01922 14.4794 0.11933 0.00015461 0.77082 0.0090512 0.010029 0.0014667 0.9859 0.99102 3.1733e-006 1.2693e-005 0.16215 0.78051 0.84348 0.001439 0.90699 0.41044 0.001937 0.41989 1.7842 1.7819 16.0181 144.9186 0.00027619 -85.3141 0.34995
7.454 0.98812 5.4732e-005 3.8183 0.011937 9.7061e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4934 0.53397 0.16335 0.019222 14.4822 0.11934 0.00015462 0.77081 0.0090516 0.010029 0.001466 0.9859 0.99102 3.1719e-006 1.2688e-005 0.16215 0.78115 0.84383 0.0014387 0.90755 0.41065 0.0019366 0.4199 1.7855 1.7833 16.0181 144.9187 0.00027564 -85.3166 0.35095
7.455 0.98812 5.4732e-005 3.8183 0.011937 9.7074e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4934 0.53401 0.16337 0.019223 14.4849 0.11935 0.00015464 0.77081 0.009052 0.01003 0.0014654 0.98591 0.99103 3.1705e-006 1.2682e-005 0.16215 0.78178 0.84419 0.0014384 0.90812 0.41085 0.0019362 0.41991 1.7869 1.7847 16.0182 144.9187 0.0002751 -85.3191 0.35195
7.456 0.98812 5.4732e-005 3.8183 0.011937 9.7087e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4935 0.53406 0.16338 0.019224 14.4877 0.11936 0.00015465 0.7708 0.0090525 0.01003 0.0014648 0.98592 0.99103 3.1691e-006 1.2677e-005 0.16216 0.78241 0.84454 0.0014381 0.90868 0.41105 0.0019358 0.41993 1.7883 1.7861 16.0182 144.9187 0.00027456 -85.3216 0.35295
7.457 0.98812 5.4732e-005 3.8183 0.011937 9.71e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4936 0.5341 0.1634 0.019225 14.4904 0.11936 0.00015466 0.77079 0.0090529 0.010031 0.0014642 0.98593 0.99104 3.1678e-006 1.2671e-005 0.16216 0.78303 0.84489 0.0014378 0.90923 0.41125 0.0019354 0.41994 1.7897 1.7875 16.0182 144.9187 0.00027402 -85.324 0.35395
7.458 0.98812 5.4732e-005 3.8183 0.011937 9.7113e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4937 0.53415 0.16341 0.019226 14.4932 0.11937 0.00015467 0.77079 0.0090533 0.010031 0.0014636 0.98594 0.99104 3.1664e-006 1.2666e-005 0.16216 0.78366 0.84524 0.0014374 0.90979 0.41146 0.001935 0.41995 1.7911 1.7889 16.0182 144.9187 0.00027348 -85.3265 0.35495
7.459 0.98812 5.4732e-005 3.8183 0.011937 9.7126e-005 0.0011695 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4938 0.53419 0.16342 0.019227 14.496 0.11938 0.00015468 0.77078 0.0090538 0.010031 0.001463 0.98594 0.99105 3.165e-006 1.266e-005 0.16217 0.78428 0.84559 0.0014371 0.91034 0.41166 0.0019346 0.41997 1.7924 1.7902 16.0182 144.9188 0.00027295 -85.3289 0.35595
7.46 0.98812 5.4732e-005 3.8183 0.011937 9.7138e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4939 0.53424 0.16344 0.019229 14.4987 0.11938 0.00015469 0.77077 0.0090542 0.010032 0.0014624 0.98595 0.99105 3.1637e-006 1.2655e-005 0.16217 0.7849 0.84593 0.0014368 0.91088 0.41186 0.0019342 0.41998 1.7938 1.7916 16.0182 144.9188 0.00027242 -85.3313 0.35695
7.461 0.98812 5.4732e-005 3.8183 0.011937 9.7151e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.494 0.53428 0.16345 0.01923 14.5015 0.11939 0.0001547 0.77076 0.0090546 0.010032 0.0014619 0.98596 0.99106 3.1623e-006 1.2649e-005 0.16217 0.78552 0.84628 0.0014365 0.91142 0.41207 0.0019338 0.41999 1.7952 1.793 16.0182 144.9188 0.00027189 -85.3337 0.35795
7.462 0.98812 5.4731e-005 3.8183 0.011937 9.7164e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4941 0.53433 0.16347 0.019231 14.5042 0.1194 0.00015471 0.77076 0.009055 0.010033 0.0014613 0.98597 0.99106 3.161e-006 1.2644e-005 0.16218 0.78614 0.84662 0.0014362 0.91196 0.41227 0.0019334 0.42001 1.7965 1.7944 16.0182 144.9188 0.00027136 -85.336 0.35895
7.463 0.98812 5.4731e-005 3.8183 0.011937 9.7177e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4942 0.53437 0.16348 0.019232 14.507 0.11941 0.00015472 0.77075 0.0090555 0.010033 0.0014607 0.98597 0.99107 3.1597e-006 1.2639e-005 0.16218 0.78675 0.84696 0.0014359 0.9125 0.41247 0.001933 0.42002 1.7979 1.7957 16.0182 144.9188 0.00027084 -85.3384 0.35995
7.464 0.98812 5.4731e-005 3.8183 0.011937 9.719e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4942 0.53442 0.16349 0.019233 14.5098 0.11941 0.00015473 0.77074 0.0090559 0.010034 0.0014601 0.98598 0.99107 3.1584e-006 1.2634e-005 0.16218 0.78737 0.8473 0.0014356 0.91303 0.41267 0.0019327 0.42003 1.7992 1.7971 16.0183 144.9188 0.00027032 -85.3407 0.36095
7.465 0.98812 5.4731e-005 3.8183 0.011937 9.7203e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4943 0.53447 0.16351 0.019234 14.5125 0.11942 0.00015474 0.77074 0.0090563 0.010034 0.0014596 0.98599 0.99108 3.1571e-006 1.2628e-005 0.16219 0.78798 0.84764 0.0014353 0.91356 0.41288 0.0019323 0.42005 1.8006 1.7984 16.0183 144.9189 0.0002698 -85.343 0.36195
7.466 0.98812 5.4731e-005 3.8183 0.011937 9.7215e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4944 0.53451 0.16352 0.019236 14.5153 0.11943 0.00015475 0.77073 0.0090567 0.010035 0.001459 0.986 0.99108 3.1558e-006 1.2623e-005 0.16219 0.78859 0.84797 0.0014351 0.91409 0.41308 0.0019319 0.42006 1.8019 1.7998 16.0183 144.9189 0.00026928 -85.3454 0.36295
7.467 0.98812 5.4731e-005 3.8183 0.011937 9.7228e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4945 0.53456 0.16354 0.019237 14.518 0.11943 0.00015476 0.77072 0.0090572 0.010035 0.0014585 0.986 0.99109 3.1545e-006 1.2618e-005 0.16219 0.78919 0.84831 0.0014348 0.91462 0.41328 0.0019315 0.42007 1.8033 1.8011 16.0183 144.9189 0.00026877 -85.3476 0.36395
7.468 0.98812 5.4731e-005 3.8183 0.011937 9.7241e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4946 0.5346 0.16355 0.019238 14.5208 0.11944 0.00015477 0.77071 0.0090576 0.010036 0.0014579 0.98601 0.99109 3.1533e-006 1.2613e-005 0.1622 0.7898 0.84864 0.0014345 0.91514 0.41348 0.0019312 0.42009 1.8046 1.8025 16.0183 144.9189 0.00026826 -85.3499 0.36495
7.469 0.98812 5.4731e-005 3.8183 0.011937 9.7254e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4947 0.53465 0.16356 0.019239 14.5236 0.11945 0.00015478 0.77071 0.009058 0.010036 0.0014574 0.98602 0.9911 3.152e-006 1.2608e-005 0.1622 0.7904 0.84897 0.0014342 0.91565 0.41369 0.0019308 0.4201 1.8059 1.8038 16.0183 144.9189 0.00026775 -85.3522 0.36595
7.47 0.98812 5.4731e-005 3.8183 0.011937 9.7267e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4948 0.53469 0.16358 0.01924 14.5263 0.11945 0.00015479 0.7707 0.0090585 0.010036 0.0014568 0.98603 0.9911 3.1508e-006 1.2603e-005 0.1622 0.79101 0.84931 0.0014339 0.91617 0.41389 0.0019304 0.42011 1.8073 1.8052 16.0183 144.9189 0.00026724 -85.3544 0.36695
7.471 0.98812 5.4731e-005 3.8183 0.011937 9.728e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4949 0.53474 0.16359 0.019242 14.5291 0.11946 0.0001548 0.77069 0.0090589 0.010037 0.0014563 0.98603 0.99111 3.1495e-006 1.2598e-005 0.16221 0.79161 0.84963 0.0014337 0.91668 0.41409 0.0019301 0.42013 1.8086 1.8065 16.0183 144.919 0.00026673 -85.3566 0.36795
7.472 0.98812 5.4731e-005 3.8183 0.011937 9.7293e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4949 0.53478 0.16361 0.019243 14.5319 0.11947 0.00015482 0.77069 0.0090593 0.010037 0.0014557 0.98604 0.99111 3.1483e-006 1.2593e-005 0.16221 0.79221 0.84996 0.0014334 0.91719 0.41429 0.0019297 0.42014 1.8099 1.8078 16.0183 144.919 0.00026623 -85.3588 0.36895
7.473 0.98812 5.4731e-005 3.8183 0.011937 9.7305e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.495 0.53483 0.16362 0.019244 14.5346 0.11948 0.00015483 0.77068 0.0090597 0.010038 0.0014552 0.98605 0.99112 3.1471e-006 1.2588e-005 0.16221 0.7928 0.85029 0.0014331 0.91769 0.4145 0.0019293 0.42015 1.8112 1.8091 16.0183 144.919 0.00026573 -85.361 0.36995
7.474 0.98812 5.473e-005 3.8183 0.011937 9.7318e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4951 0.53487 0.16363 0.019245 14.5374 0.11948 0.00015484 0.77067 0.0090602 0.010038 0.0014547 0.98605 0.99112 3.1459e-006 1.2584e-005 0.16222 0.7934 0.85061 0.0014328 0.91819 0.4147 0.001929 0.42017 1.8125 1.8105 16.0183 144.919 0.00026523 -85.3632 0.37095
7.475 0.98812 5.473e-005 3.8183 0.011937 9.7331e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4952 0.53492 0.16365 0.019246 14.5402 0.11949 0.00015485 0.77066 0.0090606 0.010039 0.0014542 0.98606 0.99113 3.1447e-006 1.2579e-005 0.16222 0.79399 0.85093 0.0014325 0.91869 0.4149 0.0019286 0.42018 1.8139 1.8118 16.0183 144.919 0.00026473 -85.3653 0.37195
7.476 0.98812 5.473e-005 3.8183 0.011937 9.7344e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4953 0.53496 0.16366 0.019247 14.5429 0.1195 0.00015486 0.77066 0.009061 0.010039 0.0014536 0.98607 0.99113 3.1435e-006 1.2574e-005 0.16222 0.79458 0.85126 0.0014323 0.91919 0.4151 0.0019283 0.42019 1.8152 1.8131 16.0184 144.9191 0.00026424 -85.3675 0.37295
7.477 0.98812 5.473e-005 3.8183 0.011937 9.7357e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4954 0.53501 0.16368 0.019249 14.5457 0.1195 0.00015487 0.77065 0.0090614 0.01004 0.0014531 0.98607 0.99113 3.1423e-006 1.2569e-005 0.16223 0.79517 0.85157 0.001432 0.91968 0.4153 0.0019279 0.42021 1.8165 1.8144 16.0184 144.9191 0.00026375 -85.3696 0.37395
7.478 0.98812 5.473e-005 3.8183 0.011937 9.737e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4955 0.53505 0.16369 0.01925 14.5485 0.11951 0.00015488 0.77064 0.0090619 0.01004 0.0014526 0.98608 0.99114 3.1411e-006 1.2565e-005 0.16223 0.79576 0.85189 0.0014317 0.92017 0.41551 0.0019276 0.42022 1.8178 1.8157 16.0184 144.9191 0.00026326 -85.3717 0.37495
7.479 0.98812 5.473e-005 3.8183 0.011937 9.7383e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4956 0.5351 0.1637 0.019251 14.5512 0.11952 0.00015489 0.77064 0.0090623 0.010041 0.0014521 0.98609 0.99114 3.14e-006 1.256e-005 0.16223 0.79634 0.85221 0.0014315 0.92066 0.41571 0.0019272 0.42023 1.8191 1.817 16.0184 144.9191 0.00026277 -85.3738 0.37595
7.48 0.98812 5.473e-005 3.8183 0.011937 9.7395e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4957 0.53515 0.16372 0.019252 14.554 0.11953 0.0001549 0.77063 0.0090627 0.010041 0.0014516 0.98609 0.99115 3.1388e-006 1.2555e-005 0.16224 0.79693 0.85253 0.0014312 0.92114 0.41591 0.0019269 0.42025 1.8204 1.8183 16.0184 144.9191 0.00026228 -85.3759 0.37695
7.481 0.98812 5.473e-005 3.8183 0.011937 9.7408e-005 0.0011696 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4957 0.53519 0.16373 0.019253 14.5568 0.11953 0.00015491 0.77062 0.0090631 0.010041 0.0014511 0.9861 0.99115 3.1377e-006 1.2551e-005 0.16224 0.79751 0.85284 0.001431 0.92162 0.41611 0.0019266 0.42026 1.8217 1.8196 16.0184 144.9192 0.0002618 -85.3779 0.37795
7.482 0.98812 5.473e-005 3.8183 0.011937 9.7421e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4958 0.53524 0.16374 0.019255 14.5595 0.11954 0.00015492 0.77062 0.0090636 0.010042 0.0014506 0.98611 0.99116 3.1365e-006 1.2546e-005 0.16224 0.79809 0.85315 0.0014307 0.9221 0.41631 0.0019262 0.42027 1.8229 1.8209 16.0184 144.9192 0.00026132 -85.38 0.37895
7.483 0.98812 5.473e-005 3.8183 0.011937 9.7434e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4959 0.53528 0.16376 0.019256 14.5623 0.11955 0.00015493 0.77061 0.009064 0.010042 0.0014501 0.98611 0.99116 3.1354e-006 1.2542e-005 0.16225 0.79867 0.85346 0.0014305 0.92257 0.41651 0.0019259 0.42029 1.8242 1.8222 16.0184 144.9192 0.00026084 -85.382 0.37995
7.484 0.98812 5.473e-005 3.8183 0.011937 9.7447e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.496 0.53533 0.16377 0.019257 14.5651 0.11955 0.00015494 0.7706 0.0090644 0.010043 0.0014496 0.98612 0.99117 3.1343e-006 1.2537e-005 0.16225 0.79924 0.85377 0.0014302 0.92305 0.41672 0.0019256 0.4203 1.8255 1.8235 16.0184 144.9192 0.00026036 -85.384 0.38095
7.485 0.98812 5.473e-005 3.8183 0.011937 9.746e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4961 0.53537 0.16379 0.019258 14.5678 0.11956 0.00015495 0.77059 0.0090648 0.010043 0.0014492 0.98613 0.99117 3.1332e-006 1.2533e-005 0.16225 0.79982 0.85408 0.0014299 0.92352 0.41692 0.0019252 0.42031 1.8268 1.8248 16.0184 144.9192 0.00025989 -85.386 0.38195
7.486 0.98812 5.473e-005 3.8183 0.011937 9.7472e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4962 0.53542 0.1638 0.019259 14.5706 0.11957 0.00015496 0.77059 0.0090653 0.010044 0.0014487 0.98613 0.99117 3.1321e-006 1.2528e-005 0.16226 0.80039 0.85439 0.0014297 0.92398 0.41712 0.0019249 0.42033 1.8281 1.8261 16.0184 144.9192 0.00025941 -85.388 0.38295
7.487 0.98812 5.4729e-005 3.8183 0.011937 9.7485e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4963 0.53546 0.16381 0.01926 14.5734 0.11957 0.00015497 0.77058 0.0090657 0.010044 0.0014482 0.98614 0.99118 3.131e-006 1.2524e-005 0.16226 0.80096 0.85469 0.0014295 0.92444 0.41732 0.0019246 0.42034 1.8293 1.8273 16.0184 144.9193 0.00025894 -85.39 0.38395
7.488 0.98812 5.4729e-005 3.8183 0.011937 9.7498e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4964 0.53551 0.16383 0.019262 14.5761 0.11958 0.00015498 0.77057 0.0090661 0.010045 0.0014477 0.98614 0.99118 3.1299e-006 1.252e-005 0.16226 0.80153 0.855 0.0014292 0.92491 0.41752 0.0019243 0.42035 1.8306 1.8286 16.0184 144.9193 0.00025848 -85.3919 0.38495
7.489 0.98812 5.4729e-005 3.8183 0.011937 9.7511e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4964 0.53555 0.16384 0.019263 14.5789 0.11959 0.000155 0.77057 0.0090666 0.010045 0.0014473 0.98615 0.99119 3.1288e-006 1.2515e-005 0.16227 0.8021 0.8553 0.001429 0.92536 0.41772 0.0019239 0.42037 1.8318 1.8299 16.0184 144.9193 0.00025801 -85.3939 0.38595
7.49 0.98812 5.4729e-005 3.8183 0.011937 9.7524e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4965 0.5356 0.16386 0.019264 14.5817 0.1196 0.00015501 0.77056 0.009067 0.010046 0.0014468 0.98616 0.99119 3.1278e-006 1.2511e-005 0.16227 0.80266 0.8556 0.0014288 0.92582 0.41792 0.0019236 0.42038 1.8331 1.8311 16.0184 144.9193 0.00025754 -85.3958 0.38695
7.491 0.98812 5.4729e-005 3.8183 0.011937 9.7537e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4966 0.53564 0.16387 0.019265 14.5844 0.1196 0.00015502 0.77055 0.0090674 0.010046 0.0014463 0.98616 0.99119 3.1267e-006 1.2507e-005 0.16227 0.80323 0.8559 0.0014285 0.92627 0.41813 0.0019233 0.4204 1.8344 1.8324 16.0184 144.9193 0.00025708 -85.3977 0.38795
7.492 0.98812 5.4729e-005 3.8183 0.011937 9.755e-005 0.0011697 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4967 0.53569 0.16388 0.019266 14.5872 0.11961 0.00015503 0.77054 0.0090678 0.010046 0.0014459 0.98617 0.9912 3.1256e-006 1.2503e-005 0.16228 0.80379 0.8562 0.0014283 0.92672 0.41833 0.001923 0.42041 1.8356 1.8337 16.0185 144.9194 0.00025662 -85.3996 0.38895
7.493 0.98812 5.4729e-005 3.8183 0.011937 9.7562e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4968 0.53573 0.1639 0.019267 14.59 0.11962 0.00015504 0.77054 0.0090683 0.010047 0.0014454 0.98618 0.9912 3.1246e-006 1.2498e-005 0.16228 0.80435 0.8565 0.0014281 0.92717 0.41853 0.0019227 0.42042 1.8369 1.8349 16.0185 144.9194 0.00025616 -85.4015 0.38995
7.494 0.98812 5.4729e-005 3.8183 0.011937 9.7575e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4969 0.53578 0.16391 0.019269 14.5928 0.11962 0.00015505 0.77053 0.0090687 0.010047 0.001445 0.98618 0.99121 3.1236e-006 1.2494e-005 0.16228 0.80491 0.8568 0.0014278 0.92761 0.41873 0.0019224 0.42044 1.8381 1.8362 16.0185 144.9194 0.00025571 -85.4034 0.39095
7.495 0.98812 5.4729e-005 3.8183 0.011937 9.7588e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.497 0.53582 0.16393 0.01927 14.5955 0.11963 0.00015506 0.77052 0.0090691 0.010048 0.0014445 0.98619 0.99121 3.1225e-006 1.249e-005 0.16229 0.80546 0.85709 0.0014276 0.92805 0.41893 0.0019221 0.42045 1.8394 1.8374 16.0185 144.9194 0.00025525 -85.4053 0.39195
7.496 0.98812 5.4729e-005 3.8183 0.011937 9.7601e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4971 0.53587 0.16394 0.019271 14.5983 0.11964 0.00015507 0.77052 0.0090695 0.010048 0.0014441 0.98619 0.99121 3.1215e-006 1.2486e-005 0.16229 0.80602 0.85738 0.0014273 0.92849 0.41913 0.0019218 0.42046 1.8406 1.8387 16.0185 144.9194 0.0002548 -85.4071 0.39295
7.497 0.98812 5.4729e-005 3.8183 0.011937 9.7614e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4971 0.53592 0.16395 0.019272 14.6011 0.11965 0.00015508 0.77051 0.00907 0.010049 0.0014436 0.9862 0.99122 3.1205e-006 1.2482e-005 0.16229 0.80657 0.85768 0.0014271 0.92893 0.41933 0.0019215 0.42048 1.8418 1.8399 16.0185 144.9194 0.00025435 -85.409 0.39395
7.498 0.98812 5.4729e-005 3.8183 0.011937 9.7627e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4972 0.53596 0.16397 0.019273 14.6038 0.11965 0.00015509 0.7705 0.0090704 0.010049 0.0014432 0.9862 0.99122 3.1195e-006 1.2478e-005 0.1623 0.80713 0.85797 0.0014269 0.92936 0.41953 0.0019212 0.42049 1.8431 1.8411 16.0185 144.9195 0.0002539 -85.4108 0.39495
7.499 0.98812 5.4728e-005 3.8183 0.011937 9.764e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4973 0.53601 0.16398 0.019274 14.6066 0.11966 0.0001551 0.7705 0.0090708 0.01005 0.0014427 0.98621 0.99122 3.1185e-006 1.2474e-005 0.1623 0.80768 0.85826 0.0014266 0.92979 0.41973 0.0019209 0.42051 1.8443 1.8424 16.0185 144.9195 0.00025345 -85.4126 0.39595
7.5 0.98812 5.4728e-005 3.8183 0.011937 9.7652e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4974 0.53605 0.164 0.019276 14.6094 0.11967 0.00015511 0.77049 0.0090712 0.01005 0.0014423 0.98622 0.99123 3.1175e-006 1.247e-005 0.1623 0.80822 0.85854 0.0014264 0.93022 0.41993 0.0019206 0.42052 1.8455 1.8436 16.0185 144.9195 0.00025301 -85.4144 0.39695
7.501 0.98812 5.4728e-005 3.8183 0.011937 9.7665e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4975 0.5361 0.16401 0.019277 14.6122 0.11967 0.00015512 0.77048 0.0090717 0.010051 0.0014419 0.98622 0.99123 3.1165e-006 1.2466e-005 0.16231 0.80877 0.85883 0.0014262 0.93064 0.42013 0.0019203 0.42053 1.8467 1.8448 16.0185 144.9195 0.00025257 -85.4162 0.39795
7.502 0.98812 5.4728e-005 3.8183 0.011937 9.7678e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4976 0.53614 0.16402 0.019278 14.6149 0.11968 0.00015513 0.77047 0.0090721 0.010051 0.0014415 0.98623 0.99124 3.1155e-006 1.2462e-005 0.16231 0.80932 0.85912 0.001426 0.93106 0.42033 0.00192 0.42055 1.8479 1.8461 16.0185 144.9195 0.00025213 -85.4179 0.39895
7.503 0.98812 5.4728e-005 3.8183 0.011937 9.7691e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4977 0.53619 0.16404 0.019279 14.6177 0.11969 0.00015514 0.77047 0.0090725 0.010051 0.001441 0.98623 0.99124 3.1146e-006 1.2458e-005 0.16231 0.80986 0.8594 0.0014258 0.93148 0.42054 0.0019197 0.42056 1.8492 1.8473 16.0185 144.9196 0.00025169 -85.4197 0.39995
7.504 0.98812 5.4728e-005 3.8183 0.011937 9.7704e-005 0.0011697 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4978 0.53623 0.16405 0.01928 14.6205 0.11969 0.00015515 0.77046 0.0090729 0.010052 0.0014406 0.98624 0.99124 3.1136e-006 1.2454e-005 0.16232 0.8104 0.85969 0.0014255 0.9319 0.42074 0.0019194 0.42057 1.8504 1.8485 16.0185 144.9196 0.00025125 -85.4214 0.40095
7.505 0.98812 5.4728e-005 3.8183 0.011937 9.7717e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4979 0.53628 0.16407 0.019282 14.6233 0.1197 0.00015516 0.77045 0.0090734 0.010052 0.0014402 0.98624 0.99125 3.1127e-006 1.2451e-005 0.16232 0.81094 0.85997 0.0014253 0.93232 0.42094 0.0019192 0.42059 1.8516 1.8497 16.0185 144.9196 0.00025081 -85.4232 0.40195
7.506 0.98812 5.4728e-005 3.8183 0.011937 9.7729e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4979 0.53632 0.16408 0.019283 14.626 0.11971 0.00015517 0.77045 0.0090738 0.010053 0.0014398 0.98625 0.99125 3.1117e-006 1.2447e-005 0.16232 0.81148 0.86025 0.0014251 0.93273 0.42114 0.0019189 0.4206 1.8528 1.8509 16.0185 144.9196 0.00025038 -85.4249 0.40295
7.507 0.98812 5.4728e-005 3.8183 0.011936 9.7742e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.498 0.53637 0.16409 0.019284 14.6288 0.11972 0.00015519 0.77044 0.0090742 0.010053 0.0014394 0.98625 0.99125 3.1108e-006 1.2443e-005 0.16233 0.81202 0.86053 0.0014249 0.93314 0.42134 0.0019186 0.42062 1.854 1.8521 16.0185 144.9196 0.00024995 -85.4266 0.40395
7.508 0.98812 5.4728e-005 3.8183 0.011936 9.7755e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4981 0.53641 0.16411 0.019285 14.6316 0.11972 0.0001552 0.77043 0.0090746 0.010054 0.001439 0.98626 0.99126 3.1098e-006 1.2439e-005 0.16233 0.81255 0.86081 0.0014247 0.93355 0.42154 0.0019183 0.42063 1.8552 1.8533 16.0185 144.9197 0.00024952 -85.4283 0.40495
7.509 0.98812 5.4728e-005 3.8183 0.011936 9.7768e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4982 0.53646 0.16412 0.019286 14.6344 0.11973 0.00015521 0.77043 0.0090751 0.010054 0.0014386 0.98626 0.99126 3.1089e-006 1.2436e-005 0.16233 0.81308 0.86108 0.0014245 0.93395 0.42174 0.0019181 0.42064 1.8564 1.8545 16.0185 144.9197 0.00024909 -85.43 0.40595
7.51 0.98812 5.4728e-005 3.8183 0.011936 9.7781e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4983 0.5365 0.16414 0.019287 14.6371 0.11974 0.00015522 0.77042 0.0090755 0.010055 0.0014382 0.98627 0.99126 3.108e-006 1.2432e-005 0.16234 0.81362 0.86136 0.0014243 0.93435 0.42194 0.0019178 0.42066 1.8576 1.8557 16.0185 144.9197 0.00024867 -85.4316 0.40695
7.511 0.98812 5.4728e-005 3.8183 0.011936 9.7794e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4984 0.53655 0.16415 0.019289 14.6399 0.11974 0.00015523 0.77041 0.0090759 0.010055 0.0014378 0.98628 0.99127 3.1071e-006 1.2428e-005 0.16234 0.81415 0.86163 0.0014241 0.93475 0.42214 0.0019175 0.42067 1.8588 1.8569 16.0185 144.9197 0.00024824 -85.4333 0.40795
7.512 0.98812 5.4727e-005 3.8183 0.011936 9.7807e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4985 0.53659 0.16416 0.01929 14.6427 0.11975 0.00015524 0.7704 0.0090763 0.010056 0.0014374 0.98628 0.99127 3.1062e-006 1.2425e-005 0.16234 0.81467 0.86191 0.0014239 0.93515 0.42234 0.0019172 0.42069 1.8599 1.8581 16.0185 144.9197 0.00024782 -85.4349 0.40895
7.513 0.98812 5.4727e-005 3.8183 0.011936 9.7819e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4986 0.53664 0.16418 0.019291 14.6455 0.11976 0.00015525 0.7704 0.0090768 0.010056 0.001437 0.98629 0.99127 3.1053e-006 1.2421e-005 0.16235 0.8152 0.86218 0.0014237 0.93554 0.42254 0.001917 0.4207 1.8611 1.8593 16.0185 144.9197 0.0002474 -85.4366 0.40995
7.514 0.98812 5.4727e-005 3.8183 0.011936 9.7832e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4986 0.53669 0.16419 0.019292 14.6482 0.11977 0.00015526 0.77039 0.0090772 0.010056 0.0014366 0.98629 0.99128 3.1044e-006 1.2418e-005 0.16235 0.81573 0.86245 0.0014235 0.93594 0.42274 0.0019167 0.42071 1.8623 1.8605 16.0185 144.9198 0.00024698 -85.4382 0.41095
7.515 0.98812 5.4727e-005 3.8183 0.011936 9.7845e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4987 0.53673 0.16421 0.019293 14.651 0.11977 0.00015527 0.77038 0.0090776 0.010057 0.0014362 0.9863 0.99128 3.1035e-006 1.2414e-005 0.16235 0.81625 0.86272 0.0014233 0.93633 0.42294 0.0019165 0.42073 1.8635 1.8617 16.0185 144.9198 0.00024657 -85.4398 0.41195
7.516 0.98812 5.4727e-005 3.8183 0.011936 9.7858e-005 0.0011698 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.4988 0.53678 0.16422 0.019294 14.6538 0.11978 0.00015528 0.77038 0.009078 0.010057 0.0014358 0.9863 0.99128 3.1026e-006 1.2411e-005 0.16236 0.81677 0.86299 0.0014231 0.93671 0.42314 0.0019162 0.42074 1.8646 1.8628 16.0185 144.9198 0.00024615 -85.4414 0.41295
7.517 0.98812 5.4727e-005 3.8183 0.011936 9.7871e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4989 0.53682 0.16423 0.019296 14.6566 0.11979 0.00015529 0.77037 0.0090784 0.010058 0.0014355 0.98631 0.99129 3.1018e-006 1.2407e-005 0.16236 0.81729 0.86326 0.0014229 0.9371 0.42334 0.0019159 0.42076 1.8658 1.864 16.0185 144.9198 0.00024574 -85.443 0.41395
7.518 0.98812 5.4727e-005 3.8183 0.011936 9.7884e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.499 0.53687 0.16425 0.019297 14.6594 0.11979 0.0001553 0.77036 0.0090789 0.010058 0.0014351 0.98631 0.99129 3.1009e-006 1.2404e-005 0.16236 0.81781 0.86352 0.0014227 0.93748 0.42354 0.0019157 0.42077 1.867 1.8652 16.0185 144.9198 0.00024533 -85.4446 0.41495
7.519 0.98812 5.4727e-005 3.8183 0.011936 9.7896e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4991 0.53691 0.16426 0.019298 14.6621 0.1198 0.00015531 0.77035 0.0090793 0.010059 0.0014347 0.98632 0.99129 3.1e-006 1.24e-005 0.16237 0.81833 0.86379 0.0014225 0.93786 0.42374 0.0019154 0.42078 1.8681 1.8664 16.0185 144.9199 0.00024492 -85.4461 0.41595
7.52 0.98812 5.4727e-005 3.8183 0.011936 9.7909e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4992 0.53696 0.16427 0.019299 14.6649 0.11981 0.00015532 0.77035 0.0090797 0.010059 0.0014343 0.98632 0.9913 3.0992e-006 1.2397e-005 0.16237 0.81884 0.86405 0.0014223 0.93824 0.42393 0.0019152 0.4208 1.8693 1.8675 16.0185 144.9199 0.00024451 -85.4477 0.41695
7.521 0.98812 5.4727e-005 3.8183 0.011936 9.7922e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4993 0.537 0.16429 0.0193 14.6677 0.11981 0.00015533 0.77034 0.0090801 0.01006 0.001434 0.98633 0.9913 3.0983e-006 1.2393e-005 0.16237 0.81936 0.86431 0.0014221 0.93862 0.42413 0.0019149 0.42081 1.8705 1.8687 16.0185 144.9199 0.0002441 -85.4492 0.41795
7.522 0.98812 5.4727e-005 3.8183 0.011936 9.7935e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4993 0.53705 0.1643 0.019301 14.6705 0.11982 0.00015534 0.77033 0.0090806 0.01006 0.0014336 0.98633 0.9913 3.0975e-006 1.239e-005 0.16238 0.81987 0.86458 0.0014219 0.93899 0.42433 0.0019147 0.42083 1.8716 1.8698 16.0185 144.9199 0.0002437 -85.4508 0.41895
7.523 0.98812 5.4727e-005 3.8183 0.011936 9.7948e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4994 0.53709 0.16432 0.019303 14.6733 0.11983 0.00015535 0.77033 0.009081 0.01006 0.0014332 0.98633 0.99131 3.0967e-006 1.2387e-005 0.16238 0.82038 0.86484 0.0014217 0.93936 0.42453 0.0019144 0.42084 1.8728 1.871 16.0185 144.9199 0.0002433 -85.4523 0.41995
7.524 0.98812 5.4726e-005 3.8183 0.011936 9.7961e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4995 0.53714 0.16433 0.019304 14.676 0.11984 0.00015536 0.77032 0.0090814 0.010061 0.0014329 0.98634 0.99131 3.0958e-006 1.2383e-005 0.16238 0.82089 0.8651 0.0014215 0.93973 0.42473 0.0019142 0.42085 1.8739 1.8721 16.0185 144.92 0.0002429 -85.4538 0.42095
7.525 0.98812 5.4726e-005 3.8183 0.011936 9.7974e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4996 0.53718 0.16434 0.019305 14.6788 0.11984 0.00015538 0.77031 0.0090818 0.010061 0.0014325 0.98634 0.99131 3.095e-006 1.238e-005 0.16239 0.82139 0.86536 0.0014213 0.94009 0.42493 0.0019139 0.42087 1.8751 1.8733 16.0185 144.92 0.0002425 -85.4553 0.42195
7.526 0.98812 5.4726e-005 3.8183 0.011936 9.7986e-005 0.0011698 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4997 0.53723 0.16436 0.019306 14.6816 0.11985 0.00015539 0.77031 0.0090823 0.010062 0.0014322 0.98635 0.99132 3.0942e-006 1.2377e-005 0.16239 0.8219 0.86561 0.0014211 0.94046 0.42513 0.0019137 0.42088 1.8762 1.8744 16.0185 144.92 0.0002421 -85.4568 0.42295
7.527 0.98812 5.4726e-005 3.8183 0.011936 9.7999e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4998 0.53727 0.16437 0.019307 14.6844 0.11986 0.0001554 0.7703 0.0090827 0.010062 0.0014318 0.98635 0.99132 3.0934e-006 1.2374e-005 0.16239 0.8224 0.86587 0.0014209 0.94082 0.42533 0.0019134 0.4209 1.8773 1.8756 16.0185 144.92 0.00024171 -85.4582 0.42395
7.528 0.98812 5.4726e-005 3.8183 0.011936 9.8012e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.4999 0.53732 0.16439 0.019309 14.6872 0.11986 0.00015541 0.77029 0.0090831 0.010063 0.0014315 0.98636 0.99132 3.0926e-006 1.237e-005 0.1624 0.82291 0.86612 0.0014208 0.94118 0.42553 0.0019132 0.42091 1.8785 1.8767 16.0185 144.92 0.00024131 -85.4597 0.42495
7.529 0.98812 5.4726e-005 3.8183 0.011936 9.8025e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5 0.53736 0.1644 0.01931 14.69 0.11987 0.00015542 0.77028 0.0090835 0.010063 0.0014311 0.98636 0.99133 3.0918e-006 1.2367e-005 0.1624 0.82341 0.86638 0.0014206 0.94154 0.42573 0.001913 0.42093 1.8796 1.8779 16.0185 144.92 0.00024092 -85.4612 0.42595
7.53 0.98812 5.4726e-005 3.8183 0.011936 9.8038e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5001 0.53741 0.16441 0.019311 14.6927 0.11988 0.00015543 0.77028 0.0090839 0.010064 0.0014308 0.98637 0.99133 3.091e-006 1.2364e-005 0.1624 0.82391 0.86663 0.0014204 0.94189 0.42593 0.0019127 0.42094 1.8807 1.879 16.0185 144.9201 0.00024053 -85.4626 0.42695
7.531 0.98812 5.4726e-005 3.8183 0.011936 9.8051e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5001 0.53746 0.16443 0.019312 14.6955 0.11989 0.00015544 0.77027 0.0090844 0.010064 0.0014304 0.98637 0.99133 3.0902e-006 1.2361e-005 0.1624 0.82441 0.86688 0.0014203 0.94225 0.42613 0.0019125 0.42095 1.8818 1.8801 16.0185 144.9201 0.00024014 -85.464 0.42795
7.532 0.98812 5.4726e-005 3.8183 0.011936 9.8063e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5002 0.5375 0.16444 0.019313 14.6983 0.11989 0.00015545 0.77026 0.0090848 0.010065 0.0014301 0.98638 0.99133 3.0894e-006 1.2358e-005 0.16241 0.8249 0.86713 0.0014201 0.9426 0.42632 0.0019123 0.42097 1.883 1.8813 16.0185 144.9201 0.00023975 -85.4655 0.42895
7.533 0.98813 5.4726e-005 3.8183 0.011936 9.8076e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5003 0.53755 0.16446 0.019314 14.7011 0.1199 0.00015546 0.77026 0.0090852 0.010065 0.0014297 0.98638 0.99134 3.0887e-006 1.2355e-005 0.16241 0.8254 0.86738 0.0014199 0.94294 0.42652 0.001912 0.42098 1.8841 1.8824 16.0185 144.9201 0.00023937 -85.4669 0.42995
7.534 0.98813 5.4726e-005 3.8183 0.011936 9.8089e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5004 0.53759 0.16447 0.019316 14.7039 0.11991 0.00015547 0.77025 0.0090856 0.010065 0.0014294 0.98638 0.99134 3.0879e-006 1.2352e-005 0.16241 0.82589 0.86763 0.0014197 0.94329 0.42672 0.0019118 0.421 1.8852 1.8835 16.0185 144.9201 0.00023898 -85.4683 0.43095
7.535 0.98813 5.4726e-005 3.8183 0.011936 9.8102e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5005 0.53764 0.16448 0.019317 14.7067 0.11991 0.00015548 0.77024 0.0090861 0.010066 0.0014291 0.98639 0.99134 3.0871e-006 1.2349e-005 0.16242 0.82638 0.86788 0.0014195 0.94363 0.42692 0.0019116 0.42101 1.8863 1.8846 16.0185 144.9202 0.0002386 -85.4697 0.43195
7.536 0.98813 5.4725e-005 3.8183 0.011936 9.8115e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5006 0.53768 0.1645 0.019318 14.7094 0.11992 0.00015549 0.77024 0.0090865 0.010066 0.0014287 0.98639 0.99135 3.0864e-006 1.2346e-005 0.16242 0.82687 0.86813 0.0014193 0.94398 0.42712 0.0019114 0.42103 1.8874 1.8857 16.0185 144.9202 0.00023822 -85.4711 0.43295
7.537 0.98813 5.4725e-005 3.8183 0.011936 9.8128e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5007 0.53773 0.16451 0.019319 14.7122 0.11993 0.0001555 0.77023 0.0090869 0.010067 0.0014284 0.9864 0.99135 3.0856e-006 1.2343e-005 0.16242 0.82736 0.86837 0.0014192 0.94432 0.42732 0.0019111 0.42104 1.8885 1.8868 16.0185 144.9202 0.00023784 -85.4724 0.43395
7.538 0.98813 5.4725e-005 3.8183 0.011936 9.8141e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5008 0.53777 0.16453 0.01932 14.715 0.11993 0.00015551 0.77022 0.0090873 0.010067 0.0014281 0.9864 0.99135 3.0849e-006 1.234e-005 0.16243 0.82785 0.86861 0.001419 0.94465 0.42752 0.0019109 0.42105 1.8896 1.888 16.0185 144.9202 0.00023746 -85.4738 0.43495
7.539 0.98813 5.4725e-005 3.8183 0.011936 9.8153e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5008 0.53782 0.16454 0.019321 14.7178 0.11994 0.00015552 0.77021 0.0090878 0.010068 0.0014278 0.98641 0.99135 3.0841e-006 1.2337e-005 0.16243 0.82833 0.86886 0.0014189 0.94499 0.42771 0.0019107 0.42107 1.8907 1.8891 16.0185 144.9202 0.00023709 -85.4752 0.43595
7.54 0.98813 5.4725e-005 3.8183 0.011936 9.8166e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5009 0.53786 0.16455 0.019323 14.7206 0.11995 0.00015553 0.77021 0.0090882 0.010068 0.0014274 0.98641 0.99136 3.0834e-006 1.2334e-005 0.16243 0.82882 0.8691 0.0014188 0.94532 0.42791 0.0019105 0.42108 1.8918 1.8902 16.0185 144.9203 0.00023671 -85.4765 0.43695
7.541 0.98813 5.4725e-005 3.8183 0.011936 9.8179e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.501 0.53791 0.16457 0.019324 14.7234 0.11996 0.00015554 0.7702 0.0090886 0.010069 0.0014271 0.98641 0.99136 3.0827e-006 1.2331e-005 0.16244 0.8293 0.86934 0.0014186 0.94566 0.42811 0.0019103 0.4211 1.8929 1.8913 16.0185 144.9203 0.00023634 -85.4778 0.43795
7.542 0.98813 5.4725e-005 3.8183 0.011936 9.8192e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5011 0.53795 0.16458 0.019325 14.7262 0.11996 0.00015555 0.77019 0.009089 0.010069 0.0014268 0.98642 0.99136 3.0819e-006 1.2328e-005 0.16244 0.82978 0.86958 0.0014184 0.94598 0.42831 0.0019101 0.42111 1.894 1.8924 16.0185 144.9203 0.00023597 -85.4792 0.43895
7.543 0.98813 5.4725e-005 3.8183 0.011936 9.8205e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5012 0.538 0.1646 0.019326 14.729 0.11997 0.00015556 0.77019 0.0090894 0.01007 0.0014265 0.98642 0.99136 3.0812e-006 1.2325e-005 0.16244 0.83026 0.86982 0.0014182 0.94631 0.42851 0.0019098 0.42112 1.8951 1.8934 16.0185 144.9203 0.0002356 -85.4805 0.43995
7.544 0.98813 5.4725e-005 3.8183 0.011936 9.8218e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5013 0.53804 0.16461 0.019327 14.7317 0.11998 0.00015558 0.77018 0.0090899 0.01007 0.0014262 0.98643 0.99137 3.0805e-006 1.2322e-005 0.16245 0.83074 0.87006 0.001418 0.94664 0.42871 0.0019096 0.42114 1.8962 1.8945 16.0185 144.9203 0.00023523 -85.4818 0.44095
7.545 0.98813 5.4725e-005 3.8183 0.011936 9.823e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5014 0.53809 0.16462 0.019328 14.7345 0.11998 0.00015559 0.77017 0.0090903 0.01007 0.0014259 0.98643 0.99137 3.0798e-006 1.2319e-005 0.16245 0.83122 0.8703 0.0014178 0.94696 0.4289 0.0019094 0.42115 1.8973 1.8956 16.0185 144.9204 0.00023487 -85.4831 0.44195
7.546 0.98813 5.4725e-005 3.8183 0.011936 9.8243e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5015 0.53813 0.16464 0.01933 14.7373 0.11999 0.0001556 0.77017 0.0090907 0.010071 0.0014256 0.98643 0.99137 3.0792e-006 1.2317e-005 0.16245 0.83169 0.87053 0.0014176 0.94728 0.4291 0.0019092 0.42117 1.8983 1.8967 16.0185 144.9204 0.0002345 -85.4844 0.44295
7.547 0.98813 5.4725e-005 3.8183 0.011936 9.8256e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5015 0.53818 0.16465 0.019331 14.7401 0.12 0.00015561 0.77016 0.0090911 0.010071 0.0014253 0.98644 0.99138 3.0784e-006 1.2314e-005 0.16246 0.83217 0.87077 0.0014175 0.9476 0.4293 0.001909 0.42118 1.8994 1.8978 16.0185 144.9204 0.00023414 -85.4856 0.44395
7.548 0.98813 5.4725e-005 3.8183 0.011936 9.8269e-005 0.0011699 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5016 0.53822 0.16466 0.019332 14.7429 0.12 0.00015562 0.77015 0.0090916 0.010072 0.001425 0.98644 0.99138 3.0777e-006 1.2311e-005 0.16246 0.83264 0.871 0.0014174 0.94792 0.4295 0.0019088 0.4212 1.9005 1.8989 16.0185 144.9204 0.00023378 -85.4869 0.44495
7.549 0.98813 5.4724e-005 3.8183 0.011936 9.8282e-005 0.00117 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5017 0.53827 0.16468 0.019333 14.7457 0.12001 0.00015563 0.77014 0.009092 0.010072 0.0014247 0.98645 0.99138 3.077e-006 1.2308e-005 0.16246 0.83311 0.87124 0.0014173 0.94823 0.42969 0.0019086 0.42121 1.9016 1.8999 16.0185 144.9204 0.00023342 -85.4882 0.44595
7.55 0.98813 5.4724e-005 3.8183 0.011936 9.8295e-005 0.00117 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5018 0.53832 0.16469 0.019334 14.7485 0.12002 0.00015564 0.77014 0.0090924 0.010073 0.0014244 0.98645 0.99138 3.0763e-006 1.2305e-005 0.16247 0.83358 0.87147 0.0014173 0.94855 0.42989 0.0019084 0.42123 1.9026 1.901 16.0185 144.9205 0.00023306 -85.4894 0.44695
7.551 0.98813 5.4724e-005 3.8183 0.011936 9.8308e-005 0.00117 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5019 0.53836 0.16471 0.019335 14.7513 0.12003 0.00015565 0.77013 0.0090928 0.010073 0.0014241 0.98645 0.99139 3.0757e-006 1.2303e-005 0.16247 0.83405 0.8717 0.0014172 0.94886 0.43009 0.0019082 0.42124 1.9037 1.9021 16.0185 144.9205 0.0002327 -85.4907 0.44795
7.552 0.98813 5.4724e-005 3.8183 0.011936 9.832e-005 0.00117 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.502 0.53841 0.16472 0.019337 14.7541 0.12003 0.00015566 0.77012 0.0090932 0.010074 0.0014238 0.98646 0.99139 3.075e-006 1.23e-005 0.16247 0.83451 0.87193 0.0014171 0.94917 0.43029 0.001908 0.42125 1.9048 1.9032 16.0185 144.9205 0.00023235 -85.4919 0.44895
7.553 0.98813 5.4724e-005 3.8183 0.011936 9.8333e-005 0.00117 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5021 0.53845 0.16473 0.019338 14.7569 0.12004 0.00015567 0.77012 0.0090937 0.010074 0.0014235 0.98646 0.99139 3.0743e-006 1.2297e-005 0.16248 0.83498 0.87216 0.0014169 0.94947 0.43049 0.0019078 0.42127 1.9058 1.9042 16.0185 144.9205 0.00023199 -85.4931 0.44995
7.554 0.98813 5.4724e-005 3.8183 0.011936 9.8346e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5022 0.5385 0.16475 0.019339 14.7596 0.12005 0.00015568 0.77011 0.0090941 0.010074 0.0014232 0.98647 0.99139 3.0737e-006 1.2295e-005 0.16248 0.83544 0.87239 0.0014167 0.94978 0.43068 0.0019076 0.42128 1.9069 1.9053 16.0185 144.9205 0.00023164 -85.4943 0.45095
7.555 0.98813 5.4724e-005 3.8183 0.011936 9.8359e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5023 0.53854 0.16476 0.01934 14.7624 0.12005 0.00015569 0.7701 0.0090945 0.010075 0.0014229 0.98647 0.9914 3.073e-006 1.2292e-005 0.16248 0.8359 0.87261 0.0014165 0.95008 0.43088 0.0019074 0.4213 1.9079 1.9063 16.0184 144.9205 0.00023129 -85.4955 0.45195
7.556 0.98813 5.4724e-005 3.8183 0.011936 9.8372e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5023 0.53859 0.16478 0.019341 14.7652 0.12006 0.0001557 0.7701 0.0090949 0.010075 0.0014226 0.98647 0.9914 3.0724e-006 1.2289e-005 0.16249 0.83636 0.87284 0.0014163 0.95039 0.43108 0.0019072 0.42131 1.909 1.9074 16.0184 144.9206 0.00023094 -85.4967 0.45295
7.557 0.98813 5.4724e-005 3.8183 0.011936 9.8385e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5024 0.53863 0.16479 0.019342 14.768 0.12007 0.00015571 0.77009 0.0090953 0.010076 0.0014224 0.98648 0.9914 3.0717e-006 1.2287e-005 0.16249 0.83682 0.87307 0.0014161 0.95068 0.43127 0.001907 0.42133 1.91 1.9084 16.0184 144.9206 0.00023059 -85.4979 0.45395
7.558 0.98813 5.4724e-005 3.8183 0.011936 9.8397e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5025 0.53868 0.1648 0.019344 14.7708 0.12007 0.00015572 0.77008 0.0090958 0.010076 0.0014221 0.98648 0.9914 3.0711e-006 1.2284e-005 0.16249 0.83728 0.87329 0.001416 0.95098 0.43147 0.0019068 0.42134 1.9111 1.9095 16.0184 144.9206 0.00023024 -85.4991 0.45495
7.559 0.98813 5.4724e-005 3.8183 0.011936 9.841e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5026 0.53872 0.16482 0.019345 14.7736 0.12008 0.00015573 0.77007 0.0090962 0.010077 0.0014218 0.98648 0.9914 3.0705e-006 1.2282e-005 0.1625 0.83774 0.87351 0.0014158 0.95128 0.43167 0.0019066 0.42135 1.9121 1.9105 16.0184 144.9206 0.0002299 -85.5003 0.45595
7.56 0.98813 5.4724e-005 3.8183 0.011936 9.8423e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5027 0.53877 0.16483 0.019346 14.7764 0.12009 0.00015574 0.77007 0.0090966 0.010077 0.0014215 0.98649 0.99141 3.0698e-006 1.2279e-005 0.1625 0.83819 0.87374 0.0014156 0.95157 0.43187 0.0019064 0.42137 1.9131 1.9116 16.0184 144.9206 0.00022955 -85.5014 0.45695
7.561 0.98813 5.4723e-005 3.8183 0.011936 9.8436e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5028 0.53881 0.16485 0.019347 14.7792 0.1201 0.00015575 0.77006 0.009097 0.010078 0.0014213 0.98649 0.99141 3.0692e-006 1.2277e-005 0.1625 0.83865 0.87396 0.0014154 0.95187 0.43206 0.0019063 0.42138 1.9142 1.9126 16.0184 144.9207 0.00022921 -85.5026 0.45795
7.562 0.98813 5.4723e-005 3.8183 0.011936 9.8449e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5029 0.53886 0.16486 0.019348 14.782 0.1201 0.00015576 0.77005 0.0090975 0.010078 0.001421 0.98649 0.99141 3.0686e-006 1.2274e-005 0.16251 0.8391 0.87418 0.0014152 0.95216 0.43226 0.0019061 0.4214 1.9152 1.9137 16.0184 144.9207 0.00022887 -85.5037 0.45895
7.563 0.98813 5.4723e-005 3.8183 0.011936 9.8462e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.503 0.5389 0.16487 0.019349 14.7848 0.12011 0.00015577 0.77005 0.0090979 0.010079 0.0014207 0.9865 0.99141 3.068e-006 1.2272e-005 0.16251 0.83955 0.8744 0.0014151 0.95244 0.43246 0.0019059 0.42141 1.9162 1.9147 16.0184 144.9207 0.00022853 -85.5049 0.45995
7.564 0.98813 5.4723e-005 3.8183 0.011936 9.8475e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.503 0.53895 0.16489 0.019351 14.7876 0.12012 0.00015579 0.77004 0.0090983 0.010079 0.0014204 0.9865 0.99142 3.0674e-006 1.2269e-005 0.16251 0.84 0.87462 0.001415 0.95273 0.43265 0.0019057 0.42143 1.9173 1.9157 16.0184 144.9207 0.00022819 -85.506 0.46095
7.565 0.98813 5.4723e-005 3.8183 0.011935 9.8487e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5031 0.53899 0.1649 0.019352 14.7904 0.12012 0.0001558 0.77003 0.0090987 0.010079 0.0014202 0.9865 0.99142 3.0668e-006 1.2267e-005 0.16252 0.84045 0.87484 0.0014148 0.95302 0.43285 0.0019055 0.42144 1.9183 1.9168 16.0184 144.9207 0.00022785 -85.5071 0.46195
7.566 0.98813 5.4723e-005 3.8183 0.011935 9.85e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5032 0.53904 0.16492 0.019353 14.7932 0.12013 0.00015581 0.77003 0.0090991 0.01008 0.0014199 0.98651 0.99142 3.0661e-006 1.2265e-005 0.16252 0.84089 0.87505 0.0014147 0.9533 0.43305 0.0019053 0.42146 1.9193 1.9178 16.0184 144.9208 0.00022752 -85.5082 0.46295
7.567 0.98813 5.4723e-005 3.8183 0.011935 9.8513e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5033 0.53908 0.16493 0.019354 14.796 0.12014 0.00015582 0.77002 0.0090996 0.01008 0.0014197 0.98651 0.99142 3.0655e-006 1.2262e-005 0.16252 0.84134 0.87527 0.0014146 0.95358 0.43324 0.0019052 0.42147 1.9203 1.9188 16.0184 144.9208 0.00022719 -85.5094 0.46395
7.568 0.98813 5.4723e-005 3.8183 0.011935 9.8526e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5034 0.53913 0.16494 0.019355 14.7988 0.12014 0.00015583 0.77001 0.0091 0.010081 0.0014194 0.98652 0.99143 3.0649e-006 1.226e-005 0.16253 0.84178 0.87548 0.0014145 0.95386 0.43344 0.001905 0.42148 1.9214 1.9198 16.0184 144.9208 0.00022685 -85.5105 0.46495
7.569 0.98813 5.4723e-005 3.8183 0.011935 9.8539e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5035 0.53918 0.16496 0.019356 14.8016 0.12015 0.00015584 0.77 0.0091004 0.010081 0.0014191 0.98652 0.99143 3.0643e-006 1.2257e-005 0.16253 0.84222 0.8757 0.0014144 0.95414 0.43364 0.0019048 0.4215 1.9224 1.9208 16.0184 144.9208 0.00022652 -85.5115 0.46595
7.57 0.98813 5.4723e-005 3.8183 0.011935 9.8552e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5036 0.53922 0.16497 0.019358 14.8044 0.12016 0.00015585 0.77 0.0091008 0.010082 0.0014189 0.98652 0.99143 3.0638e-006 1.2255e-005 0.16253 0.84267 0.87591 0.0014143 0.95441 0.43383 0.0019046 0.42151 1.9234 1.9219 16.0184 144.9208 0.00022619 -85.5126 0.46695
7.571 0.98813 5.4723e-005 3.8183 0.011935 9.8564e-005 0.00117 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5037 0.53927 0.16498 0.019359 14.8072 0.12017 0.00015586 0.76999 0.0091012 0.010082 0.0014186 0.98653 0.99143 3.0632e-006 1.2253e-005 0.16254 0.84311 0.87612 0.0014141 0.95469 0.43403 0.0019045 0.42153 1.9244 1.9229 16.0184 144.9209 0.00022586 -85.5137 0.46795
7.572 0.98813 5.4723e-005 3.8183 0.011935 9.8577e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5037 0.53931 0.165 0.01936 14.81 0.12017 0.00015587 0.76998 0.0091017 0.010083 0.0014184 0.98653 0.99143 3.0626e-006 1.225e-005 0.16254 0.84354 0.87634 0.001414 0.95496 0.43423 0.0019043 0.42154 1.9254 1.9239 16.0184 144.9209 0.00022554 -85.5148 0.46895
7.573 0.98813 5.4722e-005 3.8183 0.011935 9.859e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5038 0.53936 0.16501 0.019361 14.8128 0.12018 0.00015588 0.76998 0.0091021 0.010083 0.0014181 0.98653 0.99144 3.062e-006 1.2248e-005 0.16254 0.84398 0.87655 0.0014139 0.95523 0.43442 0.0019041 0.42156 1.9264 1.9249 16.0183 144.9209 0.00022521 -85.5158 0.46995
7.574 0.98813 5.4722e-005 3.8183 0.011935 9.8603e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5039 0.5394 0.16503 0.019362 14.8155 0.12019 0.00015589 0.76997 0.0091025 0.010083 0.0014179 0.98653 0.99144 3.0615e-006 1.2246e-005 0.16255 0.84442 0.87676 0.0014137 0.9555 0.43462 0.0019039 0.42157 1.9274 1.9259 16.0183 144.9209 0.00022489 -85.5169 0.47095
7.575 0.98813 5.4722e-005 3.8183 0.011935 9.8616e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.504 0.53945 0.16504 0.019363 14.8183 0.12019 0.0001559 0.76996 0.0091029 0.010084 0.0014176 0.98654 0.99144 3.0609e-006 1.2244e-005 0.16255 0.84485 0.87697 0.0014136 0.95577 0.43482 0.0019038 0.42159 1.9284 1.9269 16.0183 144.9209 0.00022456 -85.5179 0.47195
7.576 0.98813 5.4722e-005 3.8183 0.011935 9.8629e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5041 0.53949 0.16505 0.019365 14.8211 0.1202 0.00015591 0.76996 0.0091033 0.010084 0.0014174 0.98654 0.99144 3.0603e-006 1.2241e-005 0.16255 0.84528 0.87717 0.0014134 0.95603 0.43501 0.0019036 0.4216 1.9294 1.9279 16.0183 144.921 0.00022424 -85.519 0.47295
7.577 0.98813 5.4722e-005 3.8183 0.011935 9.8642e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5042 0.53954 0.16507 0.019366 14.8239 0.12021 0.00015592 0.76995 0.0091038 0.010085 0.0014171 0.98654 0.99144 3.0598e-006 1.2239e-005 0.16255 0.84571 0.87738 0.0014133 0.9563 0.43521 0.0019034 0.42161 1.9304 1.9289 16.0183 144.921 0.00022392 -85.52 0.47395
7.578 0.98813 5.4722e-005 3.8183 0.011935 9.8654e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5043 0.53958 0.16508 0.019367 14.8267 0.12021 0.00015593 0.76994 0.0091042 0.010085 0.0014169 0.98655 0.99145 3.0592e-006 1.2237e-005 0.16256 0.84614 0.87759 0.0014132 0.95656 0.4354 0.0019033 0.42163 1.9314 1.9299 16.0183 144.921 0.0002236 -85.521 0.47495
7.579 0.98813 5.4722e-005 3.8183 0.011935 9.8667e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5044 0.53963 0.1651 0.019368 14.8295 0.12022 0.00015594 0.76993 0.0091046 0.010086 0.0014167 0.98655 0.99145 3.0587e-006 1.2235e-005 0.16256 0.84657 0.87779 0.001413 0.95682 0.4356 0.0019031 0.42164 1.9323 1.9309 16.0183 144.921 0.00022328 -85.522 0.47595
7.58 0.98813 5.4722e-005 3.8183 0.011935 9.868e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5044 0.53967 0.16511 0.019369 14.8323 0.12023 0.00015595 0.76993 0.009105 0.010086 0.0014164 0.98655 0.99145 3.0581e-006 1.2232e-005 0.16256 0.847 0.878 0.0014129 0.95708 0.4358 0.0019029 0.42166 1.9333 1.9319 16.0183 144.921 0.00022297 -85.523 0.47695
7.581 0.98813 5.4722e-005 3.8183 0.011935 9.8693e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5045 0.53972 0.16512 0.01937 14.8351 0.12024 0.00015596 0.76992 0.0091054 0.010087 0.0014162 0.98656 0.99145 3.0576e-006 1.223e-005 0.16257 0.84743 0.8782 0.0014128 0.95734 0.43599 0.0019028 0.42167 1.9343 1.9328 16.0183 144.9211 0.00022265 -85.524 0.47795
7.582 0.98813 5.4722e-005 3.8183 0.011935 9.8706e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5046 0.53976 0.16514 0.019372 14.8379 0.12024 0.00015597 0.76991 0.0091059 0.010087 0.0014159 0.98656 0.99145 3.057e-006 1.2228e-005 0.16257 0.84785 0.87841 0.0014126 0.95759 0.43619 0.0019026 0.42169 1.9353 1.9338 16.0183 144.9211 0.00022234 -85.525 0.47895
7.583 0.98813 5.4722e-005 3.8183 0.011935 9.8719e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5047 0.53981 0.16515 0.019373 14.8408 0.12025 0.00015598 0.76991 0.0091063 0.010087 0.0014157 0.98656 0.99146 3.0565e-006 1.2226e-005 0.16257 0.84828 0.87861 0.0014125 0.95785 0.43638 0.0019025 0.4217 1.9363 1.9348 16.0183 144.9211 0.00022203 -85.526 0.47995
7.584 0.98813 5.4722e-005 3.8183 0.011935 9.8731e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5048 0.53985 0.16517 0.019374 14.8436 0.12026 0.000156 0.7699 0.0091067 0.010088 0.0014155 0.98657 0.99146 3.056e-006 1.2224e-005 0.16258 0.8487 0.87881 0.0014124 0.9581 0.43658 0.0019023 0.42172 1.9372 1.9358 16.0183 144.9211 0.00022171 -85.527 0.48095
7.585 0.98813 5.4722e-005 3.8183 0.011935 9.8744e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5049 0.5399 0.16518 0.019375 14.8464 0.12026 0.00015601 0.76989 0.0091071 0.010088 0.0014152 0.98657 0.99146 3.0555e-006 1.2222e-005 0.16258 0.84912 0.87901 0.0014123 0.95835 0.43677 0.0019021 0.42173 1.9382 1.9368 16.0183 144.9211 0.0002214 -85.528 0.48195
7.586 0.98813 5.4721e-005 3.8183 0.011935 9.8757e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.505 0.53994 0.16519 0.019376 14.8492 0.12027 0.00015602 0.76989 0.0091075 0.010089 0.001415 0.98657 0.99146 3.0549e-006 1.222e-005 0.16258 0.84954 0.87921 0.0014122 0.9586 0.43697 0.001902 0.42175 1.9392 1.9377 16.0182 144.9212 0.0002211 -85.5289 0.48295
7.587 0.98813 5.4721e-005 3.8183 0.011935 9.877e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5051 0.53999 0.16521 0.019377 14.852 0.12028 0.00015603 0.76988 0.009108 0.010089 0.0014148 0.98657 0.99146 3.0544e-006 1.2218e-005 0.16259 0.84996 0.87941 0.0014121 0.95885 0.43717 0.0019018 0.42176 1.9401 1.9387 16.0182 144.9212 0.00022079 -85.5299 0.48395
7.588 0.98813 5.4721e-005 3.8183 0.011935 9.8783e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5051 0.54003 0.16522 0.019379 14.8548 0.12028 0.00015604 0.76987 0.0091084 0.01009 0.0014146 0.98658 0.99147 3.0539e-006 1.2216e-005 0.16259 0.85037 0.87961 0.001412 0.9591 0.43736 0.0019017 0.42177 1.9411 1.9397 16.0182 144.9212 0.00022048 -85.5309 0.48495
7.589 0.98813 5.4721e-005 3.8183 0.011935 9.8796e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5052 0.54008 0.16523 0.01938 14.8576 0.12029 0.00015605 0.76986 0.0091088 0.01009 0.0014143 0.98658 0.99147 3.0534e-006 1.2213e-005 0.16259 0.85079 0.87981 0.0014119 0.95934 0.43756 0.0019015 0.42179 1.9421 1.9406 16.0182 144.9212 0.00022018 -85.5318 0.48595
7.59 0.98813 5.4721e-005 3.8183 0.011935 9.8809e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5053 0.54013 0.16525 0.019381 14.8604 0.1203 0.00015606 0.76986 0.0091092 0.010091 0.0014141 0.98658 0.99147 3.0529e-006 1.2211e-005 0.1626 0.8512 0.88 0.0014118 0.95958 0.43775 0.0019014 0.4218 1.943 1.9416 16.0182 144.9212 0.00021987 -85.5327 0.48695
7.591 0.98813 5.4721e-005 3.8183 0.011935 9.8821e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5054 0.54017 0.16526 0.019382 14.8632 0.12031 0.00015607 0.76985 0.0091096 0.010091 0.0014139 0.98659 0.99147 3.0524e-006 1.2209e-005 0.1626 0.85162 0.8802 0.0014117 0.95983 0.43795 0.0019012 0.42182 1.944 1.9426 16.0182 144.9212 0.00021957 -85.5337 0.48795
7.592 0.98813 5.4721e-005 3.8183 0.011935 9.8834e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5055 0.54022 0.16528 0.019383 14.866 0.12031 0.00015608 0.76984 0.00911 0.010091 0.0014137 0.98659 0.99147 3.0519e-006 1.2207e-005 0.1626 0.85203 0.88039 0.0014115 0.96007 0.43814 0.0019011 0.42183 1.9449 1.9435 16.0182 144.9213 0.00021927 -85.5346 0.48895
7.593 0.98813 5.4721e-005 3.8183 0.011935 9.8847e-005 0.0011701 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5056 0.54026 0.16529 0.019384 14.8688 0.12032 0.00015609 0.76984 0.0091105 0.010092 0.0014135 0.98659 0.99148 3.0514e-006 1.2205e-005 0.16261 0.85244 0.88059 0.0014114 0.9603 0.43834 0.0019009 0.42185 1.9459 1.9445 16.0182 144.9213 0.00021897 -85.5355 0.48995
7.594 0.98813 5.4721e-005 3.8183 0.011935 9.886e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5057 0.54031 0.1653 0.019386 14.8716 0.12033 0.0001561 0.76983 0.0091109 0.010092 0.0014133 0.98659 0.99148 3.0509e-006 1.2203e-005 0.16261 0.85285 0.88078 0.0014113 0.96054 0.43853 0.0019008 0.42186 1.9468 1.9454 16.0182 144.9213 0.00021867 -85.5364 0.49095
7.595 0.98813 5.4721e-005 3.8183 0.011935 9.8873e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5058 0.54035 0.16532 0.019387 14.8744 0.12033 0.00015611 0.76982 0.0091113 0.010093 0.001413 0.9866 0.99148 3.0504e-006 1.2202e-005 0.16261 0.85326 0.88097 0.0014112 0.96078 0.43873 0.0019006 0.42188 1.9478 1.9464 16.0182 144.9213 0.00021837 -85.5373 0.49195
7.596 0.98813 5.4721e-005 3.8183 0.011935 9.8886e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5058 0.5404 0.16533 0.019388 14.8772 0.12034 0.00015612 0.76982 0.0091117 0.010093 0.0014128 0.9866 0.99148 3.0499e-006 1.22e-005 0.16262 0.85366 0.88117 0.0014111 0.96101 0.43892 0.0019005 0.42189 1.9487 1.9473 16.0182 144.9213 0.00021808 -85.5382 0.49295
7.597 0.98813 5.4721e-005 3.8183 0.011935 9.8898e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5059 0.54044 0.16535 0.019389 14.88 0.12035 0.00015613 0.76981 0.0091121 0.010094 0.0014126 0.9866 0.99148 3.0494e-006 1.2198e-005 0.16262 0.85407 0.88136 0.0014109 0.96124 0.43912 0.0019003 0.42191 1.9496 1.9483 16.0181 144.9214 0.00021778 -85.5391 0.49395
7.598 0.98813 5.472e-005 3.8183 0.011935 9.8911e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.506 0.54049 0.16536 0.01939 14.8828 0.12035 0.00015614 0.7698 0.0091126 0.010094 0.0014124 0.98661 0.99148 3.0489e-006 1.2196e-005 0.16262 0.85447 0.88155 0.0014108 0.96148 0.43931 0.0019002 0.42192 1.9506 1.9492 16.0181 144.9214 0.00021749 -85.54 0.49495
7.599 0.98813 5.472e-005 3.8183 0.011935 9.8924e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5061 0.54053 0.16537 0.019391 14.8856 0.12036 0.00015615 0.76979 0.009113 0.010095 0.0014122 0.98661 0.99149 3.0485e-006 1.2194e-005 0.16263 0.85487 0.88174 0.0014107 0.96171 0.43951 0.0019001 0.42194 1.9515 1.9501 16.0181 144.9214 0.00021719 -85.5409 0.49595
7.6 0.98813 5.472e-005 3.8183 0.011935 9.8937e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5062 0.54058 0.16539 0.019393 14.8884 0.12037 0.00015616 0.76979 0.0091134 0.010095 0.001412 0.98661 0.99149 3.048e-006 1.2192e-005 0.16263 0.85528 0.88192 0.0014106 0.96193 0.4397 0.0018999 0.42195 1.9525 1.9511 16.0181 144.9214 0.0002169 -85.5418 0.49695
7.601 0.98813 5.472e-005 3.8183 0.011935 9.895e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5063 0.54062 0.1654 0.019394 14.8912 0.12038 0.00015617 0.76978 0.0091138 0.010096 0.0014118 0.98661 0.99149 3.0475e-006 1.219e-005 0.16263 0.85568 0.88211 0.0014105 0.96216 0.4399 0.0018998 0.42196 1.9534 1.952 16.0181 144.9214 0.00021661 -85.5426 0.49795
7.602 0.98813 5.472e-005 3.8183 0.011935 9.8963e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5064 0.54067 0.16542 0.019395 14.894 0.12038 0.00015618 0.76977 0.0091142 0.010096 0.0014116 0.98662 0.99149 3.0471e-006 1.2188e-005 0.16264 0.85608 0.8823 0.0014104 0.96239 0.44009 0.0018996 0.42198 1.9543 1.9529 16.0181 144.9215 0.00021632 -85.5435 0.49895
7.603 0.98813 5.472e-005 3.8183 0.011935 9.8975e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5065 0.54071 0.16543 0.019396 14.8969 0.12039 0.00015619 0.76977 0.0091146 0.010096 0.0014114 0.98662 0.99149 3.0466e-006 1.2186e-005 0.16264 0.85647 0.88249 0.0014103 0.96261 0.44028 0.0018995 0.42199 1.9552 1.9539 16.0181 144.9215 0.00021604 -85.5444 0.49995
7.604 0.98813 5.472e-005 3.8183 0.011935 9.8988e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5066 0.54076 0.16544 0.019397 14.8997 0.1204 0.0001562 0.76976 0.0091151 0.010097 0.0014112 0.98662 0.9915 3.0461e-006 1.2185e-005 0.16264 0.85687 0.88267 0.0014102 0.96283 0.44048 0.0018994 0.42201 1.9562 1.9548 16.0181 144.9215 0.00021575 -85.5452 0.50095
7.605 0.98813 5.472e-005 3.8183 0.011935 9.9001e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5066 0.5408 0.16546 0.019398 14.9025 0.1204 0.00015622 0.76975 0.0091155 0.010097 0.001411 0.98662 0.9915 3.0457e-006 1.2183e-005 0.16265 0.85727 0.88286 0.00141 0.96305 0.44067 0.0018992 0.42202 1.9571 1.9557 16.0181 144.9215 0.00021546 -85.5461 0.50195
7.606 0.98813 5.472e-005 3.8183 0.011935 9.9014e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5067 0.54085 0.16547 0.019399 14.9053 0.12041 0.00015623 0.76975 0.0091159 0.010098 0.0014108 0.98663 0.9915 3.0452e-006 1.2181e-005 0.16265 0.85766 0.88304 0.0014099 0.96327 0.44087 0.0018991 0.42204 1.958 1.9566 16.0181 144.9215 0.00021518 -85.5469 0.50295
7.607 0.98813 5.472e-005 3.8183 0.011935 9.9027e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5068 0.54089 0.16548 0.019401 14.9081 0.12042 0.00015624 0.76974 0.0091163 0.010098 0.0014106 0.98663 0.9915 3.0448e-006 1.2179e-005 0.16265 0.85805 0.88322 0.0014098 0.96349 0.44106 0.001899 0.42205 1.9589 1.9576 16.018 144.9216 0.0002149 -85.5477 0.50395
7.608 0.98813 5.472e-005 3.8183 0.011935 9.904e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5069 0.54094 0.1655 0.019402 14.9109 0.12042 0.00015625 0.76973 0.0091167 0.010099 0.0014104 0.98663 0.9915 3.0444e-006 1.2177e-005 0.16266 0.85844 0.88341 0.0014097 0.96371 0.44126 0.0018988 0.42207 1.9598 1.9585 16.018 144.9216 0.00021461 -85.5486 0.50495
7.609 0.98813 5.472e-005 3.8183 0.011935 9.9053e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.507 0.54098 0.16551 0.019403 14.9137 0.12043 0.00015626 0.76973 0.0091172 0.010099 0.0014102 0.98663 0.9915 3.0439e-006 1.2176e-005 0.16266 0.85883 0.88359 0.0014096 0.96392 0.44145 0.0018987 0.42208 1.9607 1.9594 16.018 144.9216 0.00021433 -85.5494 0.50595
7.61 0.98813 5.472e-005 3.8183 0.011935 9.9065e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5071 0.54103 0.16553 0.019404 14.9165 0.12044 0.00015627 0.76972 0.0091176 0.0101 0.00141 0.98664 0.99151 3.0435e-006 1.2174e-005 0.16266 0.85922 0.88377 0.0014095 0.96414 0.44164 0.0018986 0.4221 1.9616 1.9603 16.018 144.9216 0.00021405 -85.5502 0.50695
7.611 0.98813 5.4719e-005 3.8183 0.011935 9.9078e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5072 0.54108 0.16554 0.019405 14.9193 0.12045 0.00015628 0.76971 0.009118 0.0101 0.0014098 0.98664 0.99151 3.043e-006 1.2172e-005 0.16266 0.85961 0.88395 0.0014094 0.96435 0.44184 0.0018984 0.42211 1.9625 1.9612 16.018 144.9216 0.00021377 -85.551 0.50795
7.612 0.98813 5.4719e-005 3.8183 0.011935 9.9091e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5073 0.54112 0.16555 0.019406 14.9221 0.12045 0.00015629 0.7697 0.0091184 0.0101 0.0014096 0.98664 0.99151 3.0426e-006 1.217e-005 0.16267 0.86 0.88413 0.0014094 0.96456 0.44203 0.0018983 0.42213 1.9634 1.9621 16.018 144.9217 0.0002135 -85.5518 0.50895
7.613 0.98813 5.4719e-005 3.8183 0.011935 9.9104e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5073 0.54117 0.16557 0.019408 14.925 0.12046 0.0001563 0.7697 0.0091188 0.010101 0.0014094 0.98664 0.99151 3.0422e-006 1.2169e-005 0.16267 0.86038 0.88431 0.0014093 0.96477 0.44223 0.0018982 0.42214 1.9643 1.963 16.018 144.9217 0.00021322 -85.5526 0.50995
7.614 0.98813 5.4719e-005 3.8183 0.011935 9.9117e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5074 0.54121 0.16558 0.019409 14.9278 0.12047 0.00015631 0.76969 0.0091192 0.010101 0.0014093 0.98665 0.99151 3.0417e-006 1.2167e-005 0.16267 0.86077 0.88449 0.0014092 0.96498 0.44242 0.001898 0.42215 1.9652 1.9639 16.018 144.9217 0.00021294 -85.5534 0.51095
7.615 0.98813 5.4719e-005 3.8183 0.011935 9.913e-005 0.0011702 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5075 0.54126 0.1656 0.01941 14.9306 0.12047 0.00015632 0.76968 0.0091197 0.010102 0.0014091 0.98665 0.99151 3.0413e-006 1.2165e-005 0.16268 0.86115 0.88467 0.0014091 0.96519 0.44261 0.0018979 0.42217 1.9661 1.9648 16.018 144.9217 0.00021267 -85.5542 0.51195
7.616 0.98813 5.4719e-005 3.8183 0.011935 9.9142e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5076 0.5413 0.16561 0.019411 14.9334 0.12048 0.00015633 0.76968 0.0091201 0.010102 0.0014089 0.98665 0.99151 3.0409e-006 1.2164e-005 0.16268 0.86153 0.88484 0.001409 0.9654 0.44281 0.0018978 0.42218 1.967 1.9657 16.0179 144.9217 0.0002124 -85.555 0.51295
7.617 0.98813 5.4719e-005 3.8183 0.011935 9.9155e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5077 0.54135 0.16562 0.019412 14.9362 0.12049 0.00015634 0.76967 0.0091205 0.010103 0.0014087 0.98665 0.99152 3.0405e-006 1.2162e-005 0.16268 0.86192 0.88502 0.0014089 0.9656 0.443 0.0018977 0.4222 1.9679 1.9666 16.0179 144.9218 0.00021212 -85.5557 0.51395
7.618 0.98813 5.4719e-005 3.8183 0.011935 9.9168e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5078 0.54139 0.16564 0.019413 14.939 0.12049 0.00015635 0.76966 0.0091209 0.010103 0.0014085 0.98666 0.99152 3.0401e-006 1.216e-005 0.16269 0.8623 0.8852 0.0014088 0.9658 0.44319 0.0018975 0.42221 1.9688 1.9675 16.0179 144.9218 0.00021185 -85.5565 0.51495
7.619 0.98813 5.4719e-005 3.8183 0.011935 9.9181e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5079 0.54144 0.16565 0.019415 14.9418 0.1205 0.00015636 0.76966 0.0091213 0.010104 0.0014083 0.98666 0.99152 3.0397e-006 1.2159e-005 0.16269 0.86267 0.88537 0.0014087 0.96601 0.44339 0.0018974 0.42223 1.9697 1.9684 16.0179 144.9218 0.00021158 -85.5573 0.51595
7.62 0.98813 5.4719e-005 3.8183 0.011935 9.9194e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.508 0.54148 0.16566 0.019416 14.9446 0.12051 0.00015637 0.76965 0.0091217 0.010104 0.0014082 0.98666 0.99152 3.0393e-006 1.2157e-005 0.16269 0.86305 0.88554 0.0014086 0.96621 0.44358 0.0018973 0.42224 1.9706 1.9693 16.0179 144.9218 0.00021131 -85.558 0.51695
7.621 0.98813 5.4719e-005 3.8183 0.011935 9.9207e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.508 0.54153 0.16568 0.019417 14.9475 0.12051 0.00015638 0.76964 0.0091222 0.010104 0.001408 0.98666 0.99152 3.0388e-006 1.2155e-005 0.1627 0.86343 0.88572 0.0014085 0.96641 0.44377 0.0018972 0.42226 1.9715 1.9702 16.0179 144.9218 0.00021105 -85.5588 0.51795
7.622 0.98813 5.4719e-005 3.8183 0.011934 9.9219e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5081 0.54157 0.16569 0.019418 14.9503 0.12052 0.00015639 0.76963 0.0091226 0.010105 0.0014078 0.98667 0.99152 3.0384e-006 1.2154e-005 0.1627 0.8638 0.88589 0.0014084 0.9666 0.44397 0.0018971 0.42227 1.9723 1.971 16.0179 144.9219 0.00021078 -85.5595 0.51895
7.623 0.98813 5.4718e-005 3.8183 0.011934 9.9232e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5082 0.54162 0.16571 0.019419 14.9531 0.12053 0.0001564 0.76963 0.009123 0.010105 0.0014076 0.98667 0.99153 3.038e-006 1.2152e-005 0.1627 0.86418 0.88606 0.0014083 0.9668 0.44416 0.0018969 0.42229 1.9732 1.9719 16.0179 144.9219 0.00021051 -85.5603 0.51995
7.624 0.98813 5.4718e-005 3.8183 0.011934 9.9245e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5083 0.54166 0.16572 0.01942 14.9559 0.12054 0.00015641 0.76962 0.0091234 0.010106 0.0014075 0.98667 0.99153 3.0376e-006 1.2151e-005 0.16271 0.86455 0.88623 0.0014082 0.967 0.44435 0.0018968 0.4223 1.9741 1.9728 16.0179 144.9219 0.00021025 -85.561 0.52095
7.625 0.98813 5.4718e-005 3.8183 0.011934 9.9258e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5084 0.54171 0.16573 0.019422 14.9587 0.12054 0.00015642 0.76961 0.0091238 0.010106 0.0014073 0.98667 0.99153 3.0373e-006 1.2149e-005 0.16271 0.86492 0.8864 0.0014081 0.96719 0.44455 0.0018967 0.42232 1.975 1.9737 16.0178 144.9219 0.00020999 -85.5617 0.52195
7.626 0.98813 5.4718e-005 3.8183 0.011934 9.9271e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5085 0.54175 0.16575 0.019423 14.9615 0.12055 0.00015643 0.76961 0.0091242 0.010107 0.0014071 0.98667 0.99153 3.0369e-006 1.2147e-005 0.16271 0.86529 0.88657 0.001408 0.96739 0.44474 0.0018966 0.42233 1.9758 1.9745 16.0178 144.9219 0.00020972 -85.5625 0.52295
7.627 0.98813 5.4718e-005 3.8183 0.011934 9.9284e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5086 0.5418 0.16576 0.019424 14.9643 0.12056 0.00015645 0.7696 0.0091247 0.010107 0.001407 0.98668 0.99153 3.0365e-006 1.2146e-005 0.16272 0.86566 0.88674 0.001408 0.96758 0.44493 0.0018965 0.42234 1.9767 1.9754 16.0178 144.922 0.00020946 -85.5632 0.52395
7.628 0.98813 5.4718e-005 3.8183 0.011934 9.9297e-005 0.0011703 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5087 0.54184 0.16578 0.019425 14.9672 0.12056 0.00015646 0.76959 0.0091251 0.010108 0.0014068 0.98668 0.99153 3.0361e-006 1.2144e-005 0.16272 0.86603 0.88691 0.0014079 0.96777 0.44513 0.0018963 0.42236 1.9776 1.9763 16.0178 144.922 0.0002092 -85.5639 0.52495
7.629 0.98813 5.4718e-005 3.8183 0.011934 9.9309e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5087 0.54189 0.16579 0.019426 14.97 0.12057 0.00015647 0.76959 0.0091255 0.010108 0.0014066 0.98668 0.99153 3.0357e-006 1.2143e-005 0.16272 0.86639 0.88708 0.0014078 0.96796 0.44532 0.0018962 0.42237 1.9784 1.9772 16.0178 144.922 0.00020894 -85.5646 0.52595
7.63 0.98813 5.4718e-005 3.8183 0.011934 9.9322e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5088 0.54193 0.1658 0.019427 14.9728 0.12058 0.00015648 0.76958 0.0091259 0.010108 0.0014065 0.98668 0.99154 3.0353e-006 1.2141e-005 0.16273 0.86676 0.88725 0.0014077 0.96815 0.44551 0.0018961 0.42239 1.9793 1.978 16.0178 144.922 0.00020868 -85.5653 0.52695
7.631 0.98813 5.4718e-005 3.8183 0.011934 9.9335e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5089 0.54198 0.16582 0.019429 14.9756 0.12058 0.00015649 0.76957 0.0091263 0.010109 0.0014063 0.98669 0.99154 3.035e-006 1.214e-005 0.16273 0.86712 0.88741 0.0014076 0.96833 0.4457 0.001896 0.4224 1.9801 1.9789 16.0178 144.922 0.00020843 -85.566 0.52795
7.632 0.98813 5.4718e-005 3.8183 0.011934 9.9348e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.509 0.54202 0.16583 0.01943 14.9784 0.12059 0.0001565 0.76957 0.0091267 0.010109 0.0014061 0.98669 0.99154 3.0346e-006 1.2138e-005 0.16273 0.86749 0.88758 0.0014076 0.96852 0.4459 0.0018959 0.42242 1.981 1.9797 16.0177 144.9221 0.00020817 -85.5667 0.52895
7.633 0.98813 5.4718e-005 3.8183 0.011934 9.9361e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5091 0.54207 0.16584 0.019431 14.9813 0.1206 0.00015651 0.76956 0.0091272 0.01011 0.001406 0.98669 0.99154 3.0342e-006 1.2137e-005 0.16274 0.86785 0.88775 0.0014075 0.96871 0.44609 0.0018958 0.42243 1.9818 1.9806 16.0177 144.9221 0.00020792 -85.5674 0.52995
7.634 0.98813 5.4718e-005 3.8183 0.011934 9.9374e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5092 0.54212 0.16586 0.019432 14.9841 0.12061 0.00015652 0.76955 0.0091276 0.01011 0.0014058 0.98669 0.99154 3.0338e-006 1.2135e-005 0.16274 0.86821 0.88791 0.0014074 0.96889 0.44628 0.0018957 0.42245 1.9827 1.9815 16.0177 144.9221 0.00020766 -85.5681 0.53095
7.635 0.98813 5.4717e-005 3.8183 0.011934 9.9386e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5093 0.54216 0.16587 0.019433 14.9869 0.12061 0.00015653 0.76954 0.009128 0.010111 0.0014056 0.98669 0.99154 3.0335e-006 1.2134e-005 0.16274 0.86857 0.88807 0.0014073 0.96907 0.44647 0.0018956 0.42246 1.9835 1.9823 16.0177 144.9221 0.00020741 -85.5688 0.53195
7.636 0.98813 5.4717e-005 3.8183 0.011934 9.9399e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5094 0.54221 0.16589 0.019434 14.9897 0.12062 0.00015654 0.76954 0.0091284 0.010111 0.0014055 0.9867 0.99154 3.0331e-006 1.2132e-005 0.16275 0.86893 0.88824 0.0014072 0.96925 0.44667 0.0018955 0.42248 1.9844 1.9832 16.0177 144.9221 0.00020716 -85.5695 0.53295
7.637 0.98813 5.4717e-005 3.8183 0.011934 9.9412e-005 0.0011703 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5094 0.54225 0.1659 0.019435 14.9925 0.12063 0.00015655 0.76953 0.0091288 0.010112 0.0014053 0.9867 0.99154 3.0327e-006 1.2131e-005 0.16275 0.86929 0.8884 0.0014071 0.96943 0.44686 0.0018953 0.42249 1.9852 1.984 16.0177 144.9222 0.0002069 -85.5701 0.53395
7.638 0.98813 5.4717e-005 3.8183 0.011934 9.9425e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5095 0.5423 0.16591 0.019437 14.9954 0.12063 0.00015656 0.76952 0.0091292 0.010112 0.0014052 0.9867 0.99155 3.0324e-006 1.2129e-005 0.16275 0.86965 0.88856 0.0014071 0.96961 0.44705 0.0018952 0.42251 1.9861 1.9848 16.0177 144.9222 0.00020665 -85.5708 0.53495
7.639 0.98813 5.4717e-005 3.8183 0.011934 9.9438e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5096 0.54234 0.16593 0.019438 14.9982 0.12064 0.00015657 0.76952 0.0091297 0.010112 0.001405 0.9867 0.99155 3.032e-006 1.2128e-005 0.16275 0.87 0.88872 0.001407 0.96979 0.44724 0.0018951 0.42252 1.9869 1.9857 16.0177 144.9222 0.00020641 -85.5715 0.53595
7.64 0.98813 5.4717e-005 3.8183 0.011934 9.9451e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5097 0.54239 0.16594 0.019439 15.001 0.12065 0.00015658 0.76951 0.0091301 0.010113 0.0014049 0.9867 0.99155 3.0317e-006 1.2127e-005 0.16276 0.87036 0.88889 0.0014069 0.96997 0.44744 0.001895 0.42254 1.9878 1.9865 16.0176 144.9222 0.00020616 -85.5721 0.53695
7.641 0.98813 5.4717e-005 3.8183 0.011934 9.9463e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5098 0.54243 0.16596 0.01944 15.0038 0.12065 0.00015659 0.7695 0.0091305 0.010113 0.0014047 0.98671 0.99155 3.0313e-006 1.2125e-005 0.16276 0.87071 0.88905 0.0014068 0.97014 0.44763 0.0018949 0.42255 1.9886 1.9874 16.0176 144.9222 0.00020591 -85.5728 0.53795
7.642 0.98813 5.4717e-005 3.8183 0.011934 9.9476e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5099 0.54248 0.16597 0.019441 15.0066 0.12066 0.0001566 0.7695 0.0091309 0.010114 0.0014046 0.98671 0.99155 3.031e-006 1.2124e-005 0.16276 0.87106 0.8892 0.0014067 0.97032 0.44782 0.0018948 0.42256 1.9894 1.9882 16.0176 144.9223 0.00020566 -85.5734 0.53895
7.643 0.98813 5.4717e-005 3.8183 0.011934 9.9489e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.51 0.54252 0.16598 0.019442 15.0095 0.12067 0.00015661 0.76949 0.0091313 0.010114 0.0014044 0.98671 0.99155 3.0306e-006 1.2122e-005 0.16277 0.87141 0.88936 0.0014066 0.97049 0.44801 0.0018947 0.42258 1.9903 1.989 16.0176 144.9223 0.00020542 -85.5741 0.53995
7.644 0.98813 5.4717e-005 3.8183 0.011934 9.9502e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5101 0.54257 0.166 0.019444 15.0123 0.12067 0.00015662 0.76948 0.0091317 0.010115 0.0014043 0.98671 0.99155 3.0303e-006 1.2121e-005 0.16277 0.87176 0.88952 0.0014066 0.97066 0.4482 0.0018946 0.42259 1.9911 1.9899 16.0176 144.9223 0.00020517 -85.5747 0.54095
7.645 0.98813 5.4717e-005 3.8183 0.011934 9.9515e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5101 0.54261 0.16601 0.019445 15.0151 0.12068 0.00015663 0.76948 0.0091322 0.010115 0.0014041 0.98671 0.99155 3.0299e-006 1.212e-005 0.16277 0.87211 0.88968 0.0014065 0.97083 0.4484 0.0018945 0.42261 1.9919 1.9907 16.0176 144.9223 0.00020493 -85.5753 0.54195
7.646 0.98813 5.4717e-005 3.8183 0.011934 9.9528e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5102 0.54266 0.16603 0.019446 15.0179 0.12069 0.00015664 0.76947 0.0091326 0.010115 0.001404 0.98672 0.99156 3.0296e-006 1.2118e-005 0.16278 0.87246 0.88984 0.0014064 0.971 0.44859 0.0018944 0.42262 1.9927 1.9915 16.0176 144.9223 0.00020469 -85.576 0.54295
7.647 0.98813 5.4717e-005 3.8183 0.011934 9.9541e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5103 0.5427 0.16604 0.019447 15.0207 0.1207 0.00015665 0.76946 0.009133 0.010116 0.0014038 0.98672 0.99156 3.0293e-006 1.2117e-005 0.16278 0.87281 0.88999 0.0014063 0.97117 0.44878 0.0018943 0.42264 1.9936 1.9924 16.0175 144.9224 0.00020445 -85.5766 0.54395
7.648 0.98813 5.4716e-005 3.8183 0.011934 9.9553e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5104 0.54275 0.16605 0.019448 15.0236 0.1207 0.00015666 0.76945 0.0091334 0.010116 0.0014037 0.98672 0.99156 3.0289e-006 1.2116e-005 0.16278 0.87315 0.89015 0.0014062 0.97134 0.44897 0.0018942 0.42265 1.9944 1.9932 16.0175 144.9224 0.00020421 -85.5772 0.54495
7.649 0.98813 5.4716e-005 3.8183 0.011934 9.9566e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5105 0.54279 0.16607 0.019449 15.0264 0.12071 0.00015667 0.76945 0.0091338 0.010117 0.0014035 0.98672 0.99156 3.0286e-006 1.2114e-005 0.16279 0.8735 0.8903 0.0014062 0.97151 0.44916 0.0018941 0.42267 1.9952 1.994 16.0175 144.9224 0.00020397 -85.5778 0.54595
7.65 0.98813 5.4716e-005 3.8183 0.011934 9.9579e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5106 0.54284 0.16608 0.01945 15.0292 0.12072 0.00015668 0.76944 0.0091342 0.010117 0.0014034 0.98672 0.99156 3.0283e-006 1.2113e-005 0.16279 0.87384 0.89046 0.0014061 0.97167 0.44935 0.001894 0.42268 1.996 1.9948 16.0175 144.9224 0.00020373 -85.5785 0.54695
7.651 0.98813 5.4716e-005 3.8183 0.011934 9.9592e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5107 0.54288 0.16609 0.019452 15.032 0.12072 0.0001567 0.76943 0.0091346 0.010118 0.0014032 0.98672 0.99156 3.028e-006 1.2112e-005 0.16279 0.87418 0.89061 0.001406 0.97184 0.44955 0.0018939 0.4227 1.9968 1.9956 16.0175 144.9224 0.00020349 -85.5791 0.54795
7.652 0.98813 5.4716e-005 3.8183 0.011934 9.9605e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5108 0.54293 0.16611 0.019453 15.0349 0.12073 0.00015671 0.76943 0.0091351 0.010118 0.0014031 0.98673 0.99156 3.0276e-006 1.211e-005 0.1628 0.87452 0.89077 0.0014059 0.972 0.44974 0.0018938 0.42271 1.9976 1.9965 16.0175 144.9225 0.00020325 -85.5797 0.54895
7.653 0.98813 5.4716e-005 3.8183 0.011934 9.9618e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5108 0.54297 0.16612 0.019454 15.0377 0.12074 0.00015672 0.76942 0.0091355 0.010119 0.001403 0.98673 0.99156 3.0273e-006 1.2109e-005 0.1628 0.87486 0.89092 0.0014059 0.97217 0.44993 0.0018937 0.42273 1.9984 1.9973 16.0175 144.9225 0.00020302 -85.5803 0.54995
7.654 0.98813 5.4716e-005 3.8183 0.011934 9.963e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5109 0.54302 0.16614 0.019455 15.0405 0.12074 0.00015673 0.76941 0.0091359 0.010119 0.0014028 0.98673 0.99157 3.027e-006 1.2108e-005 0.1628 0.8752 0.89107 0.0014058 0.97233 0.45012 0.0018936 0.42274 1.9993 1.9981 16.0174 144.9225 0.00020278 -85.5809 0.55095
7.655 0.98813 5.4716e-005 3.8183 0.011934 9.9643e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.511 0.54306 0.16615 0.019456 15.0433 0.12075 0.00015674 0.76941 0.0091363 0.010119 0.0014027 0.98673 0.99157 3.0267e-006 1.2107e-005 0.16281 0.87554 0.89122 0.0014057 0.97249 0.45031 0.0018935 0.42276 2.0001 1.9989 16.0174 144.9225 0.00020255 -85.5815 0.55195
7.656 0.98813 5.4716e-005 3.8183 0.011934 9.9656e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5111 0.54311 0.16616 0.019457 15.0462 0.12076 0.00015675 0.7694 0.0091367 0.01012 0.0014025 0.98673 0.99157 3.0264e-006 1.2105e-005 0.16281 0.87588 0.89137 0.0014057 0.97265 0.4505 0.0018934 0.42277 2.0009 1.9997 16.0174 144.9225 0.00020232 -85.582 0.55295
7.657 0.98813 5.4716e-005 3.8183 0.011934 9.9669e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5112 0.54315 0.16618 0.019459 15.049 0.12076 0.00015676 0.76939 0.0091371 0.01012 0.0014024 0.98674 0.99157 3.026e-006 1.2104e-005 0.16281 0.87622 0.89152 0.0014056 0.97281 0.45069 0.0018933 0.42278 2.0017 2.0005 16.0174 144.9226 0.00020208 -85.5826 0.55395
7.658 0.98813 5.4716e-005 3.8183 0.011934 9.9682e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5113 0.5432 0.16619 0.01946 15.0518 0.12077 0.00015677 0.76938 0.0091375 0.010121 0.0014023 0.98674 0.99157 3.0257e-006 1.2103e-005 0.16282 0.87655 0.89167 0.0014055 0.97296 0.45088 0.0018932 0.4228 2.0025 2.0013 16.0174 144.9226 0.00020185 -85.5832 0.55495
7.659 0.98813 5.4716e-005 3.8183 0.011934 9.9695e-005 0.0011704 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5114 0.54324 0.1662 0.019461 15.0547 0.12078 0.00015678 0.76938 0.009138 0.010121 0.0014021 0.98674 0.99157 3.0254e-006 1.2102e-005 0.16282 0.87689 0.89182 0.0014054 0.97312 0.45107 0.0018931 0.42281 2.0033 2.0021 16.0174 144.9226 0.00020162 -85.5838 0.55595
7.66 0.98813 5.4715e-005 3.8183 0.011934 9.9707e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5115 0.54329 0.16622 0.019462 15.0575 0.12079 0.00015679 0.76937 0.0091384 0.010122 0.001402 0.98674 0.99157 3.0251e-006 1.21e-005 0.16282 0.87722 0.89197 0.0014054 0.97328 0.45127 0.0018931 0.42283 2.0041 2.0029 16.0173 144.9226 0.00020139 -85.5844 0.55695
7.661 0.98813 5.4715e-005 3.8183 0.011934 9.972e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5115 0.54334 0.16623 0.019463 15.0603 0.12079 0.0001568 0.76936 0.0091388 0.010122 0.0014019 0.98674 0.99157 3.0248e-006 1.2099e-005 0.16283 0.87755 0.89212 0.0014053 0.97343 0.45146 0.001893 0.42284 2.0048 2.0037 16.0173 144.9226 0.00020116 -85.5849 0.55795
7.662 0.98813 5.4715e-005 3.8183 0.011934 9.9733e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5116 0.54338 0.16625 0.019464 15.0631 0.1208 0.00015681 0.76936 0.0091392 0.010123 0.0014017 0.98674 0.99157 3.0245e-006 1.2098e-005 0.16283 0.87788 0.89227 0.0014052 0.97358 0.45165 0.0018929 0.42286 2.0056 2.0045 16.0173 144.9227 0.00020094 -85.5855 0.55895
7.663 0.98813 5.4715e-005 3.8183 0.011934 9.9746e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5117 0.54343 0.16626 0.019466 15.066 0.12081 0.00015682 0.76935 0.0091396 0.010123 0.0014016 0.98675 0.99158 3.0242e-006 1.2097e-005 0.16283 0.87821 0.89241 0.0014052 0.97374 0.45184 0.0018928 0.42287 2.0064 2.0053 16.0173 144.9227 0.00020071 -85.586 0.55995
7.664 0.98813 5.4715e-005 3.8183 0.011934 9.9759e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5118 0.54347 0.16627 0.019467 15.0688 0.12081 0.00015683 0.76934 0.00914 0.010123 0.0014015 0.98675 0.99158 3.0239e-006 1.2096e-005 0.16284 0.87854 0.89256 0.0014051 0.97389 0.45203 0.0018927 0.42289 2.0072 2.0061 16.0173 144.9227 0.00020048 -85.5866 0.56095
7.665 0.98813 5.4715e-005 3.8183 0.011934 9.9772e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5119 0.54352 0.16629 0.019468 15.0716 0.12082 0.00015684 0.76934 0.0091404 0.010124 0.0014013 0.98675 0.99158 3.0236e-006 1.2094e-005 0.16284 0.87887 0.89271 0.001405 0.97404 0.45222 0.0018926 0.4229 2.008 2.0069 16.0173 144.9227 0.00020026 -85.5872 0.56195
7.666 0.98813 5.4715e-005 3.8183 0.011934 9.9785e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.512 0.54356 0.1663 0.019469 15.0745 0.12083 0.00015685 0.76933 0.0091409 0.010124 0.0014012 0.98675 0.99158 3.0233e-006 1.2093e-005 0.16284 0.87919 0.89285 0.001405 0.97419 0.45241 0.0018925 0.42292 2.0088 2.0077 16.0172 144.9227 0.00020004 -85.5877 0.56295
7.667 0.98813 5.4715e-005 3.8183 0.011934 9.9797e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5121 0.54361 0.16632 0.01947 15.0773 0.12083 0.00015686 0.76932 0.0091413 0.010125 0.0014011 0.98675 0.99158 3.023e-006 1.2092e-005 0.16284 0.87952 0.893 0.0014049 0.97434 0.4526 0.0018924 0.42293 2.0096 2.0084 16.0172 144.9228 0.00019981 -85.5882 0.56395
7.668 0.98813 5.4715e-005 3.8183 0.011934 9.981e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5122 0.54365 0.16633 0.019471 15.0801 0.12084 0.00015687 0.76932 0.0091417 0.010125 0.001401 0.98675 0.99158 3.0227e-006 1.2091e-005 0.16285 0.87985 0.89314 0.0014048 0.97448 0.45279 0.0018923 0.42295 2.0103 2.0092 16.0172 144.9228 0.00019959 -85.5888 0.56495
7.669 0.98813 5.4715e-005 3.8183 0.011934 9.9823e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5122 0.5437 0.16634 0.019472 15.0829 0.12085 0.00015688 0.76931 0.0091421 0.010126 0.0014008 0.98676 0.99158 3.0225e-006 1.209e-005 0.16285 0.88017 0.89328 0.0014047 0.97463 0.45298 0.0018923 0.42296 2.0111 2.01 16.0172 144.9228 0.00019937 -85.5893 0.56595
7.67 0.98813 5.4715e-005 3.8183 0.011934 9.9836e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5123 0.54374 0.16636 0.019474 15.0858 0.12085 0.00015689 0.7693 0.0091425 0.010126 0.0014007 0.98676 0.99158 3.0222e-006 1.2089e-005 0.16285 0.88049 0.89343 0.0014047 0.97478 0.45317 0.0018922 0.42298 2.0119 2.0108 16.0172 144.9228 0.00019915 -85.5899 0.56695
7.671 0.98813 5.4715e-005 3.8183 0.011934 9.9849e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5124 0.54379 0.16637 0.019475 15.0886 0.12086 0.0001569 0.7693 0.0091429 0.010127 0.0014006 0.98676 0.99158 3.0219e-006 1.2087e-005 0.16286 0.88081 0.89357 0.0014046 0.97492 0.45336 0.0018921 0.42299 2.0127 2.0116 16.0172 144.9228 0.00019893 -85.5904 0.56795
7.672 0.98813 5.4714e-005 3.8183 0.011934 9.9862e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5125 0.54383 0.16638 0.019476 15.0914 0.12087 0.00015691 0.76929 0.0091433 0.010127 0.0014005 0.98676 0.99159 3.0216e-006 1.2086e-005 0.16286 0.88113 0.89371 0.0014045 0.97507 0.45355 0.001892 0.423 2.0134 2.0123 16.0171 144.9229 0.00019871 -85.5909 0.56895
7.673 0.98813 5.4714e-005 3.8183 0.011934 9.9874e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5126 0.54388 0.1664 0.019477 15.0943 0.12088 0.00015692 0.76928 0.0091438 0.010127 0.0014003 0.98676 0.99159 3.0213e-006 1.2085e-005 0.16286 0.88145 0.89385 0.0014045 0.97521 0.45374 0.0018919 0.42302 2.0142 2.0131 16.0171 144.9229 0.00019849 -85.5914 0.56995
7.674 0.98813 5.4714e-005 3.8183 0.011934 9.9887e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5127 0.54392 0.16641 0.019478 15.0971 0.12088 0.00015693 0.76927 0.0091442 0.010128 0.0014002 0.98676 0.99159 3.0211e-006 1.2084e-005 0.16287 0.88177 0.89399 0.0014044 0.97535 0.45393 0.0018918 0.42303 2.015 2.0139 16.0171 144.9229 0.00019827 -85.592 0.57095
7.675 0.98813 5.4714e-005 3.8183 0.011934 9.99e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5128 0.54397 0.16643 0.019479 15.0999 0.12089 0.00015694 0.76927 0.0091446 0.010128 0.0014001 0.98677 0.99159 3.0208e-006 1.2083e-005 0.16287 0.88209 0.89413 0.0014044 0.97549 0.45412 0.0018917 0.42305 2.0157 2.0146 16.0171 144.9229 0.00019806 -85.5925 0.57195
7.676 0.98813 5.4714e-005 3.8183 0.011934 9.9913e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5129 0.54401 0.16644 0.019481 15.1028 0.1209 0.00015696 0.76926 0.009145 0.010129 0.0014 0.98677 0.99159 3.0205e-006 1.2082e-005 0.16287 0.88241 0.89427 0.0014043 0.97563 0.45431 0.0018917 0.42306 2.0165 2.0154 16.0171 144.9229 0.00019784 -85.593 0.57295
7.677 0.98813 5.4714e-005 3.8183 0.011934 9.9926e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5129 0.54406 0.16645 0.019482 15.1056 0.1209 0.00015697 0.76925 0.0091454 0.010129 0.0013999 0.98677 0.99159 3.0202e-006 1.2081e-005 0.16288 0.88272 0.89441 0.0014043 0.97577 0.4545 0.0018916 0.42308 2.0173 2.0162 16.0171 144.923 0.00019763 -85.5935 0.57395
7.678 0.98813 5.4714e-005 3.8183 0.011934 9.9939e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.513 0.5441 0.16647 0.019483 15.1084 0.12091 0.00015698 0.76925 0.0091458 0.01013 0.0013997 0.98677 0.99159 3.02e-006 1.208e-005 0.16288 0.88304 0.89455 0.0014042 0.97591 0.45469 0.0018915 0.42309 2.018 2.0169 16.017 144.923 0.00019741 -85.594 0.57495
7.679 0.98813 5.4714e-005 3.8183 0.011934 9.9951e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5131 0.54415 0.16648 0.019484 15.1113 0.12092 0.00015699 0.76924 0.0091462 0.01013 0.0013996 0.98677 0.99159 3.0197e-006 1.2079e-005 0.16288 0.88335 0.89469 0.0014041 0.97605 0.45488 0.0018914 0.42311 2.0188 2.0177 16.017 144.923 0.0001972 -85.5945 0.57595
7.68 0.98813 5.4714e-005 3.8183 0.011933 9.9964e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5132 0.54419 0.1665 0.019485 15.1141 0.12092 0.000157 0.76923 0.0091466 0.010131 0.0013995 0.98677 0.99159 3.0194e-006 1.2078e-005 0.16289 0.88367 0.89483 0.001404 0.97618 0.45507 0.0018913 0.42312 2.0195 2.0184 16.017 144.923 0.00019699 -85.595 0.57695
7.681 0.98813 5.4714e-005 3.8183 0.011933 9.9977e-005 0.0011705 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5133 0.54424 0.16651 0.019486 15.1169 0.12093 0.00015701 0.76923 0.0091471 0.010131 0.0013994 0.98677 0.99159 3.0192e-006 1.2077e-005 0.16289 0.88398 0.89496 0.0014039 0.97632 0.45526 0.0018913 0.42314 2.0203 2.0192 16.017 144.923 0.00019678 -85.5955 0.57795
7.682 0.98813 5.4714e-005 3.8183 0.011933 9.999e-005 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5134 0.54428 0.16652 0.019487 15.1198 0.12094 0.00015702 0.76922 0.0091475 0.010131 0.0013993 0.98678 0.9916 3.0189e-006 1.2076e-005 0.16289 0.88429 0.8951 0.0014039 0.97646 0.45545 0.0018912 0.42315 2.021 2.02 16.017 144.9231 0.00019657 -85.596 0.57895
7.683 0.98813 5.4714e-005 3.8183 0.011933 0.0001 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5135 0.54433 0.16654 0.019489 15.1226 0.12094 0.00015703 0.76921 0.0091479 0.010132 0.0013992 0.98678 0.9916 3.0186e-006 1.2075e-005 0.1629 0.8846 0.89524 0.0014039 0.97659 0.45564 0.0018911 0.42317 2.0218 2.0207 16.017 144.9231 0.00019636 -85.5965 0.57995
7.684 0.98813 5.4714e-005 3.8183 0.011933 0.00010002 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5136 0.54437 0.16655 0.01949 15.1254 0.12095 0.00015704 0.76921 0.0091483 0.010132 0.0013991 0.98678 0.9916 3.0184e-006 1.2074e-005 0.1629 0.88491 0.89537 0.0014039 0.97672 0.45583 0.001891 0.42318 2.0225 2.0215 16.0169 144.9231 0.00019615 -85.5969 0.58095
7.685 0.98813 5.4713e-005 3.8183 0.011933 0.00010003 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5136 0.54442 0.16656 0.019491 15.1283 0.12096 0.00015705 0.7692 0.0091487 0.010133 0.001399 0.98678 0.9916 3.0181e-006 1.2073e-005 0.1629 0.88522 0.89551 0.0014039 0.97686 0.45602 0.001891 0.4232 2.0233 2.0222 16.0169 144.9231 0.00019594 -85.5974 0.58195
7.686 0.98813 5.4713e-005 3.8183 0.011933 0.00010004 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5137 0.54446 0.16658 0.019492 15.1311 0.12097 0.00015706 0.76919 0.0091491 0.010133 0.0013988 0.98678 0.9916 3.0179e-006 1.2072e-005 0.16291 0.88552 0.89564 0.0014038 0.97699 0.45621 0.0018909 0.42321 2.024 2.023 16.0169 144.9231 0.00019573 -85.5979 0.58295
7.687 0.98813 5.4713e-005 3.8183 0.011933 0.00010005 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5138 0.54451 0.16659 0.019493 15.134 0.12097 0.00015707 0.76918 0.0091495 0.010134 0.0013987 0.98678 0.9916 3.0176e-006 1.207e-005 0.16291 0.88583 0.89578 0.0014037 0.97712 0.4564 0.0018908 0.42322 2.0248 2.0237 16.0169 144.9232 0.00019553 -85.5984 0.58395
7.688 0.98813 5.4713e-005 3.8183 0.011933 0.00010007 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5139 0.54456 0.16661 0.019494 15.1368 0.12098 0.00015708 0.76918 0.00915 0.010134 0.0013986 0.98678 0.9916 3.0174e-006 1.2069e-005 0.16291 0.88613 0.89591 0.0014036 0.97725 0.45659 0.0018907 0.42324 2.0255 2.0244 16.0169 144.9232 0.00019532 -85.5988 0.58495
7.689 0.98813 5.4713e-005 3.8183 0.011933 0.00010008 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.514 0.5446 0.16662 0.019496 15.1396 0.12099 0.00015709 0.76917 0.0091504 0.010134 0.0013985 0.98679 0.9916 3.0171e-006 1.2068e-005 0.16291 0.88644 0.89604 0.0014035 0.97738 0.45677 0.0018907 0.42325 2.0262 2.0252 16.0169 144.9232 0.00019512 -85.5993 0.58595
7.69 0.98813 5.4713e-005 3.8183 0.011933 0.00010009 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5141 0.54465 0.16663 0.019497 15.1425 0.12099 0.0001571 0.76916 0.0091508 0.010135 0.0013984 0.98679 0.9916 3.0169e-006 1.2067e-005 0.16292 0.88674 0.89617 0.0014033 0.9775 0.45696 0.0018906 0.42327 2.027 2.0259 16.0168 144.9232 0.00019491 -85.5998 0.58695
7.691 0.98813 5.4713e-005 3.8183 0.011933 0.00010011 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5142 0.54469 0.16665 0.019498 15.1453 0.121 0.00015711 0.76916 0.0091512 0.010135 0.0013983 0.98679 0.9916 3.0166e-006 1.2066e-005 0.16292 0.88704 0.89631 0.0014032 0.97763 0.45715 0.0018905 0.42328 2.0277 2.0267 16.0168 144.9232 0.00019471 -85.6002 0.58795
7.692 0.98813 5.4713e-005 3.8183 0.011933 0.00010012 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5143 0.54474 0.16666 0.019499 15.1481 0.12101 0.00015712 0.76915 0.0091516 0.010136 0.0013982 0.98679 0.9916 3.0164e-006 1.2065e-005 0.16292 0.88734 0.89644 0.0014031 0.97776 0.45734 0.0018904 0.4233 2.0284 2.0274 16.0168 144.9233 0.00019451 -85.6007 0.58895
7.693 0.98813 5.4713e-005 3.8183 0.011933 0.00010013 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5143 0.54478 0.16668 0.0195 15.151 0.12101 0.00015713 0.76914 0.009152 0.010136 0.0013981 0.98679 0.99161 3.0161e-006 1.2064e-005 0.16293 0.88765 0.89657 0.0014031 0.97788 0.45753 0.0018904 0.42331 2.0292 2.0281 16.0168 144.9233 0.0001943 -85.6011 0.58995
7.694 0.98813 5.4713e-005 3.8183 0.011933 0.00010014 0.0011706 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5144 0.54483 0.16669 0.019501 15.1538 0.12102 0.00015714 0.76914 0.0091524 0.010137 0.001398 0.98679 0.99161 3.0159e-006 1.2064e-005 0.16293 0.88794 0.8967 0.001403 0.97801 0.45772 0.0018903 0.42333 2.0299 2.0289 16.0168 144.9233 0.0001941 -85.6016 0.59095
7.695 0.98813 5.4713e-005 3.8183 0.011933 0.00010016 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5145 0.54487 0.1667 0.019502 15.1567 0.12103 0.00015715 0.76913 0.0091528 0.010137 0.0013979 0.98679 0.99161 3.0157e-006 1.2063e-005 0.16293 0.88824 0.89683 0.001403 0.97813 0.45791 0.0018902 0.42334 2.0306 2.0296 16.0167 144.9233 0.0001939 -85.602 0.59195
7.696 0.98813 5.4713e-005 3.8183 0.011933 0.00010017 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5146 0.54492 0.16672 0.019504 15.1595 0.12103 0.00015716 0.76912 0.0091533 0.010138 0.0013978 0.9868 0.99161 3.0154e-006 1.2062e-005 0.16294 0.88854 0.89696 0.001403 0.97826 0.4581 0.0018901 0.42336 2.0314 2.0303 16.0167 144.9233 0.0001937 -85.6025 0.59295
7.697 0.98813 5.4712e-005 3.8183 0.011933 0.00010018 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5147 0.54496 0.16673 0.019505 15.1623 0.12104 0.00015717 0.76912 0.0091537 0.010138 0.0013977 0.9868 0.99161 3.0152e-006 1.2061e-005 0.16294 0.88884 0.89709 0.001403 0.97838 0.45828 0.0018901 0.42337 2.0321 2.031 16.0167 144.9234 0.0001935 -85.6029 0.59395
7.698 0.98813 5.4712e-005 3.8183 0.011933 0.0001002 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5148 0.54501 0.16674 0.019506 15.1652 0.12105 0.00015718 0.76911 0.0091541 0.010138 0.0013976 0.9868 0.99161 3.015e-006 1.206e-005 0.16294 0.88913 0.89721 0.001403 0.9785 0.45847 0.00189 0.42339 2.0328 2.0318 16.0167 144.9234 0.00019331 -85.6033 0.59495
7.699 0.98813 5.4712e-005 3.8183 0.011933 0.00010021 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5149 0.54505 0.16676 0.019507 15.168 0.12106 0.00015719 0.7691 0.0091545 0.010139 0.0013975 0.9868 0.99161 3.0147e-006 1.2059e-005 0.16295 0.88943 0.89734 0.001403 0.97862 0.45866 0.0018899 0.4234 2.0335 2.0325 16.0167 144.9234 0.00019311 -85.6038 0.59595
7.7 0.98813 5.4712e-005 3.8183 0.011933 0.00010022 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.515 0.5451 0.16677 0.019508 15.1709 0.12106 0.0001572 0.76909 0.0091549 0.010139 0.0013974 0.9868 0.99161 3.0145e-006 1.2058e-005 0.16295 0.88972 0.89747 0.0014029 0.97874 0.45885 0.0018899 0.42341 2.0342 2.0332 16.0167 144.9234 0.00019291 -85.6042 0.59695
7.701 0.98813 5.4712e-005 3.8183 0.011933 0.00010023 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.515 0.54514 0.16679 0.019509 15.1737 0.12107 0.00015721 0.76909 0.0091553 0.01014 0.0013973 0.9868 0.99161 3.0143e-006 1.2057e-005 0.16295 0.89002 0.8976 0.0014029 0.97886 0.45904 0.0018898 0.42343 2.035 2.0339 16.0166 144.9234 0.00019272 -85.6046 0.59795
7.702 0.98813 5.4712e-005 3.8183 0.011933 0.00010025 0.0011706 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5151 0.54519 0.1668 0.01951 15.1765 0.12108 0.00015723 0.76908 0.0091557 0.01014 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.16296 0.89031 0.89772 0.0014029 0.97898 0.45923 0.0018897 0.42344 2.0357 2.0347 16.0166 144.9235 0.00019252 -85.6051 0.59895
7.703 0.98813 5.4712e-005 3.8183 0.011933 0.00010026 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5152 0.54523 0.16681 0.019512 15.1794 0.12108 0.00015724 0.76907 0.0091561 0.010141 0.0013971 0.9868 0.99161 3.0138e-006 1.2055e-005 0.16296 0.8906 0.89785 0.0014028 0.9791 0.45941 0.0018897 0.42346 2.0364 2.0354 16.0166 144.9235 0.00019233 -85.6055 0.59995
7.704 0.98813 5.4712e-005 3.8183 0.011933 0.00010027 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5153 0.54528 0.16683 0.019513 15.1822 0.12109 0.00015725 0.76907 0.0091565 0.010141 0.001397 0.98681 0.99162 3.0136e-006 1.2054e-005 0.16296 0.89089 0.89797 0.0014028 0.97922 0.4596 0.0018896 0.42347 2.0371 2.0361 16.0166 144.9235 0.00019213 -85.6059 0.60095
7.705 0.98813 5.4712e-005 3.8183 0.011933 0.00010029 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5154 0.54532 0.16684 0.019514 15.1851 0.1211 0.00015726 0.76906 0.009157 0.010141 0.0013969 0.98681 0.99162 3.0134e-006 1.2053e-005 0.16297 0.89118 0.8981 0.0014027 0.97933 0.45979 0.0018895 0.42349 2.0378 2.0368 16.0166 144.9235 0.00019194 -85.6063 0.60195
7.706 0.98813 5.4712e-005 3.8183 0.011933 0.0001003 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5155 0.54537 0.16685 0.019515 15.1879 0.1211 0.00015727 0.76905 0.0091574 0.010142 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.16297 0.89147 0.89822 0.0014027 0.97945 0.45998 0.0018895 0.4235 2.0385 2.0375 16.0165 144.9235 0.00019175 -85.6067 0.60295
7.707 0.98813 5.4712e-005 3.8183 0.011933 0.00010031 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5156 0.54541 0.16687 0.019516 15.1908 0.12111 0.00015728 0.76905 0.0091578 0.010142 0.0013967 0.98681 0.99162 3.0129e-006 1.2052e-005 0.16297 0.89175 0.89835 0.0014026 0.97956 0.46017 0.0018894 0.42352 2.0392 2.0382 16.0165 144.9236 0.00019156 -85.6071 0.60395
7.708 0.98813 5.4712e-005 3.8183 0.011933 0.00010032 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5157 0.54546 0.16688 0.019517 15.1936 0.12112 0.00015729 0.76904 0.0091582 0.010143 0.0013966 0.98681 0.99162 3.0127e-006 1.2051e-005 0.16298 0.89204 0.89847 0.0014025 0.97968 0.46035 0.0018893 0.42353 2.0399 2.0389 16.0165 144.9236 0.00019137 -85.6075 0.60495
7.709 0.98813 5.4711e-005 3.8183 0.011933 0.00010034 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5157 0.5455 0.1669 0.019519 15.1964 0.12112 0.0001573 0.76903 0.0091586 0.010143 0.0013965 0.98681 0.99162 3.0125e-006 1.205e-005 0.16298 0.89233 0.89859 0.0014024 0.97979 0.46054 0.0018893 0.42355 2.0406 2.0396 16.0165 144.9236 0.00019118 -85.608 0.60595
7.71 0.98813 5.4711e-005 3.8183 0.011933 0.00010035 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5158 0.54555 0.16691 0.01952 15.1993 0.12113 0.00015731 0.76903 0.009159 0.010144 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.16298 0.89261 0.89872 0.0014024 0.9799 0.46073 0.0018892 0.42356 2.0413 2.0403 16.0165 144.9236 0.00019099 -85.6084 0.60695
7.711 0.98813 5.4711e-005 3.8183 0.011933 0.00010036 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5159 0.54559 0.16692 0.019521 15.2021 0.12114 0.00015732 0.76902 0.0091594 0.010144 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.16298 0.8929 0.89884 0.0014023 0.98001 0.46092 0.0018891 0.42358 2.042 2.041 16.0164 144.9236 0.0001908 -85.6088 0.60795
7.712 0.98813 5.4711e-005 3.8183 0.011933 0.00010038 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.516 0.54564 0.16694 0.019522 15.205 0.12115 0.00015733 0.76901 0.0091598 0.010145 0.0013962 0.98682 0.99162 3.0119e-006 1.2047e-005 0.16299 0.89318 0.89896 0.0014022 0.98013 0.46111 0.0018891 0.42359 2.0427 2.0417 16.0164 144.9237 0.00019061 -85.6091 0.60895
7.713 0.98813 5.4711e-005 3.8183 0.011933 0.00010039 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5161 0.54568 0.16695 0.019523 15.2078 0.12115 0.00015734 0.76901 0.0091602 0.010145 0.0013961 0.98682 0.99162 3.0117e-006 1.2047e-005 0.16299 0.89346 0.89908 0.0014022 0.98024 0.46129 0.001889 0.4236 2.0434 2.0424 16.0164 144.9237 0.00019043 -85.6095 0.60995
7.714 0.98813 5.4711e-005 3.8183 0.011933 0.0001004 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5162 0.54573 0.16697 0.019524 15.2107 0.12116 0.00015735 0.769 0.0091607 0.010145 0.001396 0.98682 0.99162 3.0115e-006 1.2046e-005 0.16299 0.89374 0.8992 0.0014022 0.98035 0.46148 0.0018889 0.42362 2.0441 2.0431 16.0164 144.9237 0.00019024 -85.6099 0.61095
7.715 0.98813 5.4711e-005 3.8183 0.011933 0.00010041 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5163 0.54577 0.16698 0.019525 15.2135 0.12117 0.00015736 0.76899 0.0091611 0.010146 0.0013959 0.98682 0.99162 3.0113e-006 1.2045e-005 0.163 0.89402 0.89932 0.0014021 0.98045 0.46167 0.0018889 0.42363 2.0448 2.0438 16.0164 144.9237 0.00019005 -85.6103 0.61195
7.716 0.98813 5.4711e-005 3.8183 0.011933 0.00010043 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5164 0.54582 0.16699 0.019527 15.2164 0.12117 0.00015737 0.76898 0.0091615 0.010146 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.163 0.8943 0.89944 0.0014021 0.98056 0.46186 0.0018888 0.42365 2.0455 2.0445 16.0163 144.9237 0.00018987 -85.6107 0.61295
7.717 0.98813 5.4711e-005 3.8183 0.011933 0.00010044 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5164 0.54586 0.16701 0.019528 15.2192 0.12118 0.00015738 0.76898 0.0091619 0.010147 0.0013958 0.98682 0.99163 3.0108e-006 1.2043e-005 0.163 0.89458 0.89956 0.0014021 0.98067 0.46204 0.0018888 0.42366 2.0462 2.0452 16.0163 144.9238 0.00018968 -85.6111 0.61395
7.718 0.98813 5.4711e-005 3.8183 0.011933 0.00010045 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5165 0.54591 0.16702 0.019529 15.2221 0.12119 0.00015739 0.76897 0.0091623 0.010147 0.0013957 0.98682 0.99163 3.0106e-006 1.2042e-005 0.16301 0.89486 0.89968 0.001402 0.98078 0.46223 0.0018887 0.42368 2.0469 2.0459 16.0163 144.9238 0.0001895 -85.6115 0.61495
7.719 0.98813 5.4711e-005 3.8183 0.011933 0.00010046 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5166 0.54596 0.16703 0.01953 15.2249 0.12119 0.0001574 0.76896 0.0091627 0.010148 0.0013956 0.98682 0.99163 3.0104e-006 1.2042e-005 0.16301 0.89514 0.8998 0.001402 0.98088 0.46242 0.0018886 0.42369 2.0475 2.0466 16.0163 144.9238 0.00018932 -85.6118 0.61595
7.72 0.98813 5.4711e-005 3.8183 0.011933 0.00010048 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5167 0.546 0.16705 0.019531 15.2278 0.1212 0.00015741 0.76896 0.0091631 0.010148 0.0013955 0.98682 0.99163 3.0102e-006 1.2041e-005 0.16301 0.89541 0.89992 0.001402 0.98099 0.4626 0.0018886 0.42371 2.0482 2.0473 16.0163 144.9238 0.00018914 -85.6122 0.61695
7.721 0.98813 5.4711e-005 3.8183 0.011933 0.00010049 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5168 0.54605 0.16706 0.019532 15.2306 0.12121 0.00015742 0.76895 0.0091635 0.010148 0.0013954 0.98683 0.99163 3.01e-006 1.204e-005 0.16302 0.89569 0.90004 0.0014019 0.98109 0.46279 0.0018885 0.42372 2.0489 2.0479 16.0162 144.9238 0.00018895 -85.6126 0.61795
7.722 0.98813 5.471e-005 3.8183 0.011933 0.0001005 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5169 0.54609 0.16708 0.019533 15.2334 0.12121 0.00015743 0.76894 0.0091639 0.010149 0.0013953 0.98683 0.99163 3.0098e-006 1.2039e-005 0.16302 0.89596 0.90015 0.0014019 0.9812 0.46298 0.0018885 0.42374 2.0496 2.0486 16.0162 144.9239 0.00018877 -85.613 0.61895
7.723 0.98813 5.471e-005 3.8183 0.011933 0.00010052 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.517 0.54614 0.16709 0.019535 15.2363 0.12122 0.00015744 0.76894 0.0091644 0.010149 0.0013952 0.98683 0.99163 3.0097e-006 1.2039e-005 0.16302 0.89624 0.90027 0.0014019 0.9813 0.46317 0.0018884 0.42375 2.0503 2.0493 16.0162 144.9239 0.00018859 -85.6133 0.61995
7.724 0.98813 5.471e-005 3.8183 0.011933 0.00010053 0.0011707 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.517 0.54618 0.1671 0.019536 15.2391 0.12123 0.00015745 0.76893 0.0091648 0.01015 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.16303 0.89651 0.90039 0.0014018 0.98141 0.46335 0.0018883 0.42377 2.0509 2.05 16.0162 144.9239 0.00018841 -85.6137 0.62095
7.725 0.98813 5.471e-005 3.8183 0.011933 0.00010054 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5171 0.54623 0.16712 0.019537 15.242 0.12123 0.00015746 0.76892 0.0091652 0.01015 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.16303 0.89678 0.9005 0.0014017 0.98151 0.46354 0.0018883 0.42378 2.0516 2.0507 16.0162 144.9239 0.00018824 -85.6141 0.62195
7.726 0.98813 5.471e-005 3.8183 0.011933 0.00010055 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5172 0.54627 0.16713 0.019538 15.2448 0.12124 0.00015747 0.76892 0.0091656 0.010151 0.001395 0.98683 0.99163 3.0091e-006 1.2036e-005 0.16303 0.89705 0.90062 0.0014017 0.98161 0.46373 0.0018882 0.42379 2.0523 2.0513 16.0161 144.9239 0.00018806 -85.6144 0.62295
7.727 0.98813 5.471e-005 3.8183 0.011933 0.00010057 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5173 0.54632 0.16714 0.019539 15.2477 0.12125 0.00015748 0.76891 0.009166 0.010151 0.0013949 0.98683 0.99163 3.0089e-006 1.2035e-005 0.16304 0.89732 0.90073 0.0014016 0.98171 0.46391 0.0018882 0.42381 2.053 2.052 16.0161 144.924 0.00018788 -85.6148 0.62395
7.728 0.98813 5.471e-005 3.8183 0.011933 0.00010058 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5174 0.54636 0.16716 0.01954 15.2505 0.12126 0.00015749 0.7689 0.0091664 0.010152 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.16304 0.89759 0.90085 0.0014016 0.98181 0.4641 0.0018881 0.42382 2.0536 2.0527 16.0161 144.924 0.0001877 -85.6151 0.62495
7.729 0.98813 5.471e-005 3.8183 0.011933 0.00010059 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5175 0.54641 0.16717 0.019541 15.2534 0.12126 0.0001575 0.7689 0.0091668 0.010152 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.16304 0.89786 0.90096 0.0014015 0.98191 0.46429 0.0018881 0.42384 2.0543 2.0534 16.0161 144.924 0.00018753 -85.6155 0.62595
7.73 0.98813 5.471e-005 3.8183 0.011933 0.00010061 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5176 0.54645 0.16719 0.019543 15.2562 0.12127 0.00015751 0.76889 0.0091672 0.010152 0.0013947 0.98684 0.99163 3.0083e-006 1.2033e-005 0.16305 0.89813 0.90107 0.0014015 0.98201 0.46447 0.001888 0.42385 2.055 2.054 16.0161 144.924 0.00018735 -85.6158 0.62695
7.731 0.98813 5.471e-005 3.8183 0.011933 0.00010062 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5177 0.5465 0.1672 0.019544 15.2591 0.12128 0.00015753 0.76888 0.0091676 0.010153 0.0013946 0.98684 0.99164 3.0081e-006 1.2032e-005 0.16305 0.89839 0.90119 0.0014014 0.98211 0.46466 0.0018879 0.42387 2.0556 2.0547 16.016 144.924 0.00018718 -85.6162 0.62795
7.732 0.98813 5.471e-005 3.8183 0.011933 0.00010063 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5177 0.54654 0.16721 0.019545 15.262 0.12128 0.00015754 0.76887 0.009168 0.010153 0.0013945 0.98684 0.99164 3.008e-006 1.2032e-005 0.16305 0.89866 0.9013 0.0014014 0.98221 0.46484 0.0018879 0.42388 2.0563 2.0554 16.016 144.9241 0.000187 -85.6165 0.62895
7.733 0.98813 5.471e-005 3.8183 0.011933 0.00010064 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5178 0.54659 0.16723 0.019546 15.2648 0.12129 0.00015755 0.76887 0.0091685 0.010154 0.0013944 0.98684 0.99164 3.0078e-006 1.2031e-005 0.16305 0.89892 0.90141 0.0014013 0.9823 0.46503 0.0018878 0.4239 2.057 2.056 16.016 144.9241 0.00018683 -85.6169 0.62995
7.734 0.98813 5.4709e-005 3.8183 0.011933 0.00010066 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5179 0.54663 0.16724 0.019547 15.2677 0.1213 0.00015756 0.76886 0.0091689 0.010154 0.0013943 0.98684 0.99164 3.0076e-006 1.203e-005 0.16306 0.89919 0.90153 0.0014013 0.9824 0.46522 0.0018878 0.42391 2.0576 2.0567 16.016 144.9241 0.00018666 -85.6172 0.63095
7.735 0.98813 5.4709e-005 3.8183 0.011933 0.00010067 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.518 0.54668 0.16725 0.019548 15.2705 0.1213 0.00015757 0.76885 0.0091693 0.010155 0.0013943 0.98684 0.99164 3.0074e-006 1.203e-005 0.16306 0.89945 0.90164 0.0014013 0.98249 0.4654 0.0018877 0.42393 2.0583 2.0573 16.0159 144.9241 0.00018649 -85.6175 0.63195
7.736 0.98813 5.4709e-005 3.8183 0.011933 0.00010068 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5181 0.54672 0.16727 0.01955 15.2734 0.12131 0.00015758 0.76885 0.0091697 0.010155 0.0013942 0.98684 0.99164 3.0072e-006 1.2029e-005 0.16306 0.89972 0.90175 0.0014012 0.98259 0.46559 0.0018877 0.42394 2.0589 2.058 16.0159 144.9242 0.00018631 -85.6179 0.63295
7.737 0.98813 5.4709e-005 3.8183 0.011932 0.0001007 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5182 0.54677 0.16728 0.019551 15.2762 0.12132 0.00015759 0.76884 0.0091701 0.010155 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.16307 0.89998 0.90186 0.0014012 0.98268 0.46578 0.0018876 0.42395 2.0596 2.0587 16.0159 144.9242 0.00018614 -85.6182 0.63395
7.738 0.98813 5.4709e-005 3.8183 0.011932 0.00010071 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5183 0.54681 0.1673 0.019552 15.2791 0.12132 0.0001576 0.76883 0.0091705 0.010156 0.001394 0.98684 0.99164 3.0069e-006 1.2027e-005 0.16307 0.90024 0.90197 0.0014012 0.98278 0.46596 0.0018876 0.42397 2.0602 2.0593 16.0159 144.9242 0.00018597 -85.6185 0.63495
7.739 0.98813 5.4709e-005 3.8183 0.011932 0.00010072 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5184 0.54686 0.16731 0.019553 15.2819 0.12133 0.00015761 0.76883 0.0091709 0.010156 0.0013939 0.98684 0.99164 3.0067e-006 1.2027e-005 0.16307 0.9005 0.90208 0.0014011 0.98287 0.46615 0.0018875 0.42398 2.0609 2.06 16.0159 144.9242 0.0001858 -85.6189 0.63595
7.74 0.98813 5.4709e-005 3.8183 0.011932 0.00010073 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5184 0.5469 0.16732 0.019554 15.2848 0.12134 0.00015762 0.76882 0.0091713 0.010157 0.0013939 0.98685 0.99164 3.0065e-006 1.2026e-005 0.16308 0.90076 0.90219 0.0014011 0.98296 0.46633 0.0018875 0.424 2.0615 2.0606 16.0158 144.9242 0.00018564 -85.6192 0.63695
7.741 0.98813 5.4709e-005 3.8183 0.011932 0.00010075 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5185 0.54695 0.16734 0.019555 15.2876 0.12134 0.00015763 0.76881 0.0091717 0.010157 0.0013938 0.98685 0.99164 3.0064e-006 1.2025e-005 0.16308 0.90102 0.9023 0.0014011 0.98306 0.46652 0.0018874 0.42401 2.0622 2.0613 16.0158 144.9243 0.00018547 -85.6195 0.63795
7.742 0.98813 5.4709e-005 3.8183 0.011932 0.00010076 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5186 0.54699 0.16735 0.019556 15.2905 0.12135 0.00015764 0.76881 0.0091721 0.010158 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.16308 0.90127 0.90241 0.001401 0.98315 0.4667 0.0018874 0.42403 2.0628 2.0619 16.0158 144.9243 0.0001853 -85.6198 0.63895
7.743 0.98813 5.4709e-005 3.8183 0.011932 0.00010077 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5187 0.54704 0.16736 0.019558 15.2933 0.12136 0.00015765 0.7688 0.0091725 0.010158 0.0013936 0.98685 0.99164 3.006e-006 1.2024e-005 0.16309 0.90153 0.90251 0.001401 0.98324 0.46689 0.0018873 0.42404 2.0635 2.0626 16.0158 144.9243 0.00018513 -85.6201 0.63995
7.744 0.98813 5.4709e-005 3.8183 0.011932 0.00010079 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5188 0.54708 0.16738 0.019559 15.2962 0.12137 0.00015766 0.76879 0.009173 0.010159 0.0013936 0.98685 0.99164 3.0059e-006 1.2023e-005 0.16309 0.90179 0.90262 0.0014009 0.98333 0.46708 0.0018873 0.42406 2.0641 2.0632 16.0158 144.9243 0.00018497 -85.6205 0.64095
7.745 0.98813 5.4709e-005 3.8183 0.011932 0.0001008 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5189 0.54713 0.16739 0.01956 15.2991 0.12137 0.00015767 0.76879 0.0091734 0.010159 0.0013935 0.98685 0.99164 3.0057e-006 1.2023e-005 0.16309 0.90204 0.90273 0.0014009 0.98342 0.46726 0.0018872 0.42407 2.0648 2.0639 16.0157 144.9243 0.0001848 -85.6208 0.64195
7.746 0.98813 5.4708e-005 3.8183 0.011932 0.00010081 0.0011708 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.519 0.54717 0.16741 0.019561 15.3019 0.12138 0.00015768 0.76878 0.0091738 0.010159 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.1631 0.9023 0.90284 0.0014008 0.98351 0.46745 0.0018872 0.42408 2.0654 2.0645 16.0157 144.9244 0.00018464 -85.6211 0.64295
7.747 0.98813 5.4708e-005 3.8183 0.011932 0.00010082 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5191 0.54722 0.16742 0.019562 15.3048 0.12139 0.00015769 0.76877 0.0091742 0.01016 0.0013934 0.98685 0.99165 3.0054e-006 1.2021e-005 0.1631 0.90255 0.90294 0.0014008 0.9836 0.46763 0.0018871 0.4241 2.0661 2.0652 16.0157 144.9244 0.00018447 -85.6214 0.64395
7.748 0.98813 5.4708e-005 3.8183 0.011932 0.00010084 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5191 0.54726 0.16743 0.019563 15.3076 0.12139 0.0001577 0.76877 0.0091746 0.01016 0.0013933 0.98685 0.99165 3.0052e-006 1.2021e-005 0.1631 0.9028 0.90305 0.0014008 0.98369 0.46782 0.0018871 0.42411 2.0667 2.0658 16.0157 144.9244 0.00018431 -85.6217 0.64495
7.749 0.98813 5.4708e-005 3.8183 0.011932 0.00010085 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5192 0.54731 0.16745 0.019564 15.3105 0.1214 0.00015771 0.76876 0.009175 0.010161 0.0013932 0.98685 0.99165 3.005e-006 1.202e-005 0.16311 0.90306 0.90316 0.0014007 0.98377 0.468 0.001887 0.42413 2.0673 2.0664 16.0156 144.9244 0.00018414 -85.622 0.64595
7.75 0.98813 5.4708e-005 3.8183 0.011932 0.00010086 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5193 0.54735 0.16746 0.019566 15.3133 0.12141 0.00015772 0.76875 0.0091754 0.010161 0.0013931 0.98686 0.99165 3.0049e-006 1.2019e-005 0.16311 0.90331 0.90326 0.0014007 0.98386 0.46819 0.001887 0.42414 2.068 2.0671 16.0156 144.9244 0.00018398 -85.6223 0.64695
7.751 0.98813 5.4708e-005 3.8183 0.011932 0.00010088 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5194 0.5474 0.16748 0.019567 15.3162 0.12141 0.00015773 0.76874 0.0091758 0.010162 0.0013931 0.98686 0.99165 3.0047e-006 1.2019e-005 0.16311 0.90356 0.90337 0.0014007 0.98395 0.46837 0.0018869 0.42416 2.0686 2.0677 16.0156 144.9245 0.00018382 -85.6226 0.64795
7.752 0.98813 5.4708e-005 3.8183 0.011932 0.00010089 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5195 0.54744 0.16749 0.019568 15.3191 0.12142 0.00015774 0.76874 0.0091762 0.010162 0.001393 0.98686 0.99165 3.0046e-006 1.2018e-005 0.16311 0.90381 0.90347 0.0014006 0.98403 0.46856 0.0018869 0.42417 2.0692 2.0683 16.0156 144.9245 0.00018366 -85.6229 0.64895
7.753 0.98813 5.4708e-005 3.8183 0.011932 0.0001009 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5196 0.54749 0.1675 0.019569 15.3219 0.12143 0.00015775 0.76873 0.0091766 0.010162 0.0013929 0.98686 0.99165 3.0044e-006 1.2017e-005 0.16312 0.90406 0.90358 0.0014006 0.98412 0.46874 0.0018868 0.42419 2.0699 2.069 16.0156 144.9245 0.0001835 -85.6232 0.64995
7.754 0.98813 5.4708e-005 3.8183 0.011932 0.00010091 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5197 0.54753 0.16752 0.01957 15.3248 0.12143 0.00015776 0.76872 0.009177 0.010163 0.0013929 0.98686 0.99165 3.0042e-006 1.2017e-005 0.16312 0.90431 0.90368 0.0014006 0.9842 0.46893 0.0018868 0.4242 2.0705 2.0696 16.0155 144.9245 0.00018334 -85.6235 0.65095
7.755 0.98813 5.4708e-005 3.8183 0.011932 0.00010093 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5198 0.54758 0.16753 0.019571 15.3276 0.12144 0.00015777 0.76872 0.0091774 0.010163 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.16312 0.90455 0.90378 0.0014005 0.98429 0.46911 0.0018867 0.42422 2.0711 2.0702 16.0155 144.9245 0.00018318 -85.6238 0.65195
7.756 0.98813 5.4708e-005 3.8183 0.011932 0.00010094 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5198 0.54763 0.16754 0.019572 15.3305 0.12145 0.00015778 0.76871 0.0091779 0.010164 0.0013927 0.98686 0.99165 3.0039e-006 1.2016e-005 0.16313 0.9048 0.90389 0.0014005 0.98437 0.4693 0.0018867 0.42423 2.0717 2.0709 16.0155 144.9246 0.00018302 -85.6241 0.65295
7.757 0.98813 5.4708e-005 3.8183 0.011932 0.00010095 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5199 0.54767 0.16756 0.019574 15.3334 0.12145 0.00015779 0.7687 0.0091783 0.010164 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.16313 0.90505 0.90399 0.0014004 0.98445 0.46948 0.0018866 0.42424 2.0724 2.0715 16.0155 144.9246 0.00018286 -85.6244 0.65395
7.758 0.98813 5.4708e-005 3.8183 0.011932 0.00010097 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.52 0.54772 0.16757 0.019575 15.3362 0.12146 0.0001578 0.7687 0.0091787 0.010165 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.16313 0.90529 0.90409 0.0014004 0.98454 0.46967 0.0018866 0.42426 2.073 2.0721 16.0154 144.9246 0.0001827 -85.6247 0.65495
7.759 0.98813 5.4707e-005 3.8183 0.011932 0.00010098 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5201 0.54776 0.16759 0.019576 15.3391 0.12147 0.00015781 0.76869 0.0091791 0.010165 0.0013925 0.98686 0.99165 3.0035e-006 1.2014e-005 0.16314 0.90554 0.90419 0.0014004 0.98462 0.46985 0.0018865 0.42427 2.0736 2.0727 16.0154 144.9246 0.00018254 -85.6249 0.65595
7.76 0.98813 5.4707e-005 3.8183 0.011932 0.00010099 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5202 0.54781 0.1676 0.019577 15.3419 0.12147 0.00015782 0.76868 0.0091795 0.010165 0.0013925 0.98686 0.99165 3.0033e-006 1.2013e-005 0.16314 0.90578 0.90429 0.0014003 0.9847 0.47004 0.0018865 0.42429 2.0742 2.0734 16.0154 144.9246 0.00018239 -85.6252 0.65695
7.761 0.98813 5.4707e-005 3.8183 0.011932 0.000101 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5203 0.54785 0.16761 0.019578 15.3448 0.12148 0.00015783 0.76868 0.0091799 0.010166 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.16314 0.90602 0.9044 0.0014003 0.98478 0.47022 0.0018864 0.4243 2.0748 2.074 16.0154 144.9247 0.00018223 -85.6255 0.65795
7.762 0.98813 5.4707e-005 3.8183 0.011932 0.00010102 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5204 0.5479 0.16763 0.019579 15.3477 0.12149 0.00015785 0.76867 0.0091803 0.010166 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.16315 0.90626 0.9045 0.0014003 0.98486 0.47041 0.0018864 0.42432 2.0755 2.0746 16.0153 144.9247 0.00018208 -85.6258 0.65895
7.763 0.98813 5.4707e-005 3.8183 0.011932 0.00010103 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5205 0.54794 0.16764 0.01958 15.3505 0.1215 0.00015786 0.76866 0.0091807 0.010167 0.0013923 0.98687 0.99165 3.0029e-006 1.2011e-005 0.16315 0.90651 0.9046 0.0014002 0.98494 0.47059 0.0018864 0.42433 2.0761 2.0752 16.0153 144.9247 0.00018192 -85.6261 0.65995
7.764 0.98813 5.4707e-005 3.8183 0.011932 0.00010104 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5205 0.54799 0.16765 0.019582 15.3534 0.1215 0.00015787 0.76866 0.0091811 0.010167 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.16315 0.90675 0.9047 0.0014002 0.98502 0.47078 0.0018863 0.42435 2.0767 2.0758 16.0153 144.9247 0.00018177 -85.6263 0.66095
7.765 0.98813 5.4707e-005 3.8183 0.011932 0.00010106 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5206 0.54803 0.16767 0.019583 15.3563 0.12151 0.00015788 0.76865 0.0091815 0.010168 0.0013921 0.98687 0.99166 3.0026e-006 1.201e-005 0.16316 0.90699 0.9048 0.0014002 0.9851 0.47096 0.0018863 0.42436 2.0773 2.0764 16.0153 144.9247 0.00018161 -85.6266 0.66195
7.766 0.98813 5.4707e-005 3.8183 0.011932 0.00010107 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5207 0.54808 0.16768 0.019584 15.3591 0.12152 0.00015789 0.76864 0.0091819 0.010168 0.0013921 0.98687 0.99166 3.0024e-006 1.201e-005 0.16316 0.90723 0.9049 0.0014001 0.98518 0.47114 0.0018862 0.42437 2.0779 2.0771 16.0153 144.9248 0.00018146 -85.6269 0.66295
7.767 0.98813 5.4707e-005 3.8183 0.011932 0.00010108 0.0011709 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5208 0.54812 0.1677 0.019585 15.362 0.12152 0.0001579 0.76864 0.0091823 0.010169 0.001392 0.98687 0.99166 3.0023e-006 1.2009e-005 0.16316 0.90746 0.905 0.0014001 0.98526 0.47133 0.0018862 0.42439 2.0785 2.0777 16.0152 144.9248 0.00018131 -85.6271 0.66395
7.768 0.98813 5.4707e-005 3.8183 0.011932 0.00010109 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5209 0.54817 0.16771 0.019586 15.3648 0.12153 0.00015791 0.76863 0.0091828 0.010169 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.16317 0.9077 0.90509 0.0014001 0.98533 0.47151 0.0018861 0.4244 2.0791 2.0783 16.0152 144.9248 0.00018115 -85.6274 0.66495
7.769 0.98813 5.4707e-005 3.8183 0.011932 0.00010111 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.521 0.54821 0.16772 0.019587 15.3677 0.12154 0.00015792 0.76862 0.0091832 0.010169 0.0013919 0.98687 0.99166 3.002e-006 1.2008e-005 0.16317 0.90794 0.90519 0.0014 0.98541 0.4717 0.0018861 0.42442 2.0797 2.0789 16.0152 144.9248 0.000181 -85.6277 0.66595
7.77 0.98813 5.4707e-005 3.8183 0.011932 0.00010112 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5211 0.54826 0.16774 0.019588 15.3706 0.12154 0.00015793 0.76861 0.0091836 0.01017 0.0013918 0.98687 0.99166 3.0019e-006 1.2007e-005 0.16317 0.90817 0.90529 0.0014 0.98549 0.47188 0.0018861 0.42443 2.0803 2.0795 16.0152 144.9248 0.00018085 -85.6279 0.66695
7.771 0.98813 5.4706e-005 3.8183 0.011932 0.00010113 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5211 0.5483 0.16775 0.01959 15.3734 0.12155 0.00015794 0.76861 0.009184 0.01017 0.0013918 0.98687 0.99166 3.0017e-006 1.2007e-005 0.16317 0.90841 0.90539 0.0014 0.98556 0.47206 0.001886 0.42445 2.081 2.0801 16.0151 144.9249 0.0001807 -85.6282 0.66795
7.772 0.98813 5.4706e-005 3.8183 0.011932 0.00010115 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5212 0.54835 0.16776 0.019591 15.3763 0.12156 0.00015795 0.7686 0.0091844 0.010171 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.16318 0.90865 0.90549 0.0014 0.98564 0.47225 0.001886 0.42446 2.0816 2.0807 16.0151 144.9249 0.00018055 -85.6285 0.66895
7.773 0.98813 5.4706e-005 3.8183 0.011932 0.00010116 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5213 0.54839 0.16778 0.019592 15.3792 0.12156 0.00015796 0.76859 0.0091848 0.010171 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.16318 0.90888 0.90558 0.0013999 0.98571 0.47243 0.0018859 0.42447 2.0822 2.0813 16.0151 144.9249 0.0001804 -85.6287 0.66995
7.774 0.98813 5.4706e-005 3.8183 0.011932 0.00010117 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5214 0.54844 0.16779 0.019593 15.382 0.12157 0.00015797 0.76859 0.0091852 0.010172 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.16318 0.90911 0.90568 0.0013999 0.98579 0.47262 0.0018859 0.42449 2.0828 2.0819 16.0151 144.9249 0.00018025 -85.629 0.67095
7.775 0.98813 5.4706e-005 3.8183 0.011932 0.00010118 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5215 0.54848 0.16781 0.019594 15.3849 0.12158 0.00015798 0.76858 0.0091856 0.010172 0.0013915 0.98688 0.99166 3.0012e-006 1.2005e-005 0.16319 0.90934 0.90577 0.0013999 0.98586 0.4728 0.0018858 0.4245 2.0834 2.0825 16.015 144.9249 0.0001801 -85.6292 0.67195
7.776 0.98813 5.4706e-005 3.8183 0.011932 0.0001012 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5216 0.54853 0.16782 0.019595 15.3878 0.12158 0.00015799 0.76857 0.009186 0.010172 0.0013915 0.98688 0.99166 3.0011e-006 1.2004e-005 0.16319 0.90958 0.90587 0.0013998 0.98593 0.47298 0.0018858 0.42452 2.0839 2.0831 16.015 144.925 0.00017996 -85.6295 0.67295
7.777 0.98813 5.4706e-005 3.8183 0.011932 0.00010121 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5217 0.54857 0.16783 0.019596 15.3906 0.12159 0.000158 0.76857 0.0091864 0.010173 0.0013914 0.98688 0.99166 3.0009e-006 1.2004e-005 0.16319 0.90981 0.90597 0.0013998 0.98601 0.47317 0.0018858 0.42453 2.0845 2.0837 16.015 144.925 0.00017981 -85.6297 0.67395
7.778 0.98813 5.4706e-005 3.8183 0.011932 0.00010122 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5218 0.54862 0.16785 0.019598 15.3935 0.1216 0.00015801 0.76856 0.0091868 0.010173 0.0013914 0.98688 0.99166 3.0008e-006 1.2003e-005 0.1632 0.91004 0.90606 0.0013998 0.98608 0.47335 0.0018857 0.42455 2.0851 2.0843 16.015 144.925 0.00017966 -85.63 0.67495
7.779 0.98813 5.4706e-005 3.8183 0.011932 0.00010124 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5218 0.54866 0.16786 0.019599 15.3964 0.1216 0.00015802 0.76855 0.0091872 0.010174 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.1632 0.91027 0.90616 0.0013997 0.98615 0.47353 0.0018857 0.42456 2.0857 2.0849 16.015 144.925 0.00017952 -85.6302 0.67595
7.78 0.98813 5.4706e-005 3.8183 0.011932 0.00010125 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5219 0.54871 0.16787 0.0196 15.3992 0.12161 0.00015803 0.76855 0.0091876 0.010174 0.0013913 0.98688 0.99166 3.0005e-006 1.2002e-005 0.1632 0.9105 0.90625 0.0013997 0.98622 0.47372 0.0018856 0.42458 2.0863 2.0855 16.0149 144.925 0.00017937 -85.6305 0.67695
7.781 0.98813 5.4706e-005 3.8183 0.011932 0.00010126 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.522 0.54875 0.16789 0.019601 15.4021 0.12162 0.00015804 0.76854 0.009188 0.010175 0.0013912 0.98688 0.99166 3.0004e-006 1.2002e-005 0.16321 0.91072 0.90634 0.0013997 0.9863 0.4739 0.0018856 0.42459 2.0869 2.0861 16.0149 144.9251 0.00017923 -85.6307 0.67795
7.782 0.98813 5.4706e-005 3.8183 0.011932 0.00010127 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5221 0.5488 0.1679 0.019602 15.405 0.12163 0.00015805 0.76853 0.0091884 0.010175 0.0013911 0.98688 0.99166 3.0003e-006 1.2001e-005 0.16321 0.91095 0.90644 0.0013996 0.98637 0.47408 0.0018856 0.4246 2.0875 2.0867 16.0149 144.9251 0.00017908 -85.631 0.67895
7.783 0.98813 5.4705e-005 3.8183 0.011932 0.00010129 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5222 0.54884 0.16792 0.019603 15.4078 0.12163 0.00015806 0.76853 0.0091889 0.010175 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.16321 0.91118 0.90653 0.0013996 0.98644 0.47427 0.0018855 0.42462 2.0881 2.0873 16.0149 144.9251 0.00017894 -85.6312 0.67995
7.784 0.98813 5.4705e-005 3.8183 0.011932 0.0001013 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5223 0.54889 0.16793 0.019604 15.4107 0.12164 0.00015807 0.76852 0.0091893 0.010176 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.16322 0.91141 0.90662 0.0013996 0.98651 0.47445 0.0018855 0.42463 2.0887 2.0879 16.0148 144.9251 0.00017879 -85.6314 0.68095
7.785 0.98813 5.4705e-005 3.8183 0.011932 0.00010131 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5224 0.54893 0.16794 0.019606 15.4136 0.12165 0.00015808 0.76851 0.0091897 0.010176 0.001391 0.98688 0.99167 2.9999e-006 1.1999e-005 0.16322 0.91163 0.90672 0.0013996 0.98658 0.47463 0.0018855 0.42465 2.0893 2.0884 16.0148 144.9251 0.00017865 -85.6317 0.68195
7.786 0.98813 5.4705e-005 3.8183 0.011932 0.00010133 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5225 0.54898 0.16796 0.019607 15.4165 0.12165 0.00015809 0.76851 0.0091901 0.010177 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.16322 0.91186 0.90681 0.0013995 0.98664 0.47481 0.0018854 0.42466 2.0898 2.089 16.0148 144.9252 0.00017851 -85.6319 0.68295
7.787 0.98813 5.4705e-005 3.8183 0.011932 0.00010134 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5225 0.54902 0.16797 0.019608 15.4193 0.12166 0.0001581 0.7685 0.0091905 0.010177 0.0013908 0.98688 0.99167 2.9996e-006 1.1998e-005 0.16322 0.91208 0.9069 0.0013995 0.98671 0.475 0.0018854 0.42468 2.0904 2.0896 16.0148 144.9252 0.00017837 -85.6321 0.68395
7.788 0.98813 5.4705e-005 3.8183 0.011932 0.00010135 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5226 0.54907 0.16798 0.019609 15.4222 0.12167 0.00015811 0.76849 0.0091909 0.010178 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.16323 0.9123 0.90699 0.0013995 0.98678 0.47518 0.0018853 0.42469 2.091 2.0902 16.0147 144.9252 0.00017823 -85.6324 0.68495
7.789 0.98813 5.4705e-005 3.8183 0.011932 0.00010136 0.001171 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5227 0.54911 0.168 0.01961 15.4251 0.12167 0.00015812 0.76848 0.0091913 0.010178 0.0013907 0.98689 0.99167 2.9994e-006 1.1997e-005 0.16323 0.91253 0.90708 0.0013994 0.98685 0.47536 0.0018853 0.4247 2.0916 2.0908 16.0147 144.9252 0.00017808 -85.6326 0.68595
7.79 0.98813 5.4705e-005 3.8183 0.011932 0.00010138 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5228 0.54916 0.16801 0.019611 15.4279 0.12168 0.00015813 0.76848 0.0091917 0.010178 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.16323 0.91275 0.90718 0.0013994 0.98691 0.47555 0.0018853 0.42472 2.0922 2.0914 16.0147 144.9252 0.00017794 -85.6328 0.68695
7.791 0.98813 5.4705e-005 3.8183 0.011932 0.00010139 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5229 0.5492 0.16803 0.019612 15.4308 0.12169 0.00015814 0.76847 0.0091921 0.010179 0.0013906 0.98689 0.99167 2.9992e-006 1.1997e-005 0.16324 0.91297 0.90727 0.0013994 0.98698 0.47573 0.0018852 0.42473 2.0927 2.0919 16.0147 144.9253 0.0001778 -85.6331 0.68795
7.792 0.98813 5.4705e-005 3.8183 0.011932 0.0001014 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.523 0.54925 0.16804 0.019614 15.4337 0.12169 0.00015815 0.76846 0.0091925 0.010179 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.16324 0.91319 0.90736 0.0013994 0.98705 0.47591 0.0018852 0.42475 2.0933 2.0925 16.0146 144.9253 0.00017767 -85.6333 0.68895
7.793 0.98813 5.4705e-005 3.8183 0.011932 0.00010141 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5231 0.54929 0.16805 0.019615 15.4366 0.1217 0.00015816 0.76846 0.0091929 0.01018 0.0013905 0.98689 0.99167 2.9989e-006 1.1996e-005 0.16324 0.91341 0.90745 0.0013993 0.98711 0.47609 0.0018852 0.42476 2.0939 2.0931 16.0146 144.9253 0.00017753 -85.6335 0.68995
7.794 0.98813 5.4705e-005 3.8183 0.011932 0.00010143 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5232 0.54934 0.16807 0.019616 15.4394 0.12171 0.00015817 0.76845 0.0091933 0.01018 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.16325 0.91363 0.90754 0.0013993 0.98718 0.47628 0.0018851 0.42478 2.0945 2.0937 16.0146 144.9253 0.00017739 -85.6337 0.69095
7.795 0.98813 5.4705e-005 3.8183 0.011931 0.00010144 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5232 0.54938 0.16808 0.019617 15.4423 0.12171 0.00015818 0.76844 0.0091937 0.010181 0.0013904 0.98689 0.99167 2.9987e-006 1.1995e-005 0.16325 0.91385 0.90763 0.0013993 0.98724 0.47646 0.0018851 0.42479 2.095 2.0942 16.0146 144.9254 0.00017725 -85.6339 0.69195
7.796 0.98813 5.4704e-005 3.8183 0.011931 0.00010145 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5233 0.54943 0.16809 0.019618 15.4452 0.12172 0.0001582 0.76844 0.0091941 0.010181 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.16325 0.91406 0.90771 0.0013993 0.98731 0.47664 0.0018851 0.4248 2.0956 2.0948 16.0145 144.9254 0.00017711 -85.6342 0.69295
7.797 0.98813 5.4704e-005 3.8183 0.011931 0.00010147 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5234 0.54947 0.16811 0.019619 15.4481 0.12173 0.00015821 0.76843 0.0091945 0.010182 0.0013903 0.98689 0.99167 2.9985e-006 1.1994e-005 0.16326 0.91428 0.9078 0.0013992 0.98737 0.47682 0.001885 0.42482 2.0962 2.0954 16.0145 144.9254 0.00017698 -85.6344 0.69395
7.798 0.98813 5.4704e-005 3.8183 0.011931 0.00010148 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5235 0.54952 0.16812 0.01962 15.4509 0.12173 0.00015822 0.76842 0.0091949 0.010182 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.16326 0.9145 0.90789 0.0013992 0.98744 0.47701 0.001885 0.42483 2.0967 2.096 16.0145 144.9254 0.00017684 -85.6346 0.69495
7.799 0.98813 5.4704e-005 3.8183 0.011931 0.00010149 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5236 0.54956 0.16814 0.019621 15.4538 0.12174 0.00015823 0.76842 0.0091954 0.010182 0.0013902 0.98689 0.99167 2.9982e-006 1.1993e-005 0.16326 0.91471 0.90798 0.0013992 0.9875 0.47719 0.001885 0.42485 2.0973 2.0965 16.0145 144.9254 0.0001767 -85.6348 0.69595
7.8 0.98813 5.4704e-005 3.8183 0.011931 0.0001015 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5237 0.54961 0.16815 0.019623 15.4567 0.12175 0.00015824 0.76841 0.0091958 0.010183 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.16327 0.91493 0.90807 0.0013991 0.98756 0.47737 0.0018849 0.42486 2.0979 2.0971 16.0144 144.9255 0.00017657 -85.635 0.69695
7.801 0.98813 5.4704e-005 3.8183 0.011931 0.00010152 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5238 0.54965 0.16816 0.019624 15.4595 0.12176 0.00015825 0.7684 0.0091962 0.010183 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.16327 0.91514 0.90815 0.0013991 0.98762 0.47755 0.0018849 0.42488 2.0984 2.0977 16.0144 144.9255 0.00017643 -85.6352 0.69795
7.802 0.98813 5.4704e-005 3.8183 0.011931 0.00010153 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5238 0.5497 0.16818 0.019625 15.4624 0.12176 0.00015826 0.7684 0.0091966 0.010184 0.0013901 0.98689 0.99167 2.9979e-006 1.1992e-005 0.16327 0.91536 0.90824 0.0013991 0.98769 0.47773 0.0018849 0.42489 2.099 2.0982 16.0144 144.9255 0.0001763 -85.6354 0.69895
7.803 0.98813 5.4704e-005 3.8183 0.011931 0.00010154 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5239 0.54974 0.16819 0.019626 15.4653 0.12177 0.00015827 0.76839 0.009197 0.010184 0.00139 0.9869 0.99167 2.9978e-006 1.1991e-005 0.16327 0.91557 0.90833 0.0013991 0.98775 0.47792 0.0018848 0.4249 2.0996 2.0988 16.0144 144.9255 0.00017617 -85.6356 0.69995
7.804 0.98813 5.4704e-005 3.8183 0.011931 0.00010156 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.524 0.54979 0.1682 0.019627 15.4682 0.12178 0.00015828 0.76838 0.0091974 0.010185 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.16328 0.91578 0.90841 0.001399 0.98781 0.4781 0.0018848 0.42492 2.1001 2.0993 16.0143 144.9255 0.00017603 -85.6359 0.70095
7.805 0.98813 5.4704e-005 3.8183 0.011931 0.00010157 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5241 0.54984 0.16822 0.019628 15.4711 0.12178 0.00015829 0.76838 0.0091978 0.010185 0.0013899 0.9869 0.99167 2.9976e-006 1.199e-005 0.16328 0.91599 0.9085 0.001399 0.98787 0.47828 0.0018848 0.42493 2.1007 2.0999 16.0143 144.9256 0.0001759 -85.6361 0.70195
7.806 0.98813 5.4704e-005 3.8183 0.011931 0.00010158 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5242 0.54988 0.16823 0.019629 15.4739 0.12179 0.0001583 0.76837 0.0091982 0.010185 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.16328 0.9162 0.90859 0.001399 0.98793 0.47846 0.0018847 0.42495 2.1012 2.1005 16.0143 144.9256 0.00017577 -85.6363 0.70295
7.807 0.98813 5.4704e-005 3.8183 0.011931 0.00010159 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5243 0.54993 0.16825 0.019631 15.4768 0.1218 0.00015831 0.76836 0.0091986 0.010186 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.16329 0.91641 0.90867 0.001399 0.98799 0.47864 0.0018847 0.42496 2.1018 2.101 16.0143 144.9256 0.00017564 -85.6365 0.70395
7.808 0.98813 5.4703e-005 3.8183 0.011931 0.00010161 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5244 0.54997 0.16826 0.019632 15.4797 0.1218 0.00015832 0.76836 0.009199 0.010186 0.0013898 0.9869 0.99168 2.9972e-006 1.1989e-005 0.16329 0.91662 0.90876 0.0013989 0.98805 0.47882 0.0018847 0.42498 2.1023 2.1016 16.0142 144.9256 0.0001755 -85.6367 0.70495
7.809 0.98813 5.4703e-005 3.8183 0.011931 0.00010162 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5245 0.55002 0.16827 0.019633 15.4826 0.12181 0.00015833 0.76835 0.0091994 0.010187 0.0013898 0.9869 0.99168 2.9971e-006 1.1988e-005 0.16329 0.91683 0.90884 0.0013989 0.98811 0.47901 0.0018846 0.42499 2.1029 2.1021 16.0142 144.9256 0.00017537 -85.6369 0.70595
7.81 0.98813 5.4703e-005 3.8183 0.011931 0.00010163 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5245 0.55006 0.16829 0.019634 15.4854 0.12182 0.00015834 0.76834 0.0091998 0.010187 0.0013897 0.9869 0.99168 2.9971e-006 1.1988e-005 0.1633 0.91704 0.90893 0.0013989 0.98817 0.47919 0.0018846 0.425 2.1034 2.1027 16.0142 144.9257 0.00017524 -85.6371 0.70695
7.811 0.98813 5.4703e-005 3.8183 0.011931 0.00010165 0.0011711 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5246 0.55011 0.1683 0.019635 15.4883 0.12182 0.00015835 0.76833 0.0092002 0.010188 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.1633 0.91725 0.90901 0.0013989 0.98823 0.47937 0.0018846 0.42502 2.104 2.1032 16.0142 144.9257 0.00017511 -85.6373 0.70795
7.812 0.98813 5.4703e-005 3.8183 0.011931 0.00010166 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5247 0.55015 0.16831 0.019636 15.4912 0.12183 0.00015836 0.76833 0.0092006 0.010188 0.0013897 0.9869 0.99168 2.9968e-006 1.1987e-005 0.1633 0.91746 0.9091 0.0013989 0.98829 0.47955 0.0018845 0.42503 2.1045 2.1038 16.0141 144.9257 0.00017498 -85.6375 0.70895
7.813 0.98813 5.4703e-005 3.8183 0.011931 0.00010167 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5248 0.5502 0.16833 0.019637 15.4941 0.12184 0.00015837 0.76832 0.009201 0.010188 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.16331 0.91766 0.90918 0.0013988 0.98834 0.47973 0.0018845 0.42505 2.1051 2.1043 16.0141 144.9257 0.00017485 -85.6377 0.70995
7.814 0.98813 5.4703e-005 3.8183 0.011931 0.00010168 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5249 0.55024 0.16834 0.019639 15.497 0.12184 0.00015838 0.76831 0.0092014 0.010189 0.0013896 0.9869 0.99168 2.9966e-006 1.1986e-005 0.16331 0.91787 0.90926 0.0013988 0.9884 0.47991 0.0018845 0.42506 2.1056 2.1049 16.0141 144.9257 0.00017472 -85.6378 0.71095
7.815 0.98813 5.4703e-005 3.8183 0.011931 0.0001017 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.525 0.55029 0.16836 0.01964 15.4998 0.12185 0.00015839 0.76831 0.0092018 0.010189 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.16331 0.91807 0.90935 0.0013988 0.98846 0.48009 0.0018844 0.42508 2.1062 2.1054 16.0141 144.9258 0.0001746 -85.638 0.71195
7.816 0.98813 5.4703e-005 3.8183 0.011931 0.00010171 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5251 0.55033 0.16837 0.019641 15.5027 0.12186 0.0001584 0.7683 0.0092022 0.01019 0.0013895 0.9869 0.99168 2.9964e-006 1.1986e-005 0.16332 0.91828 0.90943 0.0013988 0.98851 0.48028 0.0018844 0.42509 2.1067 2.106 16.014 144.9258 0.00017447 -85.6382 0.71295
7.817 0.98813 5.4703e-005 3.8183 0.011931 0.00010172 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5252 0.55038 0.16838 0.019642 15.5056 0.12186 0.00015841 0.76829 0.0092026 0.01019 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.16332 0.91848 0.90951 0.0013987 0.98857 0.48046 0.0018844 0.4251 2.1073 2.1065 16.014 144.9258 0.00017434 -85.6384 0.71395
7.818 0.98813 5.4703e-005 3.8183 0.011931 0.00010174 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5252 0.55042 0.1684 0.019643 15.5085 0.12187 0.00015842 0.76829 0.009203 0.010191 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.16332 0.91869 0.90959 0.0013987 0.98863 0.48064 0.0018843 0.42512 2.1078 2.1071 16.014 144.9258 0.00017421 -85.6386 0.71495
7.819 0.98813 5.4703e-005 3.8183 0.011931 0.00010175 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5253 0.55047 0.16841 0.019644 15.5114 0.12188 0.00015843 0.76828 0.0092034 0.010191 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.16332 0.91889 0.90967 0.0013987 0.98868 0.48082 0.0018843 0.42513 2.1084 2.1076 16.014 144.9258 0.00017409 -85.6388 0.71595
7.82 0.98813 5.4702e-005 3.8183 0.011931 0.00010176 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5254 0.55051 0.16842 0.019645 15.5142 0.12188 0.00015844 0.76827 0.0092039 0.010191 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.16333 0.91909 0.90976 0.0013987 0.98874 0.481 0.0018843 0.42515 2.1089 2.1082 16.0139 144.9259 0.00017396 -85.639 0.71695
7.821 0.98813 5.4702e-005 3.8183 0.011931 0.00010177 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5255 0.55056 0.16844 0.019647 15.5171 0.12189 0.00015845 0.76827 0.0092043 0.010192 0.0013892 0.98691 0.99168 2.9959e-006 1.1984e-005 0.16333 0.91929 0.90984 0.0013986 0.98879 0.48118 0.0018843 0.42516 2.1094 2.1087 16.0139 144.9259 0.00017384 -85.6392 0.71795
7.822 0.98813 5.4702e-005 3.8183 0.011931 0.00010179 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5256 0.5506 0.16845 0.019648 15.52 0.1219 0.00015846 0.76826 0.0092047 0.010192 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.16333 0.91949 0.90992 0.0013986 0.98885 0.48136 0.0018842 0.42518 2.11 2.1092 16.0139 144.9259 0.00017371 -85.6393 0.71895
7.823 0.98813 5.4702e-005 3.8183 0.011931 0.0001018 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5257 0.55065 0.16847 0.019649 15.5229 0.12191 0.00015847 0.76825 0.0092051 0.010193 0.0013892 0.98691 0.99168 2.9957e-006 1.1983e-005 0.16334 0.91969 0.91 0.0013986 0.9889 0.48154 0.0018842 0.42519 2.1105 2.1098 16.0138 144.9259 0.00017359 -85.6395 0.71995
7.824 0.98813 5.4702e-005 3.8183 0.011931 0.00010181 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5258 0.55069 0.16848 0.01965 15.5258 0.12191 0.00015848 0.76825 0.0092055 0.010193 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.16334 0.91989 0.91008 0.0013986 0.98895 0.48172 0.0018842 0.4252 2.111 2.1103 16.0138 144.9259 0.00017346 -85.6397 0.72095
7.825 0.98813 5.4702e-005 3.8183 0.011931 0.00010183 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5258 0.55074 0.16849 0.019651 15.5287 0.12192 0.00015849 0.76824 0.0092059 0.010194 0.0013891 0.98691 0.99168 2.9955e-006 1.1982e-005 0.16334 0.92009 0.91016 0.0013986 0.98901 0.4819 0.0018841 0.42522 2.1116 2.1108 16.0138 144.926 0.00017334 -85.6399 0.72195
7.826 0.98813 5.4702e-005 3.8183 0.011931 0.00010184 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5259 0.55078 0.16851 0.019652 15.5315 0.12193 0.0001585 0.76823 0.0092063 0.010194 0.001389 0.98691 0.99168 2.9954e-006 1.1982e-005 0.16335 0.92029 0.91024 0.0013985 0.98906 0.48208 0.0018841 0.42523 2.1121 2.1114 16.0138 144.926 0.00017322 -85.64 0.72295
7.827 0.98813 5.4702e-005 3.8183 0.011931 0.00010185 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.526 0.55083 0.16852 0.019653 15.5344 0.12193 0.00015851 0.76823 0.0092067 0.010194 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.16335 0.92049 0.91032 0.0013985 0.98911 0.48226 0.0018841 0.42525 2.1126 2.1119 16.0137 144.926 0.00017309 -85.6402 0.72395
7.828 0.98813 5.4702e-005 3.8183 0.011931 0.00010186 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5261 0.55087 0.16853 0.019654 15.5373 0.12194 0.00015852 0.76822 0.0092071 0.010195 0.0013889 0.98691 0.99168 2.9953e-006 1.1981e-005 0.16335 0.92068 0.9104 0.0013985 0.98917 0.48244 0.0018841 0.42526 2.1132 2.1124 16.0137 144.926 0.00017297 -85.6404 0.72495
7.829 0.98813 5.4702e-005 3.8183 0.011931 0.00010188 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5262 0.55092 0.16855 0.019656 15.5402 0.12195 0.00015853 0.76821 0.0092075 0.010195 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.16336 0.92088 0.91048 0.0013985 0.98922 0.48262 0.001884 0.42527 2.1137 2.113 16.0137 144.926 0.00017285 -85.6406 0.72595
7.83 0.98813 5.4702e-005 3.8183 0.011931 0.00010189 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5263 0.55096 0.16856 0.019657 15.5431 0.12195 0.00015854 0.76821 0.0092079 0.010196 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.16336 0.92108 0.91056 0.0013985 0.98927 0.4828 0.001884 0.42529 2.1142 2.1135 16.0137 144.9261 0.00017273 -85.6407 0.72695
7.831 0.98813 5.4702e-005 3.8183 0.011931 0.0001019 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5264 0.55101 0.16857 0.019658 15.546 0.12196 0.00015855 0.7682 0.0092083 0.010196 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.16336 0.92127 0.91063 0.0013984 0.98932 0.48298 0.001884 0.4253 2.1148 2.114 16.0136 144.9261 0.00017261 -85.6409 0.72795
7.832 0.98813 5.4701e-005 3.8183 0.011931 0.00010192 0.0011712 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5265 0.55105 0.16859 0.019659 15.5488 0.12197 0.00015856 0.76819 0.0092087 0.010197 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.16337 0.92147 0.91071 0.0013984 0.98937 0.48316 0.001884 0.42532 2.1153 2.1146 16.0136 144.9261 0.00017249 -85.6411 0.72895
7.833 0.98813 5.4701e-005 3.8183 0.011931 0.00010193 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5265 0.5511 0.1686 0.01966 15.5517 0.12197 0.00015857 0.76819 0.0092091 0.010197 0.0013888 0.98691 0.99168 2.9948e-006 1.1979e-005 0.16337 0.92166 0.91079 0.0013984 0.98942 0.48334 0.0018839 0.42533 2.1158 2.1151 16.0136 144.9261 0.00017237 -85.6412 0.72995
7.834 0.98813 5.4701e-005 3.8183 0.011931 0.00010194 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5266 0.55114 0.16862 0.019661 15.5546 0.12198 0.00015858 0.76818 0.0092095 0.010197 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.16337 0.92185 0.91087 0.0013984 0.98947 0.48352 0.0018839 0.42534 2.1163 2.1156 16.0136 144.9261 0.00017225 -85.6414 0.73095
7.835 0.98813 5.4701e-005 3.8183 0.011931 0.00010195 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5267 0.55119 0.16863 0.019662 15.5575 0.12199 0.00015859 0.76817 0.0092099 0.010198 0.0013887 0.98691 0.99168 2.9947e-006 1.1978e-005 0.16337 0.92205 0.91094 0.0013983 0.98952 0.4837 0.0018839 0.42536 2.1169 2.1161 16.0135 144.9262 0.00017213 -85.6416 0.73195
7.836 0.98813 5.4701e-005 3.8183 0.011931 0.00010197 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5268 0.55123 0.16864 0.019664 15.5604 0.12199 0.00015861 0.76817 0.0092103 0.010198 0.0013886 0.98691 0.99168 2.9946e-006 1.1978e-005 0.16338 0.92224 0.91102 0.0013983 0.98957 0.48388 0.0018838 0.42537 2.1174 2.1167 16.0135 144.9262 0.00017201 -85.6417 0.73295
7.837 0.98813 5.4701e-005 3.8183 0.011931 0.00010198 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5269 0.55128 0.16866 0.019665 15.5633 0.122 0.00015862 0.76816 0.0092107 0.010199 0.0013886 0.98691 0.99169 2.9945e-006 1.1978e-005 0.16338 0.92243 0.9111 0.0013983 0.98962 0.48406 0.0018838 0.42539 2.1179 2.1172 16.0135 144.9262 0.00017189 -85.6419 0.73395
7.838 0.98813 5.4701e-005 3.8183 0.011931 0.00010199 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.527 0.55132 0.16867 0.019666 15.5662 0.12201 0.00015863 0.76815 0.0092111 0.010199 0.0013886 0.98691 0.99169 2.9944e-006 1.1977e-005 0.16338 0.92262 0.91117 0.0013983 0.98967 0.48424 0.0018838 0.4254 2.1184 2.1177 16.0135 144.9262 0.00017177 -85.6421 0.73495
7.839 0.98813 5.4701e-005 3.8183 0.011931 0.00010201 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5271 0.55137 0.16868 0.019667 15.5691 0.12201 0.00015864 0.76814 0.0092115 0.0102 0.0013885 0.98691 0.99169 2.9943e-006 1.1977e-005 0.16339 0.92281 0.91125 0.0013983 0.98972 0.48442 0.0018838 0.42542 2.1189 2.1182 16.0134 144.9263 0.00017165 -85.6422 0.73595
7.84 0.98813 5.4701e-005 3.8183 0.011931 0.00010202 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5272 0.55141 0.1687 0.019668 15.5719 0.12202 0.00015865 0.76814 0.0092119 0.0102 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.16339 0.923 0.91133 0.0013982 0.98977 0.4846 0.0018837 0.42543 2.1195 2.1187 16.0134 144.9263 0.00017154 -85.6424 0.73695
7.841 0.98813 5.4701e-005 3.8183 0.011931 0.00010203 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5272 0.55146 0.16871 0.019669 15.5748 0.12203 0.00015866 0.76813 0.0092123 0.0102 0.0013885 0.98692 0.99169 2.9941e-006 1.1976e-005 0.16339 0.92319 0.9114 0.0013982 0.98982 0.48478 0.0018837 0.42544 2.12 2.1193 16.0134 144.9263 0.00017142 -85.6425 0.73795
7.842 0.98813 5.4701e-005 3.8183 0.011931 0.00010204 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5273 0.5515 0.16873 0.01967 15.5777 0.12203 0.00015867 0.76812 0.0092127 0.010201 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.1634 0.92338 0.91148 0.0013982 0.98987 0.48496 0.0018837 0.42546 2.1205 2.1198 16.0133 144.9263 0.0001713 -85.6427 0.73895
7.843 0.98813 5.4701e-005 3.8183 0.011931 0.00010206 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5274 0.55155 0.16874 0.019671 15.5806 0.12204 0.00015868 0.76812 0.0092131 0.010201 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.1634 0.92357 0.91155 0.0013982 0.98991 0.48514 0.0018837 0.42547 2.121 2.1203 16.0133 144.9263 0.00017119 -85.6429 0.73995
7.844 0.98813 5.4701e-005 3.8183 0.011931 0.00010207 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5275 0.55159 0.16875 0.019673 15.5835 0.12205 0.00015869 0.76811 0.0092135 0.010202 0.0013883 0.98692 0.99169 2.9939e-006 1.1975e-005 0.1634 0.92375 0.91163 0.0013982 0.98996 0.48532 0.0018836 0.42549 2.1215 2.1208 16.0133 144.9264 0.00017107 -85.643 0.74095
7.845 0.98813 5.47e-005 3.8183 0.011931 0.00010208 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5276 0.55164 0.16877 0.019674 15.5864 0.12205 0.0001587 0.7681 0.0092139 0.010202 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.16341 0.92394 0.9117 0.0013982 0.99001 0.4855 0.0018836 0.4255 2.122 2.1213 16.0133 144.9264 0.00017096 -85.6432 0.74195
7.846 0.98813 5.47e-005 3.8183 0.011931 0.0001021 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5277 0.55168 0.16878 0.019675 15.5893 0.12206 0.00015871 0.7681 0.0092143 0.010203 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.16341 0.92413 0.91178 0.0013981 0.99005 0.48568 0.0018836 0.42551 2.1225 2.1218 16.0132 144.9264 0.00017084 -85.6433 0.74295
7.847 0.98813 5.47e-005 3.8183 0.011931 0.00010211 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5278 0.55173 0.16879 0.019676 15.5922 0.12207 0.00015872 0.76809 0.0092147 0.010203 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16341 0.92431 0.91185 0.0013981 0.9901 0.48586 0.0018836 0.42553 2.123 2.1223 16.0132 144.9264 0.00017073 -85.6435 0.74395
7.848 0.98813 5.47e-005 3.8183 0.011931 0.00010212 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5278 0.55177 0.16881 0.019677 15.5951 0.12208 0.00015873 0.76808 0.0092151 0.010203 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16342 0.9245 0.91192 0.0013981 0.99015 0.48604 0.0018835 0.42554 2.1235 2.1228 16.0132 144.9264 0.00017062 -85.6436 0.74495
7.849 0.98813 5.47e-005 3.8183 0.011931 0.00010213 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5279 0.55182 0.16882 0.019678 15.598 0.12208 0.00015874 0.76808 0.0092155 0.010204 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.16342 0.92468 0.912 0.0013981 0.99019 0.48622 0.0018835 0.42556 2.1241 2.1234 16.0132 144.9265 0.0001705 -85.6438 0.74595
7.85 0.98813 5.47e-005 3.8183 0.011931 0.00010215 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.528 0.55186 0.16884 0.019679 15.6008 0.12209 0.00015875 0.76807 0.0092159 0.010204 0.0013881 0.98692 0.99169 2.9934e-006 1.1974e-005 0.16342 0.92487 0.91207 0.0013981 0.99024 0.4864 0.0018835 0.42557 2.1246 2.1239 16.0131 144.9265 0.00017039 -85.6439 0.74695
7.851 0.98813 5.47e-005 3.8183 0.011931 0.00010216 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5281 0.55191 0.16885 0.019681 15.6037 0.1221 0.00015876 0.76806 0.0092163 0.010205 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.16342 0.92505 0.91214 0.001398 0.99028 0.48657 0.0018835 0.42558 2.1251 2.1244 16.0131 144.9265 0.00017028 -85.6441 0.74795
7.852 0.98813 5.47e-005 3.8183 0.01193 0.00010217 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5282 0.55195 0.16886 0.019682 15.6066 0.1221 0.00015877 0.76806 0.0092168 0.010205 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.16343 0.92523 0.91222 0.001398 0.99033 0.48675 0.0018834 0.4256 2.1256 2.1249 16.0131 144.9265 0.00017016 -85.6442 0.74895
7.853 0.98813 5.47e-005 3.8183 0.01193 0.00010218 0.0011713 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5283 0.552 0.16888 0.019683 15.6095 0.12211 0.00015878 0.76805 0.0092172 0.010206 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.16343 0.92541 0.91229 0.001398 0.99037 0.48693 0.0018834 0.42561 2.1261 2.1254 16.013 144.9265 0.00017005 -85.6444 0.74995
7.854 0.98813 5.47e-005 3.8183 0.01193 0.0001022 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5284 0.55204 0.16889 0.019684 15.6124 0.12212 0.00015879 0.76804 0.0092176 0.010206 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.16343 0.9256 0.91236 0.001398 0.99042 0.48711 0.0018834 0.42563 2.1266 2.1259 16.013 144.9266 0.00016994 -85.6445 0.75095
7.855 0.98813 5.47e-005 3.8183 0.01193 0.00010221 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5285 0.55209 0.1689 0.019685 15.6153 0.12212 0.0001588 0.76804 0.009218 0.010206 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.16344 0.92578 0.91243 0.001398 0.99046 0.48729 0.0018834 0.42564 2.1271 2.1264 16.013 144.9266 0.00016983 -85.6446 0.75195
7.856 0.98813 5.47e-005 3.8183 0.01193 0.00010222 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5285 0.55213 0.16892 0.019686 15.6182 0.12213 0.00015881 0.76803 0.0092184 0.010207 0.0013879 0.98692 0.99169 2.9929e-006 1.1972e-005 0.16344 0.92596 0.9125 0.001398 0.9905 0.48747 0.0018834 0.42565 2.1276 2.1269 16.013 144.9266 0.00016972 -85.6448 0.75295
7.857 0.98813 5.4699e-005 3.8183 0.01193 0.00010224 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5286 0.55218 0.16893 0.019687 15.6211 0.12214 0.00015882 0.76802 0.0092188 0.010207 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.16344 0.92614 0.91258 0.0013979 0.99055 0.48765 0.0018833 0.42567 2.1281 2.1274 16.0129 144.9266 0.00016961 -85.6449 0.75395
7.858 0.98813 5.4699e-005 3.8183 0.01193 0.00010225 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5287 0.55222 0.16895 0.019688 15.624 0.12214 0.00015883 0.76802 0.0092192 0.010208 0.0013878 0.98692 0.99169 2.9928e-006 1.1971e-005 0.16345 0.92632 0.91265 0.0013979 0.99059 0.48783 0.0018833 0.42568 2.1286 2.1279 16.0129 144.9266 0.0001695 -85.6451 0.75495
7.859 0.98813 5.4699e-005 3.8183 0.01193 0.00010226 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5288 0.55227 0.16896 0.01969 15.6269 0.12215 0.00015884 0.76801 0.0092196 0.010208 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.16345 0.9265 0.91272 0.0013979 0.99063 0.488 0.0018833 0.4257 2.1291 2.1284 16.0129 144.9267 0.00016939 -85.6452 0.75595
7.86 0.98813 5.4699e-005 3.8183 0.01193 0.00010227 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5289 0.55231 0.16897 0.019691 15.6298 0.12216 0.00015885 0.768 0.00922 0.010209 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.16345 0.92667 0.91279 0.0013979 0.99068 0.48818 0.0018833 0.42571 2.1296 2.1289 16.0129 144.9267 0.00016928 -85.6453 0.75695
7.861 0.98813 5.4699e-005 3.8183 0.01193 0.00010229 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.529 0.55236 0.16899 0.019692 15.6327 0.12216 0.00015886 0.768 0.0092204 0.010209 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.16346 0.92685 0.91286 0.0013979 0.99072 0.48836 0.0018832 0.42572 2.13 2.1294 16.0128 144.9267 0.00016917 -85.6455 0.75795
7.862 0.98813 5.4699e-005 3.8183 0.01193 0.0001023 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5291 0.5524 0.169 0.019693 15.6356 0.12217 0.00015887 0.76799 0.0092208 0.010209 0.0013877 0.98693 0.99169 2.9925e-006 1.197e-005 0.16346 0.92703 0.91293 0.0013979 0.99076 0.48854 0.0018832 0.42574 2.1305 2.1299 16.0128 144.9267 0.00016906 -85.6456 0.75895
7.863 0.98813 5.4699e-005 3.8183 0.01193 0.00010231 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5291 0.55245 0.16901 0.019694 15.6385 0.12218 0.00015888 0.76798 0.0092212 0.01021 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.16346 0.92721 0.913 0.0013978 0.9908 0.48872 0.0018832 0.42575 2.131 2.1304 16.0128 144.9267 0.00016895 -85.6458 0.75995
7.864 0.98813 5.4699e-005 3.8183 0.01193 0.00010233 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5292 0.55249 0.16903 0.019695 15.6414 0.12218 0.00015889 0.76798 0.0092216 0.01021 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.16346 0.92738 0.91307 0.0013978 0.99084 0.48889 0.0018832 0.42577 2.1315 2.1308 16.0127 144.9268 0.00016885 -85.6459 0.76095
7.865 0.98813 5.4699e-005 3.8183 0.01193 0.00010234 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5293 0.55254 0.16904 0.019696 15.6443 0.12219 0.0001589 0.76797 0.009222 0.010211 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.16347 0.92756 0.91314 0.0013978 0.99088 0.48907 0.0018832 0.42578 2.132 2.1313 16.0127 144.9268 0.00016874 -85.646 0.76195
7.866 0.98813 5.4699e-005 3.8183 0.01193 0.00010235 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5294 0.55258 0.16905 0.019698 15.6472 0.1222 0.00015891 0.76796 0.0092224 0.010211 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.16347 0.92773 0.91321 0.0013978 0.99092 0.48925 0.0018831 0.42579 2.1325 2.1318 16.0127 144.9268 0.00016863 -85.6462 0.76295
7.867 0.98813 5.4699e-005 3.8183 0.01193 0.00010236 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5295 0.55263 0.16907 0.019699 15.6501 0.1222 0.00015892 0.76796 0.0092228 0.010212 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.16347 0.92791 0.91328 0.0013978 0.99097 0.48943 0.0018831 0.42581 2.133 2.1323 16.0127 144.9268 0.00016853 -85.6463 0.76395
7.868 0.98813 5.4699e-005 3.8183 0.01193 0.00010238 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5296 0.55267 0.16908 0.0197 15.653 0.12221 0.00015893 0.76795 0.0092232 0.010212 0.0013875 0.98693 0.99169 2.9921e-006 1.1968e-005 0.16348 0.92808 0.91335 0.0013978 0.99101 0.48961 0.0018831 0.42582 2.1335 2.1328 16.0126 144.9268 0.00016842 -85.6464 0.76495
7.869 0.98813 5.4698e-005 3.8183 0.01193 0.00010239 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5297 0.55272 0.1691 0.019701 15.6559 0.12222 0.00015894 0.76794 0.0092236 0.010212 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16348 0.92825 0.91341 0.0013977 0.99105 0.48978 0.0018831 0.42584 2.134 2.1333 16.0126 144.9269 0.00016832 -85.6465 0.76595
7.87 0.98813 5.4698e-005 3.8183 0.01193 0.0001024 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5298 0.55276 0.16911 0.019702 15.6588 0.12222 0.00015895 0.76793 0.009224 0.010213 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.16348 0.92843 0.91348 0.0013977 0.99109 0.48996 0.0018831 0.42585 2.1344 2.1338 16.0126 144.9269 0.00016821 -85.6467 0.76695
7.871 0.98813 5.4698e-005 3.8183 0.01193 0.00010242 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5298 0.55281 0.16912 0.019703 15.6617 0.12223 0.00015896 0.76793 0.0092244 0.010213 0.0013875 0.98693 0.99169 2.9919e-006 1.1967e-005 0.16349 0.9286 0.91355 0.0013977 0.99113 0.49014 0.001883 0.42586 2.1349 2.1343 16.0125 144.9269 0.0001681 -85.6468 0.76795
7.872 0.98813 5.4698e-005 3.8183 0.01193 0.00010243 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5299 0.55285 0.16914 0.019704 15.6646 0.12224 0.00015897 0.76792 0.0092248 0.010214 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.16349 0.92877 0.91362 0.0013977 0.99116 0.49032 0.001883 0.42588 2.1354 2.1347 16.0125 144.9269 0.000168 -85.6469 0.76895
7.873 0.98813 5.4698e-005 3.8183 0.01193 0.00010244 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.53 0.5529 0.16915 0.019705 15.6675 0.12224 0.00015898 0.76791 0.0092252 0.010214 0.0013874 0.98693 0.9917 2.9917e-006 1.1967e-005 0.16349 0.92894 0.91369 0.0013977 0.9912 0.4905 0.001883 0.42589 2.1359 2.1352 16.0125 144.9269 0.0001679 -85.6471 0.76995
7.874 0.98813 5.4698e-005 3.8183 0.01193 0.00010245 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5301 0.55294 0.16916 0.019707 15.6703 0.12225 0.00015899 0.76791 0.0092256 0.010215 0.0013874 0.98693 0.9917 2.9917e-006 1.1967e-005 0.1635 0.92911 0.91375 0.0013977 0.99124 0.49067 0.001883 0.42591 2.1364 2.1357 16.0125 144.927 0.00016779 -85.6472 0.77095
7.875 0.98813 5.4698e-005 3.8183 0.01193 0.00010247 0.0011714 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5302 0.55299 0.16918 0.019708 15.6733 0.12226 0.000159 0.7679 0.009226 0.010215 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.1635 0.92928 0.91382 0.0013976 0.99128 0.49085 0.001883 0.42592 2.1369 2.1362 16.0124 144.927 0.00016769 -85.6473 0.77195
7.876 0.98813 5.4698e-005 3.8183 0.01193 0.00010248 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5303 0.55303 0.16919 0.019709 15.6762 0.12226 0.00015901 0.76789 0.0092264 0.010215 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.1635 0.92945 0.91389 0.0013976 0.99132 0.49103 0.0018829 0.42593 2.1373 2.1367 16.0124 144.927 0.00016759 -85.6474 0.77295
7.877 0.98813 5.4698e-005 3.8183 0.01193 0.00010249 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5304 0.55308 0.16921 0.01971 15.6791 0.12227 0.00015902 0.76789 0.0092268 0.010216 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.1635 0.92962 0.91395 0.0013976 0.99136 0.4912 0.0018829 0.42595 2.1378 2.1372 16.0124 144.927 0.00016748 -85.6475 0.77395
7.878 0.98813 5.4698e-005 3.8183 0.01193 0.00010251 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5305 0.55312 0.16922 0.019711 15.682 0.12228 0.00015903 0.76788 0.0092272 0.010216 0.0013872 0.98693 0.9917 2.9914e-006 1.1966e-005 0.16351 0.92979 0.91402 0.0013976 0.9914 0.49138 0.0018829 0.42596 2.1383 2.1376 16.0123 144.9271 0.00016738 -85.6477 0.77495
7.879 0.98813 5.4698e-005 3.8183 0.01193 0.00010252 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5305 0.55317 0.16923 0.019712 15.6849 0.12229 0.00015904 0.76787 0.0092276 0.010217 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16351 0.92996 0.91408 0.0013976 0.99143 0.49156 0.0018829 0.42598 2.1388 2.1381 16.0123 144.9271 0.00016728 -85.6478 0.77595
7.88 0.98813 5.4698e-005 3.8183 0.01193 0.00010253 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5306 0.55321 0.16925 0.019713 15.6878 0.12229 0.00015905 0.76787 0.009228 0.010217 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16351 0.93012 0.91415 0.0013976 0.99147 0.49174 0.0018829 0.42599 2.1392 2.1386 16.0123 144.9271 0.00016718 -85.6479 0.77695
7.881 0.98813 5.4698e-005 3.8183 0.01193 0.00010254 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5307 0.55326 0.16926 0.019714 15.6907 0.1223 0.00015906 0.76786 0.0092284 0.010218 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.16352 0.93029 0.91422 0.0013976 0.99151 0.49191 0.0018828 0.426 2.1397 2.1391 16.0123 144.9271 0.00016708 -85.648 0.77795
7.882 0.98813 5.4697e-005 3.8183 0.01193 0.00010256 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5308 0.5533 0.16927 0.019716 15.6936 0.12231 0.00015907 0.76785 0.0092288 0.010218 0.0013871 0.98693 0.9917 2.9912e-006 1.1965e-005 0.16352 0.93046 0.91428 0.0013975 0.99154 0.49209 0.0018828 0.42602 2.1402 2.1395 16.0122 144.9271 0.00016697 -85.6481 0.77895
7.883 0.98813 5.4697e-005 3.8183 0.01193 0.00010257 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5309 0.55335 0.16929 0.019717 15.6965 0.12231 0.00015909 0.76785 0.0092292 0.010218 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.16352 0.93062 0.91435 0.0013975 0.99158 0.49227 0.0018828 0.42603 2.1406 2.14 16.0122 144.9272 0.00016687 -85.6483 0.77995
7.884 0.98813 5.4697e-005 3.8183 0.01193 0.00010258 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.531 0.55339 0.1693 0.019718 15.6994 0.12232 0.0001591 0.76784 0.0092296 0.010219 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16353 0.93079 0.91441 0.0013975 0.99162 0.49244 0.0018828 0.42605 2.1411 2.1405 16.0122 144.9272 0.00016677 -85.6484 0.78095
7.885 0.98813 5.4697e-005 3.8183 0.01193 0.0001026 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5311 0.55344 0.16931 0.019719 15.7023 0.12233 0.00015911 0.76783 0.00923 0.010219 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16353 0.93095 0.91448 0.0013975 0.99165 0.49262 0.0018828 0.42606 2.1416 2.1409 16.0121 144.9272 0.00016667 -85.6485 0.78195
7.886 0.98813 5.4697e-005 3.8183 0.01193 0.00010261 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5311 0.55348 0.16933 0.01972 15.7052 0.12233 0.00015912 0.76783 0.0092304 0.01022 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.16353 0.93112 0.91454 0.0013975 0.99169 0.4928 0.0018827 0.42607 2.1421 2.1414 16.0121 144.9272 0.00016657 -85.6486 0.78295
7.887 0.98813 5.4697e-005 3.8183 0.01193 0.00010262 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5312 0.55353 0.16934 0.019721 15.7081 0.12234 0.00015913 0.76782 0.0092308 0.01022 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.16354 0.93128 0.9146 0.0013975 0.99173 0.49297 0.0018827 0.42609 2.1425 2.1419 16.0121 144.9272 0.00016648 -85.6487 0.78395
7.888 0.98813 5.4697e-005 3.8183 0.01193 0.00010263 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5313 0.55358 0.16936 0.019722 15.711 0.12235 0.00015914 0.76781 0.0092312 0.010221 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.16354 0.93145 0.91467 0.0013975 0.99176 0.49315 0.0018827 0.4261 2.143 2.1424 16.0121 144.9273 0.00016638 -85.6488 0.78495
7.889 0.98813 5.4697e-005 3.8183 0.01193 0.00010265 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5314 0.55362 0.16937 0.019724 15.7139 0.12235 0.00015915 0.76781 0.0092316 0.010221 0.001387 0.98693 0.9917 2.9907e-006 1.1963e-005 0.16354 0.93161 0.91473 0.0013974 0.9918 0.49333 0.0018827 0.42611 2.1435 2.1428 16.012 144.9273 0.00016628 -85.6489 0.78595
7.89 0.98813 5.4697e-005 3.8183 0.01193 0.00010266 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5315 0.55367 0.16938 0.019725 15.7168 0.12236 0.00015916 0.7678 0.009232 0.010221 0.0013869 0.98694 0.9917 2.9907e-006 1.1963e-005 0.16355 0.93177 0.9148 0.0013974 0.99183 0.4935 0.0018827 0.42613 2.1439 2.1433 16.012 144.9273 0.00016618 -85.6491 0.78695
7.891 0.98813 5.4697e-005 3.8183 0.01193 0.00010267 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5316 0.55371 0.1694 0.019726 15.7197 0.12237 0.00015917 0.76779 0.0092324 0.010222 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16355 0.93193 0.91486 0.0013974 0.99187 0.49368 0.0018827 0.42614 2.1444 2.1438 16.012 144.9273 0.00016608 -85.6492 0.78795
7.892 0.98813 5.4697e-005 3.8183 0.01193 0.00010269 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5317 0.55376 0.16941 0.019727 15.7226 0.12237 0.00015918 0.76779 0.0092328 0.010222 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16355 0.93209 0.91492 0.0013974 0.9919 0.49386 0.0018826 0.42616 2.1448 2.1442 16.0119 144.9273 0.00016598 -85.6493 0.78895
7.893 0.98813 5.4697e-005 3.8183 0.01193 0.0001027 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5318 0.5538 0.16942 0.019728 15.7255 0.12238 0.00015919 0.76778 0.0092332 0.010223 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16355 0.93225 0.91499 0.0013974 0.99193 0.49403 0.0018826 0.42617 2.1453 2.1447 16.0119 144.9274 0.00016589 -85.6494 0.78995
7.894 0.98813 5.4696e-005 3.8183 0.01193 0.00010271 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5318 0.55385 0.16944 0.019729 15.7284 0.12239 0.0001592 0.76777 0.0092336 0.010223 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16356 0.93241 0.91505 0.0013974 0.99197 0.49421 0.0018826 0.42618 2.1458 2.1451 16.0119 144.9274 0.00016579 -85.6495 0.79095
7.895 0.98813 5.4696e-005 3.8183 0.01193 0.00010272 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5319 0.55389 0.16945 0.01973 15.7313 0.12239 0.00015921 0.76777 0.009234 0.010224 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.16356 0.93257 0.91511 0.0013974 0.992 0.49439 0.0018826 0.4262 2.1462 2.1456 16.0119 144.9274 0.00016569 -85.6496 0.79195
7.896 0.98813 5.4696e-005 3.8183 0.01193 0.00010274 0.0011715 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.532 0.55394 0.16947 0.019731 15.7342 0.1224 0.00015922 0.76776 0.0092344 0.010224 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16356 0.93273 0.91517 0.0013974 0.99204 0.49456 0.0018826 0.42621 2.1467 2.1461 16.0118 144.9274 0.0001656 -85.6497 0.79295
7.897 0.98813 5.4696e-005 3.8183 0.01193 0.00010275 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5321 0.55398 0.16948 0.019733 15.7371 0.12241 0.00015923 0.76775 0.0092348 0.010224 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16357 0.93289 0.91523 0.0013973 0.99207 0.49474 0.0018826 0.42622 2.1471 2.1465 16.0118 144.9274 0.0001655 -85.6498 0.79395
7.898 0.98813 5.4696e-005 3.8183 0.01193 0.00010276 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5322 0.55403 0.16949 0.019734 15.74 0.12241 0.00015924 0.76775 0.0092352 0.010225 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16357 0.93305 0.9153 0.0013973 0.9921 0.49491 0.0018825 0.42624 2.1476 2.147 16.0118 144.9275 0.00016541 -85.6499 0.79495
7.899 0.98813 5.4696e-005 3.8183 0.01193 0.00010278 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5323 0.55407 0.16951 0.019735 15.743 0.12242 0.00015925 0.76774 0.0092356 0.010225 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16357 0.93321 0.91536 0.0013973 0.99214 0.49509 0.0018825 0.42625 2.1481 2.1474 16.0117 144.9275 0.00016531 -85.65 0.79595
7.9 0.98813 5.4696e-005 3.8183 0.01193 0.00010279 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5324 0.55412 0.16952 0.019736 15.7459 0.12243 0.00015926 0.76773 0.009236 0.010226 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.16358 0.93337 0.91542 0.0013973 0.99217 0.49527 0.0018825 0.42627 2.1485 2.1479 16.0117 144.9275 0.00016522 -85.6501 0.79695
7.901 0.98813 5.4696e-005 3.8183 0.01193 0.0001028 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5324 0.55416 0.16953 0.019737 15.7488 0.12243 0.00015927 0.76773 0.0092364 0.010226 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.16358 0.93352 0.91548 0.0013973 0.9922 0.49544 0.0018825 0.42628 2.149 2.1484 16.0117 144.9275 0.00016512 -85.6502 0.79795
7.902 0.98813 5.4696e-005 3.8183 0.01193 0.00010281 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5325 0.55421 0.16955 0.019738 15.7517 0.12244 0.00015928 0.76772 0.0092368 0.010226 0.0013867 0.98694 0.9917 2.99e-006 1.196e-005 0.16358 0.93368 0.91554 0.0013973 0.99223 0.49562 0.0018825 0.42629 2.1494 2.1488 16.0117 144.9275 0.00016503 -85.6503 0.79895
7.903 0.98813 5.4696e-005 3.8183 0.01193 0.00010283 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5326 0.55425 0.16956 0.019739 15.7546 0.12245 0.00015929 0.76771 0.0092372 0.010227 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.16359 0.93383 0.9156 0.0013973 0.99227 0.49579 0.0018825 0.42631 2.1499 2.1493 16.0116 144.9276 0.00016493 -85.6504 0.79995
7.904 0.98813 5.4696e-005 3.8183 0.01193 0.00010284 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5327 0.5543 0.16957 0.01974 15.7575 0.12245 0.0001593 0.76771 0.0092376 0.010227 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.16359 0.93399 0.91566 0.0013973 0.9923 0.49597 0.0018824 0.42632 2.1503 2.1497 16.0116 144.9276 0.00016484 -85.6505 0.80095
7.905 0.98813 5.4696e-005 3.8183 0.01193 0.00010285 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5328 0.55434 0.16959 0.019742 15.7604 0.12246 0.00015931 0.7677 0.009238 0.010228 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.16359 0.93415 0.91572 0.0013972 0.99233 0.49615 0.0018824 0.42634 2.1508 2.1502 16.0116 144.9276 0.00016475 -85.6506 0.80195
7.906 0.98813 5.4695e-005 3.8183 0.01193 0.00010286 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5329 0.55439 0.1696 0.019743 15.7633 0.12247 0.00015932 0.76769 0.0092384 0.010228 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.16359 0.9343 0.91578 0.0013972 0.99236 0.49632 0.0018824 0.42635 2.1512 2.1506 16.0115 144.9276 0.00016465 -85.6507 0.80295
7.907 0.98813 5.4695e-005 3.8183 0.01193 0.00010288 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.533 0.55443 0.16962 0.019744 15.7662 0.12247 0.00015933 0.76769 0.0092388 0.010229 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.1636 0.93445 0.91584 0.0013972 0.99239 0.4965 0.0018824 0.42636 2.1517 2.1511 16.0115 144.9276 0.00016456 -85.6508 0.80395
7.908 0.98813 5.4695e-005 3.8183 0.01193 0.00010289 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5331 0.55448 0.16963 0.019745 15.7691 0.12248 0.00015934 0.76768 0.0092392 0.010229 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.1636 0.93461 0.9159 0.0013972 0.99242 0.49667 0.0018824 0.42638 2.1521 2.1515 16.0115 144.9277 0.00016447 -85.6509 0.80495
7.909 0.98813 5.4695e-005 3.8183 0.011929 0.0001029 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5331 0.55452 0.16964 0.019746 15.7721 0.12249 0.00015935 0.76767 0.0092396 0.010229 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.1636 0.93476 0.91596 0.0013972 0.99245 0.49685 0.0018824 0.42639 2.1526 2.152 16.0114 144.9277 0.00016438 -85.651 0.80595
7.91 0.98813 5.4695e-005 3.8183 0.011929 0.00010292 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5332 0.55457 0.16966 0.019747 15.775 0.12249 0.00015936 0.76766 0.00924 0.01023 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16361 0.93491 0.91602 0.0013972 0.99248 0.49702 0.0018823 0.4264 2.153 2.1524 16.0114 144.9277 0.00016429 -85.6511 0.80695
7.911 0.98813 5.4695e-005 3.8183 0.011929 0.00010293 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5333 0.55461 0.16967 0.019748 15.7779 0.1225 0.00015937 0.76766 0.0092404 0.01023 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16361 0.93506 0.91608 0.0013972 0.99252 0.4972 0.0018823 0.42642 2.1535 2.1529 16.0114 144.9277 0.0001642 -85.6512 0.80795
7.912 0.98813 5.4695e-005 3.8183 0.011929 0.00010294 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5334 0.55466 0.16968 0.019749 15.7808 0.12251 0.00015938 0.76765 0.0092408 0.010231 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16361 0.93522 0.91614 0.0013972 0.99255 0.49737 0.0018823 0.42643 2.1539 2.1533 16.0114 144.9277 0.0001641 -85.6513 0.80895
7.913 0.98813 5.4695e-005 3.8183 0.011929 0.00010295 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5335 0.5547 0.1697 0.019751 15.7837 0.12251 0.00015939 0.76764 0.0092412 0.010231 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16362 0.93537 0.9162 0.0013971 0.99258 0.49755 0.0018823 0.42645 2.1544 2.1538 16.0113 144.9278 0.00016401 -85.6514 0.80995
7.914 0.98813 5.4695e-005 3.8183 0.011929 0.00010297 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5336 0.55475 0.16971 0.019752 15.7866 0.12252 0.0001594 0.76764 0.0092416 0.010232 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.16362 0.93552 0.91626 0.0013971 0.99261 0.49772 0.0018823 0.42646 2.1548 2.1542 16.0113 144.9278 0.00016392 -85.6515 0.81095
7.915 0.98813 5.4695e-005 3.8183 0.011929 0.00010298 0.0011716 0.23374 0.00065931 0.23439 0.2163 0 0.032257 0.0389 0 1.5337 0.55479 0.16973 0.019753 15.7895 0.12253 0.00015941 0.76763 0.009242 0.010232 0.0013864 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16362 0.93567 0.91631 0.0013971 0.99264 0.4979 0.0018823 0.42647 2.1552 2.1546 16.0113 144.9278 0.00016383 -85.6516 0.81195
7.916 0.98813 5.4695e-005 3.8183 0.011929 0.00010299 0.0011716 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5337 0.55484 0.16974 0.019754 15.7924 0.12253 0.00015942 0.76762 0.0092424 0.010232 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16363 0.93582 0.91637 0.0013971 0.99266 0.49807 0.0018823 0.42649 2.1557 2.1551 16.0112 144.9278 0.00016374 -85.6517 0.81295
7.917 0.98813 5.4695e-005 3.8183 0.011929 0.00010301 0.0011716 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5338 0.55488 0.16975 0.019755 15.7954 0.12254 0.00015943 0.76762 0.0092428 0.010233 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16363 0.93597 0.91643 0.0013971 0.99269 0.49825 0.0018822 0.4265 2.1561 2.1555 16.0112 144.9279 0.00016365 -85.6517 0.81395
7.918 0.98813 5.4694e-005 3.8183 0.011929 0.00010302 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5339 0.55493 0.16977 0.019756 15.7983 0.12255 0.00015944 0.76761 0.0092432 0.010233 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16363 0.93611 0.91649 0.0013971 0.99272 0.49842 0.0018822 0.42651 2.1566 2.156 16.0112 144.9279 0.00016357 -85.6518 0.81495
7.919 0.98813 5.4694e-005 3.8183 0.011929 0.00010303 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.534 0.55497 0.16978 0.019757 15.8012 0.12255 0.00015945 0.7676 0.0092436 0.010234 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16363 0.93626 0.91654 0.0013971 0.99275 0.4986 0.0018822 0.42653 2.157 2.1564 16.0111 144.9279 0.00016348 -85.6519 0.81595
7.92 0.98813 5.4694e-005 3.8183 0.011929 0.00010304 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5341 0.55502 0.16979 0.019758 15.8041 0.12256 0.00015946 0.7676 0.009244 0.010234 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.16364 0.93641 0.9166 0.0013971 0.99278 0.49877 0.0018822 0.42654 2.1574 2.1568 16.0111 144.9279 0.00016339 -85.652 0.81695
7.921 0.98813 5.4694e-005 3.8183 0.011929 0.00010306 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5342 0.55506 0.16981 0.01976 15.807 0.12257 0.00015947 0.76759 0.0092443 0.010235 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.16364 0.93656 0.91666 0.0013971 0.99281 0.49895 0.0018822 0.42655 2.1579 2.1573 16.0111 144.9279 0.0001633 -85.6521 0.81795
7.922 0.98813 5.4694e-005 3.8183 0.011929 0.00010307 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5343 0.55511 0.16982 0.019761 15.8099 0.12258 0.00015948 0.76758 0.0092447 0.010235 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16364 0.9367 0.91672 0.001397 0.99284 0.49912 0.0018822 0.42657 2.1583 2.1577 16.0111 144.928 0.00016321 -85.6522 0.81895
7.923 0.98813 5.4694e-005 3.8183 0.011929 0.00010308 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5344 0.55515 0.16983 0.019762 15.8129 0.12258 0.00015949 0.76758 0.0092451 0.010235 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16365 0.93685 0.91677 0.001397 0.99287 0.4993 0.0018822 0.42658 2.1587 2.1582 16.011 144.928 0.00016313 -85.6523 0.81995
7.924 0.98813 5.4694e-005 3.8183 0.011929 0.0001031 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5344 0.5552 0.16985 0.019763 15.8158 0.12259 0.0001595 0.76757 0.0092455 0.010236 0.0013862 0.98695 0.99171 2.9889e-006 1.1956e-005 0.16365 0.937 0.91683 0.001397 0.99289 0.49947 0.0018821 0.4266 2.1592 2.1586 16.011 144.928 0.00016304 -85.6524 0.82095
7.925 0.98813 5.4694e-005 3.8183 0.011929 0.00010311 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5345 0.55524 0.16986 0.019764 15.8187 0.1226 0.00015951 0.76756 0.0092459 0.010236 0.0013862 0.98695 0.99171 2.9889e-006 1.1955e-005 0.16365 0.93714 0.91688 0.001397 0.99292 0.49964 0.0018821 0.42661 2.1596 2.159 16.011 144.928 0.00016295 -85.6524 0.82195
7.926 0.98813 5.4694e-005 3.8183 0.011929 0.00010312 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5346 0.55529 0.16988 0.019765 15.8216 0.1226 0.00015952 0.76756 0.0092463 0.010237 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16366 0.93729 0.91694 0.001397 0.99295 0.49982 0.0018821 0.42662 2.16 2.1595 16.0109 144.928 0.00016286 -85.6525 0.82295
7.927 0.98813 5.4694e-005 3.8183 0.011929 0.00010313 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5347 0.55533 0.16989 0.019766 15.8245 0.12261 0.00015953 0.76755 0.0092467 0.010237 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16366 0.93743 0.917 0.001397 0.99298 0.49999 0.0018821 0.42664 2.1605 2.1599 16.0109 144.9281 0.00016278 -85.6526 0.82395
7.928 0.98813 5.4694e-005 3.8183 0.011929 0.00010315 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5348 0.55538 0.1699 0.019767 15.8274 0.12262 0.00015954 0.76754 0.0092471 0.010237 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16366 0.93758 0.91705 0.001397 0.993 0.50017 0.0018821 0.42665 2.1609 2.1603 16.0109 144.9281 0.00016269 -85.6527 0.82495
7.929 0.98813 5.4694e-005 3.8183 0.011929 0.00010316 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5349 0.55542 0.16992 0.019769 15.8304 0.12262 0.00015955 0.76754 0.0092475 0.010238 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16366 0.93772 0.91711 0.001397 0.99303 0.50034 0.0018821 0.42666 2.1613 2.1608 16.0108 144.9281 0.00016261 -85.6528 0.82595
7.93 0.98813 5.4694e-005 3.8183 0.011929 0.00010317 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.535 0.55547 0.16993 0.01977 15.8333 0.12263 0.00015956 0.76753 0.0092479 0.010238 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16367 0.93786 0.91716 0.001397 0.99306 0.50052 0.0018821 0.42668 2.1618 2.1612 16.0108 144.9281 0.00016252 -85.6529 0.82695
7.931 0.98813 5.4693e-005 3.8183 0.011929 0.00010319 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.535 0.55551 0.16994 0.019771 15.8362 0.12264 0.00015957 0.76752 0.0092483 0.010239 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16367 0.93801 0.91722 0.001397 0.99309 0.50069 0.0018821 0.42669 2.1622 2.1616 16.0108 144.9281 0.00016244 -85.6529 0.82795
7.932 0.98813 5.4693e-005 3.8183 0.011929 0.0001032 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5351 0.55556 0.16996 0.019772 15.8391 0.12264 0.00015958 0.76752 0.0092487 0.010239 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16367 0.93815 0.91727 0.0013969 0.99311 0.50086 0.001882 0.4267 2.1626 2.162 16.0108 144.9282 0.00016235 -85.653 0.82895
7.933 0.98813 5.4693e-005 3.8183 0.011929 0.00010321 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5352 0.5556 0.16997 0.019773 15.842 0.12265 0.00015959 0.76751 0.0092491 0.01024 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16368 0.93829 0.91733 0.0013969 0.99314 0.50104 0.001882 0.42672 2.163 2.1625 16.0107 144.9282 0.00016227 -85.6531 0.82995
7.934 0.98813 5.4693e-005 3.8183 0.011929 0.00010322 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5353 0.55565 0.16998 0.019774 15.845 0.12266 0.0001596 0.7675 0.0092495 0.01024 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16368 0.93843 0.91738 0.0013969 0.99316 0.50121 0.001882 0.42673 2.1635 2.1629 16.0107 144.9282 0.00016218 -85.6532 0.83095
7.935 0.98813 5.4693e-005 3.8183 0.011929 0.00010324 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5354 0.55569 0.17 0.019775 15.8479 0.12266 0.00015961 0.7675 0.0092499 0.01024 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16368 0.93857 0.91744 0.0013969 0.99319 0.50139 0.001882 0.42675 2.1639 2.1633 16.0107 144.9282 0.0001621 -85.6533 0.83195
7.936 0.98813 5.4693e-005 3.8183 0.011929 0.00010325 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5355 0.55574 0.17001 0.019776 15.8508 0.12267 0.00015962 0.76749 0.0092503 0.010241 0.0013859 0.98695 0.99171 2.9884e-006 1.1954e-005 0.16369 0.93871 0.91749 0.0013969 0.99322 0.50156 0.001882 0.42676 2.1643 2.1637 16.0106 144.9282 0.00016201 -85.6533 0.83295
7.937 0.98813 5.4693e-005 3.8183 0.011929 0.00010326 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5356 0.55578 0.17003 0.019778 15.8537 0.12268 0.00015963 0.76748 0.0092507 0.010241 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.16369 0.93885 0.91754 0.0013969 0.99324 0.50173 0.001882 0.42677 2.1647 2.1642 16.0106 144.9283 0.00016193 -85.6534 0.83395
7.938 0.98813 5.4693e-005 3.8183 0.011929 0.00010328 0.0011717 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5357 0.55583 0.17004 0.019779 15.8566 0.12268 0.00015964 0.76748 0.0092511 0.010242 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16369 0.93899 0.9176 0.0013969 0.99327 0.50191 0.001882 0.42679 2.1652 2.1646 16.0106 144.9283 0.00016185 -85.6535 0.83495
7.939 0.98813 5.4693e-005 3.8183 0.011929 0.00010329 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5357 0.55587 0.17005 0.01978 15.8596 0.12269 0.00015965 0.76747 0.0092515 0.010242 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.1637 0.93913 0.91765 0.0013969 0.99329 0.50208 0.001882 0.4268 2.1656 2.165 16.0105 144.9283 0.00016177 -85.6536 0.83595
7.94 0.98813 5.4693e-005 3.8183 0.011929 0.0001033 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5358 0.55592 0.17007 0.019781 15.8625 0.1227 0.00015966 0.76746 0.0092519 0.010243 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.1637 0.93927 0.9177 0.0013969 0.99332 0.50225 0.0018819 0.42681 2.166 2.1654 16.0105 144.9283 0.00016168 -85.6537 0.83695
7.941 0.98813 5.4693e-005 3.8183 0.011929 0.00010331 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5359 0.55596 0.17008 0.019782 15.8654 0.1227 0.00015967 0.76746 0.0092523 0.010243 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.1637 0.93941 0.91776 0.0013969 0.99334 0.50243 0.0018819 0.42683 2.1664 2.1659 16.0105 144.9283 0.0001616 -85.6537 0.83795
7.942 0.98813 5.4693e-005 3.8183 0.011929 0.00010333 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.536 0.55601 0.17009 0.019783 15.8683 0.12271 0.00015968 0.76745 0.0092527 0.010243 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.1637 0.93955 0.91781 0.0013969 0.99337 0.5026 0.0018819 0.42684 2.1668 2.1663 16.0105 144.9284 0.00016152 -85.6538 0.83895
7.943 0.98813 5.4692e-005 3.8183 0.011929 0.00010334 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5361 0.55605 0.17011 0.019784 15.8713 0.12272 0.00015969 0.76744 0.0092531 0.010244 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16371 0.93968 0.91786 0.0013968 0.99339 0.50277 0.0018819 0.42685 2.1673 2.1667 16.0104 144.9284 0.00016144 -85.6539 0.83995
7.944 0.98813 5.4692e-005 3.8183 0.011929 0.00010335 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5362 0.5561 0.17012 0.019785 15.8742 0.12272 0.0001597 0.76744 0.0092535 0.010244 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16371 0.93982 0.91792 0.0013968 0.99342 0.50295 0.0018819 0.42687 2.1677 2.1671 16.0104 144.9284 0.00016136 -85.6539 0.84095
7.945 0.98813 5.4692e-005 3.8183 0.011929 0.00010337 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5363 0.55614 0.17013 0.019787 15.8771 0.12273 0.00015972 0.76743 0.0092539 0.010245 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16371 0.93996 0.91797 0.0013968 0.99344 0.50312 0.0018819 0.42688 2.1681 2.1675 16.0104 144.9284 0.00016127 -85.654 0.84195
7.946 0.98813 5.4692e-005 3.8183 0.011929 0.00010338 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5363 0.55619 0.17015 0.019788 15.88 0.12274 0.00015973 0.76742 0.0092543 0.010245 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16372 0.94009 0.91802 0.0013968 0.99347 0.50329 0.0018819 0.42689 2.1685 2.168 16.0103 144.9284 0.00016119 -85.6541 0.84295
7.947 0.98813 5.4692e-005 3.8183 0.011929 0.00010339 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5364 0.55623 0.17016 0.019789 15.8829 0.12274 0.00015974 0.76742 0.0092547 0.010246 0.0013857 0.98695 0.99171 2.988e-006 1.1952e-005 0.16372 0.94023 0.91807 0.0013968 0.99349 0.50347 0.0018819 0.42691 2.1689 2.1684 16.0103 144.9285 0.00016111 -85.6542 0.84395
7.948 0.98813 5.4692e-005 3.8183 0.011929 0.0001034 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5365 0.55628 0.17018 0.01979 15.8859 0.12275 0.00015975 0.76741 0.0092551 0.010246 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.16372 0.94037 0.91812 0.0013968 0.99351 0.50364 0.0018818 0.42692 2.1693 2.1688 16.0103 144.9285 0.00016103 -85.6542 0.84495
7.949 0.98813 5.4692e-005 3.8183 0.011929 0.00010342 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5366 0.55632 0.17019 0.019791 15.8888 0.12276 0.00015976 0.7674 0.0092555 0.010246 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.16373 0.9405 0.91818 0.0013968 0.99354 0.50381 0.0018818 0.42694 2.1698 2.1692 16.0102 144.9285 0.00016095 -85.6543 0.84595
7.95 0.98813 5.4692e-005 3.8183 0.011929 0.00010343 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5367 0.55637 0.1702 0.019792 15.8917 0.12276 0.00015977 0.7674 0.0092559 0.010247 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.16373 0.94063 0.91823 0.0013968 0.99356 0.50399 0.0018818 0.42695 2.1702 2.1696 16.0102 144.9285 0.00016087 -85.6544 0.84695
7.951 0.98813 5.4692e-005 3.8183 0.011929 0.00010344 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5368 0.55641 0.17022 0.019793 15.8946 0.12277 0.00015978 0.76739 0.0092563 0.010247 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16373 0.94077 0.91828 0.0013968 0.99359 0.50416 0.0018818 0.42696 2.1706 2.17 16.0102 144.9286 0.00016079 -85.6544 0.84795
7.952 0.98813 5.4692e-005 3.8183 0.011929 0.00010345 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5369 0.55646 0.17023 0.019794 15.8976 0.12278 0.00015979 0.76738 0.0092567 0.010248 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16374 0.9409 0.91833 0.0013968 0.99361 0.50433 0.0018818 0.42698 2.171 2.1704 16.0101 144.9286 0.00016072 -85.6545 0.84895
7.953 0.98813 5.4692e-005 3.8183 0.011929 0.00010347 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5369 0.5565 0.17024 0.019796 15.9005 0.12278 0.0001598 0.76738 0.009257 0.010248 0.0013856 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16374 0.94104 0.91838 0.0013968 0.99363 0.5045 0.0018818 0.42699 2.1714 2.1709 16.0101 144.9286 0.00016064 -85.6546 0.84995
7.954 0.98813 5.4692e-005 3.8183 0.011929 0.00010348 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.537 0.55655 0.17026 0.019797 15.9034 0.12279 0.00015981 0.76737 0.0092574 0.010248 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16374 0.94117 0.91843 0.0013967 0.99366 0.50468 0.0018818 0.427 2.1718 2.1713 16.0101 144.9286 0.00016056 -85.6547 0.85095
7.955 0.98813 5.4691e-005 3.8183 0.011929 0.00010349 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5371 0.55659 0.17027 0.019798 15.9064 0.1228 0.00015982 0.76736 0.0092578 0.010249 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16374 0.9413 0.91848 0.0013967 0.99368 0.50485 0.0018818 0.42702 2.1722 2.1717 16.01 144.9286 0.00016048 -85.6547 0.85195
7.956 0.98813 5.4691e-005 3.8183 0.011929 0.00010351 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5372 0.55664 0.17028 0.019799 15.9093 0.1228 0.00015983 0.76736 0.0092582 0.010249 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16375 0.94143 0.91853 0.0013967 0.9937 0.50502 0.0018818 0.42703 2.1726 2.1721 16.01 144.9287 0.0001604 -85.6548 0.85295
7.957 0.98813 5.4691e-005 3.8183 0.011929 0.00010352 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5373 0.55668 0.1703 0.0198 15.9122 0.12281 0.00015984 0.76735 0.0092586 0.01025 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16375 0.94156 0.91858 0.0013967 0.99372 0.50519 0.0018817 0.42704 2.173 2.1725 16.01 144.9287 0.00016032 -85.6549 0.85395
7.958 0.98813 5.4691e-005 3.8183 0.011929 0.00010353 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5374 0.55673 0.17031 0.019801 15.9151 0.12282 0.00015985 0.76734 0.009259 0.01025 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16375 0.9417 0.91863 0.0013967 0.99375 0.50537 0.0018817 0.42706 2.1734 2.1729 16.01 144.9287 0.00016025 -85.6549 0.85495
7.959 0.98813 5.4691e-005 3.8183 0.011929 0.00010354 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5375 0.55677 0.17033 0.019802 15.9181 0.12282 0.00015986 0.76734 0.0092594 0.010251 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.16376 0.94183 0.91868 0.0013967 0.99377 0.50554 0.0018817 0.42707 2.1739 2.1733 16.0099 144.9287 0.00016017 -85.655 0.85595
7.96 0.98813 5.4691e-005 3.8183 0.011929 0.00010356 0.0011718 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5376 0.55682 0.17034 0.019803 15.921 0.12283 0.00015987 0.76733 0.0092598 0.010251 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.16376 0.94196 0.91873 0.0013967 0.99379 0.50571 0.0018817 0.42708 2.1743 2.1737 16.0099 144.9287 0.00016009 -85.6551 0.85695
7.961 0.98813 5.4691e-005 3.8183 0.011929 0.00010357 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5376 0.55686 0.17035 0.019804 15.9239 0.12284 0.00015988 0.76732 0.0092602 0.010251 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.16376 0.94209 0.91878 0.0013967 0.99381 0.50588 0.0018817 0.4271 2.1747 2.1741 16.0099 144.9288 0.00016001 -85.6551 0.85795
7.962 0.98813 5.4691e-005 3.8183 0.011929 0.00010358 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5377 0.55691 0.17037 0.019806 15.9269 0.12284 0.00015989 0.76732 0.0092606 0.010252 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.16377 0.94222 0.91883 0.0013967 0.99383 0.50606 0.0018817 0.42711 2.1751 2.1745 16.0098 144.9288 0.00015994 -85.6552 0.85895
7.963 0.98813 5.4691e-005 3.8183 0.011929 0.0001036 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5378 0.55695 0.17038 0.019807 15.9298 0.12285 0.0001599 0.76731 0.009261 0.010252 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.16377 0.94235 0.91888 0.0013967 0.99386 0.50623 0.0018817 0.42712 2.1755 2.1749 16.0098 144.9288 0.00015986 -85.6552 0.85995
7.964 0.98813 5.4691e-005 3.8183 0.011929 0.00010361 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5379 0.557 0.17039 0.019808 15.9327 0.12286 0.00015991 0.7673 0.0092614 0.010253 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.16377 0.94247 0.91893 0.0013967 0.99388 0.5064 0.0018817 0.42714 2.1759 2.1753 16.0098 144.9288 0.00015979 -85.6553 0.86095
7.965 0.98813 5.4691e-005 3.8183 0.011929 0.00010362 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.538 0.55704 0.17041 0.019809 15.9356 0.12286 0.00015992 0.7673 0.0092618 0.010253 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16377 0.9426 0.91898 0.0013967 0.9939 0.50657 0.0018817 0.42715 2.1763 2.1757 16.0097 144.9288 0.00015971 -85.6554 0.86195
7.966 0.98813 5.4691e-005 3.8183 0.011928 0.00010363 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5381 0.55709 0.17042 0.01981 15.9386 0.12287 0.00015993 0.76729 0.0092622 0.010254 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16378 0.94273 0.91903 0.0013967 0.99392 0.50674 0.0018817 0.42716 2.1767 2.1761 16.0097 144.9289 0.00015963 -85.6554 0.86295
7.967 0.98813 5.469e-005 3.8183 0.011928 0.00010365 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5382 0.55713 0.17043 0.019811 15.9415 0.12288 0.00015994 0.76728 0.0092626 0.010254 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16378 0.94286 0.91908 0.0013966 0.99394 0.50691 0.0018816 0.42718 2.1771 2.1765 16.0097 144.9289 0.00015956 -85.6555 0.86395
7.968 0.98813 5.469e-005 3.8183 0.011928 0.00010366 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5382 0.55718 0.17045 0.019812 15.9444 0.12288 0.00015995 0.76728 0.009263 0.010254 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16378 0.94298 0.91912 0.0013966 0.99396 0.50709 0.0018816 0.42719 2.1775 2.1769 16.0096 144.9289 0.00015948 -85.6556 0.86495
7.969 0.98813 5.469e-005 3.8183 0.011928 0.00010367 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5383 0.55722 0.17046 0.019813 15.9474 0.12289 0.00015996 0.76727 0.0092634 0.010255 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16379 0.94311 0.91917 0.0013966 0.99398 0.50726 0.0018816 0.4272 2.1779 2.1773 16.0096 144.9289 0.00015941 -85.6556 0.86595
7.97 0.98813 5.469e-005 3.8183 0.011928 0.00010369 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5384 0.55727 0.17048 0.019815 15.9503 0.1229 0.00015997 0.76726 0.0092638 0.010255 0.0013854 0.98696 0.99171 2.9872e-006 1.1949e-005 0.16379 0.94324 0.91922 0.0013966 0.994 0.50743 0.0018816 0.42722 2.1783 2.1777 16.0096 144.9289 0.00015934 -85.6557 0.86695
7.971 0.98813 5.469e-005 3.8183 0.011928 0.0001037 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5385 0.55731 0.17049 0.019816 15.9532 0.1229 0.00015998 0.76726 0.0092642 0.010256 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16379 0.94336 0.91927 0.0013966 0.99402 0.5076 0.0018816 0.42723 2.1787 2.1781 16.0095 144.929 0.00015926 -85.6557 0.86795
7.972 0.98813 5.469e-005 3.8183 0.011928 0.00010371 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5386 0.55736 0.1705 0.019817 15.9562 0.12291 0.00015999 0.76725 0.0092646 0.010256 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.1638 0.94349 0.91932 0.0013966 0.99405 0.50777 0.0018816 0.42724 2.1791 2.1785 16.0095 144.929 0.00015919 -85.6558 0.86895
7.973 0.98813 5.469e-005 3.8183 0.011928 0.00010372 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5387 0.5574 0.17052 0.019818 15.9591 0.12292 0.00016 0.76724 0.009265 0.010256 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.1638 0.94361 0.91936 0.0013966 0.99407 0.50794 0.0018816 0.42726 2.1795 2.1789 16.0095 144.929 0.00015911 -85.6559 0.86995
7.974 0.98813 5.469e-005 3.8183 0.011928 0.00010374 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5388 0.55745 0.17053 0.019819 15.962 0.12292 0.00016001 0.76724 0.0092653 0.010257 0.0013853 0.98696 0.99171 2.9871e-006 1.1948e-005 0.1638 0.94374 0.91941 0.0013966 0.99409 0.50812 0.0018816 0.42727 2.1799 2.1793 16.0095 144.929 0.00015904 -85.6559 0.87095
7.975 0.98813 5.469e-005 3.8183 0.011928 0.00010375 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5389 0.55749 0.17054 0.01982 15.965 0.12293 0.00016002 0.76723 0.0092657 0.010257 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16381 0.94386 0.91946 0.0013966 0.99411 0.50829 0.0018816 0.42728 2.1802 2.1797 16.0094 144.929 0.00015897 -85.656 0.87195
7.976 0.98813 5.469e-005 3.8183 0.011928 0.00010376 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5389 0.55753 0.17056 0.019821 15.9679 0.12294 0.00016003 0.76722 0.0092661 0.010258 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16381 0.94399 0.91951 0.0013966 0.99413 0.50846 0.0018816 0.4273 2.1806 2.1801 16.0094 144.9291 0.00015889 -85.656 0.87295
7.977 0.98813 5.469e-005 3.8183 0.011928 0.00010378 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.539 0.55758 0.17057 0.019822 15.9708 0.12294 0.00016004 0.76722 0.0092665 0.010258 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16381 0.94411 0.91955 0.0013966 0.99415 0.50863 0.0018815 0.42731 2.181 2.1805 16.0094 144.9291 0.00015882 -85.6561 0.87395
7.978 0.98813 5.469e-005 3.8183 0.011928 0.00010379 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5391 0.55762 0.17058 0.019823 15.9738 0.12295 0.00016005 0.76721 0.0092669 0.010259 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16381 0.94423 0.9196 0.0013966 0.99417 0.5088 0.0018815 0.42732 2.1814 2.1809 16.0093 144.9291 0.00015875 -85.6561 0.87495
7.979 0.98813 5.4689e-005 3.8183 0.011928 0.0001038 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5392 0.55767 0.1706 0.019825 15.9767 0.12296 0.00016006 0.7672 0.0092673 0.010259 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16382 0.94436 0.91965 0.0013966 0.99418 0.50897 0.0018815 0.42734 2.1818 2.1813 16.0093 144.9291 0.00015868 -85.6562 0.87595
7.98 0.98813 5.4689e-005 3.8183 0.011928 0.00010381 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5393 0.55771 0.17061 0.019826 15.9796 0.12296 0.00016007 0.7672 0.0092677 0.010259 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16382 0.94448 0.91969 0.0013966 0.9942 0.50914 0.0018815 0.42735 2.1822 2.1817 16.0093 144.9291 0.00015861 -85.6562 0.87695
7.981 0.98813 5.4689e-005 3.8183 0.011928 0.00010383 0.0011719 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5394 0.55776 0.17063 0.019827 15.9826 0.12297 0.00016008 0.76719 0.0092681 0.01026 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16382 0.9446 0.91974 0.0013965 0.99422 0.50931 0.0018815 0.42736 2.1826 2.1821 16.0092 144.9292 0.00015853 -85.6563 0.87795
7.982 0.98813 5.4689e-005 3.8183 0.011928 0.00010384 0.001172 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5395 0.5578 0.17064 0.019828 15.9855 0.12298 0.00016009 0.76718 0.0092685 0.01026 0.0013853 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16383 0.94472 0.91978 0.0013965 0.99424 0.50949 0.0018815 0.42738 2.183 2.1825 16.0092 144.9292 0.00015846 -85.6564 0.87895
7.983 0.98813 5.4689e-005 3.8183 0.011928 0.00010385 0.001172 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5395 0.55785 0.17065 0.019829 15.9884 0.12298 0.0001601 0.76718 0.0092689 0.010261 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16383 0.94485 0.91983 0.0013965 0.99426 0.50966 0.0018815 0.42739 2.1834 2.1829 16.0092 144.9292 0.00015839 -85.6564 0.87995
7.984 0.98813 5.4689e-005 3.8183 0.011928 0.00010387 0.001172 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5396 0.55789 0.17067 0.01983 15.9914 0.12299 0.00016011 0.76717 0.0092693 0.010261 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16383 0.94497 0.91988 0.0013965 0.99428 0.50983 0.0018815 0.4274 2.1838 2.1832 16.0091 144.9292 0.00015832 -85.6565 0.88095
7.985 0.98813 5.4689e-005 3.8183 0.011928 0.00010388 0.001172 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5397 0.55794 0.17068 0.019831 15.9943 0.123 0.00016012 0.76716 0.0092697 0.010261 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16384 0.94509 0.91992 0.0013965 0.9943 0.51 0.0018815 0.42742 2.1842 2.1836 16.0091 144.9293 0.00015825 -85.6565 0.88195
7.986 0.98813 5.4689e-005 3.8183 0.011928 0.00010389 0.001172 0.23374 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5398 0.55798 0.17069 0.019832 15.9973 0.123 0.00016013 0.76716 0.0092701 0.010262 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16384 0.94521 0.91997 0.0013965 0.99432 0.51017 0.0018815 0.42743 2.1845 2.184 16.0091 144.9293 0.00015818 -85.6566 0.88295
7.987 0.98813 5.4689e-005 3.8183 0.011928 0.0001039 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5399 0.55803 0.17071 0.019834 16.0002 0.12301 0.00016014 0.76715 0.0092705 0.010262 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16384 0.94533 0.92001 0.0013965 0.99434 0.51034 0.0018815 0.42744 2.1849 2.1844 16.009 144.9293 0.00015811 -85.6566 0.88395
7.988 0.98813 5.4689e-005 3.8183 0.011928 0.00010392 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.54 0.55807 0.17072 0.019835 16.0031 0.12302 0.00016015 0.76714 0.0092709 0.010263 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16384 0.94545 0.92006 0.0013965 0.99436 0.51051 0.0018815 0.42746 2.1853 2.1848 16.009 144.9293 0.00015804 -85.6567 0.88495
7.989 0.98813 5.4689e-005 3.8183 0.011928 0.00010393 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5401 0.55812 0.17073 0.019836 16.0061 0.12302 0.00016016 0.76714 0.0092713 0.010263 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16385 0.94556 0.9201 0.0013965 0.99437 0.51068 0.0018814 0.42747 2.1857 2.1852 16.009 144.9293 0.00015797 -85.6567 0.88595
7.99 0.98813 5.4689e-005 3.8183 0.011928 0.00010394 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5401 0.55816 0.17075 0.019837 16.009 0.12303 0.00016017 0.76713 0.0092717 0.010264 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16385 0.94568 0.92015 0.0013965 0.99439 0.51085 0.0018814 0.42748 2.1861 2.1856 16.0089 144.9294 0.0001579 -85.6568 0.88695
7.991 0.98813 5.4689e-005 3.8183 0.011928 0.00010396 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5402 0.55821 0.17076 0.019838 16.012 0.12304 0.00016018 0.76712 0.009272 0.010264 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16385 0.9458 0.92019 0.0013965 0.99441 0.51102 0.0018814 0.4275 2.1865 2.1859 16.0089 144.9294 0.00015783 -85.6568 0.88795
7.992 0.98813 5.4688e-005 3.8183 0.011928 0.00010397 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5403 0.55825 0.17078 0.019839 16.0149 0.12304 0.00016019 0.76712 0.0092724 0.010264 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16386 0.94592 0.92024 0.0013965 0.99443 0.51119 0.0018814 0.42751 2.1868 2.1863 16.0089 144.9294 0.00015776 -85.6569 0.88895
7.993 0.98813 5.4688e-005 3.8183 0.011928 0.00010398 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5404 0.5583 0.17079 0.01984 16.0178 0.12305 0.0001602 0.76711 0.0092728 0.010265 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16386 0.94604 0.92028 0.0013965 0.99445 0.51136 0.0018814 0.42752 2.1872 2.1867 16.0088 144.9294 0.00015769 -85.6569 0.88995
7.994 0.98813 5.4688e-005 3.8183 0.011928 0.00010399 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5405 0.55834 0.1708 0.019841 16.0208 0.12306 0.00016021 0.7671 0.0092732 0.010265 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16386 0.94615 0.92033 0.0013965 0.99446 0.51153 0.0018814 0.42754 2.1876 2.1871 16.0088 144.9294 0.00015762 -85.657 0.89095
7.995 0.98813 5.4688e-005 3.8183 0.011928 0.00010401 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5406 0.55839 0.17082 0.019842 16.0237 0.12306 0.00016022 0.7671 0.0092736 0.010266 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16387 0.94627 0.92037 0.0013965 0.99448 0.5117 0.0018814 0.42755 2.188 2.1875 16.0088 144.9295 0.00015756 -85.657 0.89195
7.996 0.98813 5.4688e-005 3.8183 0.011928 0.00010402 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5407 0.55843 0.17083 0.019844 16.0267 0.12307 0.00016023 0.76709 0.009274 0.010266 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.16387 0.94639 0.92041 0.0013965 0.9945 0.51187 0.0018814 0.42756 2.1884 2.1879 16.0088 144.9295 0.00015749 -85.6571 0.89295
7.997 0.98813 5.4688e-005 3.8183 0.011928 0.00010403 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5408 0.55848 0.17084 0.019845 16.0296 0.12308 0.00016024 0.76708 0.0092744 0.010266 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.16387 0.9465 0.92046 0.0013964 0.99452 0.51204 0.0018814 0.42758 2.1887 2.1882 16.0087 144.9295 0.00015742 -85.6571 0.89395
7.998 0.98813 5.4688e-005 3.8183 0.011928 0.00010404 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5408 0.55852 0.17086 0.019846 16.0325 0.12308 0.00016025 0.76708 0.0092748 0.010267 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.16388 0.94662 0.9205 0.0013964 0.99453 0.51221 0.0018814 0.42759 2.1891 2.1886 16.0087 144.9295 0.00015735 -85.6572 0.89495
7.999 0.98813 5.4688e-005 3.8183 0.011928 0.00010406 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5409 0.55857 0.17087 0.019847 16.0355 0.12309 0.00016026 0.76707 0.0092752 0.010267 0.0013851 0.98696 0.99171 2.9864e-006 1.1945e-005 0.16388 0.94674 0.92054 0.0013964 0.99455 0.51238 0.0018814 0.4276 2.1895 2.189 16.0087 144.9295 0.00015728 -85.6572 0.89595
8 0.98813 5.4688e-005 3.8183 0.011928 0.00010407 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.541 0.55861 0.17088 0.019848 16.0384 0.1231 0.00016027 0.76706 0.0092756 0.010268 0.0013851 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16388 0.94685 0.92059 0.0013964 0.99457 0.51255 0.0018814 0.42762 2.1899 2.1894 16.0086 144.9296 0.00015722 -85.6573 0.89695
8.001 0.98813 5.4688e-005 3.8183 0.011928 0.00010408 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5411 0.55866 0.1709 0.019849 16.0414 0.1231 0.00016028 0.76706 0.009276 0.010268 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16388 0.94696 0.92063 0.0013964 0.99458 0.51272 0.0018814 0.42763 2.1903 2.1897 16.0086 144.9296 0.00015715 -85.6573 0.89795
8.002 0.98813 5.4688e-005 3.8183 0.011928 0.0001041 0.001172 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5412 0.5587 0.17091 0.01985 16.0443 0.12311 0.00016029 0.76705 0.0092764 0.010269 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16389 0.94708 0.92067 0.0013964 0.9946 0.51289 0.0018813 0.42764 2.1906 2.1901 16.0086 144.9296 0.00015708 -85.6574 0.89895
8.003 0.98813 5.4688e-005 3.8183 0.011928 0.00010411 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5413 0.55875 0.17092 0.019851 16.0472 0.12312 0.0001603 0.76704 0.0092768 0.010269 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16389 0.94719 0.92072 0.0013964 0.99462 0.51306 0.0018813 0.42766 2.191 2.1905 16.0085 144.9296 0.00015702 -85.6574 0.89995
8.004 0.98813 5.4687e-005 3.8183 0.011928 0.00010412 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5414 0.55879 0.17094 0.019853 16.0502 0.12312 0.00016031 0.76704 0.0092772 0.010269 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16389 0.94731 0.92076 0.0013964 0.99463 0.51323 0.0018813 0.42767 2.1914 2.1909 16.0085 144.9296 0.00015695 -85.6575 0.90095
8.005 0.98813 5.4687e-005 3.8183 0.011928 0.00010413 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5414 0.55884 0.17095 0.019854 16.0531 0.12313 0.00016032 0.76703 0.0092775 0.01027 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.1639 0.94742 0.9208 0.0013964 0.99465 0.5134 0.0018813 0.42768 2.1917 2.1912 16.0085 144.9297 0.00015688 -85.6575 0.90195
8.006 0.98813 5.4687e-005 3.8183 0.011928 0.00010415 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5415 0.55888 0.17097 0.019855 16.0561 0.12314 0.00016033 0.76702 0.0092779 0.01027 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.1639 0.94753 0.92085 0.0013964 0.99467 0.51357 0.0018813 0.4277 2.1921 2.1916 16.0084 144.9297 0.00015682 -85.6575 0.90295
8.007 0.98813 5.4687e-005 3.8183 0.011928 0.00010416 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5416 0.55893 0.17098 0.019856 16.059 0.12314 0.00016034 0.76702 0.0092783 0.010271 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.1639 0.94765 0.92089 0.0013964 0.99468 0.51374 0.0018813 0.42771 2.1925 2.192 16.0084 144.9297 0.00015675 -85.6576 0.90395
8.008 0.98813 5.4687e-005 3.8183 0.011928 0.00010417 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5417 0.55897 0.17099 0.019857 16.062 0.12315 0.00016035 0.76701 0.0092787 0.010271 0.001385 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16391 0.94776 0.92093 0.0013964 0.9947 0.51391 0.0018813 0.42772 2.1929 2.1924 16.0084 144.9297 0.00015669 -85.6576 0.90495
8.009 0.98813 5.4687e-005 3.8183 0.011928 0.00010419 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5418 0.55902 0.17101 0.019858 16.0649 0.12316 0.00016036 0.767 0.0092791 0.010272 0.001385 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16391 0.94787 0.92097 0.0013964 0.99472 0.51408 0.0018813 0.42774 2.1932 2.1927 16.0083 144.9297 0.00015662 -85.6577 0.90595
8.01 0.98813 5.4687e-005 3.8183 0.011928 0.0001042 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5419 0.55906 0.17102 0.019859 16.0679 0.12316 0.00016037 0.767 0.0092795 0.010272 0.001385 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16391 0.94798 0.92101 0.0013964 0.99473 0.51425 0.0018813 0.42775 2.1936 2.1931 16.0083 144.9298 0.00015656 -85.6577 0.90695
8.011 0.98813 5.4687e-005 3.8183 0.011928 0.00010421 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.542 0.55911 0.17103 0.01986 16.0708 0.12317 0.00016038 0.76699 0.0092799 0.010272 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16391 0.94809 0.92106 0.0013964 0.99475 0.51442 0.0018813 0.42776 2.194 2.1935 16.0083 144.9298 0.00015649 -85.6578 0.90795
8.012 0.98813 5.4687e-005 3.8183 0.011928 0.00010422 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.542 0.55915 0.17105 0.019861 16.0738 0.12318 0.00016039 0.76698 0.0092803 0.010273 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16392 0.9482 0.9211 0.0013964 0.99476 0.51459 0.0018813 0.42778 2.1943 2.1939 16.0082 144.9298 0.00015643 -85.6578 0.90895
8.013 0.98813 5.4687e-005 3.8183 0.011928 0.00010424 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5421 0.5592 0.17106 0.019863 16.0767 0.12318 0.0001604 0.76698 0.0092807 0.010273 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16392 0.94831 0.92114 0.0013964 0.99478 0.51476 0.0018813 0.42779 2.1947 2.1942 16.0082 144.9298 0.00015636 -85.6578 0.90995
8.014 0.98813 5.4687e-005 3.8183 0.011928 0.00010425 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5422 0.55924 0.17107 0.019864 16.0796 0.12319 0.00016041 0.76697 0.0092811 0.010274 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16392 0.94842 0.92118 0.0013964 0.99479 0.51493 0.0018813 0.4278 2.1951 2.1946 16.0082 144.9298 0.0001563 -85.6579 0.91095
8.015 0.98813 5.4687e-005 3.8183 0.011928 0.00010426 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5423 0.55929 0.17109 0.019865 16.0826 0.1232 0.00016042 0.76696 0.0092815 0.010274 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16393 0.94853 0.92122 0.0013963 0.99481 0.51509 0.0018813 0.42782 2.1954 2.195 16.0081 144.9299 0.00015624 -85.6579 0.91195
8.016 0.98813 5.4686e-005 3.8183 0.011928 0.00010428 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5424 0.55933 0.1711 0.019866 16.0855 0.1232 0.00016043 0.76696 0.0092819 0.010274 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16393 0.94864 0.92126 0.0013963 0.99483 0.51526 0.0018812 0.42783 2.1958 2.1953 16.0081 144.9299 0.00015617 -85.658 0.91295
8.017 0.98813 5.4686e-005 3.8183 0.011928 0.00010429 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5425 0.55938 0.17112 0.019867 16.0885 0.12321 0.00016044 0.76695 0.0092823 0.010275 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16393 0.94875 0.9213 0.0013963 0.99484 0.51543 0.0018812 0.42784 2.1962 2.1957 16.0081 144.9299 0.00015611 -85.658 0.91395
8.018 0.98813 5.4686e-005 3.8183 0.011928 0.0001043 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5426 0.55942 0.17113 0.019868 16.0914 0.12322 0.00016045 0.76694 0.0092826 0.010275 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16394 0.94886 0.92134 0.0013963 0.99486 0.5156 0.0018812 0.42785 2.1965 2.1961 16.008 144.9299 0.00015605 -85.6581 0.91495
8.019 0.98813 5.4686e-005 3.8183 0.011928 0.00010431 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5427 0.55947 0.17114 0.019869 16.0944 0.12322 0.00016046 0.76694 0.009283 0.010276 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16394 0.94897 0.92138 0.0013963 0.99487 0.51577 0.0018812 0.42787 2.1969 2.1964 16.008 144.93 0.00015598 -85.6581 0.91595
8.02 0.98813 5.4686e-005 3.8183 0.011928 0.00010433 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032257 0.0389 0 1.5427 0.55951 0.17116 0.01987 16.0973 0.12323 0.00016047 0.76693 0.0092834 0.010276 0.0013849 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16394 0.94908 0.92143 0.0013963 0.99489 0.51594 0.0018812 0.42788 2.1973 2.1968 16.008 144.93 0.00015592 -85.6581 0.91695
8.021 0.98813 5.4686e-005 3.8183 0.011928 0.00010434 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5428 0.55956 0.17117 0.019871 16.1003 0.12324 0.00016048 0.76692 0.0092838 0.010277 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16394 0.94918 0.92147 0.0013963 0.9949 0.51611 0.0018812 0.42789 2.1976 2.1972 16.0079 144.93 0.00015586 -85.6582 0.91795
8.022 0.98813 5.4686e-005 3.8183 0.011928 0.00010435 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5429 0.5596 0.17118 0.019873 16.1032 0.12324 0.00016049 0.76692 0.0092842 0.010277 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16395 0.94929 0.92151 0.0013963 0.99492 0.51628 0.0018812 0.42791 2.198 2.1975 16.0079 144.93 0.00015579 -85.6582 0.91895
8.023 0.98813 5.4686e-005 3.8183 0.011927 0.00010437 0.0011721 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.543 0.55965 0.1712 0.019874 16.1062 0.12325 0.0001605 0.76691 0.0092846 0.010277 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16395 0.9494 0.92155 0.0013963 0.99493 0.51644 0.0018812 0.42792 2.1984 2.1979 16.0079 144.93 0.00015573 -85.6582 0.91995
8.024 0.98813 5.4686e-005 3.8183 0.011927 0.00010438 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5431 0.55969 0.17121 0.019875 16.1091 0.12326 0.00016051 0.7669 0.009285 0.010278 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16395 0.94951 0.92159 0.0013963 0.99495 0.51661 0.0018812 0.42793 2.1987 2.1982 16.0078 144.9301 0.00015567 -85.6583 0.92095
8.025 0.98813 5.4686e-005 3.8183 0.011927 0.00010439 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5432 0.55974 0.17122 0.019876 16.1121 0.12326 0.00016052 0.7669 0.0092854 0.010278 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16396 0.94961 0.92163 0.0013963 0.99496 0.51678 0.0018812 0.42795 2.1991 2.1986 16.0078 144.9301 0.00015561 -85.6583 0.92195
8.026 0.98813 5.4686e-005 3.8183 0.011927 0.0001044 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5433 0.55978 0.17124 0.019877 16.115 0.12327 0.00016053 0.76689 0.0092858 0.010279 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16396 0.94972 0.92167 0.0013963 0.99497 0.51695 0.0018812 0.42796 2.1994 2.199 16.0078 144.9301 0.00015555 -85.6584 0.92295
8.027 0.98813 5.4686e-005 3.8183 0.011927 0.00010442 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5433 0.55983 0.17125 0.019878 16.118 0.12328 0.00016054 0.76688 0.0092862 0.010279 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16396 0.94982 0.92171 0.0013963 0.99499 0.51712 0.0018812 0.42797 2.1998 2.1993 16.0077 144.9301 0.00015549 -85.6584 0.92395
8.028 0.98813 5.4685e-005 3.8183 0.011927 0.00010443 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5434 0.55987 0.17126 0.019879 16.1209 0.12328 0.00016055 0.76688 0.0092866 0.010279 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16397 0.94993 0.92174 0.0013963 0.995 0.51729 0.0018812 0.42799 2.2002 2.1997 16.0077 144.9301 0.00015543 -85.6584 0.92495
8.029 0.98813 5.4685e-005 3.8183 0.011927 0.00010444 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5435 0.55992 0.17128 0.01988 16.1239 0.12329 0.00016056 0.76687 0.009287 0.01028 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16397 0.95003 0.92178 0.0013963 0.99502 0.51745 0.0018812 0.428 2.2005 2.2 16.0077 144.9302 0.00015536 -85.6585 0.92595
8.03 0.98813 5.4685e-005 3.8183 0.011927 0.00010446 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5436 0.55996 0.17129 0.019881 16.1268 0.1233 0.00016057 0.76686 0.0092873 0.01028 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16397 0.95014 0.92182 0.0013963 0.99503 0.51762 0.0018812 0.42801 2.2009 2.2004 16.0076 144.9302 0.0001553 -85.6585 0.92695
8.031 0.98813 5.4685e-005 3.8183 0.011927 0.00010447 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5437 0.56001 0.17131 0.019883 16.1298 0.1233 0.00016058 0.76686 0.0092877 0.010281 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16397 0.95024 0.92186 0.0013963 0.99504 0.51779 0.0018812 0.42802 2.2012 2.2008 16.0076 144.9302 0.00015524 -85.6585 0.92795
8.032 0.98813 5.4685e-005 3.8183 0.011927 0.00010448 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5438 0.56005 0.17132 0.019884 16.1327 0.12331 0.00016059 0.76685 0.0092881 0.010281 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16398 0.95035 0.9219 0.0013963 0.99506 0.51796 0.0018812 0.42804 2.2016 2.2011 16.0076 144.9302 0.00015518 -85.6586 0.92895
8.033 0.98813 5.4685e-005 3.8183 0.011927 0.00010449 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5439 0.5601 0.17133 0.019885 16.1357 0.12332 0.0001606 0.76684 0.0092885 0.010282 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16398 0.95045 0.92194 0.0013963 0.99507 0.51813 0.0018811 0.42805 2.202 2.2015 16.0075 144.9302 0.00015512 -85.6586 0.92995
8.034 0.98813 5.4685e-005 3.8183 0.011927 0.00010451 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5439 0.56014 0.17135 0.019886 16.1387 0.12332 0.00016061 0.76684 0.0092889 0.010282 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16398 0.95055 0.92198 0.0013963 0.99509 0.51829 0.0018811 0.42806 2.2023 2.2018 16.0075 144.9303 0.00015506 -85.6587 0.93095
8.035 0.98813 5.4685e-005 3.8183 0.011927 0.00010452 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.544 0.56019 0.17136 0.019887 16.1416 0.12333 0.00016062 0.76683 0.0092893 0.010282 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16399 0.95066 0.92202 0.0013963 0.9951 0.51846 0.0018811 0.42808 2.2027 2.2022 16.0075 144.9303 0.000155 -85.6587 0.93195
8.036 0.98813 5.4685e-005 3.8183 0.011927 0.00010453 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5441 0.56023 0.17137 0.019888 16.1446 0.12334 0.00016063 0.76682 0.0092897 0.010283 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16399 0.95076 0.92206 0.0013963 0.99511 0.51863 0.0018811 0.42809 2.203 2.2025 16.0074 144.9303 0.00015494 -85.6587 0.93295
8.037 0.98813 5.4685e-005 3.8183 0.011927 0.00010455 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5442 0.56028 0.17139 0.019889 16.1475 0.12334 0.00016064 0.76682 0.0092901 0.010283 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16399 0.95086 0.92209 0.0013962 0.99513 0.5188 0.0018811 0.4281 2.2034 2.2029 16.0074 144.9303 0.00015488 -85.6588 0.93395
8.038 0.98813 5.4685e-005 3.8183 0.011927 0.00010456 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5443 0.56032 0.1714 0.01989 16.1505 0.12335 0.00016065 0.76681 0.0092905 0.010284 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.164 0.95096 0.92213 0.0013962 0.99514 0.51897 0.0018811 0.42812 2.2037 2.2033 16.0074 144.9303 0.00015483 -85.6588 0.93495
8.039 0.98813 5.4685e-005 3.8183 0.011927 0.00010457 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5444 0.56037 0.17141 0.019891 16.1534 0.12336 0.00016066 0.7668 0.0092909 0.010284 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.164 0.95107 0.92217 0.0013962 0.99515 0.51913 0.0018811 0.42813 2.2041 2.2036 16.0073 144.9304 0.00015477 -85.6588 0.93595
8.04 0.98813 5.4685e-005 3.8183 0.011927 0.00010458 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5445 0.56041 0.17143 0.019893 16.1564 0.12336 0.00016067 0.7668 0.0092913 0.010284 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.164 0.95117 0.92221 0.0013962 0.99517 0.5193 0.0018811 0.42814 2.2044 2.204 16.0073 144.9304 0.00015471 -85.6589 0.93695
8.041 0.98813 5.4684e-005 3.8183 0.011927 0.0001046 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5446 0.56046 0.17144 0.019894 16.1593 0.12337 0.00016068 0.76679 0.0092916 0.010285 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.164 0.95127 0.92224 0.0013962 0.99518 0.51947 0.0018811 0.42815 2.2048 2.2043 16.0073 144.9304 0.00015465 -85.6589 0.93795
8.042 0.98813 5.4684e-005 3.8183 0.011927 0.00010461 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5446 0.5605 0.17145 0.019895 16.1623 0.12338 0.00016069 0.76678 0.009292 0.010285 0.0013846 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16401 0.95137 0.92228 0.0013962 0.99519 0.51964 0.0018811 0.42817 2.2051 2.2047 16.0072 144.9304 0.00015459 -85.6589 0.93895
8.043 0.98813 5.4684e-005 3.8183 0.011927 0.00010462 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5447 0.56055 0.17147 0.019896 16.1653 0.12338 0.0001607 0.76678 0.0092924 0.010286 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.16401 0.95147 0.92232 0.0013962 0.9952 0.5198 0.0018811 0.42818 2.2055 2.205 16.0072 144.9304 0.00015453 -85.659 0.93995
8.044 0.98813 5.4684e-005 3.8183 0.011927 0.00010463 0.0011722 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5448 0.56059 0.17148 0.019897 16.1682 0.12339 0.00016071 0.76677 0.0092928 0.010286 0.0013846 0.98696 0.99172 2.9854e-006 1.1942e-005 0.16401 0.95157 0.92236 0.0013962 0.99522 0.51997 0.0018811 0.42819 2.2058 2.2054 16.0072 144.9305 0.00015447 -85.659 0.94095
8.045 0.98813 5.4684e-005 3.8183 0.011927 0.00010465 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5449 0.56064 0.1715 0.019898 16.1712 0.1234 0.00016072 0.76676 0.0092932 0.010286 0.0013846 0.98697 0.99172 2.9854e-006 1.1942e-005 0.16402 0.95167 0.92239 0.0013962 0.99523 0.52014 0.0018811 0.42821 2.2062 2.2057 16.0071 144.9305 0.00015442 -85.659 0.94195
8.046 0.98813 5.4684e-005 3.8183 0.011927 0.00010466 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.545 0.56068 0.17151 0.019899 16.1741 0.1234 0.00016073 0.76676 0.0092936 0.010287 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16402 0.95177 0.92243 0.0013962 0.99524 0.52031 0.0018811 0.42822 2.2065 2.2061 16.0071 144.9305 0.00015436 -85.659 0.94295
8.047 0.98813 5.4684e-005 3.8183 0.011927 0.00010467 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5451 0.56073 0.17152 0.0199 16.1771 0.12341 0.00016074 0.76675 0.009294 0.010287 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16402 0.95187 0.92247 0.0013962 0.99526 0.52047 0.0018811 0.42823 2.2069 2.2064 16.0071 144.9305 0.0001543 -85.6591 0.94395
8.048 0.98813 5.4684e-005 3.8183 0.011927 0.00010469 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5452 0.56077 0.17154 0.019901 16.18 0.12342 0.00016075 0.76674 0.0092944 0.010288 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16403 0.95197 0.92251 0.0013962 0.99527 0.52064 0.0018811 0.42825 2.2072 2.2068 16.007 144.9305 0.00015424 -85.6591 0.94495
8.049 0.98813 5.4684e-005 3.8183 0.011927 0.0001047 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5452 0.56082 0.17155 0.019903 16.183 0.12342 0.00016076 0.76674 0.0092948 0.010288 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16403 0.95207 0.92254 0.0013962 0.99528 0.52081 0.0018811 0.42826 2.2076 2.2071 16.007 144.9306 0.00015419 -85.6591 0.94595
8.05 0.98813 5.4684e-005 3.8183 0.011927 0.00010471 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5453 0.56086 0.17156 0.019904 16.186 0.12343 0.00016077 0.76673 0.0092952 0.010289 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16403 0.95217 0.92258 0.0013962 0.99529 0.52097 0.0018811 0.42827 2.2079 2.2075 16.007 144.9306 0.00015413 -85.6592 0.94695
8.051 0.98813 5.4684e-005 3.8183 0.011927 0.00010472 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5454 0.56091 0.17158 0.019905 16.1889 0.12344 0.00016078 0.76672 0.0092955 0.010289 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16404 0.95226 0.92262 0.0013962 0.9953 0.52114 0.0018811 0.42828 2.2083 2.2078 16.0069 144.9306 0.00015407 -85.6592 0.94795
8.052 0.98813 5.4684e-005 3.8183 0.011927 0.00010474 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5455 0.56095 0.17159 0.019906 16.1919 0.12344 0.00016079 0.76672 0.0092959 0.010289 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16404 0.95236 0.92265 0.0013962 0.99532 0.52131 0.001881 0.4283 2.2086 2.2081 16.0069 144.9306 0.00015402 -85.6592 0.94895
8.053 0.98813 5.4683e-005 3.8183 0.011927 0.00010475 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5456 0.561 0.1716 0.019907 16.1948 0.12345 0.0001608 0.76671 0.0092963 0.01029 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16404 0.95246 0.92269 0.0013962 0.99533 0.52147 0.001881 0.42831 2.2089 2.2085 16.0069 144.9307 0.00015396 -85.6593 0.94995
8.054 0.98813 5.4683e-005 3.8183 0.011927 0.00010476 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5457 0.56104 0.17162 0.019908 16.1978 0.12346 0.00016081 0.7667 0.0092967 0.01029 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16404 0.95256 0.92272 0.0013962 0.99534 0.52164 0.001881 0.42832 2.2093 2.2088 16.0068 144.9307 0.00015391 -85.6593 0.95095
8.055 0.98813 5.4683e-005 3.8183 0.011927 0.00010478 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5458 0.56109 0.17163 0.019909 16.2008 0.12346 0.00016082 0.7667 0.0092971 0.010291 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16405 0.95265 0.92276 0.0013962 0.99535 0.52181 0.001881 0.42834 2.2096 2.2092 16.0068 144.9307 0.00015385 -85.6593 0.95195
8.056 0.98813 5.4683e-005 3.8183 0.011927 0.00010479 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5458 0.56113 0.17164 0.01991 16.2037 0.12347 0.00016083 0.76669 0.0092975 0.010291 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16405 0.95275 0.9228 0.0013962 0.99536 0.52197 0.001881 0.42835 2.21 2.2095 16.0068 144.9307 0.00015379 -85.6594 0.95295
8.057 0.98813 5.4683e-005 3.8183 0.011927 0.0001048 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5459 0.56118 0.17166 0.019911 16.2067 0.12348 0.00016084 0.76668 0.0092979 0.010291 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16405 0.95284 0.92283 0.0013962 0.99538 0.52214 0.001881 0.42836 2.2103 2.2099 16.0067 144.9307 0.00015374 -85.6594 0.95395
8.058 0.98813 5.4683e-005 3.8183 0.011927 0.00010481 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.546 0.56122 0.17167 0.019913 16.2096 0.12348 0.00016085 0.76668 0.0092983 0.010292 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16406 0.95294 0.92287 0.0013962 0.99539 0.52231 0.001881 0.42837 2.2107 2.2102 16.0067 144.9308 0.00015368 -85.6594 0.95495
8.059 0.98813 5.4683e-005 3.8183 0.011927 0.00010483 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5461 0.56126 0.17169 0.019914 16.2126 0.12349 0.00016086 0.76667 0.0092987 0.010292 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16406 0.95304 0.9229 0.0013962 0.9954 0.52247 0.001881 0.42839 2.211 2.2106 16.0067 144.9308 0.00015363 -85.6594 0.95595
8.06 0.98813 5.4683e-005 3.8183 0.011927 0.00010484 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5462 0.56131 0.1717 0.019915 16.2156 0.1235 0.00016087 0.76666 0.0092991 0.010293 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16406 0.95313 0.92294 0.0013962 0.99541 0.52264 0.001881 0.4284 2.2113 2.2109 16.0066 144.9308 0.00015357 -85.6595 0.95695
8.061 0.98813 5.4683e-005 3.8183 0.011927 0.00010485 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5463 0.56135 0.17171 0.019916 16.2185 0.1235 0.00016088 0.76666 0.0092994 0.010293 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16407 0.95323 0.92297 0.0013962 0.99542 0.52281 0.001881 0.42841 2.2117 2.2112 16.0066 144.9308 0.00015352 -85.6595 0.95795
8.062 0.98813 5.4683e-005 3.8183 0.011927 0.00010487 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5464 0.5614 0.17173 0.019917 16.2215 0.12351 0.00016089 0.76665 0.0092998 0.010294 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16407 0.95332 0.92301 0.0013962 0.99543 0.52297 0.001881 0.42843 2.212 2.2116 16.0066 144.9308 0.00015346 -85.6595 0.95895
8.063 0.98813 5.4683e-005 3.8183 0.011927 0.00010488 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5464 0.56144 0.17174 0.019918 16.2245 0.12352 0.0001609 0.76664 0.0093002 0.010294 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16407 0.95342 0.92304 0.0013962 0.99545 0.52314 0.001881 0.42844 2.2124 2.2119 16.0065 144.9309 0.00015341 -85.6595 0.95995
8.064 0.98813 5.4683e-005 3.8183 0.011927 0.00010489 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5465 0.56149 0.17175 0.019919 16.2274 0.12352 0.00016091 0.76664 0.0093006 0.010294 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16407 0.95351 0.92308 0.0013961 0.99546 0.5233 0.001881 0.42845 2.2127 2.2123 16.0065 144.9309 0.00015336 -85.6596 0.96095
8.065 0.98813 5.4682e-005 3.8183 0.011927 0.0001049 0.0011723 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5466 0.56153 0.17177 0.01992 16.2304 0.12353 0.00016092 0.76663 0.009301 0.010295 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16408 0.9536 0.92311 0.0013961 0.99547 0.52347 0.001881 0.42846 2.213 2.2126 16.0065 144.9309 0.0001533 -85.6596 0.96195
8.066 0.98813 5.4682e-005 3.8183 0.011927 0.00010492 0.0011724 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5467 0.56158 0.17178 0.019921 16.2333 0.12354 0.00016093 0.76662 0.0093014 0.010295 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16408 0.9537 0.92315 0.0013961 0.99548 0.52364 0.001881 0.42848 2.2134 2.2129 16.0064 144.9309 0.00015325 -85.6596 0.96295
8.067 0.98813 5.4682e-005 3.8183 0.011927 0.00010493 0.0011724 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5468 0.56162 0.17179 0.019923 16.2363 0.12354 0.00016094 0.76662 0.0093018 0.010296 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16408 0.95379 0.92318 0.0013961 0.99549 0.5238 0.001881 0.42849 2.2137 2.2133 16.0064 144.9309 0.00015319 -85.6596 0.96395
8.068 0.98813 5.4682e-005 3.8183 0.011927 0.00010494 0.0011724 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.5469 0.56167 0.17181 0.019924 16.2393 0.12355 0.00016095 0.76661 0.0093022 0.010296 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16409 0.95388 0.92322 0.0013961 0.9955 0.52397 0.001881 0.4285 2.214 2.2136 16.0064 144.931 0.00015314 -85.6597 0.96495
8.069 0.98813 5.4682e-005 3.8183 0.011927 0.00010496 0.0011724 0.23373 0.00065931 0.23439 0.21629 0 0.032258 0.0389 0 1.547 0.56171 0.17182 0.019925 16.2422 0.12356 0.00016096 0.7666 0.0093026 0.010296 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16409 0.95398 0.92325 0.0013961 0.99551 0.52413 0.001881 0.42852 2.2144 2.2139 16.0063 144.931 0.00015309 -85.6597 0.96595
8.07 0.98813 5.4682e-005 3.8183 0.011927 0.00010497 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5471 0.56176 0.17183 0.019926 16.2452 0.12356 0.00016097 0.7666 0.0093029 0.010297 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16409 0.95407 0.92329 0.0013961 0.99552 0.5243 0.001881 0.42853 2.2147 2.2143 16.0063 144.931 0.00015304 -85.6597 0.96695
8.071 0.98813 5.4682e-005 3.8183 0.011927 0.00010498 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5471 0.5618 0.17185 0.019927 16.2482 0.12357 0.00016098 0.76659 0.0093033 0.010297 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.1641 0.95416 0.92332 0.0013961 0.99553 0.52447 0.001881 0.42854 2.2151 2.2146 16.0063 144.931 0.00015298 -85.6598 0.96795
8.072 0.98813 5.4682e-005 3.8183 0.011927 0.00010499 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5472 0.56185 0.17186 0.019928 16.2511 0.12358 0.00016099 0.76658 0.0093037 0.010298 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.1641 0.95425 0.92335 0.0013961 0.99554 0.52463 0.001881 0.42855 2.2154 2.2149 16.0062 144.931 0.00015293 -85.6598 0.96895
8.073 0.98813 5.4682e-005 3.8183 0.011927 0.00010501 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5473 0.56189 0.17188 0.019929 16.2541 0.12358 0.000161 0.76658 0.0093041 0.010298 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.1641 0.95434 0.92339 0.0013961 0.99555 0.5248 0.001881 0.42857 2.2157 2.2153 16.0062 144.9311 0.00015288 -85.6598 0.96995
8.074 0.98813 5.4682e-005 3.8183 0.011927 0.00010502 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5474 0.56194 0.17189 0.01993 16.2571 0.12359 0.00016101 0.76657 0.0093045 0.010298 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.1641 0.95444 0.92342 0.0013961 0.99556 0.52496 0.001881 0.42858 2.2161 2.2156 16.0062 144.9311 0.00015282 -85.6598 0.97095
8.075 0.98813 5.4682e-005 3.8183 0.011927 0.00010503 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5475 0.56198 0.1719 0.019931 16.26 0.1236 0.00016102 0.76656 0.0093049 0.010299 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.16411 0.95453 0.92345 0.0013961 0.99558 0.52513 0.0018809 0.42859 2.2164 2.2159 16.0061 144.9311 0.00015277 -85.6598 0.97195
8.076 0.98813 5.4682e-005 3.8183 0.011927 0.00010505 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5476 0.56203 0.17192 0.019933 16.263 0.1236 0.00016103 0.76656 0.0093053 0.010299 0.0013844 0.98697 0.99172 2.985e-006 1.194e-005 0.16411 0.95462 0.92349 0.0013961 0.99559 0.52529 0.0018809 0.42861 2.2167 2.2163 16.0061 144.9311 0.00015272 -85.6599 0.97295
8.077 0.98813 5.4681e-005 3.8183 0.011927 0.00010506 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5477 0.56207 0.17193 0.019934 16.266 0.12361 0.00016104 0.76655 0.0093057 0.0103 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16411 0.95471 0.92352 0.0013961 0.9956 0.52546 0.0018809 0.42862 2.2171 2.2166 16.0061 144.9311 0.00015267 -85.6599 0.97395
8.078 0.98813 5.4681e-005 3.8183 0.011927 0.00010507 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5477 0.56212 0.17194 0.019935 16.2689 0.12362 0.00016105 0.76654 0.009306 0.0103 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16412 0.9548 0.92355 0.0013961 0.99561 0.52562 0.0018809 0.42863 2.2174 2.2169 16.006 144.9312 0.00015262 -85.6599 0.97495
8.079 0.98813 5.4681e-005 3.8183 0.011926 0.00010508 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5478 0.56216 0.17196 0.019936 16.2719 0.12362 0.00016106 0.76654 0.0093064 0.010301 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16412 0.95489 0.92359 0.0013961 0.99562 0.52579 0.0018809 0.42864 2.2177 2.2173 16.006 144.9312 0.00015257 -85.6599 0.97595
8.08 0.98813 5.4681e-005 3.8183 0.011926 0.0001051 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5479 0.56221 0.17197 0.019937 16.2749 0.12363 0.00016107 0.76653 0.0093068 0.010301 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16412 0.95498 0.92362 0.0013961 0.99563 0.52596 0.0018809 0.42866 2.218 2.2176 16.006 144.9312 0.00015251 -85.66 0.97695
8.081 0.98813 5.4681e-005 3.8183 0.011926 0.00010511 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.548 0.56225 0.17198 0.019938 16.2779 0.12364 0.00016108 0.76653 0.0093072 0.010301 0.0013844 0.98697 0.99172 2.9849e-006 1.194e-005 0.16412 0.95507 0.92365 0.0013961 0.99564 0.52612 0.0018809 0.42867 2.2184 2.2179 16.0059 144.9312 0.00015246 -85.66 0.97795
8.082 0.98813 5.4681e-005 3.8183 0.011926 0.00010512 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5481 0.5623 0.172 0.019939 16.2808 0.12364 0.00016109 0.76652 0.0093076 0.010302 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16413 0.95515 0.92369 0.0013961 0.99565 0.52629 0.0018809 0.42868 2.2187 2.2183 16.0059 144.9312 0.00015241 -85.66 0.97895
8.083 0.98813 5.4681e-005 3.8183 0.011926 0.00010513 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5482 0.56234 0.17201 0.01994 16.2838 0.12365 0.0001611 0.76651 0.009308 0.010302 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16413 0.95524 0.92372 0.0013961 0.99566 0.52645 0.0018809 0.4287 2.219 2.2186 16.0059 144.9313 0.00015236 -85.66 0.97995
8.084 0.98813 5.4681e-005 3.8183 0.011926 0.00010515 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5483 0.56239 0.17202 0.019941 16.2868 0.12366 0.00016111 0.76651 0.0093084 0.010303 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16413 0.95533 0.92375 0.0013961 0.99567 0.52662 0.0018809 0.42871 2.2194 2.2189 16.0058 144.9313 0.00015231 -85.6601 0.98095
8.085 0.98813 5.4681e-005 3.8183 0.011926 0.00010516 0.0011724 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5483 0.56243 0.17204 0.019942 16.2897 0.12366 0.00016112 0.7665 0.0093088 0.010303 0.0013844 0.98697 0.99172 2.9849e-006 1.1939e-005 0.16414 0.95542 0.92378 0.0013961 0.99568 0.52678 0.0018809 0.42872 2.2197 2.2193 16.0058 144.9313 0.00015226 -85.6601 0.98195
8.086 0.98813 5.4681e-005 3.8183 0.011926 0.00010517 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5484 0.56248 0.17205 0.019944 16.2927 0.12367 0.00016113 0.76649 0.0093092 0.010303 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16414 0.95551 0.92382 0.0013961 0.99569 0.52695 0.0018809 0.42873 2.22 2.2196 16.0058 144.9313 0.00015221 -85.6601 0.98295
8.087 0.98813 5.4681e-005 3.8183 0.011926 0.00010519 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5485 0.56252 0.17207 0.019945 16.2957 0.12368 0.00016114 0.76649 0.0093095 0.010304 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16414 0.9556 0.92385 0.0013961 0.9957 0.52711 0.0018809 0.42875 2.2203 2.2199 16.0057 144.9314 0.00015216 -85.6601 0.98395
8.088 0.98813 5.4681e-005 3.8183 0.011926 0.0001052 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5486 0.56257 0.17208 0.019946 16.2986 0.12368 0.00016115 0.76648 0.0093099 0.010304 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16415 0.95568 0.92388 0.0013961 0.99571 0.52727 0.0018809 0.42876 2.2207 2.2202 16.0057 144.9314 0.00015211 -85.6601 0.98495
8.089 0.98813 5.468e-005 3.8183 0.011926 0.00010521 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5487 0.56261 0.17209 0.019947 16.3016 0.12369 0.00016116 0.76647 0.0093103 0.010305 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16415 0.95577 0.92391 0.0013961 0.99571 0.52744 0.0018809 0.42877 2.221 2.2206 16.0057 144.9314 0.00015206 -85.6602 0.98595
8.09 0.98813 5.468e-005 3.8183 0.011926 0.00010522 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5488 0.56266 0.17211 0.019948 16.3046 0.1237 0.00016117 0.76647 0.0093107 0.010305 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16415 0.95586 0.92395 0.0013961 0.99572 0.5276 0.0018809 0.42878 2.2213 2.2209 16.0056 144.9314 0.00015201 -85.6602 0.98695
8.091 0.98813 5.468e-005 3.8183 0.011926 0.00010524 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5489 0.5627 0.17212 0.019949 16.3076 0.1237 0.00016118 0.76646 0.0093111 0.010305 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16415 0.95594 0.92398 0.0013961 0.99573 0.52777 0.0018809 0.4288 2.2216 2.2212 16.0056 144.9314 0.00015196 -85.6602 0.98795
8.092 0.98813 5.468e-005 3.8183 0.011926 0.00010525 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5489 0.56275 0.17213 0.01995 16.3105 0.12371 0.00016119 0.76645 0.0093115 0.010306 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16416 0.95603 0.92401 0.0013961 0.99574 0.52793 0.0018809 0.42881 2.222 2.2215 16.0056 144.9315 0.00015191 -85.6602 0.98895
8.093 0.98813 5.468e-005 3.8183 0.011926 0.00010526 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.549 0.56279 0.17215 0.019951 16.3135 0.12372 0.0001612 0.76645 0.0093119 0.010306 0.0013844 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16416 0.95612 0.92404 0.0013961 0.99575 0.5281 0.0018809 0.42882 2.2223 2.2219 16.0055 144.9315 0.00015186 -85.6602 0.98995
8.094 0.98813 5.468e-005 3.8183 0.011926 0.00010528 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5491 0.56284 0.17216 0.019952 16.3165 0.12372 0.00016121 0.76644 0.0093123 0.010307 0.0013843 0.98697 0.99172 2.9848e-006 1.1939e-005 0.16416 0.9562 0.92407 0.0013961 0.99576 0.52826 0.0018809 0.42883 2.2226 2.2222 16.0055 144.9315 0.00015181 -85.6603 0.99095
8.095 0.98813 5.468e-005 3.8183 0.011926 0.00010529 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5492 0.56288 0.17217 0.019954 16.3195 0.12373 0.00016122 0.76643 0.0093126 0.010307 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16417 0.95629 0.9241 0.0013961 0.99577 0.52843 0.0018809 0.42885 2.2229 2.2225 16.0055 144.9315 0.00015176 -85.6603 0.99195
8.096 0.98813 5.468e-005 3.8183 0.011926 0.0001053 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5493 0.56293 0.17219 0.019955 16.3224 0.12374 0.00016123 0.76643 0.009313 0.010308 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16417 0.95637 0.92414 0.0013961 0.99578 0.52859 0.0018809 0.42886 2.2233 2.2228 16.0054 144.9315 0.00015172 -85.6603 0.99295
8.097 0.98813 5.468e-005 3.8183 0.011926 0.00010531 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5494 0.56297 0.1722 0.019956 16.3254 0.12374 0.00016124 0.76642 0.0093134 0.010308 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16417 0.95646 0.92417 0.0013961 0.99579 0.52875 0.0018809 0.42887 2.2236 2.2232 16.0054 144.9316 0.00015167 -85.6603 0.99395
8.098 0.98813 5.468e-005 3.8183 0.011926 0.00010533 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5495 0.56302 0.17221 0.019957 16.3284 0.12375 0.00016125 0.76641 0.0093138 0.010308 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16418 0.95654 0.9242 0.0013961 0.9958 0.52892 0.0018809 0.42889 2.2239 2.2235 16.0053 144.9316 0.00015162 -85.6603 0.99495
8.099 0.98813 5.468e-005 3.8183 0.011926 0.00010534 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5495 0.56306 0.17223 0.019958 16.3314 0.12375 0.00016126 0.76641 0.0093142 0.010309 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16418 0.95663 0.92423 0.0013961 0.99581 0.52908 0.0018809 0.4289 2.2242 2.2238 16.0053 144.9316 0.00015157 -85.6604 0.99595
8.1 0.98813 5.468e-005 3.8183 0.011926 0.00010535 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5496 0.56311 0.17224 0.019959 16.3343 0.12376 0.00016127 0.7664 0.0093146 0.010309 0.0013843 0.98697 0.99172 2.9847e-006 1.1939e-005 0.16418 0.95671 0.92426 0.001396 0.99582 0.52925 0.0018809 0.42891 2.2245 2.2241 16.0053 144.9316 0.00015152 -85.6593 0.99695
8.101 0.98813 5.468e-005 3.8183 0.011926 0.00010537 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5497 0.56315 0.17225 0.01996 16.3373 0.12377 0.00016128 0.76639 0.009315 0.01031 0.0064769 0.98322 0.99099 1.4526e-005 5.3364e-005 0.16418 0.95674 0.92429 0.0027739 0.99581 0.52939 0.0023959 0.42887 2.2249 2.2244 16.0052 144.9316 0.00015148 -76.1571 0.99795
8.102 0.98813 5.4679e-005 3.8183 0.011926 0.00010538 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5498 0.5632 0.17227 0.019961 16.3403 0.12377 0.00016129 0.76639 0.0093153 0.01031 0.026234 0.9717 0.98766 6.602e-005 0.00022964 0.16419 0.95656 0.92432 0.0053019 0.99576 0.52951 0.0033368 0.42875 2.2252 2.2248 16.0052 144.9316 0.00015147 -67.1434 0.99895
8.103 0.98813 5.4679e-005 3.8183 0.011926 0.00010539 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5499 0.56324 0.17228 0.019962 16.3433 0.12378 0.0001613 0.76638 0.0093157 0.01031 0.094919 0.9472 0.97732 0.00028456 0.0009136 0.16419 0.95582 0.92435 0.0092494 0.9955 0.52962 0.0044256 0.42859 2.2255 2.2251 16.0051 144.9316 0.00015147 -58.0116 0.99995
8.104 0.98813 5.4679e-005 3.8183 0.011926 0.0001054 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.55 0.56329 0.1723 0.019963 16.3462 0.12379 0.00016131 0.76637 0.0093161 0.010311 0.48858 0.85611 0.93869 0.0021831 0.0054838 0.16419 0.95382 0.92438 0.015757 0.99138 0.52967 0.0056246 0.4284 2.2258 2.2254 16.0058 144.9316 0.00015151 -37.1877 0.1555
8.105 0.98813 5.4679e-005 3.8183 0.011926 0.00010542 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5501 0.56333 0.17231 0.019965 16.3492 0.12379 0.00016132 0.76637 0.0093165 0.010311 0.99964 0.0021578 0.71203 0.94373 0.99666 0.1642 0.92053 0.92131 0.33599 0.96397 0.51803 0.044552 0.4282 2.1678 0.9776 16.0097 144.9312 0.00024928 25.2483 0.0019412
8.106 0.98813 5.4679e-005 3.8183 0.011926 0.00010543 0.0011725 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5501 0.56337 0.17232 0.019966 16.3522 0.1238 0.00016133 0.76636 0.0093169 0.010312 0.99955 1.2919e-006 0.52805 0.99838 0.99962 0.1642 0.88064 0.90277 0.63018 0.93682 0.50352 0.1014 0.42799 1.9507 0.6242 16.0093 144.9298 0.0003687 22.4714 0.0029412
8.107 0.98814 5.4679e-005 3.8183 0.011926 0.00010544 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5502 0.56342 0.17234 0.019967 16.3552 0.12381 0.00016134 0.76635 0.0093173 0.010312 0.99924 -1.7322e-009 0.39184 0.99691 0.99914 0.1642 0.84281 0.87868 0.75939 0.91043 0.48953 0.14621 0.42779 1.7488 0.61105 16.009 144.928 0.00044724 17.632 0.0039412
8.108 0.98814 5.4679e-005 3.8183 0.011926 0.00010546 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5503 0.56346 0.17235 0.019968 16.3582 0.12381 0.00016135 0.76635 0.0093177 0.010312 0.9989 2.2068e-010 0.29101 0.99436 0.99843 0.16421 0.80733 0.85155 0.81607 0.88479 0.47614 0.18171 0.42758 1.5819 0.66103 16.0086 144.9261 0.00050754 14.2457 0.0049412
8.109 0.98814 5.4679e-005 3.8183 0.011926 0.00010547 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5504 0.56351 0.17236 0.019969 16.3611 0.12382 0.00016136 0.76634 0.0093181 0.010313 0.9986 -9.1268e-011 0.2163 0.99145 0.99763 0.16421 0.77416 0.82265 0.84109 0.85987 0.46336 0.21158 0.42738 1.45 0.7309 16.0083 144.9242 0.00055476 12.0042 0.0059412
8.11 0.98814 5.4679e-005 3.8183 0.011926 0.00010548 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5505 0.56355 0.17238 0.01997 16.3641 0.12383 0.00016137 0.76633 0.0093184 0.010313 0.99832 -7.5582e-011 0.16087 0.98837 0.9968 0.16421 0.74311 0.7929 0.85059 0.83566 0.45117 0.23765 0.42718 1.3495 0.80464 16.0079 144.9224 0.00059144 10.333 0.0069412
8.111 0.98814 5.4679e-005 3.8183 0.011926 0.00010549 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5506 0.5636 0.17239 0.019971 16.3671 0.12383 0.00016138 0.76633 0.0093188 0.010314 0.99805 -4.2269e-010 0.11973 0.98508 0.9959 0.16421 0.71399 0.76298 0.85168 0.81213 0.43953 0.26083 0.42697 1.2752 0.87375 16.0076 144.9207 0.00061968 8.9313 0.0079412
8.112 0.98814 5.4679e-005 3.8183 0.011926 0.00010551 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5507 0.56364 0.1724 0.019972 16.3701 0.12384 0.00016139 0.76632 0.0093192 0.010314 0.99776 -2.7277e-012 0.089164 0.98145 0.99489 0.16422 0.68668 0.73339 0.8478 0.78927 0.42844 0.28162 0.42677 1.2222 0.9336 16.0073 144.919 0.00064143 7.6592 0.0089412
8.113 0.98814 5.4679e-005 3.8183 0.011926 0.00010552 0.0011726 0.23373 0.00065931 0.23438 0.21629 0 0.032258 0.0389 0 1.5508 0.56369 0.17242 0.019973 16.373 0.12385 0.0001614 0.76631 0.0093196 0.010315 0.99744 1.0049e-010 0.066447 0.97734 0.99371 0.16422 0.66107 0.7045 0.84075 0.76705 0.41789 0.30034 0.42657 1.1856 0.98239 16.007 144.9174 0.00065835 6.4487 0.0099412
8.114 0.98814 5.4678e-005 3.8183 0.011926 0.00010553 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5508 0.56373 0.17243 0.019975 16.376 0.12385 0.00016141 0.76631 0.00932 0.010315 0.99709 -3.9379e-011 0.049554 0.97258 0.99233 0.16422 0.63709 0.67655 0.83149 0.74546 0.40788 0.31718 0.42637 1.1611 1.0204 16.0067 144.9158 0.0006718 5.263 0.010941
8.115 0.98814 5.4678e-005 3.8183 0.011926 0.00010555 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5509 0.56378 0.17244 0.019976 16.379 0.12386 0.00016142 0.7663 0.0093204 0.010315 0.99669 4.1807e-012 0.036986 0.967 0.99068 0.16423 0.61465 0.64974 0.82055 0.72449 0.39842 0.33232 0.42616 1.1454 1.0489 16.0064 144.9144 0.00068277 4.0796 0.011941
8.116 0.98814 5.4678e-005 3.8183 0.011926 0.00010556 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.551 0.56382 0.17246 0.019977 16.382 0.12387 0.00016143 0.76629 0.0093208 0.010316 0.99622 -5.0358e-012 0.027631 0.96041 0.98867 0.16423 0.59372 0.62416 0.8082 0.7041 0.38952 0.34589 0.42596 1.1358 1.0699 16.0061 144.913 0.00069196 2.882 0.012941
8.117 0.98814 5.4678e-005 3.8183 0.011926 0.00010557 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5511 0.56387 0.17247 0.019978 16.385 0.12387 0.00016144 0.76629 0.0093211 0.010316 0.99568 -5.9048e-014 0.020664 0.95255 0.98621 0.16423 0.57423 0.59993 0.79458 0.6843 0.3812 0.35798 0.42576 1.1305 1.0852 16.0059 144.9117 0.00069985 1.6551 0.013941
8.118 0.98814 5.4678e-005 3.8183 0.011926 0.00010558 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5512 0.56391 0.17248 0.019979 16.388 0.12388 0.00016145 0.76628 0.0093215 0.010317 0.99503 7.5132e-013 0.015472 0.9431 0.98318 0.16424 0.55615 0.5771 0.77971 0.66506 0.37346 0.36868 0.42555 1.1279 1.0964 16.0056 144.9105 0.00070674 0.3833 0.014941
8.119 0.98814 5.4678e-005 3.8183 0.011926 0.0001056 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5513 0.56396 0.1725 0.01998 16.3909 0.12389 0.00016146 0.76627 0.0093219 0.010317 0.99425 -9.7915e-013 0.011601 0.93165 0.97938 0.16424 0.53944 0.55576 0.76352 0.64637 0.36634 0.37805 0.42535 1.1272 1.1047 16.0053 144.9094 0.00071283 -0.95241 0.015941
8.12 0.98814 5.4678e-005 3.8183 0.011926 0.00010561 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5514 0.564 0.17251 0.019981 16.3939 0.12389 0.00016147 0.76627 0.0093223 0.010317 0.99327 8.363e-013 0.0087135 0.91765 0.97454 0.16424 0.5241 0.53597 0.74591 0.62821 0.35984 0.38615 0.42515 1.1278 1.1111 16.0051 144.9083 0.00071823 -2.3766 0.016941
8.121 0.98814 5.4678e-005 3.8183 0.011926 0.00010562 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5514 0.56405 0.17253 0.019982 16.3969 0.1239 0.00016148 0.76626 0.0093227 0.010318 0.99201 -1.7283e-012 0.0065583 0.90033 0.96829 0.16424 0.5101 0.5178 0.72668 0.61058 0.354 0.393 0.42495 1.1291 1.1162 16.0048 144.9073 0.000723 -3.9226 0.017941
8.122 0.98814 5.4678e-005 3.8183 0.011926 0.00010563 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5515 0.56409 0.17254 0.019983 16.3999 0.12391 0.00016149 0.76626 0.0093231 0.010318 0.99034 9.7168e-013 0.0049493 0.87863 0.96003 0.16425 0.49747 0.50137 0.70557 0.59346 0.34885 0.39862 0.42474 1.1309 1.1204 16.0046 144.9064 0.00072714 -5.6373 0.018941
8.123 0.98814 5.4678e-005 3.8183 0.011926 0.00010565 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5516 0.56414 0.17255 0.019984 16.4029 0.12391 0.0001615 0.76625 0.0093235 0.010319 0.98801 3.7377e-013 0.0037479 0.85098 0.94886 0.16425 0.48623 0.48677 0.68225 0.57684 0.34442 0.40301 0.42454 1.1331 1.124 16.0044 144.9055 0.00073066 -7.5869 0.019941
8.124 0.98814 5.4678e-005 3.8183 0.011926 0.00010566 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5517 0.56418 0.17257 0.019986 16.4059 0.12392 0.00016151 0.76624 0.0093238 0.010319 0.98454 -1.6362e-012 0.0028514 0.81512 0.93331 0.16425 0.47642 0.47415 0.65628 0.56073 0.34074 0.40616 0.42434 1.1354 1.1274 16.0041 144.9047 0.00073349 -9.8658 0.020941
8.125 0.98814 5.4678e-005 3.8183 0.011926 0.00010567 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5518 0.56423 0.17258 0.019987 16.4088 0.12393 0.00016152 0.76624 0.0093242 0.010319 0.97903 3.2207e-012 0.0021841 0.76773 0.91099 0.16426 0.4681 0.46367 0.62722 0.54514 0.33783 0.40803 0.42414 1.1379 1.1304 16.0039 144.904 0.00073557 -12.604 0.021941
8.126 0.98814 5.4677e-005 3.8183 0.011926 0.00010569 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5519 0.56427 0.17259 0.019988 16.4118 0.12393 0.00016153 0.76623 0.0093246 0.01032 0.96949 -6.8037e-013 0.00169 0.70406 0.87803 0.16426 0.46131 0.45546 0.59468 0.53009 0.33567 0.40863 0.42394 1.1405 1.1334 16.0037 144.9034 0.00073679 -15.9661 0.022941
8.127 0.98814 5.4677e-005 3.8183 0.011926 0.0001057 0.0011726 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.552 0.56432 0.17261 0.019989 16.4148 0.12394 0.00016154 0.76622 0.009325 0.01032 0.95154 4.018e-013 0.0013286 0.61796 0.82824 0.16426 0.45605 0.44959 0.55857 0.51569 0.33421 0.40799 0.42374 1.1431 1.1363 16.0036 144.9029 0.00073702 -20.1115 0.023941
8.128 0.98814 5.4677e-005 3.8183 0.011926 0.00010571 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.552 0.56436 0.17262 0.01999 16.4178 0.12395 0.00016155 0.76622 0.0093254 0.010321 0.91601 2.8781e-013 0.0010706 0.50382 0.75292 0.16426 0.45215 0.4459 0.5191 0.50219 0.33332 0.40624 0.42354 1.1457 1.1391 16.0034 144.9024 0.00073625 -25.0649 0.024941
8.129 0.98814 5.4677e-005 3.8183 0.011926 0.00010572 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5521 0.56441 0.17263 0.019991 16.4208 0.12395 0.00016156 0.76621 0.0093258 0.010321 0.84806 -1.2136e-013 0.00089326 0.36361 0.64351 0.16427 0.44935 0.44391 0.47618 0.49018 0.33283 0.40348 0.42334 1.1484 1.1418 16.0033 144.9021 0.00073462 -30.5066 0.025941
8.13 0.98814 5.4677e-005 3.8183 0.011926 0.00010574 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5522 0.56445 0.17265 0.019992 16.4238 0.12396 0.00016157 0.7662 0.0093262 0.010321 0.73845 2.3066e-014 0.00077566 0.21823 0.50067 0.16427 0.44731 0.44292 0.42847 0.48082 0.33261 0.39967 0.42314 1.1511 1.1446 16.0032 144.9018 0.00073249 -35.779 0.026941
8.131 0.98814 5.4677e-005 3.8183 0.011926 0.00010575 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5523 0.5645 0.17266 0.019993 16.4267 0.12397 0.00016158 0.7662 0.0093265 0.010322 0.60203 3.3236e-005 0.00070568 0.10302 0.34392 0.16427 0.44579 0.44256 0.37418 0.47528 0.33255 0.39452 0.42294 1.1538 1.1473 16.0031 144.9015 0.00073018 -40.3755 0.027941
8.132 0.98814 5.4677e-005 3.8183 0.011926 0.00010576 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5524 0.56454 0.17267 0.019994 16.4297 0.12397 0.00016159 0.76619 0.0093269 0.010322 0.46839 0.00051689 0.00084335 0.037436 0.20432 0.16428 0.44466 0.44303 0.31346 0.47354 0.33259 0.38764 0.42274 1.1564 1.15 16.0031 144.9013 0.0007278 -44.211 0.028941
8.133 0.98814 5.4677e-005 3.8183 0.011926 0.00010578 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5525 0.56459 0.17269 0.019995 16.4327 0.12398 0.0001616 0.76618 0.0093273 0.010323 0.35811 0.0013022 0.0012172 0.0111 0.10426 0.16428 0.44386 0.44462 0.24954 0.47424 0.33268 0.37869 0.42255 1.1591 1.1527 16.003 144.9012 0.00072537 -47.3717 0.029941
8.134 0.98814 5.4677e-005 3.8183 0.011926 0.00010579 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5526 0.56463 0.1727 0.019997 16.4357 0.12399 0.00016161 0.76618 0.0093277 0.010323 0.27602 0.0025004 0.001857 0.0034067 0.046397 0.16428 0.44336 0.44725 0.18792 0.47601 0.33281 0.36751 0.42236 1.1618 1.1554 16.003 144.9011 0.0007229 -49.9633 0.030941
8.135 0.98814 5.4677e-005 3.8183 0.011926 0.0001058 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5526 0.56468 0.17271 0.019998 16.4387 0.12399 0.00016162 0.76617 0.0093281 0.010324 0.21747 0.0041925 0.0027796 0.0015142 0.018989 0.16429 0.44312 0.45052 0.13417 0.47808 0.33295 0.35413 0.42217 1.1645 1.1581 16.003 144.901 0.00072041 -52.0949 0.031941
8.136 0.98814 5.4677e-005 3.8183 0.011925 0.00010581 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5527 0.56472 0.17273 0.019999 16.4417 0.124 0.00016163 0.76616 0.0093285 0.010324 0.17566 0.0064387 0.0039911 0.00095428 0.0080026 0.16429 0.44309 0.45407 0.091702 0.48016 0.33311 0.33874 0.42199 1.1672 1.1608 16.003 144.9009 0.0007179 -53.8756 0.032941
8.137 0.98814 5.4677e-005 3.8183 0.011925 0.00010583 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5528 0.56477 0.17274 0.02 16.4447 0.12401 0.00016164 0.76616 0.0093289 0.010324 0.14494 0.0092877 0.0054934 0.00069492 0.0040175 0.16429 0.44324 0.45772 0.061111 0.48215 0.33327 0.32161 0.42181 1.1699 1.1635 16.003 144.9009 0.00071538 -55.4037 0.033941
8.138 0.98814 5.4676e-005 3.8183 0.011925 0.00010584 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5529 0.56481 0.17276 0.020001 16.4477 0.12401 0.00016165 0.76615 0.0093292 0.010325 0.12148 0.012789 0.0072901 0.0005347 0.0025324 0.16429 0.44355 0.46136 0.04079 0.48403 0.33343 0.30305 0.42163 1.1725 1.1662 16.003 144.9008 0.00071285 -56.7587 0.034941
8.139 0.98814 5.4676e-005 3.8183 0.011925 0.00010585 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.553 0.56486 0.17277 0.020002 16.4506 0.12402 0.00016166 0.76614 0.0093296 0.010325 0.1029 0.017002 0.0093896 0.00042356 0.0018574 0.1643 0.44399 0.46498 0.028161 0.4858 0.3336 0.28333 0.42145 1.1752 1.1689 16.003 144.9008 0.00071031 -57.9984 0.035941
8.14 0.98814 5.4676e-005 3.8183 0.011925 0.00010587 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5531 0.5649 0.17278 0.020003 16.4536 0.12402 0.00016167 0.76614 0.00933 0.010326 0.087749 0.022003 0.011806 0.00034162 0.0014573 0.1643 0.44456 0.46857 0.020665 0.48747 0.33376 0.26275 0.42128 1.1779 1.1716 16.003 144.9008 0.00070776 -59.1609 0.036941
8.141 0.98814 5.4676e-005 3.8183 0.011925 0.00010588 0.0011727 0.23373 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5532 0.56495 0.1728 0.020004 16.4566 0.12403 0.00016168 0.76613 0.0093304 0.010326 0.075158 0.027883 0.01456 0.00027942 0.0011753 0.1643 0.44523 0.47212 0.016277 0.48906 0.33393 0.24156 0.42111 1.1806 1.1743 16.0031 144.9007 0.00070521 -60.2694 0.037941
8.142 0.98814 5.4676e-005 3.8183 0.011925 0.00010589 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5532 0.56499 0.17281 0.020005 16.4596 0.12404 0.00016169 0.76612 0.0093308 0.010326 0.064575 0.034749 0.017674 0.00022964 0.00096076 0.16431 0.446 0.47563 0.013623 0.49056 0.3341 0.22004 0.42094 1.1832 1.177 16.0031 144.9007 0.00070266 -61.3372 0.038941
8.143 0.98814 5.4676e-005 3.8183 0.011925 0.0001059 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5533 0.56503 0.17282 0.020006 16.4626 0.12404 0.0001617 0.76612 0.0093312 0.010327 0.055624 0.042721 0.021175 0.00019059 0.00079227 0.16431 0.44687 0.4791 0.011882 0.49201 0.33427 0.19848 0.42077 1.1859 1.1797 16.0031 144.9007 0.0007001 -62.3715 0.039941
8.144 0.98814 5.4676e-005 3.8183 0.011925 0.00010592 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5534 0.56508 0.17284 0.020008 16.4656 0.12405 0.00016171 0.76611 0.0093315 0.010327 0.048027 0.051923 0.025092 0.00015889 0.00065789 0.16431 0.44781 0.48254 0.010615 0.49339 0.33444 0.17717 0.42061 1.1886 1.1824 16.0032 144.9007 0.00069754 -63.376 0.040941
8.145 0.98814 5.4676e-005 3.8183 0.011925 0.00010593 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5535 0.56512 0.17285 0.020009 16.4686 0.12406 0.00016172 0.7661 0.0093319 0.010328 0.041564 0.062491 0.029458 0.00013324 0.00054963 0.16432 0.44883 0.48594 0.0096054 0.49473 0.3346 0.1564 0.42046 1.1912 1.1851 16.0032 144.9006 0.00069498 -64.3531 0.041941
8.146 0.98814 5.4676e-005 3.8183 0.011925 0.00010594 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5536 0.56517 0.17286 0.02001 16.4716 0.12406 0.00016173 0.7661 0.0093323 0.010328 0.036059 0.074558 0.034304 0.00011231 0.00046174 0.16432 0.44991 0.4893 0.0087541 0.49603 0.33477 0.13645 0.4203 1.1939 1.1877 16.0033 144.9006 0.00069242 -65.3039 0.042941
8.147 0.98814 5.4676e-005 3.8183 0.011925 0.00010596 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5537 0.56521 0.17288 0.020011 16.4746 0.12407 0.00016174 0.76609 0.0093327 0.010328 0.03136 0.08826 0.039667 9.5096e-005 0.00038993 0.16432 0.45105 0.49262 0.0080152 0.4973 0.33494 0.11759 0.42016 1.1966 1.1904 16.0033 144.9006 0.00068986 -66.2294 0.043941
8.148 0.98814 5.4676e-005 3.8183 0.011925 0.00010597 0.0011727 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5538 0.56526 0.17289 0.020012 16.4776 0.12408 0.00016175 0.76608 0.0093331 0.010329 0.027345 0.10373 0.045586 8.0896e-005 0.00033095 0.16432 0.45224 0.49591 0.0073645 0.49854 0.33511 0.10005 0.42001 1.1992 1.1931 16.0034 144.9005 0.00068731 -67.1301 0.044941
8.149 0.98814 5.4676e-005 3.8183 0.011925 0.00010598 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5538 0.5653 0.1729 0.020013 16.4806 0.12408 0.00016176 0.76608 0.0093335 0.010329 0.023909 0.12108 0.052103 6.916e-005 0.00028225 0.16433 0.45348 0.49915 0.0067873 0.49978 0.33528 0.084021 0.41987 1.2019 1.1958 16.0035 144.9005 0.00068475 -68.0063 0.045941
8.15 0.98814 5.4675e-005 3.8183 0.011925 0.00010599 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5539 0.56535 0.17292 0.020014 16.4835 0.12409 0.00016177 0.76607 0.0093338 0.01033 0.020964 0.14043 0.059262 5.9369e-005 0.00024188 0.16433 0.45476 0.50237 0.0062733 0.501 0.33545 0.069633 0.41974 1.2045 1.1984 16.0036 144.9005 0.00068219 -68.8581 0.046941
8.151 0.98814 5.4675e-005 3.8183 0.011925 0.00010601 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.554 0.56539 0.17293 0.020015 16.4865 0.1241 0.00016178 0.76606 0.0093342 0.01033 0.018438 0.16185 0.067115 5.1213e-005 0.00020825 0.16433 0.45608 0.50554 0.0058139 0.50222 0.33562 0.056961 0.41961 1.2072 1.2011 16.0036 144.9005 0.00067963 -69.6853 0.047941
8.152 0.98814 5.4675e-005 3.8183 0.011925 0.00010602 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5541 0.56544 0.17294 0.020016 16.4895 0.1241 0.00016179 0.76606 0.0093346 0.01033 0.016267 0.1854 0.075713 4.4363e-005 0.00018016 0.16434 0.45743 0.50869 0.0054024 0.50344 0.33579 0.046019 0.41948 1.2098 1.2038 16.0037 144.9004 0.00067708 -70.4876 0.048941
8.153 0.98814 5.4675e-005 3.8183 0.011925 0.00010603 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5542 0.56548 0.17296 0.020017 16.4925 0.12411 0.0001618 0.76605 0.009335 0.010331 0.0144 0.21111 0.085113 3.8617e-005 0.0001566 0.16434 0.4588 0.51179 0.0050333 0.50467 0.33596 0.036763 0.41936 1.2125 1.2065 16.0038 144.9004 0.00067453 -71.2644 0.049941
8.154 0.98814 5.4675e-005 3.8183 0.011925 0.00010605 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5543 0.56553 0.17297 0.020019 16.4955 0.12412 0.00016181 0.76605 0.0093354 0.010331 0.012793 0.23894 0.095373 3.3795e-005 0.0001368 0.16434 0.4602 0.51486 0.0047017 0.50591 0.33613 0.029094 0.41924 1.2151 1.2091 16.0039 144.9004 0.00067199 -72.015 0.050941
8.155 0.98814 5.4675e-005 3.8183 0.011925 0.00010606 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5544 0.56557 0.17298 0.02002 16.4985 0.12412 0.00016182 0.76604 0.0093358 0.010332 0.011408 0.26882 0.10655 2.9686e-005 0.00012009 0.16434 0.46162 0.5179 0.0044036 0.50717 0.33631 0.022875 0.41913 1.2178 1.2118 16.004 144.9003 0.00066944 -72.7386 0.051941
8.156 0.98814 5.4675e-005 3.8183 0.011925 0.00010607 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5544 0.56562 0.173 0.020021 16.5015 0.12413 0.00016183 0.76603 0.0093361 0.010332 0.010213 0.30063 0.1187 2.6218e-005 0.00010596 0.16435 0.46306 0.5209 0.0041354 0.50846 0.33648 0.017938 0.41903 1.2204 1.2144 16.0041 144.9003 0.00066691 -73.4344 0.052941
8.157 0.98814 5.4675e-005 3.8183 0.011925 0.00010608 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5545 0.56566 0.17301 0.020022 16.5045 0.12414 0.00016184 0.76603 0.0093365 0.010333 0.0091824 0.33418 0.13186 2.3284e-005 9.3991e-005 0.16435 0.46451 0.52387 0.0038941 0.50976 0.33666 0.014101 0.41893 1.2231 1.2171 16.0042 144.9003 0.00066437 -74.1015 0.053941
8.158 0.98814 5.4675e-005 3.8183 0.011925 0.0001061 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5546 0.56571 0.17303 0.020023 16.5075 0.12414 0.00016185 0.76602 0.0093369 0.010333 0.0082914 0.36922 0.14608 2.0777e-005 8.3822e-005 0.16435 0.46597 0.52681 0.0036771 0.5111 0.33683 0.011177 0.41883 1.2257 1.2197 16.0043 144.9003 0.00066185 -74.7391 0.054941
8.159 0.98814 5.4675e-005 3.8183 0.011925 0.00010611 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5547 0.56575 0.17304 0.020024 16.5105 0.12415 0.00016186 0.76601 0.0093373 0.010333 0.007521 0.40547 0.16136 1.865e-005 7.5163e-005 0.16436 0.46745 0.52972 0.0034819 0.51247 0.33701 0.0089914 0.41874 1.2283 1.2224 16.0044 144.9002 0.00065933 -75.3465 0.055941
8.16 0.98814 5.4675e-005 3.8183 0.011925 0.00010612 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5548 0.5658 0.17305 0.020025 16.5135 0.12416 0.00016187 0.76601 0.0093377 0.010334 0.0068539 0.44257 0.17772 1.6829e-005 6.7775e-005 0.16436 0.46894 0.53259 0.0033065 0.51387 0.33719 0.0073826 0.41866 1.231 1.225 16.0045 144.9002 0.00065681 -75.9233 0.056941
8.161 0.98814 5.4675e-005 3.8183 0.011925 0.00010613 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5549 0.56584 0.17307 0.020026 16.5165 0.12416 0.00016188 0.766 0.0093381 0.010334 0.0062757 0.48015 0.19512 1.5264e-005 6.1456e-005 0.16436 0.47043 0.53544 0.0031488 0.51531 0.33738 0.006213 0.41858 1.2336 1.2277 16.0046 144.9002 0.0006543 -76.4692 0.057941
8.162 0.98814 5.4674e-005 3.8183 0.011925 0.00010615 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.555 0.56589 0.17308 0.020027 16.5195 0.12417 0.00016189 0.76599 0.0093384 0.010335 0.0057743 0.51781 0.21351 1.3931e-005 5.6039e-005 0.16437 0.47193 0.53825 0.0030071 0.51678 0.33756 0.0053686 0.4185 1.2362 1.2303 16.0047 144.9002 0.0006518 -76.984 0.058941
8.163 0.98814 5.4674e-005 3.8183 0.011925 0.00010616 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.555 0.56593 0.17309 0.020028 16.5225 0.12418 0.0001619 0.76599 0.0093388 0.010335 0.0053386 0.55515 0.23283 1.2784e-005 5.1386e-005 0.16437 0.47343 0.54103 0.0028799 0.51829 0.33774 0.0047592 0.41843 1.2389 1.233 16.0048 144.9001 0.00064931 -77.4679 0.059941
8.164 0.98814 5.4674e-005 3.8183 0.011925 0.00010617 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5551 0.56598 0.17311 0.020029 16.5255 0.12418 0.00016191 0.76598 0.0093392 0.010335 0.004959 0.59176 0.25299 1.1785e-005 4.7377e-005 0.16437 0.47494 0.54378 0.0027656 0.51985 0.33793 0.0043163 0.41837 1.2415 1.2356 16.0049 144.9001 0.00064683 -77.9214 0.060941
8.165 0.98814 5.4674e-005 3.8183 0.011925 0.00010619 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5552 0.56602 0.17312 0.020031 16.5285 0.12419 0.00016192 0.76597 0.0093396 0.010336 0.0046289 0.62729 0.27387 1.0934e-005 4.3916e-005 0.16437 0.47645 0.5465 0.0026631 0.52144 0.33812 0.0039893 0.4183 1.2441 1.2383 16.005 144.9001 0.00064435 -78.345 0.061941
8.166 0.98814 5.4674e-005 3.8183 0.011925 0.0001062 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5553 0.56607 0.17313 0.020032 16.5315 0.1242 0.00016193 0.76597 0.00934 0.010336 0.0043404 0.66139 0.29535 1.0193e-005 4.0921e-005 0.16438 0.47796 0.5492 0.0025711 0.52307 0.33831 0.0037423 0.41824 1.2467 1.2409 16.0051 144.9001 0.00064189 -78.7397 0.062941
8.167 0.98814 5.4674e-005 3.8183 0.011925 0.00010621 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5554 0.56611 0.17315 0.020033 16.5345 0.1242 0.00016194 0.76596 0.0093404 0.010337 0.0040881 0.6938 0.31731 9.548e-006 3.8323e-005 0.16438 0.47948 0.55186 0.0024885 0.52474 0.3385 0.0035506 0.41819 1.2493 1.2435 16.0052 144.9001 0.00063943 -79.1063 0.063941
8.168 0.98814 5.4674e-005 3.8183 0.011925 0.00010622 0.0011728 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5555 0.56616 0.17316 0.020034 16.5375 0.12421 0.00016195 0.76595 0.0093407 0.010337 0.0038673 0.72428 0.33961 8.9884e-006 3.6063e-005 0.16438 0.48099 0.5545 0.0024144 0.52645 0.33869 0.0033976 0.41814 1.2519 1.2461 16.0054 144.9 0.00063699 -79.4461 0.064941
8.169 0.98814 5.4674e-005 3.8183 0.011925 0.00010624 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5556 0.5662 0.17317 0.020035 16.5405 0.12421 0.00016196 0.76595 0.0093411 0.010337 0.0036734 0.75268 0.36213 8.5004e-006 3.4093e-005 0.16439 0.48251 0.55711 0.0023479 0.52819 0.33889 0.003272 0.41809 1.2545 1.2488 16.0055 144.9 0.00063455 -79.7603 0.065941
8.17 0.98814 5.4674e-005 3.8183 0.011925 0.00010625 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5556 0.56625 0.17319 0.020036 16.5435 0.12422 0.00016197 0.76594 0.0093415 0.010338 0.0035028 0.77889 0.38473 8.0726e-006 3.237e-005 0.16439 0.48402 0.55969 0.0022881 0.52997 0.33908 0.0031664 0.41805 1.2571 1.2514 16.0056 144.9 0.00063213 -80.0503 0.066941
8.171 0.98814 5.4674e-005 3.8183 0.011925 0.00010626 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5557 0.56629 0.1732 0.020037 16.5465 0.12423 0.00016198 0.76593 0.0093419 0.010338 0.0033527 0.80287 0.40731 7.6979e-006 3.0861e-005 0.16439 0.48553 0.56224 0.0022345 0.53178 0.33928 0.0030758 0.418 1.2597 1.254 16.0057 144.9 0.00062971 -80.3175 0.067941
8.172 0.98814 5.4674e-005 3.8183 0.011925 0.00010628 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5558 0.56634 0.17321 0.020038 16.5495 0.12423 0.00016199 0.76593 0.0093423 0.010339 0.0032201 0.82463 0.42975 7.3692e-006 2.9535e-005 0.16439 0.48704 0.56477 0.0021863 0.53362 0.33948 0.002997 0.41796 1.2623 1.2566 16.0058 144.9 0.00062731 -80.5632 0.068941
8.173 0.98814 5.4674e-005 3.8183 0.011925 0.00010629 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5559 0.56638 0.17323 0.020039 16.5525 0.12424 0.000162 0.76592 0.0093427 0.010339 0.0031028 0.84422 0.45195 7.0794e-006 2.8367e-005 0.1644 0.48855 0.56727 0.0021429 0.53549 0.33967 0.002928 0.41793 1.2649 1.2592 16.006 144.9 0.00062492 -80.789 0.069941
8.174 0.98814 5.4674e-005 3.8183 0.011925 0.0001063 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.556 0.56642 0.17324 0.02004 16.5555 0.12425 0.00016201 0.76591 0.009343 0.010339 0.0029988 0.86173 0.47384 6.823e-006 2.7336e-005 0.1644 0.49006 0.56974 0.0021039 0.53738 0.33987 0.0028669 0.41789 1.2675 1.2619 16.0061 144.9 0.00062254 -80.9963 0.070941
8.175 0.98814 5.4673e-005 3.8183 0.011925 0.00010631 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5561 0.56647 0.17325 0.020042 16.5585 0.12425 0.00016202 0.76591 0.0093434 0.01034 0.0029064 0.87728 0.49534 6.5961e-006 2.6424e-005 0.1644 0.49156 0.57219 0.0020687 0.5393 0.34007 0.0028127 0.41786 1.2701 1.2645 16.0062 144.8999 0.00062018 -81.1863 0.071941
8.176 0.98814 5.4673e-005 3.8183 0.011925 0.00010633 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5562 0.56651 0.17327 0.020043 16.5615 0.12426 0.00016203 0.7659 0.0093438 0.01034 0.0028243 0.89099 0.51637 6.3954e-006 2.5615e-005 0.16441 0.49306 0.57462 0.002037 0.54125 0.34028 0.0027643 0.41783 1.2727 1.2671 16.0063 144.8999 0.00061782 -81.3605 0.072941
8.177 0.98814 5.4673e-005 3.8183 0.011925 0.00010634 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5562 0.56656 0.17328 0.020044 16.5645 0.12427 0.00016204 0.76589 0.0093442 0.010341 0.002751 0.90302 0.53691 6.2167e-006 2.4895e-005 0.16441 0.49456 0.57702 0.0020084 0.54321 0.34048 0.002721 0.4178 1.2753 1.2697 16.0064 144.8999 0.00061548 -81.5202 0.073941
8.178 0.98814 5.4673e-005 3.8183 0.011925 0.00010635 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5563 0.5666 0.1733 0.020045 16.5675 0.12427 0.00016205 0.76589 0.0093446 0.010341 0.0026853 0.91352 0.55689 6.0568e-006 2.4254e-005 0.16441 0.49606 0.57939 0.0019826 0.54519 0.34068 0.0026821 0.41777 1.2779 1.2723 16.0066 144.8999 0.00061315 -81.6664 0.074941
8.179 0.98814 5.4673e-005 3.8183 0.011925 0.00010637 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5564 0.56665 0.17331 0.020046 16.5705 0.12428 0.00016206 0.76588 0.009345 0.010341 0.0026266 0.92264 0.57628 5.9139e-006 2.3681e-005 0.16442 0.49755 0.58174 0.0019592 0.54719 0.34089 0.0026472 0.41775 1.2805 1.2749 16.0067 144.8999 0.00061083 -81.8005 0.075941
8.18 0.98814 5.4673e-005 3.8183 0.011925 0.00010638 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5565 0.56669 0.17332 0.020047 16.5735 0.12429 0.00016207 0.76588 0.0093453 0.010342 0.002574 0.93053 0.59507 5.7865e-006 2.3167e-005 0.16442 0.49904 0.58407 0.001938 0.5492 0.34109 0.0026158 0.41772 1.283 1.2775 16.0068 144.8999 0.00060852 -81.9233 0.076941
8.181 0.98814 5.4673e-005 3.8183 0.011925 0.00010639 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5566 0.56674 0.17334 0.020048 16.5765 0.12429 0.00016208 0.76587 0.0093457 0.010342 0.0025268 0.93733 0.61324 5.673e-006 2.2706e-005 0.16442 0.50052 0.58637 0.0019187 0.55122 0.34129 0.0025874 0.4177 1.2856 1.28 16.0069 144.8999 0.00060623 -82.036 0.077941
8.182 0.98814 5.4673e-005 3.8183 0.011925 0.0001064 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5567 0.56678 0.17335 0.020049 16.5795 0.1243 0.00016209 0.76586 0.0093461 0.010343 0.0024838 0.94317 0.63076 5.5695e-006 2.2291e-005 0.16442 0.50201 0.58865 0.0019013 0.55325 0.3415 0.0025617 0.41768 1.2882 1.2826 16.007 144.8999 0.00060395 -82.1394 0.078941
8.183 0.98814 5.4673e-005 3.8183 0.011925 0.00010642 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5568 0.56683 0.17336 0.02005 16.5825 0.12431 0.0001621 0.76586 0.0093465 0.010343 0.0024449 0.94818 0.64765 5.4755e-006 2.1917e-005 0.16443 0.50348 0.59091 0.0018854 0.5553 0.34171 0.0025384 0.41766 1.2908 1.2852 16.0072 144.8999 0.00060168 -82.2345 0.079941
8.184 0.98814 5.4673e-005 3.8183 0.011925 0.00010643 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5568 0.56687 0.17338 0.020051 16.5855 0.12431 0.00016211 0.76585 0.0093469 0.010343 0.0024098 0.95246 0.66389 5.3906e-006 2.1578e-005 0.16443 0.50496 0.59315 0.0018709 0.55735 0.34191 0.0025173 0.41764 1.2933 1.2878 16.0073 144.8999 0.00059942 -82.3219 0.080941
8.185 0.98814 5.4673e-005 3.8183 0.011925 0.00010644 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5569 0.56692 0.17339 0.020053 16.5885 0.12432 0.00016212 0.76584 0.0093472 0.010344 0.0023781 0.95611 0.6795 5.315e-006 2.1271e-005 0.16443 0.50643 0.59536 0.0018576 0.55941 0.34212 0.0024981 0.41762 1.2959 1.2904 16.0074 144.8999 0.00059718 -82.4024 0.081941
8.186 0.98814 5.4673e-005 3.8183 0.011925 0.00010646 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.557 0.56696 0.1734 0.020054 16.5915 0.12433 0.00016213 0.76584 0.0093476 0.010344 0.0023492 0.95922 0.69447 5.2454e-006 2.0991e-005 0.16444 0.5079 0.59755 0.0018454 0.56147 0.34233 0.0024806 0.4176 1.2984 1.2929 16.0075 144.8999 0.00059495 -82.4767 0.082941
8.187 0.98814 5.4672e-005 3.8183 0.011925 0.00010647 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5571 0.56701 0.17342 0.020055 16.5945 0.12433 0.00016214 0.76583 0.009348 0.010345 0.0023226 0.96187 0.70882 5.1814e-006 2.0736e-005 0.16444 0.50936 0.59972 0.0018343 0.56353 0.34254 0.0024646 0.41758 1.301 1.2955 16.0076 144.8999 0.00059273 -82.5453 0.083941
8.188 0.98814 5.4672e-005 3.8183 0.011925 0.00010648 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5572 0.56705 0.17343 0.020056 16.5975 0.12434 0.00016215 0.76582 0.0093484 0.010345 0.0022982 0.96413 0.72256 5.1229e-006 2.0502e-005 0.16444 0.51082 0.60187 0.001824 0.5656 0.34274 0.0024499 0.41757 1.3035 1.2981 16.0078 144.8999 0.00059053 -82.6089 0.084941
8.189 0.98814 5.4672e-005 3.8183 0.011925 0.00010649 0.0011729 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5573 0.5671 0.17344 0.020057 16.6005 0.12435 0.00016216 0.76582 0.0093488 0.010346 0.002276 0.96605 0.73571 5.0699e-006 2.0288e-005 0.16444 0.51228 0.60399 0.0018146 0.56768 0.34295 0.0024364 0.41755 1.3061 1.3007 16.0079 144.8999 0.00058833 -82.6679 0.085941
8.19 0.98814 5.4672e-005 3.8183 0.011925 0.00010651 0.001173 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5574 0.56714 0.17346 0.020058 16.6035 0.12435 0.00016217 0.76581 0.0093492 0.010346 0.0022555 0.96769 0.74827 5.021e-006 2.0091e-005 0.16445 0.51373 0.6061 0.0018058 0.56975 0.34316 0.002424 0.41753 1.3086 1.3032 16.008 144.8999 0.00058615 -82.7227 0.086941
8.191 0.98814 5.4672e-005 3.8183 0.011925 0.00010652 0.001173 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5574 0.56719 0.17347 0.020059 16.6065 0.12436 0.00016218 0.7658 0.0093495 0.010346 0.0022364 0.96909 0.76027 4.9755e-006 1.9909e-005 0.16445 0.51517 0.60819 0.0017977 0.57182 0.34337 0.0024125 0.41752 1.3112 1.3058 16.0081 144.8999 0.00058398 -82.7738 0.087941
8.192 0.98814 5.4672e-005 3.8183 0.011925 0.00010653 0.001173 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5575 0.56723 0.17348 0.02006 16.6095 0.12437 0.00016219 0.7658 0.0093499 0.010347 0.0022188 0.97028 0.77173 4.9336e-006 1.9741e-005 0.16445 0.51662 0.61025 0.0017902 0.57389 0.34358 0.0024019 0.41751 1.3137 1.3083 16.0082 144.8999 0.00058183 -82.8215 0.088941
8.193 0.98814 5.4672e-005 3.8183 0.011924 0.00010654 0.001173 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5576 0.56728 0.1735 0.020061 16.6125 0.12437 0.0001622 0.76579 0.0093503 0.010347 0.0022025 0.9713 0.78266 4.8948e-006 1.9585e-005 0.16446 0.51806 0.6123 0.0017831 0.57596 0.34379 0.002392 0.41749 1.3162 1.3109 16.0083 144.8999 0.00057968 -82.8662 0.089941
8.194 0.98814 5.4672e-005 3.8183 0.011924 0.00010656 0.001173 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5577 0.56732 0.17351 0.020062 16.6155 0.12438 0.00016221 0.76578 0.0093507 0.010348 0.0021873 0.97218 0.79308 4.8585e-006 1.9439e-005 0.16446 0.51949 0.61432 0.0017765 0.57803 0.344 0.0023829 0.41748 1.3188 1.3134 16.0085 144.8999 0.00057755 -82.9081 0.090941
8.195 0.98814 5.4672e-005 3.8183 0.011924 0.00010657 0.001173 0.23372 0.00065931 0.23438 0.21628 0 0.032258 0.0389 0 1.5578 0.56737 0.17352 0.020063 16.6186 0.12438 0.00016222 0.76578 0.0093511 0.010348 0.002173 0.97293 0.80301 4.8245e-006 1.9303e-005 0.16446 0.52092 0.61633 0.0017704 0.5801 0.34421 0.0023743 0.41747 1.3213 1.316 16.0086 144.8999 0.00057543 -82.9476 0.091941
8.196 0.98814 5.4672e-005 3.8183 0.011924 0.00010658 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5579 0.56741 0.17354 0.020065 16.6216 0.12439 0.00016223 0.76577 0.0093514 0.010348 0.0021596 0.97358 0.81246 4.7927e-006 1.9176e-005 0.16447 0.52235 0.61832 0.0017646 0.58217 0.34442 0.0023662 0.41745 1.3238 1.3185 16.0087 144.8999 0.00057332 -82.9849 0.092941
8.197 0.98814 5.4672e-005 3.8183 0.011924 0.0001066 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.558 0.56746 0.17355 0.020066 16.6246 0.1244 0.00016224 0.76576 0.0093518 0.010349 0.0021471 0.97415 0.82147 4.7629e-006 1.9056e-005 0.16447 0.52377 0.62028 0.0017591 0.58423 0.34463 0.0023587 0.41744 1.3264 1.3211 16.0088 144.8999 0.00057123 -83.0202 0.093941
8.198 0.98814 5.4672e-005 3.8183 0.011924 0.00010661 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.558 0.5675 0.17356 0.020067 16.6276 0.1244 0.00016225 0.76576 0.0093522 0.010349 0.0021353 0.97464 0.83003 4.7348e-006 1.8943e-005 0.16447 0.52519 0.62223 0.001754 0.58629 0.34484 0.0023516 0.41743 1.3289 1.3236 16.0089 144.8999 0.00056915 -83.0536 0.094941
8.199 0.98814 5.4671e-005 3.8183 0.011924 0.00010662 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5581 0.56755 0.17358 0.020068 16.6306 0.12441 0.00016226 0.76575 0.0093526 0.01035 0.0021239 0.97507 0.83819 4.708e-006 1.8836e-005 0.16447 0.5266 0.62416 0.0017491 0.58834 0.34505 0.0023449 0.41742 1.3314 1.3261 16.009 144.8999 0.00056708 -83.0854 0.095941
8.2 0.98814 5.4671e-005 3.8183 0.011924 0.00010663 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5582 0.56759 0.17359 0.020069 16.6336 0.12442 0.00016227 0.76574 0.009353 0.01035 0.0021133 0.97545 0.84594 4.6827e-006 1.8735e-005 0.16448 0.52801 0.62608 0.0017444 0.59039 0.34526 0.0023385 0.41741 1.3339 1.3286 16.0091 144.8999 0.00056502 -83.1158 0.096941
8.201 0.98814 5.4671e-005 3.8183 0.011924 0.00010665 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5583 0.56763 0.17361 0.02007 16.6366 0.12442 0.00016228 0.76574 0.0093534 0.01035 0.0021032 0.97578 0.85331 4.6588e-006 1.8639e-005 0.16448 0.52942 0.62797 0.00174 0.59244 0.34547 0.0023324 0.4174 1.3364 1.3312 16.0092 144.8999 0.00056297 -83.1448 0.097941
8.202 0.98814 5.4671e-005 3.8183 0.011924 0.00010666 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5584 0.56768 0.17362 0.020071 16.6396 0.12443 0.00016229 0.76573 0.0093537 0.010351 0.0020936 0.97608 0.86032 4.6359e-006 1.8547e-005 0.16448 0.53082 0.62985 0.0017357 0.59448 0.34568 0.0023267 0.41739 1.3389 1.3337 16.0094 144.8999 0.00056093 -83.1726 0.098941
8.203 0.98814 5.4671e-005 3.8183 0.011924 0.00010667 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5585 0.56772 0.17363 0.020072 16.6426 0.12444 0.0001623 0.76573 0.0093541 0.010351 0.0020843 0.97635 0.86697 4.614e-006 1.8459e-005 0.16449 0.53222 0.63171 0.0017316 0.59652 0.34589 0.0023212 0.41738 1.3414 1.3362 16.0095 144.8999 0.00055891 -83.1993 0.099941
8.204 0.98814 5.4671e-005 3.8183 0.011924 0.00010669 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5586 0.56777 0.17365 0.020073 16.6456 0.12444 0.00016231 0.76572 0.0093545 0.010352 0.0020755 0.97659 0.8733 4.593e-006 1.8375e-005 0.16449 0.53361 0.63355 0.0017277 0.59855 0.3461 0.0023159 0.41737 1.3439 1.3387 16.0096 144.8999 0.00055689 -83.225 0.10094
8.205 0.98814 5.4671e-005 3.8183 0.011924 0.0001067 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5586 0.56781 0.17366 0.020074 16.6486 0.12445 0.00016232 0.76571 0.0093549 0.010352 0.0020669 0.97681 0.8793 4.5729e-006 1.8294e-005 0.16449 0.535 0.63538 0.001724 0.60058 0.34631 0.0023108 0.41736 1.3464 1.3412 16.0097 144.8999 0.00055489 -83.2498 0.10194
8.206 0.98814 5.4671e-005 3.8183 0.011924 0.00010671 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5587 0.56786 0.17367 0.020075 16.6517 0.12446 0.00016233 0.76571 0.0093553 0.010352 0.0020587 0.97701 0.88501 4.5535e-006 1.8217e-005 0.16449 0.53639 0.63719 0.0017203 0.6026 0.34652 0.0023059 0.41735 1.3489 1.3437 16.0098 144.8999 0.0005529 -83.2738 0.10294
8.207 0.98814 5.4671e-005 3.8183 0.011924 0.00010672 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5588 0.5679 0.17369 0.020077 16.6547 0.12446 0.00016234 0.7657 0.0093556 0.010353 0.0020508 0.97719 0.89042 4.5347e-006 1.8142e-005 0.1645 0.53777 0.63898 0.0017168 0.60461 0.34673 0.0023012 0.41734 1.3514 1.3462 16.0099 144.8999 0.00055093 -83.2971 0.10394
8.208 0.98814 5.4671e-005 3.8183 0.011924 0.00010674 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5589 0.56795 0.1737 0.020078 16.6577 0.12447 0.00016235 0.76569 0.009356 0.010353 0.0020431 0.97736 0.89556 4.5166e-006 1.8069e-005 0.1645 0.53914 0.64075 0.0017134 0.60662 0.34694 0.0022967 0.41733 1.3539 1.3488 16.01 144.8999 0.00054896 -83.3197 0.10494
8.209 0.98814 5.4671e-005 3.8183 0.011924 0.00010675 0.001173 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.559 0.56799 0.17371 0.020079 16.6607 0.12448 0.00016236 0.76569 0.0093564 0.010354 0.0020357 0.97751 0.90044 4.4991e-006 1.7999e-005 0.1645 0.54052 0.64251 0.0017101 0.60863 0.34716 0.0022923 0.41733 1.3564 1.3512 16.0101 144.8999 0.000547 -83.3416 0.10594
8.21 0.98814 5.4671e-005 3.8183 0.011924 0.00010676 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5591 0.56804 0.17373 0.02008 16.6637 0.12448 0.00016237 0.76568 0.0093568 0.010354 0.0020285 0.97766 0.90507 4.4821e-006 1.7931e-005 0.16451 0.54189 0.64426 0.0017069 0.61062 0.34737 0.002288 0.41732 1.3588 1.3537 16.0102 144.8999 0.00054506 -83.363 0.10694
8.211 0.98814 5.467e-005 3.8183 0.011924 0.00010678 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5592 0.56808 0.17374 0.020081 16.6667 0.12449 0.00016238 0.76567 0.0093572 0.010354 0.0020215 0.9778 0.90946 4.4656e-006 1.7865e-005 0.16451 0.54325 0.64598 0.0017038 0.61261 0.34758 0.0022839 0.41731 1.3613 1.3562 16.0103 144.8999 0.00054312 -83.3839 0.10794
8.212 0.98814 5.467e-005 3.8183 0.011924 0.00010679 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5592 0.56813 0.17375 0.020082 16.6697 0.1245 0.00016239 0.76567 0.0093575 0.010355 0.0020147 0.97793 0.91363 4.4495e-006 1.78e-005 0.16451 0.54461 0.6477 0.0017008 0.6146 0.34779 0.0022798 0.4173 1.3638 1.3587 16.0104 144.8999 0.0005412 -83.4043 0.10894
8.213 0.98814 5.467e-005 3.8183 0.011924 0.0001068 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5593 0.56817 0.17377 0.020083 16.6727 0.1245 0.0001624 0.76566 0.0093579 0.010355 0.002008 0.97805 0.91758 4.4338e-006 1.7737e-005 0.16452 0.54597 0.64939 0.0016978 0.61658 0.348 0.0022759 0.41729 1.3662 1.3612 16.0105 144.9 0.00053929 -83.4242 0.10994
8.214 0.98814 5.467e-005 3.8183 0.011924 0.00010681 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5594 0.56822 0.17378 0.020084 16.6758 0.12451 0.00016241 0.76565 0.0093583 0.010356 0.0020016 0.97817 0.92133 4.4185e-006 1.7676e-005 0.16452 0.54732 0.65108 0.0016949 0.61855 0.34821 0.002272 0.41729 1.3687 1.3637 16.0106 144.9 0.00053739 -83.4437 0.11094
8.215 0.98814 5.467e-005 3.8183 0.011924 0.00010683 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5595 0.56826 0.17379 0.020085 16.6788 0.12452 0.00016242 0.76565 0.0093587 0.010356 0.0019952 0.97829 0.92488 4.4035e-006 1.7616e-005 0.16452 0.54867 0.65274 0.0016921 0.62052 0.34842 0.0022683 0.41728 1.3712 1.3662 16.0107 144.9 0.0005355 -83.4629 0.11194
8.216 0.98814 5.467e-005 3.8183 0.011924 0.00010684 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5596 0.56831 0.17381 0.020086 16.6818 0.12452 0.00016243 0.76564 0.0093591 0.010356 0.001989 0.97839 0.92825 4.3889e-006 1.7558e-005 0.16452 0.55001 0.65439 0.0016893 0.62247 0.34864 0.0022646 0.41727 1.3736 1.3686 16.0108 144.9 0.00053362 -83.4817 0.11294
8.217 0.98814 5.467e-005 3.8183 0.011924 0.00010685 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5597 0.56835 0.17382 0.020087 16.6848 0.12453 0.00016244 0.76563 0.0093594 0.010357 0.0019829 0.9785 0.93145 4.3746e-006 1.75e-005 0.16453 0.55135 0.65603 0.0016865 0.62443 0.34885 0.002261 0.41727 1.3761 1.3711 16.0109 144.9 0.00053175 -83.5002 0.11394
8.218 0.98814 5.467e-005 3.8183 0.011924 0.00010687 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5598 0.5684 0.17383 0.020089 16.6878 0.12453 0.00016245 0.76563 0.0093598 0.010357 0.001977 0.9786 0.93448 4.3605e-006 1.7444e-005 0.16453 0.55269 0.65765 0.0016839 0.62637 0.34906 0.0022574 0.41726 1.3785 1.3736 16.011 144.9 0.00052989 -83.5184 0.11494
8.219 0.98814 5.467e-005 3.8183 0.011924 0.00010688 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5598 0.56844 0.17385 0.02009 16.6908 0.12454 0.00016246 0.76562 0.0093602 0.010358 0.0019711 0.9787 0.93735 4.3467e-006 1.7389e-005 0.16453 0.55402 0.65926 0.0016812 0.62831 0.34927 0.002254 0.41726 1.381 1.376 16.0111 144.9 0.00052804 -83.5362 0.11594
8.22 0.98814 5.467e-005 3.8183 0.011924 0.00010689 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5599 0.56849 0.17386 0.020091 16.6938 0.12455 0.00016246 0.76561 0.0093606 0.010358 0.0019654 0.97879 0.94007 4.3332e-006 1.7335e-005 0.16454 0.55535 0.66086 0.0016786 0.63024 0.34948 0.0022506 0.41725 1.3834 1.3785 16.0112 144.9 0.0005262 -83.5539 0.11694
8.221 0.98814 5.467e-005 3.8183 0.011924 0.0001069 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.56 0.56853 0.17387 0.020092 16.6969 0.12455 0.00016247 0.76561 0.009361 0.010358 0.0019597 0.97888 0.94265 4.3199e-006 1.7281e-005 0.16454 0.55667 0.66244 0.0016761 0.63217 0.3497 0.0022472 0.41724 1.3858 1.3809 16.0113 144.9 0.00052437 -83.5712 0.11794
8.222 0.98814 5.467e-005 3.8183 0.011924 0.00010692 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5601 0.56858 0.17389 0.020093 16.6999 0.12456 0.00016248 0.7656 0.0093613 0.010359 0.0019542 0.97897 0.94509 4.3068e-006 1.7229e-005 0.16454 0.55799 0.664 0.0016736 0.63409 0.34991 0.0022439 0.41724 1.3883 1.3834 16.0114 144.9 0.00052256 -83.5883 0.11894
8.223 0.98814 5.4669e-005 3.8183 0.011924 0.00010693 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5602 0.56862 0.1739 0.020094 16.7029 0.12457 0.00016249 0.76559 0.0093617 0.010359 0.0019487 0.97906 0.9474 4.294e-006 1.7178e-005 0.16454 0.55931 0.66556 0.0016711 0.636 0.35012 0.0022406 0.41723 1.3907 1.3858 16.0115 144.9 0.00052075 -83.6052 0.11994
8.224 0.98814 5.4669e-005 3.8183 0.011924 0.00010694 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5603 0.56867 0.17391 0.020095 16.7059 0.12457 0.0001625 0.76559 0.0093621 0.01036 0.0019433 0.97914 0.9496 4.2813e-006 1.7127e-005 0.16455 0.56062 0.6671 0.0016687 0.63791 0.35033 0.0022374 0.41723 1.3931 1.3883 16.0116 144.9 0.00051895 -83.6219 0.12094
8.225 0.98814 5.4669e-005 3.8183 0.011924 0.00010695 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5604 0.56871 0.17393 0.020096 16.7089 0.12458 0.00016251 0.76558 0.0093625 0.01036 0.001938 0.97922 0.95168 4.2689e-006 1.7077e-005 0.16455 0.56193 0.66862 0.0016663 0.6398 0.35054 0.0022343 0.41722 1.3956 1.3907 16.0117 144.9 0.00051717 -83.6383 0.12194
8.226 0.98814 5.4669e-005 3.8183 0.011924 0.00010697 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5604 0.56875 0.17394 0.020097 16.712 0.12459 0.00016252 0.76558 0.0093629 0.01036 0.0019328 0.97931 0.95365 4.2566e-006 1.7028e-005 0.16455 0.56323 0.67014 0.0016639 0.64169 0.35076 0.0022312 0.41722 1.398 1.3931 16.0118 144.9 0.00051539 -83.6546 0.12294
8.227 0.98814 5.4669e-005 3.8183 0.011924 0.00010698 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5605 0.5688 0.17396 0.020098 16.715 0.12459 0.00016253 0.76557 0.0093632 0.010361 0.0019276 0.97938 0.95551 4.2445e-006 1.698e-005 0.16456 0.56453 0.67164 0.0016616 0.64358 0.35097 0.0022281 0.41722 1.4004 1.3956 16.0119 144.9 0.00051362 -83.6707 0.12394
8.228 0.98814 5.4669e-005 3.8183 0.011924 0.00010699 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5606 0.56884 0.17397 0.020099 16.718 0.1246 0.00016254 0.76556 0.0093636 0.010361 0.0019226 0.97946 0.95728 4.2326e-006 1.6932e-005 0.16456 0.56583 0.67312 0.0016592 0.64546 0.35118 0.0022251 0.41721 1.4028 1.398 16.012 144.9 0.00051186 -83.6866 0.12494
8.229 0.98814 5.4669e-005 3.8183 0.011924 0.00010701 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5607 0.56889 0.17398 0.020101 16.721 0.12461 0.00016255 0.76556 0.009364 0.010362 0.0019176 0.97954 0.95895 4.2208e-006 1.6885e-005 0.16456 0.56712 0.6746 0.001657 0.64733 0.35139 0.0022221 0.41721 1.4052 1.4004 16.0121 144.9 0.00051012 -83.7023 0.12594
8.23 0.98814 5.4669e-005 3.8183 0.011924 0.00010702 0.0011731 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5608 0.56893 0.174 0.020102 16.724 0.12461 0.00016256 0.76555 0.0093644 0.010362 0.0019126 0.97962 0.96054 4.2092e-006 1.6838e-005 0.16456 0.56841 0.67606 0.0016547 0.64919 0.3516 0.0022191 0.4172 1.4076 1.4028 16.0122 144.9 0.00050838 -83.7178 0.12694
8.231 0.98814 5.4669e-005 3.8183 0.011924 0.00010703 0.0011732 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.5609 0.56898 0.17401 0.020103 16.727 0.12462 0.00016257 0.76554 0.0093648 0.010362 0.0019077 0.97969 0.96204 4.1978e-006 1.6793e-005 0.16457 0.56969 0.67751 0.0016525 0.65104 0.35182 0.0022162 0.4172 1.41 1.4052 16.0123 144.9 0.00050665 -83.7332 0.12794
8.232 0.98814 5.4669e-005 3.8183 0.011924 0.00010704 0.0011732 0.23372 0.00065931 0.23437 0.21628 0 0.032258 0.0389 0 1.561 0.56902 0.17402 0.020104 16.7301 0.12463 0.00016258 0.76554 0.0093651 0.010363 0.0019029 0.97976 0.96346 4.1865e-006 1.6747e-005 0.16457 0.57098 0.67895 0.0016503 0.65289 0.35203 0.0022133 0.4172 1.4124 1.4077 16.0124 144.9001 0.00050493 -83.7484 0.12894
8.233 0.98814 5.4669e-005 3.8183 0.011924 0.00010706 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.561 0.56907 0.17404 0.020105 16.7331 0.12463 0.00016259 0.76553 0.0093655 0.010363 0.0018982 0.97983 0.96481 4.1753e-006 1.6703e-005 0.16457 0.57225 0.68038 0.0016481 0.65473 0.35224 0.0022105 0.41719 1.4148 1.4101 16.0125 144.9001 0.00050322 -83.7635 0.12994
8.234 0.98814 5.4669e-005 3.8183 0.011924 0.00010707 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5611 0.56911 0.17405 0.020106 16.7361 0.12464 0.0001626 0.76552 0.0093659 0.010364 0.0018935 0.9799 0.96608 4.1643e-006 1.6659e-005 0.16458 0.57352 0.68179 0.001646 0.65657 0.35245 0.0022077 0.41719 1.4172 1.4125 16.0126 144.9001 0.00050152 -83.7785 0.13094
8.235 0.98814 5.4668e-005 3.8183 0.011924 0.00010708 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5612 0.56916 0.17406 0.020107 16.7391 0.12465 0.00016261 0.76552 0.0093663 0.010364 0.0018888 0.97997 0.96729 4.1534e-006 1.6615e-005 0.16458 0.57479 0.68319 0.0016438 0.6584 0.35267 0.0022049 0.41719 1.4196 1.4149 16.0126 144.9001 0.00049983 -83.7932 0.13194
8.236 0.98814 5.4668e-005 3.8183 0.011924 0.0001071 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5613 0.5692 0.17408 0.020108 16.7421 0.12465 0.00016262 0.76551 0.0093666 0.010364 0.0018842 0.98004 0.96844 4.1426e-006 1.6572e-005 0.16458 0.57606 0.68458 0.0016417 0.66022 0.35288 0.0022021 0.41718 1.422 1.4173 16.0127 144.9001 0.00049815 -83.8079 0.13294
8.237 0.98814 5.4668e-005 3.8183 0.011924 0.00010711 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5614 0.56925 0.17409 0.020109 16.7452 0.12466 0.00016263 0.7655 0.009367 0.010365 0.0018797 0.98011 0.96952 4.132e-006 1.6529e-005 0.16459 0.57732 0.68596 0.0016396 0.66203 0.35309 0.0021994 0.41718 1.4243 1.4197 16.0128 144.9001 0.00049648 -83.8224 0.13394
8.238 0.98814 5.4668e-005 3.8183 0.011924 0.00010712 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5615 0.56929 0.1741 0.02011 16.7482 0.12467 0.00016264 0.7655 0.0093674 0.010365 0.0018752 0.98018 0.97055 4.1215e-006 1.6488e-005 0.16459 0.57858 0.68733 0.0016376 0.66384 0.3533 0.0021967 0.41718 1.4267 1.422 16.0129 144.9001 0.00049481 -83.8368 0.13494
8.239 0.98814 5.4668e-005 3.8183 0.011924 0.00010713 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5616 0.56934 0.17412 0.020111 16.7512 0.12467 0.00016265 0.76549 0.0093678 0.010366 0.0018708 0.98024 0.97152 4.1112e-006 1.6446e-005 0.16459 0.57983 0.68869 0.0016355 0.66563 0.35352 0.002194 0.41718 1.4291 1.4244 16.013 144.9001 0.00049316 -83.851 0.13594
8.24 0.98814 5.4668e-005 3.8183 0.011924 0.00010715 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5616 0.56938 0.17413 0.020113 16.7542 0.12468 0.00016266 0.76548 0.0093682 0.010366 0.0018664 0.98031 0.97244 4.1009e-006 1.6405e-005 0.16459 0.58108 0.69003 0.0016335 0.66743 0.35373 0.0021914 0.41717 1.4314 1.4268 16.0131 144.9001 0.00049152 -83.8651 0.13694
8.241 0.98814 5.4668e-005 3.8183 0.011924 0.00010716 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5617 0.56943 0.17414 0.020114 16.7573 0.12468 0.00016267 0.76548 0.0093685 0.010366 0.0018621 0.98037 0.97331 4.0908e-006 1.6364e-005 0.1646 0.58233 0.69137 0.0016315 0.66921 0.35394 0.0021888 0.41717 1.4338 1.4292 16.0132 144.9001 0.00048988 -83.8791 0.13794
8.242 0.98814 5.4668e-005 3.8183 0.011924 0.00010717 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5618 0.56947 0.17416 0.020115 16.7603 0.12469 0.00016268 0.76547 0.0093689 0.010367 0.0018578 0.98044 0.97414 4.0808e-006 1.6324e-005 0.1646 0.58357 0.69269 0.0016295 0.67099 0.35415 0.0021862 0.41717 1.4362 1.4316 16.0133 144.9001 0.00048825 -83.893 0.13894
8.243 0.98814 5.4668e-005 3.8183 0.011924 0.00010719 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5619 0.56952 0.17417 0.020116 16.7633 0.1247 0.00016269 0.76547 0.0093693 0.010367 0.0018536 0.9805 0.97492 4.0709e-006 1.6285e-005 0.1646 0.58481 0.694 0.0016276 0.67276 0.35437 0.0021836 0.41717 1.4385 1.4339 16.0134 144.9001 0.00048664 -83.9067 0.13994
8.244 0.98814 5.4668e-005 3.8183 0.011924 0.0001072 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.562 0.56956 0.17418 0.020117 16.7663 0.1247 0.0001627 0.76546 0.0093697 0.010368 0.0018494 0.98056 0.97566 4.0611e-006 1.6245e-005 0.16461 0.58604 0.69531 0.0016257 0.67452 0.35458 0.0021811 0.41717 1.4409 1.4363 16.0134 144.9001 0.00048503 -83.9203 0.14094
8.245 0.98814 5.4668e-005 3.8183 0.011924 0.00010721 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5621 0.56961 0.1742 0.020118 16.7694 0.12471 0.00016271 0.76545 0.0093701 0.010368 0.0018453 0.98062 0.97636 4.0514e-006 1.6207e-005 0.16461 0.58727 0.6966 0.0016237 0.67628 0.35479 0.0021786 0.41716 1.4432 1.4386 16.0135 144.9001 0.00048343 -83.9338 0.14194
8.246 0.98814 5.4668e-005 3.8183 0.011924 0.00010722 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5622 0.56965 0.17421 0.020119 16.7724 0.12472 0.00016272 0.76545 0.0093704 0.010369 0.0018412 0.98068 0.97703 4.0418e-006 1.6168e-005 0.16461 0.5885 0.69788 0.0016218 0.67803 0.355 0.0021761 0.41716 1.4455 1.441 16.0136 144.9002 0.00048184 -83.9472 0.14294
8.247 0.98814 5.4667e-005 3.8183 0.011924 0.00010724 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5622 0.5697 0.17422 0.02012 16.7754 0.12472 0.00016273 0.76544 0.0093708 0.010369 0.0018371 0.98074 0.97766 4.0323e-006 1.613e-005 0.16461 0.58972 0.69915 0.0016199 0.67977 0.35522 0.0021736 0.41716 1.4479 1.4433 16.0137 144.9002 0.00048025 -83.9604 0.14394
8.248 0.98814 5.4667e-005 3.8183 0.011924 0.00010725 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5623 0.56974 0.17424 0.020121 16.7784 0.12473 0.00016274 0.76543 0.0093712 0.010369 0.0018331 0.9808 0.97825 4.0229e-006 1.6093e-005 0.16462 0.59094 0.70041 0.0016181 0.6815 0.35543 0.0021712 0.41716 1.4502 1.4457 16.0138 144.9002 0.00047868 -83.9736 0.14494
8.249 0.98814 5.4667e-005 3.8183 0.011923 0.00010726 0.0011732 0.23372 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5624 0.56978 0.17425 0.020122 16.7815 0.12474 0.00016275 0.76543 0.0093716 0.01037 0.0018292 0.98086 0.97882 4.0137e-006 1.6056e-005 0.16462 0.59216 0.70166 0.0016162 0.68323 0.35564 0.0021688 0.41716 1.4525 1.448 16.0139 144.9002 0.00047711 -83.9866 0.14594
8.25 0.98814 5.4667e-005 3.8183 0.011923 0.00010728 0.0011732 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5625 0.56983 0.17426 0.020123 16.7845 0.12474 0.00016276 0.76542 0.0093719 0.01037 0.0018252 0.98091 0.97935 4.0045e-006 1.6019e-005 0.16462 0.59337 0.70291 0.0016144 0.68495 0.35585 0.0021664 0.41716 1.4549 1.4504 16.0139 144.9002 0.00047556 -83.9996 0.14694
8.251 0.98814 5.4667e-005 3.8183 0.011923 0.00010729 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5626 0.56987 0.17428 0.020125 16.7875 0.12475 0.00016277 0.76541 0.0093723 0.010371 0.0018214 0.98097 0.97986 3.9954e-006 1.5983e-005 0.16463 0.59458 0.70414 0.0016126 0.68666 0.35607 0.002164 0.41716 1.4572 1.4527 16.014 144.9002 0.00047401 -84.0124 0.14794
8.252 0.98814 5.4667e-005 3.8183 0.011923 0.0001073 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5627 0.56992 0.17429 0.020126 16.7905 0.12476 0.00016278 0.76541 0.0093727 0.010371 0.0018175 0.98103 0.98034 3.9864e-006 1.5947e-005 0.16463 0.59579 0.70536 0.0016108 0.68837 0.35628 0.0021617 0.41716 1.4595 1.455 16.0141 144.9002 0.00047247 -84.0251 0.14894
8.253 0.98814 5.4667e-005 3.8183 0.011923 0.00010731 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5628 0.56996 0.1743 0.020127 16.7936 0.12476 0.00016279 0.7654 0.0093731 0.010371 0.0018137 0.98108 0.9808 3.9776e-006 1.5911e-005 0.16463 0.59699 0.70657 0.001609 0.69006 0.35649 0.0021594 0.41716 1.4618 1.4574 16.0142 144.9002 0.00047093 -84.0377 0.14994
8.254 0.98814 5.4667e-005 3.8183 0.011923 0.00010733 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5628 0.57001 0.17432 0.020128 16.7966 0.12477 0.0001628 0.76539 0.0093735 0.010372 0.00181 0.98114 0.98123 3.9688e-006 1.5876e-005 0.16463 0.59819 0.70778 0.0016073 0.69175 0.35671 0.0021571 0.41716 1.4641 1.4597 16.0143 144.9002 0.00046941 -84.0502 0.15094
8.255 0.98814 5.4667e-005 3.8183 0.011923 0.00010734 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5629 0.57005 0.17433 0.020129 16.7996 0.12478 0.00016281 0.76539 0.0093738 0.010372 0.0018062 0.98119 0.98164 3.9601e-006 1.5841e-005 0.16464 0.59938 0.70897 0.0016055 0.69344 0.35692 0.0021548 0.41716 1.4664 1.462 16.0143 144.9002 0.00046789 -84.0626 0.15194
8.256 0.98814 5.4667e-005 3.8183 0.011923 0.00010735 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.563 0.5701 0.17434 0.02013 16.8026 0.12478 0.00016282 0.76538 0.0093742 0.010373 0.0018025 0.98124 0.98203 3.9515e-006 1.5807e-005 0.16464 0.60057 0.71016 0.0016038 0.69512 0.35713 0.0021525 0.41716 1.4687 1.4643 16.0144 144.9002 0.00046639 -84.0749 0.15294
8.257 0.98814 5.4667e-005 3.8183 0.011923 0.00010736 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5631 0.57014 0.17436 0.020131 16.8057 0.12479 0.00016283 0.76537 0.0093746 0.010373 0.0017989 0.9813 0.98239 3.9429e-006 1.5773e-005 0.16464 0.60176 0.71133 0.0016021 0.69678 0.35734 0.0021503 0.41716 1.471 1.4666 16.0145 144.9002 0.00046489 -84.0871 0.15394
8.258 0.98814 5.4667e-005 3.8183 0.011923 0.00010738 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5632 0.57019 0.17437 0.020132 16.8087 0.12479 0.00016284 0.76537 0.009375 0.010373 0.0017953 0.98135 0.98274 3.9345e-006 1.5739e-005 0.16465 0.60294 0.7125 0.0016004 0.69845 0.35756 0.0021481 0.41716 1.4733 1.4689 16.0146 144.9003 0.0004634 -84.0992 0.15494
8.259 0.98814 5.4667e-005 3.8183 0.011923 0.00010739 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5633 0.57023 0.17439 0.020133 16.8117 0.1248 0.00016285 0.76536 0.0093753 0.010374 0.0017917 0.9814 0.98307 3.9262e-006 1.5706e-005 0.16465 0.60412 0.71365 0.0015987 0.7001 0.35777 0.0021459 0.41716 1.4756 1.4712 16.0147 144.9003 0.00046191 -84.1111 0.15594
8.26 0.98814 5.4666e-005 3.8183 0.011923 0.0001074 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5634 0.57028 0.1744 0.020134 16.8148 0.12481 0.00016286 0.76536 0.0093757 0.010374 0.0017882 0.98145 0.98339 3.9179e-006 1.5673e-005 0.16465 0.60529 0.7148 0.0015971 0.70175 0.35798 0.0021437 0.41716 1.4779 1.4735 16.0147 144.9003 0.00046044 -84.123 0.15694
8.261 0.98814 5.4666e-005 3.8183 0.011923 0.00010742 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5634 0.57032 0.17441 0.020135 16.8178 0.12481 0.00016287 0.76535 0.0093761 0.010375 0.0017847 0.9815 0.98368 3.9098e-006 1.564e-005 0.16466 0.60647 0.71594 0.0015954 0.70339 0.3582 0.0021416 0.41716 1.4802 1.4758 16.0148 144.9003 0.00045897 -84.1348 0.15794
8.262 0.98814 5.4666e-005 3.8183 0.011923 0.00010743 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5635 0.57037 0.17443 0.020136 16.8208 0.12482 0.00016288 0.76534 0.0093765 0.010375 0.0017812 0.98155 0.98397 3.9017e-006 1.5608e-005 0.16466 0.60764 0.71708 0.0015938 0.70502 0.35841 0.0021394 0.41716 1.4824 1.4781 16.0149 144.9003 0.00045751 -84.1465 0.15894
8.263 0.98814 5.4666e-005 3.8183 0.011923 0.00010744 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5636 0.57041 0.17444 0.020138 16.8238 0.12483 0.00016289 0.76534 0.0093769 0.010375 0.0017778 0.9816 0.98423 3.8937e-006 1.5576e-005 0.16466 0.6088 0.7182 0.0015922 0.70665 0.35862 0.0021373 0.41716 1.4847 1.4804 16.015 144.9003 0.00045606 -84.1581 0.15994
8.264 0.98814 5.4666e-005 3.8183 0.011923 0.00010745 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5637 0.57046 0.17445 0.020139 16.8269 0.12483 0.0001629 0.76533 0.0093772 0.010376 0.0017744 0.98165 0.98449 3.8858e-006 1.5544e-005 0.16466 0.60996 0.71931 0.0015906 0.70827 0.35883 0.0021352 0.41716 1.487 1.4827 16.015 144.9003 0.00045461 -84.1696 0.16094
8.265 0.98814 5.4666e-005 3.8183 0.011923 0.00010747 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5638 0.5705 0.17447 0.02014 16.8299 0.12484 0.00016291 0.76532 0.0093776 0.010376 0.001771 0.9817 0.98473 3.8779e-006 1.5513e-005 0.16467 0.61112 0.72042 0.001589 0.70988 0.35905 0.0021331 0.41717 1.4892 1.485 16.0151 144.9003 0.00045318 -84.1811 0.16194
8.266 0.98814 5.4666e-005 3.8183 0.011923 0.00010748 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032258 0.0389 0 1.5639 0.57055 0.17448 0.020141 16.8329 0.12485 0.00016292 0.76532 0.009378 0.010377 0.0017677 0.98175 0.98496 3.8702e-006 1.5482e-005 0.16467 0.61228 0.72152 0.0015874 0.71149 0.35926 0.0021311 0.41717 1.4915 1.4872 16.0152 144.9003 0.00045175 -84.1924 0.16294
8.267 0.98814 5.4666e-005 3.8183 0.011923 0.00010749 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.564 0.57059 0.17449 0.020142 16.836 0.12485 0.00016293 0.76531 0.0093784 0.010377 0.0017644 0.98179 0.98518 3.8625e-006 1.5451e-005 0.16467 0.61343 0.72261 0.0015858 0.71308 0.35947 0.0021291 0.41717 1.4937 1.4895 16.0153 144.9003 0.00045033 -84.2036 0.16394
8.268 0.98814 5.4666e-005 3.8183 0.011923 0.00010751 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.564 0.57064 0.17451 0.020143 16.839 0.12486 0.00016294 0.7653 0.0093787 0.010377 0.0017611 0.98184 0.98538 3.8549e-006 1.542e-005 0.16468 0.61457 0.72369 0.0015843 0.71467 0.35969 0.002127 0.41717 1.496 1.4918 16.0153 144.9003 0.00044891 -84.2147 0.16494
8.269 0.98814 5.4666e-005 3.8183 0.011923 0.00010752 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5641 0.57068 0.17452 0.020144 16.842 0.12487 0.00016295 0.7653 0.0093791 0.010378 0.0017579 0.98189 0.98558 3.8473e-006 1.539e-005 0.16468 0.61572 0.72476 0.0015828 0.71626 0.3599 0.002125 0.41717 1.4982 1.494 16.0154 144.9004 0.00044751 -84.2258 0.16594
8.27 0.98814 5.4666e-005 3.8183 0.011923 0.00010753 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5642 0.57073 0.17453 0.020145 16.8451 0.12487 0.00016296 0.76529 0.0093795 0.010378 0.0017547 0.98193 0.98577 3.8399e-006 1.536e-005 0.16468 0.61686 0.72583 0.0015813 0.71783 0.36011 0.002123 0.41717 1.5005 1.4963 16.0155 144.9004 0.00044611 -84.2367 0.16694
8.271 0.98814 5.4666e-005 3.8183 0.011923 0.00010754 0.0011733 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5643 0.57077 0.17455 0.020146 16.8481 0.12488 0.00016297 0.76528 0.0093799 0.010379 0.0017516 0.98198 0.98595 3.8325e-006 1.5331e-005 0.16468 0.618 0.72689 0.0015798 0.7194 0.36032 0.0021211 0.41718 1.5027 1.4985 16.0155 144.9004 0.00044472 -84.2476 0.16794
8.272 0.98814 5.4665e-005 3.8183 0.011923 0.00010756 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5644 0.57081 0.17456 0.020147 16.8511 0.12489 0.00016298 0.76528 0.0093802 0.010379 0.0017484 0.98202 0.98611 3.8252e-006 1.5302e-005 0.16469 0.61913 0.72794 0.0015783 0.72097 0.36054 0.0021191 0.41718 1.505 1.5008 16.0156 144.9004 0.00044333 -84.2584 0.16894
8.273 0.98814 5.4665e-005 3.8183 0.011923 0.00010757 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5645 0.57086 0.17457 0.020148 16.8542 0.12489 0.00016299 0.76527 0.0093806 0.010379 0.0017453 0.98207 0.98628 3.818e-006 1.5273e-005 0.16469 0.62026 0.72898 0.0015768 0.72252 0.36075 0.0021172 0.41718 1.5072 1.503 16.0157 144.9004 0.00044195 -84.2691 0.16994
8.274 0.98814 5.4665e-005 3.8183 0.011923 0.00010758 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5646 0.5709 0.17459 0.020149 16.8572 0.1249 0.000163 0.76526 0.009381 0.01038 0.0017423 0.98211 0.98643 3.8108e-006 1.5244e-005 0.16469 0.62139 0.73001 0.0015753 0.72407 0.36096 0.0021153 0.41718 1.5094 1.5053 16.0158 144.9004 0.00044058 -84.2797 0.17094
8.275 0.98814 5.4665e-005 3.8183 0.011923 0.0001076 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5646 0.57095 0.1746 0.020151 16.8602 0.1249 0.00016301 0.76526 0.0093814 0.01038 0.0017392 0.98215 0.98657 3.8037e-006 1.5216e-005 0.1647 0.62251 0.73104 0.0015739 0.72561 0.36118 0.0021134 0.41719 1.5116 1.5075 16.0158 144.9004 0.00043922 -84.2902 0.17194
8.276 0.98814 5.4665e-005 3.8183 0.011923 0.00010761 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5647 0.57099 0.17461 0.020152 16.8633 0.12491 0.00016302 0.76525 0.0093818 0.010381 0.0017362 0.9822 0.98671 3.7967e-006 1.5188e-005 0.1647 0.62363 0.73206 0.0015724 0.72714 0.36139 0.0021115 0.41719 1.5138 1.5097 16.0159 144.9004 0.00043787 -84.3007 0.17294
8.277 0.98814 5.4665e-005 3.8183 0.011923 0.00010762 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5648 0.57104 0.17463 0.020153 16.8663 0.12492 0.00016303 0.76525 0.0093821 0.010381 0.0017331 0.98224 0.98685 3.7897e-006 1.516e-005 0.1647 0.62474 0.73307 0.001571 0.72867 0.3616 0.0021097 0.41719 1.516 1.5119 16.016 144.9004 0.00043652 -84.311 0.17394
8.278 0.98814 5.4665e-005 3.8183 0.011923 0.00010763 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5649 0.57108 0.17464 0.020154 16.8693 0.12492 0.00016304 0.76524 0.0093825 0.010381 0.0017302 0.98228 0.98697 3.7828e-006 1.5132e-005 0.1647 0.62586 0.73408 0.0015696 0.73019 0.36182 0.0021078 0.41719 1.5183 1.5142 16.016 144.9004 0.00043518 -84.3213 0.17494
8.279 0.98814 5.4665e-005 3.8183 0.011923 0.00010765 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.565 0.57113 0.17465 0.020155 16.8724 0.12493 0.00016305 0.76523 0.0093829 0.010382 0.0017273 0.98232 0.98709 3.776e-006 1.5105e-005 0.16471 0.62697 0.73508 0.0015682 0.7317 0.36203 0.002106 0.4172 1.5205 1.5164 16.0161 144.9005 0.00043384 -84.3315 0.17594
8.28 0.98814 5.4665e-005 3.8183 0.011923 0.00010766 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5651 0.57117 0.17467 0.020156 16.8754 0.12494 0.00016306 0.76523 0.0093833 0.010382 0.0017244 0.98236 0.98721 3.7693e-006 1.5078e-005 0.16471 0.62807 0.73607 0.0015668 0.73321 0.36224 0.0021042 0.4172 1.5227 1.5186 16.0162 144.9005 0.00043252 -84.3416 0.17694
8.281 0.98814 5.4665e-005 3.8183 0.011923 0.00010767 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5652 0.57122 0.17468 0.020157 16.8784 0.12494 0.00016307 0.76522 0.0093836 0.010383 0.0017216 0.98241 0.98732 3.7626e-006 1.5051e-005 0.16471 0.62918 0.73705 0.0015654 0.73471 0.36245 0.0021024 0.4172 1.5249 1.5208 16.0162 144.9005 0.0004312 -84.3516 0.17794
8.282 0.98814 5.4665e-005 3.8183 0.011923 0.00010769 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5652 0.57126 0.17469 0.020158 16.8815 0.12495 0.00016308 0.76521 0.009384 0.010383 0.0017188 0.98245 0.98742 3.756e-006 1.5025e-005 0.16472 0.63027 0.73803 0.0015641 0.7362 0.36267 0.0021006 0.41721 1.527 1.523 16.0163 144.9005 0.00042988 -84.3616 0.17894
8.283 0.98814 5.4665e-005 3.8183 0.011923 0.0001077 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5653 0.57131 0.17471 0.020159 16.8845 0.12496 0.00016308 0.76521 0.0093844 0.010383 0.001716 0.98249 0.98752 3.7495e-006 1.4999e-005 0.16472 0.63137 0.739 0.0015627 0.73768 0.36288 0.0020988 0.41721 1.5292 1.5252 16.0164 144.9005 0.00042858 -84.3714 0.17994
8.284 0.98814 5.4664e-005 3.8183 0.011923 0.00010771 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5654 0.57135 0.17472 0.02016 16.8876 0.12496 0.00016309 0.7652 0.0093848 0.010384 0.0017132 0.98253 0.98761 3.743e-006 1.4973e-005 0.16472 0.63246 0.73996 0.0015614 0.73916 0.36309 0.0020971 0.41721 1.5314 1.5274 16.0164 144.9005 0.00042728 -84.3812 0.18094
8.285 0.98814 5.4664e-005 3.8183 0.011923 0.00010772 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5655 0.5714 0.17473 0.020161 16.8906 0.12497 0.0001631 0.76519 0.0093851 0.010384 0.0017103 0.98256 0.98771 3.7365e-006 1.4947e-005 0.16472 0.63355 0.74092 0.0015601 0.74063 0.36331 0.0020953 0.41722 1.5336 1.5296 16.0165 144.9005 0.00042599 -84.3909 0.18194
8.286 0.98814 5.4664e-005 3.8183 0.011923 0.00010774 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5656 0.57144 0.17475 0.020163 16.8936 0.12498 0.00016311 0.76519 0.0093855 0.010385 0.0017075 0.9826 0.98779 3.7301e-006 1.4921e-005 0.16473 0.63464 0.74187 0.0015587 0.7421 0.36352 0.0020936 0.41722 1.5358 1.5318 16.0166 144.9005 0.0004247 -84.4006 0.18294
8.287 0.98814 5.4664e-005 3.8183 0.011923 0.00010775 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5657 0.57149 0.17476 0.020164 16.8967 0.12498 0.00016312 0.76518 0.0093859 0.010385 0.0017047 0.98264 0.98788 3.7237e-006 1.4896e-005 0.16473 0.63572 0.74281 0.0015574 0.74355 0.36373 0.0020919 0.41723 1.5379 1.5339 16.0166 144.9005 0.00042342 -84.4101 0.18394
8.288 0.98814 5.4664e-005 3.8183 0.011923 0.00010776 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5657 0.57153 0.17477 0.020165 16.8997 0.12499 0.00016313 0.76517 0.0093863 0.010385 0.0017019 0.98268 0.98796 3.7174e-006 1.4871e-005 0.16473 0.6368 0.74375 0.0015561 0.74501 0.36394 0.0020902 0.41723 1.5401 1.5361 16.0167 144.9006 0.00042215 -84.4196 0.18494
8.289 0.98814 5.4664e-005 3.8183 0.011923 0.00010777 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5658 0.57158 0.17479 0.020166 16.9027 0.125 0.00016314 0.76517 0.0093866 0.010386 0.0016992 0.98272 0.98803 3.7112e-006 1.4846e-005 0.16474 0.63788 0.74468 0.0015548 0.74645 0.36416 0.0020886 0.41723 1.5422 1.5383 16.0168 144.9006 0.00042088 -84.429 0.18594
8.29 0.98814 5.4664e-005 3.8183 0.011923 0.00010779 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5659 0.57162 0.1748 0.020167 16.9058 0.125 0.00016315 0.76516 0.009387 0.010386 0.0016966 0.98275 0.9881 3.7051e-006 1.4821e-005 0.16474 0.63895 0.74561 0.0015536 0.74788 0.36437 0.0020869 0.41724 1.5444 1.5405 16.0168 144.9006 0.00041962 -84.4383 0.18694
8.291 0.98814 5.4664e-005 3.8183 0.011923 0.0001078 0.0011734 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.566 0.57166 0.17481 0.020168 16.9088 0.12501 0.00016316 0.76515 0.0093874 0.010387 0.0016941 0.98279 0.98818 3.6991e-006 1.4797e-005 0.16474 0.64002 0.74652 0.0015523 0.74931 0.36458 0.0020853 0.41724 1.5465 1.5426 16.0169 144.9006 0.00041837 -84.4476 0.18794
8.292 0.98814 5.4664e-005 3.8183 0.011923 0.00010781 0.0011735 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5661 0.57171 0.17483 0.020169 16.9119 0.12501 0.00016317 0.76515 0.0093878 0.010387 0.0016916 0.98283 0.98824 3.6932e-006 1.4773e-005 0.16474 0.64108 0.74744 0.0015511 0.75074 0.3648 0.0020836 0.41725 1.5487 1.5448 16.0169 144.9006 0.00041712 -84.4568 0.18894
8.293 0.98814 5.4664e-005 3.8183 0.011923 0.00010783 0.0011735 0.23371 0.00065931 0.23437 0.21627 0 0.032259 0.0389 0 1.5662 0.57175 0.17484 0.02017 16.9149 0.12502 0.00016318 0.76514 0.0093881 0.010387 0.0016891 0.98286 0.98831 3.6873e-006 1.475e-005 0.16475 0.64215 0.74834 0.0015499 0.75215 0.36501 0.002082 0.41725 1.5508 1.5469 16.017 144.9006 0.00041588 -84.4659 0.18994
8.294 0.98814 5.4664e-005 3.8183 0.011923 0.00010784 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5663 0.5718 0.17485 0.020171 16.9179 0.12503 0.00016319 0.76514 0.0093885 0.010388 0.0016866 0.9829 0.98837 3.6814e-006 1.4726e-005 0.16475 0.64321 0.74924 0.0015486 0.75356 0.36522 0.0020804 0.41726 1.553 1.5491 16.0171 144.9006 0.00041465 -84.4749 0.19094
8.295 0.98814 5.4664e-005 3.8183 0.011923 0.00010785 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5663 0.57184 0.17487 0.020172 16.921 0.12503 0.0001632 0.76513 0.0093889 0.010388 0.0016841 0.98293 0.98843 3.6756e-006 1.4703e-005 0.16475 0.64426 0.75013 0.0015474 0.75496 0.36543 0.0020788 0.41726 1.5551 1.5512 16.0171 144.9006 0.00041342 -84.4839 0.19194
8.296 0.98814 5.4663e-005 3.8183 0.011923 0.00010786 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5664 0.57189 0.17488 0.020173 16.924 0.12504 0.00016321 0.76512 0.0093893 0.010389 0.0016816 0.98297 0.98849 3.6698e-006 1.468e-005 0.16476 0.64532 0.75102 0.0015462 0.75636 0.36565 0.0020772 0.41727 1.5572 1.5534 16.0172 144.9006 0.0004122 -84.4928 0.19294
8.297 0.98814 5.4663e-005 3.8183 0.011923 0.00010788 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5665 0.57193 0.1749 0.020174 16.9271 0.12505 0.00016322 0.76512 0.0093896 0.010389 0.0016792 0.983 0.98854 3.6641e-006 1.4657e-005 0.16476 0.64637 0.7519 0.001545 0.75775 0.36586 0.0020757 0.41727 1.5594 1.5555 16.0173 144.9007 0.00041099 -84.5016 0.19394
8.298 0.98814 5.4663e-005 3.8183 0.011923 0.00010789 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5666 0.57198 0.17491 0.020176 16.9301 0.12505 0.00016323 0.76511 0.00939 0.010389 0.0016767 0.98304 0.98859 3.6584e-006 1.4634e-005 0.16476 0.64741 0.75277 0.0015439 0.75913 0.36607 0.0020741 0.41728 1.5615 1.5576 16.0173 144.9007 0.00040978 -84.5104 0.19494
8.299 0.98814 5.4663e-005 3.8183 0.011923 0.0001079 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5667 0.57202 0.17492 0.020177 16.9332 0.12506 0.00016324 0.7651 0.0093904 0.01039 0.0016743 0.98307 0.98864 3.6528e-006 1.4612e-005 0.16477 0.64846 0.75364 0.0015427 0.76051 0.36629 0.0020726 0.41728 1.5636 1.5598 16.0174 144.9007 0.00040858 -84.519 0.19594
8.3 0.98814 5.4663e-005 3.8183 0.011923 0.00010792 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5668 0.57207 0.17494 0.020178 16.9362 0.12507 0.00016325 0.7651 0.0093908 0.01039 0.0016719 0.98311 0.98869 3.6472e-006 1.4589e-005 0.16477 0.6495 0.75451 0.0015415 0.76187 0.3665 0.0020711 0.41729 1.5657 1.5619 16.0174 144.9007 0.00040738 -84.5277 0.19694
8.301 0.98814 5.4663e-005 3.8183 0.011923 0.00010793 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5669 0.57211 0.17495 0.020179 16.9392 0.12507 0.00016326 0.76509 0.0093912 0.01039 0.0016695 0.98314 0.98874 3.6417e-006 1.4567e-005 0.16477 0.65053 0.75536 0.0015404 0.76324 0.36671 0.0020696 0.41729 1.5678 1.564 16.0175 144.9007 0.00040619 -84.5362 0.19794
8.302 0.98814 5.4663e-005 3.8183 0.011923 0.00010794 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5669 0.57216 0.17496 0.02018 16.9423 0.12508 0.00016327 0.76508 0.0093915 0.010391 0.0016671 0.98317 0.98879 3.6362e-006 1.4545e-005 0.16477 0.65157 0.75622 0.0015392 0.76459 0.36692 0.0020681 0.4173 1.5699 1.5661 16.0175 144.9007 0.00040501 -84.5447 0.19894
8.303 0.98814 5.4663e-005 3.8183 0.011923 0.00010795 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.567 0.5722 0.17498 0.020181 16.9453 0.12509 0.00016328 0.76508 0.0093919 0.010391 0.0016648 0.9832 0.98883 3.6308e-006 1.4524e-005 0.16478 0.6526 0.75706 0.0015381 0.76594 0.36714 0.0020666 0.4173 1.572 1.5682 16.0176 144.9007 0.00040383 -84.5531 0.19994
8.304 0.98814 5.4663e-005 3.8183 0.011923 0.00010797 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5671 0.57225 0.17499 0.020182 16.9484 0.12509 0.00016329 0.76507 0.0093923 0.010392 0.0016625 0.98324 0.98887 3.6254e-006 1.4502e-005 0.16478 0.65363 0.7579 0.0015369 0.76728 0.36735 0.0020651 0.41731 1.5741 1.5703 16.0177 144.9007 0.00040266 -84.5615 0.20094
8.305 0.98814 5.4663e-005 3.8183 0.011923 0.00010798 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5672 0.57229 0.175 0.020183 16.9514 0.1251 0.0001633 0.76506 0.0093927 0.010392 0.0016602 0.98327 0.98892 3.6201e-006 1.4481e-005 0.16478 0.65465 0.75874 0.0015358 0.76862 0.36756 0.0020637 0.41731 1.5762 1.5724 16.0177 144.9008 0.00040149 -84.5698 0.20194
8.306 0.98814 5.4663e-005 3.8183 0.011922 0.00010799 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5673 0.57234 0.17502 0.020184 16.9545 0.12511 0.00016331 0.76506 0.009393 0.010392 0.0016579 0.9833 0.98896 3.6148e-006 1.446e-005 0.16479 0.65567 0.75957 0.0015347 0.76994 0.36777 0.0020622 0.41732 1.5783 1.5745 16.0178 144.9008 0.00040033 -84.578 0.20294
8.307 0.98814 5.4663e-005 3.8183 0.011922 0.00010801 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5674 0.57238 0.17503 0.020185 16.9575 0.12511 0.00016332 0.76505 0.0093934 0.010393 0.0016557 0.98333 0.98899 3.6096e-006 1.4439e-005 0.16479 0.65669 0.76039 0.0015336 0.77127 0.36799 0.0020608 0.41733 1.5803 1.5766 16.0178 144.9008 0.00039918 -84.5861 0.20394
8.308 0.98814 5.4662e-005 3.8183 0.011922 0.00010802 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5675 0.57243 0.17504 0.020186 16.9605 0.12512 0.00016333 0.76505 0.0093938 0.010393 0.0016534 0.98336 0.98903 3.6045e-006 1.4418e-005 0.16479 0.6577 0.76121 0.0015325 0.77258 0.3682 0.0020594 0.41733 1.5824 1.5787 16.0179 144.9008 0.00039803 -84.5942 0.20494
8.309 0.98814 5.4662e-005 3.8183 0.011922 0.00010803 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5675 0.57247 0.17506 0.020187 16.9636 0.12512 0.00016334 0.76504 0.0093941 0.010394 0.0016512 0.98339 0.98907 3.5993e-006 1.4398e-005 0.16479 0.65872 0.76202 0.0015315 0.77389 0.36841 0.002058 0.41734 1.5845 1.5808 16.0179 144.9008 0.00039689 -84.6022 0.20594
8.31 0.98814 5.4662e-005 3.8183 0.011922 0.00010804 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5676 0.57251 0.17507 0.020188 16.9666 0.12513 0.00016335 0.76503 0.0093945 0.010394 0.0016491 0.98342 0.9891 3.5943e-006 1.4378e-005 0.1648 0.65973 0.76283 0.0015304 0.77519 0.36863 0.0020566 0.41734 1.5866 1.5829 16.018 144.9008 0.00039575 -84.6102 0.20694
8.311 0.98814 5.4662e-005 3.8183 0.011922 0.00010806 0.0011735 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5677 0.57256 0.17508 0.02019 16.9697 0.12514 0.00016336 0.76503 0.0093949 0.010394 0.0016469 0.98345 0.98914 3.5893e-006 1.4358e-005 0.1648 0.66073 0.76363 0.0015294 0.77649 0.36884 0.0020552 0.41735 1.5886 1.5849 16.018 144.9008 0.00039462 -84.6181 0.20794
8.312 0.98814 5.4662e-005 3.8183 0.011922 0.00010807 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5678 0.5726 0.1751 0.020191 16.9727 0.12514 0.00016337 0.76502 0.0093953 0.010395 0.0016448 0.98348 0.98917 3.5843e-006 1.4338e-005 0.1648 0.66173 0.76443 0.0015283 0.77778 0.36905 0.0020538 0.41736 1.5907 1.587 16.0181 144.9008 0.0003935 -84.626 0.20894
8.313 0.98814 5.4662e-005 3.8183 0.011922 0.00010808 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5679 0.57265 0.17511 0.020192 16.9758 0.12515 0.00016338 0.76501 0.0093956 0.010395 0.0016426 0.98351 0.9892 3.5794e-006 1.4318e-005 0.16481 0.66273 0.76522 0.0015273 0.77906 0.36926 0.0020525 0.41736 1.5927 1.5891 16.0182 144.9009 0.00039238 -84.6337 0.20994
8.314 0.98814 5.4662e-005 3.8183 0.011922 0.0001081 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.568 0.57269 0.17512 0.020193 16.9788 0.12516 0.00016339 0.76501 0.009396 0.010396 0.0016405 0.98354 0.98923 3.5745e-006 1.4298e-005 0.16481 0.66373 0.76601 0.0015262 0.78034 0.36948 0.0020511 0.41737 1.5948 1.5911 16.0182 144.9009 0.00039126 -84.6415 0.21094
8.315 0.98814 5.4662e-005 3.8183 0.011922 0.00010811 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5681 0.57274 0.17514 0.020194 16.9819 0.12516 0.0001634 0.765 0.0093964 0.010396 0.0016384 0.98357 0.98927 3.5696e-006 1.4279e-005 0.16481 0.66472 0.76679 0.0015252 0.78161 0.36969 0.0020498 0.41738 1.5968 1.5932 16.0183 144.9009 0.00039016 -84.6491 0.21194
8.316 0.98814 5.4662e-005 3.8183 0.011922 0.00010812 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5681 0.57278 0.17515 0.020195 16.9849 0.12517 0.00016341 0.76499 0.0093968 0.010396 0.0016364 0.9836 0.98929 3.5648e-006 1.426e-005 0.16481 0.66571 0.76757 0.0015242 0.78287 0.3699 0.0020485 0.41738 1.5989 1.5952 16.0183 144.9009 0.00038905 -84.6567 0.21294
8.317 0.98814 5.4662e-005 3.8183 0.011922 0.00010813 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5682 0.57283 0.17516 0.020196 16.988 0.12518 0.00016342 0.76499 0.0093971 0.010397 0.0016343 0.98363 0.98932 3.5601e-006 1.4241e-005 0.16482 0.6667 0.76834 0.0015232 0.78413 0.37011 0.0020471 0.41739 1.6009 1.5973 16.0184 144.9009 0.00038796 -84.6643 0.21394
8.318 0.98814 5.4662e-005 3.8183 0.011922 0.00010815 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5683 0.57287 0.17518 0.020197 16.991 0.12518 0.00016343 0.76498 0.0093975 0.010397 0.0016323 0.98366 0.98935 3.5554e-006 1.4222e-005 0.16482 0.66768 0.76911 0.0015222 0.78538 0.37033 0.0020458 0.4174 1.6029 1.5993 16.0184 144.9009 0.00038687 -84.6717 0.21494
8.319 0.98814 5.4662e-005 3.8183 0.011922 0.00010816 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5684 0.57292 0.17519 0.020198 16.9941 0.12519 0.00016344 0.76497 0.0093979 0.010398 0.0016303 0.98368 0.98938 3.5507e-006 1.4203e-005 0.16482 0.66867 0.76988 0.0015212 0.78662 0.37054 0.0020445 0.4174 1.6049 1.6014 16.0185 144.9009 0.00038578 -84.6792 0.21594
8.32 0.98814 5.4661e-005 3.8183 0.011922 0.00010817 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5685 0.57296 0.1752 0.020199 16.9971 0.1252 0.00016345 0.76497 0.0093983 0.010398 0.0016283 0.98371 0.98941 3.5461e-006 1.4185e-005 0.16483 0.66964 0.77063 0.0015202 0.78786 0.37075 0.0020433 0.41741 1.607 1.6034 16.0185 144.9009 0.0003847 -84.6865 0.21694
8.321 0.98814 5.4661e-005 3.8183 0.011922 0.00010818 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5686 0.57301 0.17522 0.0202 17.0002 0.1252 0.00016346 0.76496 0.0093986 0.010398 0.0016263 0.98374 0.98943 3.5415e-006 1.4166e-005 0.16483 0.67062 0.77139 0.0015193 0.78909 0.37096 0.002042 0.41742 1.609 1.6054 16.0186 144.901 0.00038363 -84.6938 0.21794
8.322 0.98814 5.4661e-005 3.8183 0.011922 0.0001082 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5687 0.57305 0.17523 0.020201 17.0032 0.12521 0.00016347 0.76496 0.009399 0.010399 0.0016243 0.98377 0.98946 3.537e-006 1.4148e-005 0.16483 0.67159 0.77214 0.0015183 0.79031 0.37118 0.0020407 0.41742 1.611 1.6075 16.0186 144.901 0.00038256 -84.7011 0.21894
8.323 0.98814 5.4661e-005 3.8183 0.011922 0.00010821 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5687 0.5731 0.17524 0.020203 17.0063 0.12521 0.00016348 0.76495 0.0093994 0.010399 0.0016224 0.98379 0.98948 3.5325e-006 1.413e-005 0.16483 0.67256 0.77288 0.0015173 0.79153 0.37139 0.0020395 0.41743 1.613 1.6095 16.0187 144.901 0.0003815 -84.7083 0.21994
8.324 0.98814 5.4661e-005 3.8183 0.011922 0.00010822 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5688 0.57314 0.17526 0.020204 17.0093 0.12522 0.00016349 0.76494 0.0093998 0.0104 0.0016205 0.98382 0.98951 3.528e-006 1.4112e-005 0.16484 0.67353 0.77362 0.0015164 0.79275 0.3716 0.0020382 0.41744 1.615 1.6115 16.0187 144.901 0.00038044 -84.7154 0.22094
8.325 0.98814 5.4661e-005 3.8183 0.011922 0.00010824 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5689 0.57319 0.17527 0.020205 17.0124 0.12523 0.0001635 0.76494 0.0094001 0.0104 0.0016185 0.98385 0.98953 3.5236e-006 1.4095e-005 0.16484 0.67449 0.77435 0.0015154 0.79395 0.37181 0.002037 0.41745 1.617 1.6135 16.0188 144.901 0.00037938 -84.7225 0.22194
8.326 0.98814 5.4661e-005 3.8183 0.011922 0.00010825 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.569 0.57323 0.17528 0.020206 17.0154 0.12523 0.00016351 0.76493 0.0094005 0.0104 0.0016166 0.98387 0.98955 3.5192e-006 1.4077e-005 0.16484 0.67545 0.77508 0.0015145 0.79515 0.37203 0.0020358 0.41745 1.619 1.6155 16.0188 144.901 0.00037834 -84.7295 0.22294
8.327 0.98814 5.4661e-005 3.8183 0.011922 0.00010826 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5691 0.57328 0.1753 0.020207 17.0185 0.12524 0.00016352 0.76492 0.0094009 0.010401 0.0016147 0.9839 0.98958 3.5148e-006 1.406e-005 0.16485 0.67641 0.77581 0.0015136 0.79635 0.37224 0.0020346 0.41746 1.621 1.6175 16.0189 144.901 0.00037729 -84.7365 0.22394
8.328 0.98814 5.4661e-005 3.8183 0.011922 0.00010827 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5692 0.57332 0.17531 0.020208 17.0215 0.12525 0.00016353 0.76492 0.0094013 0.010401 0.0016129 0.98392 0.9896 3.5105e-006 1.4043e-005 0.16485 0.67736 0.77653 0.0015127 0.79753 0.37245 0.0020334 0.41747 1.623 1.6195 16.0189 144.901 0.00037626 -84.7434 0.22494
8.329 0.98814 5.4661e-005 3.8183 0.011922 0.00010829 0.0011736 0.23371 0.00065931 0.23436 0.21627 0 0.032259 0.0389 0 1.5692 0.57336 0.17532 0.020209 17.0246 0.12525 0.00016354 0.76491 0.0094016 0.010402 0.001611 0.98395 0.98962 3.5063e-006 1.4026e-005 0.16485 0.67831 0.77725 0.0015118 0.79871 0.37266 0.0020322 0.41748 1.625 1.6215 16.019 144.9011 0.00037522 -84.7503 0.22594
8.33 0.98814 5.4661e-005 3.8183 0.011922 0.0001083 0.0011736 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5693 0.57341 0.17534 0.02021 17.0276 0.12526 0.00016355 0.7649 0.009402 0.010402 0.0016092 0.98397 0.98964 3.502e-006 1.4009e-005 0.16485 0.67926 0.77796 0.0015109 0.79989 0.37287 0.002031 0.41748 1.6269 1.6235 16.019 144.9011 0.0003742 -84.7571 0.22694
8.331 0.98814 5.4661e-005 3.8183 0.011922 0.00010831 0.0011736 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5694 0.57345 0.17535 0.020211 17.0307 0.12527 0.00016355 0.7649 0.0094024 0.010402 0.0016074 0.984 0.98966 3.4979e-006 1.3992e-005 0.16486 0.68021 0.77867 0.00151 0.80106 0.37309 0.0020299 0.41749 1.6289 1.6255 16.0191 144.9011 0.00037318 -84.7639 0.22794
8.332 0.98814 5.466e-005 3.8183 0.011922 0.00010833 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5695 0.5735 0.17536 0.020212 17.0337 0.12527 0.00016356 0.76489 0.0094028 0.010403 0.0016056 0.98402 0.98969 3.4937e-006 1.3975e-005 0.16486 0.68115 0.77937 0.0015091 0.80222 0.3733 0.0020287 0.4175 1.6309 1.6274 16.0191 144.9011 0.00037216 -84.7706 0.22894
8.333 0.98814 5.466e-005 3.8183 0.011922 0.00010834 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5696 0.57354 0.17538 0.020213 17.0368 0.12528 0.00016357 0.76488 0.0094031 0.010403 0.0016039 0.98405 0.98971 3.4896e-006 1.3959e-005 0.16486 0.68209 0.78007 0.0015082 0.80338 0.37351 0.0020276 0.41751 1.6328 1.6294 16.0191 144.9011 0.00037115 -84.7772 0.22994
8.334 0.98814 5.466e-005 3.8183 0.011922 0.00010835 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5697 0.57359 0.17539 0.020214 17.0398 0.12529 0.00016358 0.76488 0.0094035 0.010404 0.0016021 0.98407 0.98973 3.4855e-006 1.3943e-005 0.16487 0.68303 0.78077 0.0015073 0.80453 0.37372 0.0020264 0.41752 1.6348 1.6314 16.0192 144.9011 0.00037014 -84.7838 0.23094
8.335 0.98814 5.466e-005 3.8183 0.011922 0.00010836 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5698 0.57363 0.1754 0.020215 17.0429 0.12529 0.00016359 0.76487 0.0094039 0.010404 0.0016004 0.9841 0.98975 3.4815e-006 1.3926e-005 0.16487 0.68396 0.78146 0.0015065 0.80567 0.37394 0.0020253 0.41752 1.6367 1.6334 16.0192 144.9011 0.00036914 -84.7904 0.23194
8.336 0.98814 5.466e-005 3.8183 0.011922 0.00010838 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5698 0.57368 0.17542 0.020217 17.0459 0.1253 0.0001636 0.76487 0.0094042 0.010404 0.0015986 0.98412 0.98976 3.4775e-006 1.391e-005 0.16487 0.68489 0.78214 0.0015056 0.80681 0.37415 0.0020242 0.41753 1.6387 1.6353 16.0193 144.9012 0.00036814 -84.7969 0.23294
8.337 0.98814 5.466e-005 3.8183 0.011922 0.00010839 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5699 0.57372 0.17543 0.020218 17.049 0.1253 0.00016361 0.76486 0.0094046 0.010405 0.0015969 0.98414 0.98978 3.4735e-006 1.3894e-005 0.16487 0.68582 0.78283 0.0015048 0.80795 0.37436 0.0020231 0.41754 1.6406 1.6373 16.0193 144.9012 0.00036715 -84.8033 0.23394
8.338 0.98814 5.466e-005 3.8183 0.011922 0.0001084 0.0011737 0.23371 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.57 0.57377 0.17544 0.020219 17.0521 0.12531 0.00016362 0.76485 0.009405 0.010405 0.0015952 0.98417 0.9898 3.4696e-006 1.3879e-005 0.16488 0.68675 0.7835 0.0015039 0.80907 0.37457 0.002022 0.41755 1.6426 1.6392 16.0194 144.9012 0.00036616 -84.8097 0.23494
8.339 0.98814 5.466e-005 3.8183 0.011922 0.00010842 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5701 0.57381 0.17546 0.02022 17.0551 0.12532 0.00016363 0.76485 0.0094054 0.010406 0.0015935 0.98419 0.98982 3.4657e-006 1.3863e-005 0.16488 0.68767 0.78418 0.0015031 0.81019 0.37478 0.0020209 0.41756 1.6445 1.6412 16.0194 144.9012 0.00036518 -84.8161 0.23594
8.34 0.98814 5.466e-005 3.8183 0.011922 0.00010843 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5702 0.57386 0.17547 0.020221 17.0582 0.12532 0.00016364 0.76484 0.0094057 0.010406 0.0015919 0.98421 0.98984 3.4618e-006 1.3848e-005 0.16488 0.68859 0.78485 0.0015023 0.81131 0.375 0.0020198 0.41757 1.6464 1.6431 16.0195 144.9012 0.00036421 -84.8224 0.23694
8.341 0.98814 5.466e-005 3.8183 0.011922 0.00010844 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5703 0.5739 0.17548 0.020222 17.0612 0.12533 0.00016365 0.76483 0.0094061 0.010406 0.0015902 0.98424 0.98986 3.458e-006 1.3832e-005 0.16489 0.68951 0.78552 0.0015014 0.81242 0.37521 0.0020187 0.41757 1.6484 1.645 16.0195 144.9012 0.00036323 -84.8287 0.23794
8.342 0.98814 5.466e-005 3.8183 0.011922 0.00010845 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5704 0.57395 0.1755 0.020223 17.0643 0.12534 0.00016366 0.76483 0.0094065 0.010407 0.0015885 0.98426 0.98987 3.4542e-006 1.3817e-005 0.16489 0.69042 0.78618 0.0015006 0.81352 0.37542 0.0020176 0.41758 1.6503 1.647 16.0195 144.9012 0.00036227 -84.8349 0.23894
8.343 0.98814 5.466e-005 3.8183 0.011922 0.00010847 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5704 0.57399 0.17551 0.020224 17.0673 0.12534 0.00016367 0.76482 0.0094069 0.010407 0.0015869 0.98428 0.98989 3.4504e-006 1.3802e-005 0.16489 0.69133 0.78684 0.0014998 0.81462 0.37563 0.0020166 0.41759 1.6522 1.6489 16.0196 144.9013 0.0003613 -84.841 0.23994
8.344 0.98814 5.4659e-005 3.8183 0.011922 0.00010848 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5705 0.57404 0.17552 0.020225 17.0704 0.12535 0.00016368 0.76481 0.0094072 0.010408 0.0015853 0.9843 0.98991 3.4467e-006 1.3787e-005 0.16489 0.69224 0.78749 0.001499 0.81571 0.37584 0.0020155 0.4176 1.6541 1.6508 16.0196 144.9013 0.00036035 -84.8471 0.24094
8.345 0.98814 5.4659e-005 3.8183 0.011922 0.00010849 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5706 0.57408 0.17554 0.020226 17.0735 0.12536 0.00016369 0.76481 0.0094076 0.010408 0.0015837 0.98432 0.98993 3.443e-006 1.3772e-005 0.1649 0.69314 0.78814 0.0014982 0.81679 0.37605 0.0020145 0.41761 1.656 1.6528 16.0197 144.9013 0.00035939 -84.8532 0.24194
8.346 0.98814 5.4659e-005 3.8183 0.011922 0.00010851 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5707 0.57412 0.17555 0.020227 17.0765 0.12536 0.0001637 0.7648 0.009408 0.010408 0.0015821 0.98435 0.98994 3.4393e-006 1.3758e-005 0.1649 0.69405 0.78879 0.0014974 0.81787 0.37627 0.0020135 0.41762 1.6579 1.6547 16.0197 144.9013 0.00035845 -84.8592 0.24294
8.347 0.98814 5.4659e-005 3.8183 0.011922 0.00010852 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5708 0.57417 0.17556 0.020228 17.0796 0.12537 0.00016371 0.76479 0.0094083 0.010409 0.0015806 0.98437 0.98996 3.4357e-006 1.3743e-005 0.1649 0.69495 0.78943 0.0014966 0.81895 0.37648 0.0020124 0.41763 1.6598 1.6566 16.0198 144.9013 0.0003575 -84.8652 0.24394
8.348 0.98814 5.4659e-005 3.8183 0.011922 0.00010853 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5709 0.57421 0.17558 0.020229 17.0826 0.12538 0.00016372 0.76479 0.0094087 0.010409 0.001579 0.98439 0.98997 3.4321e-006 1.3729e-005 0.16491 0.69584 0.79007 0.0014959 0.82002 0.37669 0.0020114 0.41764 1.6617 1.6585 16.0198 144.9013 0.00035656 -84.8711 0.24494
8.349 0.98814 5.4659e-005 3.8183 0.011922 0.00010854 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.571 0.57426 0.17559 0.020231 17.0857 0.12538 0.00016373 0.76478 0.0094091 0.01041 0.0015774 0.98441 0.98999 3.4285e-006 1.3714e-005 0.16491 0.69674 0.79071 0.0014951 0.82108 0.3769 0.0020104 0.41764 1.6636 1.6604 16.0198 144.9013 0.00035563 -84.877 0.24594
8.35 0.98814 5.4659e-005 3.8183 0.011922 0.00010856 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.571 0.5743 0.1756 0.020232 17.0887 0.12539 0.00016374 0.76478 0.0094095 0.01041 0.0015759 0.98443 0.99001 3.425e-006 1.37e-005 0.16491 0.69763 0.79134 0.0014943 0.82213 0.37711 0.0020094 0.41765 1.6655 1.6623 16.0199 144.9014 0.0003547 -84.8828 0.24694
8.351 0.98814 5.4659e-005 3.8183 0.011922 0.00010857 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5711 0.57435 0.17562 0.020233 17.0918 0.12539 0.00016375 0.76477 0.0094098 0.01041 0.0015744 0.98445 0.99002 3.4215e-006 1.3686e-005 0.16491 0.69852 0.79197 0.0014936 0.82319 0.37733 0.0020084 0.41766 1.6674 1.6642 16.0199 144.9014 0.00035377 -84.8886 0.24794
8.352 0.98814 5.4659e-005 3.8183 0.011922 0.00010858 0.0011737 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5712 0.57439 0.17563 0.020234 17.0949 0.1254 0.00016376 0.76476 0.0094102 0.010411 0.0015729 0.98447 0.99004 3.418e-006 1.3672e-005 0.16492 0.69941 0.7926 0.0014928 0.82423 0.37754 0.0020074 0.41767 1.6693 1.6661 16.02 144.9014 0.00035285 -84.8944 0.24894
8.353 0.98814 5.4659e-005 3.8183 0.011922 0.00010859 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5713 0.57444 0.17564 0.020235 17.0979 0.12541 0.00016377 0.76476 0.0094106 0.010411 0.0015714 0.98449 0.99005 3.4145e-006 1.3659e-005 0.16492 0.70029 0.79322 0.0014921 0.82527 0.37775 0.0020065 0.41768 1.6711 1.6679 16.02 144.9014 0.00035194 -84.9001 0.24994
8.354 0.98814 5.4659e-005 3.8183 0.011922 0.00010861 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5714 0.57448 0.17566 0.020236 17.101 0.12541 0.00016378 0.76475 0.0094109 0.010411 0.0015699 0.98451 0.99007 3.4111e-006 1.3645e-005 0.16492 0.70117 0.79383 0.0014913 0.8263 0.37796 0.0020055 0.41769 1.673 1.6698 16.02 144.9014 0.00035103 -84.9057 0.25094
8.355 0.98814 5.4659e-005 3.8183 0.011922 0.00010862 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5715 0.57453 0.17567 0.020237 17.104 0.12542 0.00016379 0.76474 0.0094113 0.010412 0.0015684 0.98453 0.99008 3.4077e-006 1.3631e-005 0.16493 0.70205 0.79445 0.0014906 0.82733 0.37817 0.0020045 0.4177 1.6749 1.6717 16.0201 144.9014 0.00035012 -84.9114 0.25194
8.356 0.98814 5.4659e-005 3.8183 0.011922 0.00010863 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5716 0.57457 0.17568 0.020238 17.1071 0.12543 0.0001638 0.76474 0.0094117 0.010412 0.001567 0.98455 0.99009 3.4044e-006 1.3618e-005 0.16493 0.70292 0.79506 0.0014899 0.82836 0.37838 0.0020036 0.41771 1.6767 1.6736 16.0201 144.9014 0.00034922 -84.9169 0.25294
8.357 0.98814 5.4658e-005 3.8183 0.011922 0.00010865 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5716 0.57462 0.1757 0.020239 17.1102 0.12543 0.00016381 0.76473 0.0094121 0.010413 0.0015655 0.98457 0.99011 3.4011e-006 1.3605e-005 0.16493 0.7038 0.79567 0.0014892 0.82937 0.37859 0.0020027 0.41772 1.6786 1.6754 16.0202 144.9015 0.00034832 -84.9225 0.25394
8.358 0.98814 5.4658e-005 3.8183 0.011922 0.00010866 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5717 0.57466 0.17571 0.02024 17.1132 0.12544 0.00016382 0.76472 0.0094124 0.010413 0.0015641 0.98459 0.99012 3.3977e-006 1.3591e-005 0.16493 0.70467 0.79627 0.0014884 0.83038 0.37881 0.0020017 0.41773 1.6804 1.6773 16.0202 144.9015 0.00034743 -84.928 0.25494
8.359 0.98814 5.4658e-005 3.8183 0.011922 0.00010867 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5718 0.57471 0.17572 0.020241 17.1163 0.12545 0.00016383 0.76472 0.0094128 0.010413 0.0015627 0.98461 0.99014 3.3945e-006 1.3578e-005 0.16494 0.70553 0.79687 0.0014877 0.83139 0.37902 0.0020008 0.41774 1.6823 1.6791 16.0202 144.9015 0.00034654 -84.9334 0.25594
8.36 0.98814 5.4658e-005 3.8183 0.011922 0.00010868 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5719 0.57475 0.17574 0.020242 17.1194 0.12545 0.00016384 0.76471 0.0094132 0.010414 0.0015613 0.98463 0.99015 3.3912e-006 1.3565e-005 0.16494 0.7064 0.79747 0.001487 0.83239 0.37923 0.0019999 0.41775 1.6841 1.681 16.0203 144.9015 0.00034565 -84.9388 0.25694
8.361 0.98814 5.4658e-005 3.8183 0.011922 0.0001087 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.572 0.5748 0.17575 0.020243 17.1224 0.12546 0.00016385 0.7647 0.0094136 0.010414 0.0015599 0.98465 0.99016 3.388e-006 1.3552e-005 0.16494 0.70726 0.79806 0.0014863 0.83339 0.37944 0.001999 0.41776 1.6859 1.6828 16.0203 144.9015 0.00034477 -84.9442 0.25794
8.362 0.98814 5.4658e-005 3.8183 0.011921 0.00010871 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5721 0.57484 0.17576 0.020245 17.1255 0.12547 0.00016386 0.7647 0.0094139 0.010415 0.0015585 0.98467 0.99018 3.3848e-006 1.354e-005 0.16495 0.70812 0.79865 0.0014856 0.83438 0.37965 0.0019981 0.41777 1.6878 1.6847 16.0203 144.9015 0.00034389 -84.9495 0.25894
8.363 0.98814 5.4658e-005 3.8183 0.011921 0.00010872 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5721 0.57488 0.17578 0.020246 17.1285 0.12547 0.00016387 0.76469 0.0094143 0.010415 0.0015572 0.98469 0.99019 3.3817e-006 1.3527e-005 0.16495 0.70898 0.79924 0.001485 0.83536 0.37986 0.0019972 0.41778 1.6896 1.6865 16.0204 144.9016 0.00034302 -84.9548 0.25994
8.364 0.98814 5.4658e-005 3.8183 0.011921 0.00010874 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5722 0.57493 0.17579 0.020247 17.1316 0.12548 0.00016388 0.76469 0.0094147 0.010415 0.0015558 0.9847 0.9902 3.3785e-006 1.3514e-005 0.16495 0.70983 0.79982 0.0014843 0.83634 0.38007 0.0019963 0.41779 1.6914 1.6884 16.0204 144.9016 0.00034215 -84.96 0.26094
8.365 0.98814 5.4658e-005 3.8183 0.011921 0.00010875 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5723 0.57497 0.17581 0.020248 17.1347 0.12548 0.00016389 0.76468 0.009415 0.010416 0.0015544 0.98472 0.99022 3.3754e-006 1.3502e-005 0.16495 0.71068 0.8004 0.0014836 0.83731 0.38028 0.0019954 0.4178 1.6932 1.6902 16.0204 144.9016 0.00034129 -84.9652 0.26194
8.366 0.98814 5.4658e-005 3.8183 0.011921 0.00010876 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5724 0.57502 0.17582 0.020249 17.1377 0.12549 0.0001639 0.76467 0.0094154 0.010416 0.0015531 0.98474 0.99023 3.3723e-006 1.349e-005 0.16496 0.71153 0.80098 0.0014829 0.83828 0.3805 0.0019945 0.41781 1.6951 1.692 16.0205 144.9016 0.00034043 -84.9704 0.26294
8.367 0.98814 5.4658e-005 3.8183 0.011921 0.00010877 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5725 0.57506 0.17583 0.02025 17.1408 0.1255 0.00016391 0.76467 0.0094158 0.010417 0.0015518 0.98476 0.99024 3.3693e-006 1.3477e-005 0.16496 0.71238 0.80155 0.0014823 0.83924 0.38071 0.0019936 0.41782 1.6969 1.6938 16.0205 144.9016 0.00033957 -84.9755 0.26394
8.368 0.98814 5.4658e-005 3.8183 0.011921 0.00010879 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5726 0.57511 0.17585 0.020251 17.1439 0.1255 0.00016392 0.76466 0.0094162 0.010417 0.0015505 0.98478 0.99025 3.3662e-006 1.3465e-005 0.16496 0.71322 0.80213 0.0014816 0.8402 0.38092 0.0019928 0.41783 1.6987 1.6957 16.0206 144.9016 0.00033872 -84.9806 0.26494
8.369 0.98814 5.4657e-005 3.8183 0.011921 0.0001088 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5727 0.57515 0.17586 0.020252 17.1469 0.12551 0.00016393 0.76465 0.0094165 0.010417 0.0015492 0.98479 0.99027 3.3632e-006 1.3453e-005 0.16497 0.71406 0.80269 0.001481 0.84115 0.38113 0.0019919 0.41784 1.7005 1.6975 16.0206 144.9016 0.00033788 -84.9856 0.26594
8.37 0.98814 5.4657e-005 3.8183 0.011921 0.00010881 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5727 0.5752 0.17587 0.020253 17.15 0.12552 0.00016394 0.76465 0.0094169 0.010418 0.0015479 0.98481 0.99028 3.3603e-006 1.3441e-005 0.16497 0.7149 0.80326 0.0014803 0.8421 0.38134 0.0019911 0.41785 1.7023 1.6993 16.0206 144.9017 0.00033703 -84.9906 0.26694
8.371 0.98814 5.4657e-005 3.8183 0.011921 0.00010883 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5728 0.57524 0.17589 0.020254 17.1531 0.12552 0.00016394 0.76464 0.0094173 0.010418 0.0015466 0.98483 0.99029 3.3573e-006 1.343e-005 0.16497 0.71574 0.80382 0.0014797 0.84304 0.38155 0.0019902 0.41786 1.7041 1.7011 16.0207 144.9017 0.00033619 -84.9956 0.26794
8.372 0.98814 5.4657e-005 3.8183 0.011921 0.00010884 0.0011738 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5729 0.57529 0.1759 0.020255 17.1561 0.12553 0.00016395 0.76463 0.0094176 0.010419 0.0015453 0.98485 0.9903 3.3544e-006 1.3418e-005 0.16497 0.71657 0.80438 0.001479 0.84398 0.38176 0.0019894 0.41787 1.7059 1.7029 16.0207 144.9017 0.00033536 -85.0005 0.26894
8.373 0.98814 5.4657e-005 3.8183 0.011921 0.00010885 0.0011739 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.573 0.57533 0.17591 0.020256 17.1592 0.12554 0.00016396 0.76463 0.009418 0.010419 0.0015441 0.98486 0.99032 3.3515e-006 1.3406e-005 0.16498 0.7174 0.80493 0.0014784 0.84491 0.38197 0.0019886 0.41788 1.7076 1.7047 16.0207 144.9017 0.00033453 -85.0054 0.26994
8.374 0.98814 5.4657e-005 3.8183 0.011921 0.00010886 0.0011739 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5731 0.57538 0.17593 0.020257 17.1623 0.12554 0.00016397 0.76462 0.0094184 0.010419 0.0015428 0.98488 0.99033 3.3486e-006 1.3395e-005 0.16498 0.71823 0.80548 0.0014778 0.84584 0.38218 0.0019877 0.41789 1.7094 1.7065 16.0208 144.9017 0.0003337 -85.0103 0.27094
8.375 0.98814 5.4657e-005 3.8183 0.011921 0.00010888 0.0011739 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5732 0.57542 0.17594 0.020259 17.1653 0.12555 0.00016398 0.76462 0.0094188 0.01042 0.0015416 0.9849 0.99034 3.3457e-006 1.3383e-005 0.16498 0.71905 0.80603 0.0014771 0.84676 0.38239 0.0019869 0.4179 1.7112 1.7082 16.0208 144.9017 0.00033288 -85.0151 0.27194
8.376 0.98814 5.4657e-005 3.8183 0.011921 0.00010889 0.0011739 0.2337 0.00065931 0.23436 0.21626 0 0.032259 0.0389 0 1.5733 0.57547 0.17595 0.02026 17.1684 0.12555 0.00016399 0.76461 0.0094191 0.01042 0.0015403 0.98491 0.99035 3.3429e-006 1.3372e-005 0.16499 0.71988 0.80658 0.0014765 0.84767 0.38261 0.0019861 0.41791 1.713 1.71 16.0208 144.9017 0.00033206 -85.0199 0.27294
8.377 0.98814 5.4657e-005 3.8183 0.011921 0.0001089 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5733 0.57551 0.17597 0.020261 17.1715 0.12556 0.000164 0.7646 0.0094195 0.010421 0.0015391 0.98493 0.99036 3.3401e-006 1.3361e-005 0.16499 0.7207 0.80712 0.0014759 0.84858 0.38282 0.0019853 0.41792 1.7147 1.7118 16.0208 144.9018 0.00033125 -85.0246 0.27394
8.378 0.98814 5.4657e-005 3.8183 0.011921 0.00010891 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5734 0.57555 0.17598 0.020262 17.1745 0.12557 0.00016401 0.7646 0.0094199 0.010421 0.0015379 0.98494 0.99037 3.3373e-006 1.335e-005 0.16499 0.72151 0.80766 0.0014753 0.84949 0.38303 0.0019845 0.41793 1.7165 1.7136 16.0209 144.9018 0.00033043 -85.0293 0.27494
8.379 0.98814 5.4657e-005 3.8183 0.011921 0.00010893 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5735 0.5756 0.17599 0.020263 17.1776 0.12557 0.00016402 0.76459 0.0094202 0.010421 0.0015367 0.98496 0.99038 3.3346e-006 1.3339e-005 0.16499 0.72233 0.8082 0.0014747 0.85039 0.38324 0.0019837 0.41794 1.7182 1.7153 16.0209 144.9018 0.00032963 -85.034 0.27594
8.38 0.98814 5.4657e-005 3.8183 0.011921 0.00010894 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5736 0.57564 0.17601 0.020264 17.1807 0.12558 0.00016403 0.76458 0.0094206 0.010422 0.0015355 0.98498 0.9904 3.3318e-006 1.3328e-005 0.165 0.72314 0.80874 0.0014741 0.85128 0.38345 0.001983 0.41795 1.72 1.7171 16.0209 144.9018 0.00032882 -85.0387 0.27694
8.381 0.98814 5.4656e-005 3.8183 0.011921 0.00010895 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5737 0.57569 0.17602 0.020265 17.1837 0.12559 0.00016404 0.76458 0.009421 0.010422 0.0015343 0.98499 0.99041 3.3291e-006 1.3317e-005 0.165 0.72395 0.80927 0.0014735 0.85217 0.38366 0.0019822 0.41796 1.7217 1.7189 16.021 144.9018 0.00032803 -85.0433 0.27794
8.382 0.98814 5.4656e-005 3.8183 0.011921 0.00010897 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5738 0.57573 0.17603 0.020266 17.1868 0.12559 0.00016405 0.76457 0.0094213 0.010423 0.0015332 0.98501 0.99042 3.3264e-006 1.3306e-005 0.165 0.72476 0.8098 0.0014729 0.85306 0.38387 0.0019814 0.41797 1.7235 1.7206 16.021 144.9018 0.00032723 -85.0478 0.27894
8.383 0.98814 5.4656e-005 3.8183 0.011921 0.00010898 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5738 0.57578 0.17605 0.020267 17.1899 0.1256 0.00016406 0.76456 0.0094217 0.010423 0.001532 0.98502 0.99043 3.3238e-006 1.3295e-005 0.16501 0.72557 0.81032 0.0014723 0.85394 0.38408 0.0019806 0.41798 1.7252 1.7224 16.021 144.9019 0.00032644 -85.0524 0.27994
8.384 0.98814 5.4656e-005 3.8183 0.011921 0.00010899 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5739 0.57582 0.17606 0.020268 17.193 0.12561 0.00016407 0.76456 0.0094221 0.010423 0.0015309 0.98504 0.99044 3.3211e-006 1.3285e-005 0.16501 0.72637 0.81084 0.0014717 0.85481 0.38429 0.0019799 0.418 1.727 1.7241 16.0211 144.9019 0.00032565 -85.0569 0.28094
8.385 0.98814 5.4656e-005 3.8183 0.011921 0.000109 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.574 0.57587 0.17607 0.020269 17.196 0.12561 0.00016408 0.76455 0.0094225 0.010424 0.0015297 0.98505 0.99045 3.3185e-006 1.3274e-005 0.16501 0.72717 0.81137 0.0014712 0.85569 0.3845 0.0019791 0.41801 1.7287 1.7258 16.0211 144.9019 0.00032487 -85.0613 0.28194
8.386 0.98814 5.4656e-005 3.8183 0.011921 0.00010902 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5741 0.57591 0.17609 0.02027 17.1991 0.12562 0.00016409 0.76455 0.0094228 0.010424 0.0015286 0.98507 0.99046 3.3159e-006 1.3264e-005 0.16501 0.72797 0.81188 0.0014706 0.85655 0.38471 0.0019784 0.41802 1.7304 1.7276 16.0211 144.9019 0.00032409 -85.0658 0.28294
8.387 0.98814 5.4656e-005 3.8183 0.011921 0.00010903 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5742 0.57596 0.1761 0.020271 17.2022 0.12563 0.0001641 0.76454 0.0094232 0.010424 0.0015275 0.98509 0.99047 3.3133e-006 1.3253e-005 0.16502 0.72876 0.8124 0.00147 0.85741 0.38492 0.0019776 0.41803 1.7321 1.7293 16.0212 144.9019 0.00032331 -85.0702 0.28394
8.388 0.98814 5.4656e-005 3.8183 0.011921 0.00010904 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5743 0.576 0.17611 0.020272 17.2052 0.12563 0.00016411 0.76453 0.0094236 0.010425 0.0015264 0.9851 0.99048 3.3107e-006 1.3243e-005 0.16502 0.72956 0.81291 0.0014695 0.85827 0.38513 0.0019769 0.41804 1.7339 1.731 16.0212 144.9019 0.00032254 -85.0745 0.28494
8.389 0.98814 5.4656e-005 3.8183 0.011921 0.00010906 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5744 0.57605 0.17613 0.020274 17.2083 0.12564 0.00016412 0.76453 0.0094239 0.010425 0.0015253 0.98511 0.99049 3.3082e-006 1.3233e-005 0.16502 0.73035 0.81342 0.0014689 0.85912 0.38534 0.0019762 0.41805 1.7356 1.7328 16.0212 144.902 0.00032177 -85.0789 0.28594
8.39 0.98814 5.4656e-005 3.8183 0.011921 0.00010907 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5744 0.57609 0.17614 0.020275 17.2114 0.12564 0.00016413 0.76452 0.0094243 0.010426 0.0015242 0.98513 0.9905 3.3057e-006 1.3223e-005 0.16503 0.73113 0.81393 0.0014684 0.85996 0.38555 0.0019755 0.41806 1.7373 1.7345 16.0212 144.902 0.000321 -85.0832 0.28694
8.391 0.98814 5.4656e-005 3.8183 0.011921 0.00010908 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5745 0.57614 0.17615 0.020276 17.2145 0.12565 0.00016414 0.76451 0.0094247 0.010426 0.0015231 0.98514 0.99051 3.3032e-006 1.3213e-005 0.16503 0.73192 0.81443 0.0014678 0.86081 0.38576 0.0019747 0.41807 1.739 1.7362 16.0213 144.902 0.00032024 -85.0874 0.28794
8.392 0.98814 5.4656e-005 3.8183 0.011921 0.00010909 0.0011739 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5746 0.57618 0.17617 0.020277 17.2175 0.12566 0.00016415 0.76451 0.009425 0.010426 0.001522 0.98516 0.99052 3.3007e-006 1.3203e-005 0.16503 0.7327 0.81493 0.0014673 0.86164 0.38597 0.001974 0.41808 1.7407 1.7379 16.0213 144.902 0.00031948 -85.0917 0.28894
8.393 0.98814 5.4655e-005 3.8183 0.011921 0.00010911 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5747 0.57623 0.17618 0.020278 17.2206 0.12566 0.00016416 0.7645 0.0094254 0.010427 0.001521 0.98517 0.99053 3.2983e-006 1.3193e-005 0.16503 0.73348 0.81543 0.0014667 0.86247 0.38618 0.0019733 0.4181 1.7424 1.7396 16.0213 144.902 0.00031873 -85.0959 0.28994
8.394 0.98814 5.4655e-005 3.8183 0.011921 0.00010912 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5748 0.57627 0.17619 0.020279 17.2237 0.12567 0.00016417 0.76449 0.0094258 0.010427 0.0015199 0.98519 0.99054 3.2958e-006 1.3184e-005 0.16504 0.73426 0.81593 0.0014662 0.8633 0.38639 0.0019726 0.41811 1.7441 1.7413 16.0213 144.902 0.00031798 -85.1 0.29094
8.395 0.98814 5.4655e-005 3.8183 0.011921 0.00010913 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5749 0.57631 0.17621 0.02028 17.2267 0.12568 0.00016418 0.76449 0.0094262 0.010428 0.0015189 0.9852 0.99055 3.2934e-006 1.3174e-005 0.16504 0.73504 0.81642 0.0014657 0.86412 0.3866 0.0019719 0.41812 1.7458 1.743 16.0214 144.9021 0.00031723 -85.1042 0.29194
8.396 0.98814 5.4655e-005 3.8183 0.011921 0.00010915 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.575 0.57636 0.17622 0.020281 17.2298 0.12568 0.00016419 0.76448 0.0094265 0.010428 0.0015178 0.98521 0.99056 3.291e-006 1.3164e-005 0.16504 0.73581 0.81691 0.0014652 0.86494 0.38681 0.0019712 0.41813 1.7474 1.7447 16.0214 144.9021 0.00031648 -85.1083 0.29294
8.397 0.98814 5.4655e-005 3.8183 0.011921 0.00010916 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.575 0.5764 0.17623 0.020282 17.2329 0.12569 0.0001642 0.76448 0.0094269 0.010428 0.0015168 0.98523 0.99057 3.2886e-006 1.3155e-005 0.16505 0.73658 0.8174 0.0014646 0.86575 0.38702 0.0019706 0.41814 1.7491 1.7464 16.0214 144.9021 0.00031574 -85.1124 0.29394
8.398 0.98814 5.4655e-005 3.8183 0.011921 0.00010917 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5751 0.57645 0.17625 0.020283 17.236 0.1257 0.00016421 0.76447 0.0094273 0.010429 0.0015158 0.98524 0.99058 3.2863e-006 1.3145e-005 0.16505 0.73735 0.81788 0.0014641 0.86656 0.38723 0.0019699 0.41815 1.7508 1.7481 16.0215 144.9021 0.00031501 -85.1164 0.29494
8.399 0.98814 5.4655e-005 3.8183 0.011921 0.00010918 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5752 0.57649 0.17626 0.020284 17.239 0.1257 0.00016422 0.76446 0.0094276 0.010429 0.0015148 0.98526 0.99059 3.284e-006 1.3136e-005 0.16505 0.73812 0.81837 0.0014636 0.86736 0.38744 0.0019692 0.41816 1.7525 1.7497 16.0215 144.9021 0.00031427 -85.1204 0.29594
8.4 0.98814 5.4655e-005 3.8183 0.011921 0.0001092 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5753 0.57654 0.17627 0.020285 17.2421 0.12571 0.00016423 0.76446 0.009428 0.01043 0.0015138 0.98527 0.9906 3.2816e-006 1.3127e-005 0.16505 0.73888 0.81885 0.0014631 0.86816 0.38765 0.0019685 0.41818 1.7541 1.7514 16.0215 144.9021 0.00031354 -85.1244 0.29694
8.401 0.98814 5.4655e-005 3.8183 0.011921 0.00010921 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5754 0.57658 0.17629 0.020286 17.2452 0.12571 0.00016424 0.76445 0.0094284 0.01043 0.0015128 0.98528 0.9906 3.2793e-006 1.3118e-005 0.16506 0.73964 0.81933 0.0014626 0.86896 0.38786 0.0019679 0.41819 1.7558 1.7531 16.0215 144.9022 0.00031282 -85.1284 0.29794
8.402 0.98814 5.4655e-005 3.8183 0.011921 0.00010922 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5755 0.57663 0.1763 0.020287 17.2483 0.12572 0.00016425 0.76444 0.0094287 0.01043 0.0015118 0.9853 0.99061 3.2771e-006 1.3108e-005 0.16506 0.7404 0.8198 0.0014621 0.86975 0.38807 0.0019672 0.4182 1.7574 1.7547 16.0216 144.9022 0.00031209 -85.1323 0.29894
8.403 0.98814 5.4655e-005 3.8183 0.011921 0.00010924 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5756 0.57667 0.17631 0.020289 17.2514 0.12573 0.00016426 0.76444 0.0094291 0.010431 0.0015108 0.98531 0.99062 3.2748e-006 1.3099e-005 0.16506 0.74116 0.82028 0.0014616 0.87053 0.38828 0.0019666 0.41821 1.7591 1.7564 16.0216 144.9022 0.00031138 -85.1362 0.29994
8.404 0.98814 5.4655e-005 3.8183 0.011921 0.00010925 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5756 0.57672 0.17633 0.02029 17.2544 0.12573 0.00016427 0.76443 0.0094295 0.010431 0.0015098 0.98532 0.99063 3.2726e-006 1.309e-005 0.16507 0.74191 0.82075 0.0014611 0.87131 0.38849 0.0019659 0.41822 1.7607 1.7581 16.0216 144.9022 0.00031066 -85.1401 0.30094
8.405 0.98814 5.4654e-005 3.8183 0.011921 0.00010926 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5757 0.57676 0.17634 0.020291 17.2575 0.12574 0.00016428 0.76442 0.0094299 0.010432 0.0015089 0.98534 0.99064 3.2703e-006 1.3082e-005 0.16507 0.74267 0.82122 0.0014606 0.87209 0.3887 0.0019653 0.41824 1.7624 1.7597 16.0216 144.9022 0.00030995 -85.1439 0.30194
8.406 0.98814 5.4654e-005 3.8183 0.011921 0.00010927 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5758 0.57681 0.17635 0.020292 17.2606 0.12575 0.00016428 0.76442 0.0094302 0.010432 0.0015079 0.98535 0.99065 3.2681e-006 1.3073e-005 0.16507 0.74342 0.82168 0.0014601 0.87286 0.38891 0.0019646 0.41825 1.764 1.7614 16.0217 144.9022 0.00030924 -85.1477 0.30294
8.407 0.98814 5.4654e-005 3.8183 0.011921 0.00010929 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5759 0.57685 0.17637 0.020293 17.2637 0.12575 0.00016429 0.76441 0.0094306 0.010432 0.001507 0.98536 0.99066 3.266e-006 1.3064e-005 0.16507 0.74416 0.82215 0.0014596 0.87363 0.38912 0.001964 0.41826 1.7657 1.763 16.0217 144.9022 0.00030853 -85.1515 0.30394
8.408 0.98814 5.4654e-005 3.8183 0.011921 0.0001093 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.576 0.5769 0.17638 0.020294 17.2667 0.12576 0.0001643 0.7644 0.009431 0.010433 0.001506 0.98537 0.99067 3.2638e-006 1.3055e-005 0.16508 0.74491 0.82261 0.0014592 0.87439 0.38933 0.0019634 0.41827 1.7673 1.7647 16.0217 144.9023 0.00030783 -85.1553 0.30494
8.409 0.98814 5.4654e-005 3.8183 0.011921 0.00010931 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5761 0.57694 0.17639 0.020295 17.2698 0.12577 0.00016431 0.7644 0.0094313 0.010433 0.0015051 0.98539 0.99067 3.2616e-006 1.3047e-005 0.16508 0.74565 0.82307 0.0014587 0.87515 0.38954 0.0019628 0.41828 1.7689 1.7663 16.0217 144.9023 0.00030713 -85.159 0.30594
8.41 0.98814 5.4654e-005 3.8183 0.011921 0.00010932 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5761 0.57698 0.17641 0.020296 17.2729 0.12577 0.00016432 0.76439 0.0094317 0.010433 0.0015042 0.9854 0.99068 3.2595e-006 1.3038e-005 0.16508 0.74639 0.82352 0.0014582 0.87591 0.38975 0.0019621 0.41829 1.7705 1.7679 16.0217 144.9023 0.00030643 -85.1627 0.30694
8.411 0.98814 5.4654e-005 3.8183 0.011921 0.00010934 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5762 0.57703 0.17642 0.020297 17.276 0.12578 0.00016433 0.76439 0.0094321 0.010434 0.0015032 0.98541 0.99069 3.2574e-006 1.303e-005 0.16509 0.74713 0.82398 0.0014577 0.87665 0.38996 0.0019615 0.41831 1.7722 1.7695 16.0218 144.9023 0.00030574 -85.1663 0.30794
8.412 0.98814 5.4654e-005 3.8183 0.011921 0.00010935 0.001174 0.2337 0.00065931 0.23435 0.21626 0 0.032259 0.0389 0 1.5763 0.57707 0.17643 0.020298 17.2791 0.12578 0.00016434 0.76438 0.0094324 0.010434 0.0015023 0.98542 0.9907 3.2553e-006 1.3021e-005 0.16509 0.74787 0.82443 0.0014573 0.8774 0.39017 0.0019609 0.41832 1.7738 1.7712 16.0218 144.9023 0.00030505 -85.17 0.30894
8.413 0.98814 5.4654e-005 3.8183 0.011921 0.00010936 0.0011741 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5764 0.57712 0.17645 0.020299 17.2821 0.12579 0.00016435 0.76437 0.0094328 0.010435 0.0015014 0.98543 0.99071 3.2532e-006 1.3013e-005 0.16509 0.7486 0.82488 0.0014568 0.87814 0.39038 0.0019603 0.41833 1.7754 1.7728 16.0218 144.9024 0.00030436 -85.1736 0.30994
8.414 0.98814 5.4654e-005 3.8183 0.011921 0.00010938 0.0011741 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5765 0.57716 0.17646 0.0203 17.2852 0.1258 0.00016436 0.76437 0.0094332 0.010435 0.0015005 0.98545 0.99072 3.2511e-006 1.3005e-005 0.16509 0.74933 0.82533 0.0014563 0.87888 0.39058 0.0019597 0.41834 1.777 1.7744 16.0218 144.9024 0.00030368 -85.1772 0.31094
8.415 0.98814 5.4654e-005 3.8183 0.011921 0.00010939 0.0011741 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5766 0.57721 0.17647 0.020301 17.2883 0.1258 0.00016437 0.76436 0.0094335 0.010435 0.0014996 0.98546 0.99072 3.2491e-006 1.2997e-005 0.1651 0.75006 0.82577 0.0014559 0.87961 0.39079 0.0019591 0.41836 1.7786 1.776 16.0219 144.9024 0.000303 -85.1808 0.31194
8.416 0.98814 5.4654e-005 3.8183 0.011921 0.0001094 0.0011741 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5767 0.57725 0.17649 0.020302 17.2914 0.12581 0.00016438 0.76435 0.0094339 0.010436 0.0014987 0.98547 0.99073 3.2471e-006 1.2988e-005 0.1651 0.75079 0.82622 0.0014554 0.88034 0.391 0.0019585 0.41837 1.7802 1.7776 16.0219 144.9024 0.00030232 -85.1843 0.31294
8.417 0.98814 5.4653e-005 3.8183 0.011921 0.00010941 0.0011741 0.2337 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5767 0.5773 0.1765 0.020303 17.2945 0.12582 0.00016439 0.76435 0.0094343 0.010436 0.0014979 0.98548 0.99074 3.245e-006 1.298e-005 0.1651 0.75151 0.82666 0.001455 0.88106 0.39121 0.001958 0.41838 1.7818 1.7792 16.0219 144.9024 0.00030165 -85.1878 0.31394
8.418 0.98814 5.4653e-005 3.8183 0.01192 0.00010943 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5768 0.57734 0.17651 0.020305 17.2975 0.12582 0.0001644 0.76434 0.0094346 0.010437 0.001497 0.98549 0.99075 3.243e-006 1.2972e-005 0.16511 0.75224 0.8271 0.0014546 0.88178 0.39142 0.0019574 0.41839 1.7834 1.7808 16.0219 144.9024 0.00030098 -85.1913 0.31494
8.419 0.98814 5.4653e-005 3.8183 0.01192 0.00010944 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5769 0.57739 0.17653 0.020306 17.3006 0.12583 0.00016441 0.76433 0.009435 0.010437 0.0014961 0.9855 0.99075 3.2411e-006 1.2964e-005 0.16511 0.75296 0.82753 0.0014541 0.8825 0.39163 0.0019568 0.4184 1.785 1.7824 16.0219 144.9025 0.00030031 -85.1947 0.31594
8.42 0.98814 5.4653e-005 3.8183 0.01192 0.00010945 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.577 0.57743 0.17654 0.020307 17.3037 0.12584 0.00016442 0.76433 0.0094354 0.010437 0.0014953 0.98552 0.99076 3.2391e-006 1.2957e-005 0.16511 0.75368 0.82797 0.0014537 0.88321 0.39184 0.0019562 0.41842 1.7865 1.784 16.022 144.9025 0.00029965 -85.1982 0.31694
8.421 0.98814 5.4653e-005 3.8183 0.01192 0.00010947 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5771 0.57748 0.17655 0.020308 17.3068 0.12584 0.00016443 0.76432 0.0094358 0.010438 0.0014944 0.98553 0.99077 3.2371e-006 1.2949e-005 0.16511 0.75439 0.8284 0.0014532 0.88392 0.39205 0.0019557 0.41843 1.7881 1.7856 16.022 144.9025 0.00029899 -85.2016 0.31794
8.422 0.98814 5.4653e-005 3.8183 0.01192 0.00010948 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5772 0.57752 0.17657 0.020309 17.3099 0.12585 0.00016444 0.76432 0.0094361 0.010438 0.0014936 0.98554 0.99078 3.2352e-006 1.2941e-005 0.16512 0.75511 0.82883 0.0014528 0.88462 0.39226 0.0019551 0.41844 1.7897 1.7872 16.022 144.9025 0.00029833 -85.2049 0.31894
8.423 0.98814 5.4653e-005 3.8183 0.01192 0.00010949 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5773 0.57756 0.17658 0.02031 17.313 0.12585 0.00016445 0.76431 0.0094365 0.010439 0.0014927 0.98555 0.99078 3.2333e-006 1.2933e-005 0.16512 0.75582 0.82926 0.0014524 0.88532 0.39246 0.0019545 0.41845 1.7912 1.7887 16.022 144.9025 0.00029767 -85.2083 0.31994
8.424 0.98814 5.4653e-005 3.8183 0.01192 0.0001095 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5773 0.57761 0.17659 0.020311 17.316 0.12586 0.00016446 0.7643 0.0094369 0.010439 0.0014919 0.98556 0.99079 3.2314e-006 1.2926e-005 0.16512 0.75653 0.82968 0.001452 0.88601 0.39267 0.001954 0.41847 1.7928 1.7903 16.022 144.9025 0.00029702 -85.2116 0.32094
8.425 0.98814 5.4653e-005 3.8183 0.01192 0.00010952 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5774 0.57765 0.17661 0.020312 17.3191 0.12587 0.00016447 0.7643 0.0094372 0.010439 0.0014911 0.98557 0.9908 3.2295e-006 1.2918e-005 0.16513 0.75723 0.83011 0.0014515 0.8867 0.39288 0.0019534 0.41848 1.7944 1.7919 16.0221 144.9026 0.00029637 -85.2149 0.32194
8.426 0.98814 5.4653e-005 3.8183 0.01192 0.00010953 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5775 0.5777 0.17662 0.020313 17.3222 0.12587 0.00016448 0.76429 0.0094376 0.01044 0.0014903 0.98558 0.99081 3.2276e-006 1.2911e-005 0.16513 0.75794 0.83053 0.0014511 0.88739 0.39309 0.0019529 0.41849 1.7959 1.7934 16.0221 144.9026 0.00029573 -85.2182 0.32294
8.427 0.98814 5.4653e-005 3.8183 0.01192 0.00010954 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5776 0.57774 0.17663 0.020314 17.3253 0.12588 0.00016449 0.76428 0.009438 0.01044 0.0014895 0.98559 0.99081 3.2258e-006 1.2903e-005 0.16513 0.75864 0.83095 0.0014507 0.88807 0.3933 0.0019524 0.4185 1.7975 1.795 16.0221 144.9026 0.00029508 -85.2215 0.32394
8.428 0.98814 5.4653e-005 3.8183 0.01192 0.00010956 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5777 0.57779 0.17665 0.020315 17.3284 0.12589 0.0001645 0.76428 0.0094383 0.010441 0.0014887 0.9856 0.99082 3.2239e-006 1.2896e-005 0.16513 0.75934 0.83136 0.0014503 0.88875 0.39351 0.0019518 0.41852 1.799 1.7966 16.0221 144.9026 0.00029444 -85.2247 0.32494
8.429 0.98814 5.4652e-005 3.8183 0.01192 0.00010957 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5778 0.57783 0.17666 0.020316 17.3315 0.12589 0.00016451 0.76427 0.0094387 0.010441 0.0014879 0.98561 0.99083 3.2221e-006 1.2889e-005 0.16514 0.76004 0.83178 0.0014499 0.88943 0.39372 0.0019513 0.41853 1.8006 1.7981 16.0221 144.9026 0.00029381 -85.2279 0.32594
8.43 0.98814 5.4652e-005 3.8183 0.01192 0.00010958 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5778 0.57788 0.17667 0.020317 17.3346 0.1259 0.00016452 0.76427 0.0094391 0.010441 0.0014871 0.98563 0.99084 3.2203e-006 1.2881e-005 0.16514 0.76074 0.83219 0.0014495 0.8901 0.39392 0.0019508 0.41854 1.8021 1.7997 16.0222 144.9026 0.00029317 -85.2311 0.32694
8.431 0.98814 5.4652e-005 3.8183 0.01192 0.00010959 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.032259 0.0389 0 1.5779 0.57792 0.17669 0.020318 17.3376 0.12591 0.00016453 0.76426 0.0094394 0.010442 0.0014863 0.98564 0.99084 3.2185e-006 1.2874e-005 0.16514 0.76143 0.8326 0.0014491 0.89077 0.39413 0.0019502 0.41855 1.8036 1.8012 16.0222 144.9027 0.00029254 -85.2342 0.32794
8.432 0.98814 5.4652e-005 3.8183 0.01192 0.00010961 0.0011741 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.578 0.57797 0.1767 0.02032 17.3407 0.12591 0.00016454 0.76425 0.0094398 0.010442 0.0014855 0.98565 0.99085 3.2167e-006 1.2867e-005 0.16514 0.76212 0.83301 0.0014487 0.89143 0.39434 0.0019497 0.41857 1.8052 1.8027 16.0222 144.9027 0.00029191 -85.2374 0.32894
8.433 0.98814 5.4652e-005 3.8183 0.01192 0.00010962 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5781 0.57801 0.17671 0.020321 17.3438 0.12592 0.00016455 0.76425 0.0094402 0.010442 0.0014848 0.98566 0.99086 3.2149e-006 1.286e-005 0.16515 0.76281 0.83342 0.0014483 0.89209 0.39455 0.0019492 0.41858 1.8067 1.8043 16.0222 144.9027 0.00029129 -85.2405 0.32994
8.434 0.98814 5.4652e-005 3.8183 0.01192 0.00010963 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5782 0.57806 0.17673 0.020322 17.3469 0.12592 0.00016456 0.76424 0.0094405 0.010443 0.001484 0.98567 0.99086 3.2132e-006 1.2853e-005 0.16515 0.7635 0.83383 0.0014479 0.89274 0.39476 0.0019487 0.41859 1.8082 1.8058 16.0222 144.9027 0.00029067 -85.2436 0.33094
8.435 0.98814 5.4652e-005 3.8183 0.01192 0.00010964 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5783 0.5781 0.17674 0.020323 17.35 0.12593 0.00016457 0.76423 0.0094409 0.010443 0.0014832 0.98568 0.99087 3.2114e-006 1.2846e-005 0.16515 0.76418 0.83423 0.0014475 0.89339 0.39497 0.0019482 0.41861 1.8097 1.8073 16.0222 144.9027 0.00029005 -85.2466 0.33194
8.436 0.98814 5.4652e-005 3.8183 0.01192 0.00010966 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5784 0.57815 0.17675 0.020324 17.3531 0.12594 0.00016458 0.76423 0.0094413 0.010444 0.0014825 0.98569 0.99088 3.2097e-006 1.2839e-005 0.16516 0.76487 0.83463 0.0014471 0.89404 0.39517 0.0019477 0.41862 1.8113 1.8089 16.0223 144.9027 0.00028943 -85.2497 0.33294
8.437 0.98814 5.4652e-005 3.8183 0.01192 0.00010967 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5784 0.57819 0.17677 0.020325 17.3562 0.12594 0.00016459 0.76422 0.0094416 0.010444 0.0014817 0.9857 0.99088 3.208e-006 1.2832e-005 0.16516 0.76555 0.83503 0.0014467 0.89468 0.39538 0.0019472 0.41863 1.8128 1.8104 16.0223 144.9028 0.00028882 -85.2527 0.33394
8.438 0.98814 5.4652e-005 3.8183 0.01192 0.00010968 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5785 0.57823 0.17678 0.020326 17.3592 0.12595 0.00016459 0.76421 0.009442 0.010444 0.001481 0.98571 0.99089 3.2063e-006 1.2825e-005 0.16516 0.76623 0.83543 0.0014463 0.89532 0.39559 0.0019467 0.41864 1.8143 1.8119 16.0223 144.9028 0.0002882 -85.2557 0.33494
8.439 0.98814 5.4652e-005 3.8183 0.01192 0.0001097 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5786 0.57828 0.17679 0.020327 17.3623 0.12596 0.0001646 0.76421 0.0094424 0.010445 0.0014802 0.98572 0.9909 3.2046e-006 1.2819e-005 0.16516 0.76691 0.83582 0.001446 0.89596 0.3958 0.0019462 0.41866 1.8158 1.8134 16.0223 144.9028 0.0002876 -85.2587 0.33594
8.44 0.98814 5.4652e-005 3.8183 0.01192 0.00010971 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5787 0.57832 0.17681 0.020328 17.3654 0.12596 0.00016461 0.7642 0.0094427 0.010445 0.0014795 0.98573 0.9909 3.2029e-006 1.2812e-005 0.16517 0.76758 0.83622 0.0014456 0.89659 0.39601 0.0019457 0.41867 1.8173 1.8149 16.0223 144.9028 0.00028699 -85.2616 0.33694
8.441 0.98814 5.4651e-005 3.8183 0.01192 0.00010972 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5788 0.57837 0.17682 0.020329 17.3685 0.12597 0.00016462 0.7642 0.0094431 0.010446 0.0014788 0.98573 0.99091 3.2013e-006 1.2805e-005 0.16517 0.76825 0.83661 0.0014452 0.89722 0.39621 0.0019452 0.41868 1.8188 1.8164 16.0223 144.9028 0.00028639 -85.2645 0.33794
8.442 0.98814 5.4651e-005 3.8183 0.01192 0.00010973 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5789 0.57841 0.17683 0.02033 17.3716 0.12598 0.00016463 0.76419 0.0094435 0.010446 0.0014781 0.98574 0.99091 3.1996e-006 1.2799e-005 0.16517 0.76892 0.837 0.0014449 0.89785 0.39642 0.0019447 0.4187 1.8203 1.8179 16.0224 144.9028 0.00028579 -85.2675 0.33894
8.443 0.98814 5.4651e-005 3.8183 0.01192 0.00010975 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.579 0.57846 0.17684 0.020331 17.3747 0.12598 0.00016464 0.76418 0.0094438 0.010446 0.0014774 0.98575 0.99092 3.198e-006 1.2792e-005 0.16518 0.76959 0.83739 0.0014445 0.89847 0.39663 0.0019443 0.41871 1.8217 1.8194 16.0224 144.9029 0.00028519 -85.2703 0.33994
8.444 0.98814 5.4651e-005 3.8183 0.01192 0.00010976 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.579 0.5785 0.17686 0.020332 17.3778 0.12599 0.00016465 0.76418 0.0094442 0.010447 0.0014767 0.98576 0.99093 3.1964e-006 1.2786e-005 0.16518 0.77026 0.83777 0.0014441 0.89908 0.39684 0.0019438 0.41872 1.8232 1.8209 16.0224 144.9029 0.0002846 -85.2732 0.34094
8.445 0.98814 5.4651e-005 3.8183 0.01192 0.00010977 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5791 0.57855 0.17687 0.020333 17.3809 0.12599 0.00016466 0.76417 0.0094446 0.010447 0.001476 0.98577 0.99093 3.1948e-006 1.2779e-005 0.16518 0.77092 0.83816 0.0014438 0.8997 0.39704 0.0019433 0.41874 1.8247 1.8224 16.0224 144.9029 0.00028401 -85.276 0.34194
8.446 0.98814 5.4651e-005 3.8183 0.01192 0.00010979 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5792 0.57859 0.17688 0.020334 17.384 0.126 0.00016467 0.76416 0.0094449 0.010448 0.0014753 0.98578 0.99094 3.1932e-006 1.2773e-005 0.16518 0.77159 0.83854 0.0014434 0.90031 0.39725 0.0019429 0.41875 1.8262 1.8239 16.0224 144.9029 0.00028342 -85.2789 0.34294
8.447 0.98814 5.4651e-005 3.8183 0.01192 0.0001098 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5793 0.57864 0.1769 0.020336 17.3871 0.12601 0.00016468 0.76416 0.0094453 0.010448 0.0014746 0.98579 0.99095 3.1916e-006 1.2766e-005 0.16519 0.77225 0.83892 0.0014431 0.90091 0.39746 0.0019424 0.41876 1.8277 1.8253 16.0224 144.9029 0.00028283 -85.2817 0.34394
8.448 0.98814 5.4651e-005 3.8183 0.01192 0.00010981 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5794 0.57868 0.17691 0.020337 17.3901 0.12601 0.00016469 0.76415 0.0094457 0.010448 0.0014739 0.9858 0.99095 3.19e-006 1.276e-005 0.16519 0.7729 0.8393 0.0014427 0.90152 0.39767 0.0019419 0.41877 1.8291 1.8268 16.0224 144.903 0.00028225 -85.2845 0.34494
8.449 0.98814 5.4651e-005 3.8183 0.01192 0.00010982 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5795 0.57873 0.17692 0.020338 17.3932 0.12602 0.0001647 0.76414 0.009446 0.010449 0.0014732 0.98581 0.99096 3.1884e-006 1.2754e-005 0.16519 0.77356 0.83968 0.0014424 0.90211 0.39787 0.0019415 0.41879 1.8306 1.8283 16.0225 144.903 0.00028167 -85.2872 0.34594
8.45 0.98814 5.4651e-005 3.8183 0.01192 0.00010984 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5795 0.57877 0.17694 0.020339 17.3963 0.12603 0.00016471 0.76414 0.0094464 0.010449 0.0014725 0.98582 0.99096 3.1869e-006 1.2748e-005 0.1652 0.77422 0.84005 0.001442 0.90271 0.39808 0.001941 0.4188 1.832 1.8298 16.0225 144.903 0.00028109 -85.29 0.34694
8.451 0.98814 5.4651e-005 3.8183 0.01192 0.00010985 0.0011742 0.23369 0.00065931 0.23435 0.21625 0 0.03226 0.0389 0 1.5796 0.57881 0.17695 0.02034 17.3994 0.12603 0.00016472 0.76413 0.0094468 0.010449 0.0014719 0.98583 0.99097 3.1854e-006 1.2742e-005 0.1652 0.77487 0.84043 0.0014417 0.9033 0.39829 0.0019406 0.41881 1.8335 1.8312 16.0225 144.903 0.00028051 -85.2927 0.34794
8.452 0.98814 5.4651e-005 3.8183 0.01192 0.00010986 0.0011742 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5797 0.57886 0.17696 0.020341 17.4025 0.12604 0.00016473 0.76413 0.0094471 0.01045 0.0014712 0.98584 0.99098 3.1838e-006 1.2735e-005 0.1652 0.77552 0.8408 0.0014413 0.90389 0.3985 0.0019401 0.41883 1.8349 1.8327 16.0225 144.903 0.00027994 -85.2954 0.34894
8.453 0.98814 5.465e-005 3.8183 0.01192 0.00010988 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5798 0.5789 0.17698 0.020342 17.4056 0.12605 0.00016474 0.76412 0.0094475 0.01045 0.0014706 0.98584 0.99098 3.1823e-006 1.2729e-005 0.1652 0.77617 0.84117 0.001441 0.90448 0.3987 0.0019397 0.41884 1.8364 1.8341 16.0225 144.903 0.00027937 -85.2981 0.34994
8.454 0.98814 5.465e-005 3.8183 0.01192 0.00010989 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5799 0.57895 0.17699 0.020343 17.4087 0.12605 0.00016475 0.76411 0.0094479 0.010451 0.0014699 0.98585 0.99099 3.1808e-006 1.2723e-005 0.16521 0.77681 0.84154 0.0014407 0.90506 0.39891 0.0019392 0.41885 1.8378 1.8356 16.0225 144.9031 0.0002788 -85.3007 0.35094
8.455 0.98814 5.465e-005 3.8183 0.01192 0.0001099 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.58 0.57899 0.177 0.020344 17.4118 0.12606 0.00016476 0.76411 0.0094482 0.010451 0.0014693 0.98586 0.99099 3.1794e-006 1.2717e-005 0.16521 0.77746 0.8419 0.0014403 0.90563 0.39912 0.0019388 0.41887 1.8393 1.837 16.0225 144.9031 0.00027824 -85.3034 0.35194
8.456 0.98814 5.465e-005 3.8183 0.01192 0.00010991 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5801 0.57904 0.17702 0.020345 17.4149 0.12606 0.00016477 0.7641 0.0094486 0.010451 0.0014686 0.98587 0.991 3.1779e-006 1.2712e-005 0.16521 0.7781 0.84227 0.00144 0.90621 0.39932 0.0019384 0.41888 1.8407 1.8385 16.0226 144.9031 0.00027767 -85.306 0.35294
8.457 0.98814 5.465e-005 3.8183 0.01192 0.00010993 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5801 0.57908 0.17703 0.020346 17.418 0.12607 0.00016478 0.76409 0.009449 0.010452 0.001468 0.98588 0.991 3.1764e-006 1.2706e-005 0.16522 0.77874 0.84263 0.0014397 0.90678 0.39953 0.001938 0.41889 1.8421 1.8399 16.0226 144.9031 0.00027711 -85.3086 0.35394
8.458 0.98814 5.465e-005 3.8183 0.01192 0.00010994 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5802 0.57913 0.17704 0.020347 17.4211 0.12608 0.00016479 0.76409 0.0094493 0.010452 0.0014673 0.98589 0.99101 3.175e-006 1.27e-005 0.16522 0.77938 0.84299 0.0014393 0.90735 0.39974 0.0019375 0.41891 1.8436 1.8413 16.0226 144.9031 0.00027656 -85.3112 0.35494
8.459 0.98814 5.465e-005 3.8183 0.01192 0.00010995 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5803 0.57917 0.17706 0.020348 17.4242 0.12608 0.0001648 0.76408 0.0094497 0.010453 0.0014667 0.98589 0.99102 3.1735e-006 1.2694e-005 0.16522 0.78001 0.84335 0.001439 0.90791 0.39995 0.0019371 0.41892 1.845 1.8428 16.0226 144.9031 0.000276 -85.3137 0.35594
8.46 0.98814 5.465e-005 3.8183 0.01192 0.00010996 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5804 0.57922 0.17707 0.020349 17.4273 0.12609 0.00016481 0.76407 0.0094501 0.010453 0.0014661 0.9859 0.99102 3.1721e-006 1.2688e-005 0.16522 0.78065 0.84371 0.0014387 0.90847 0.40015 0.0019367 0.41893 1.8464 1.8442 16.0226 144.9032 0.00027545 -85.3163 0.35694
8.461 0.98814 5.465e-005 3.8183 0.01192 0.00010998 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5805 0.57926 0.17708 0.02035 17.4304 0.1261 0.00016482 0.76407 0.0094504 0.010453 0.0014655 0.98591 0.99103 3.1707e-006 1.2683e-005 0.16523 0.78128 0.84407 0.0014384 0.90903 0.40036 0.0019363 0.41895 1.8478 1.8456 16.0226 144.9032 0.0002749 -85.3188 0.35794
8.462 0.98814 5.465e-005 3.8183 0.01192 0.00010999 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5806 0.57931 0.1771 0.020351 17.4335 0.1261 0.00016483 0.76406 0.0094508 0.010454 0.0014649 0.98592 0.99103 3.1693e-006 1.2677e-005 0.16523 0.78191 0.84442 0.0014381 0.90958 0.40057 0.0019359 0.41896 1.8492 1.8471 16.0226 144.9032 0.00027435 -85.3213 0.35894
8.463 0.98814 5.465e-005 3.8183 0.01192 0.00011 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5806 0.57935 0.17711 0.020353 17.4366 0.12611 0.00016484 0.76406 0.0094512 0.010454 0.0014643 0.98593 0.99104 3.1679e-006 1.2672e-005 0.16523 0.78254 0.84478 0.0014378 0.91013 0.40077 0.0019354 0.41897 1.8507 1.8485 16.0226 144.9032 0.00027381 -85.3238 0.35994
8.464 0.98814 5.465e-005 3.8183 0.01192 0.00011002 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5807 0.57939 0.17712 0.020354 17.4397 0.12612 0.00016485 0.76405 0.0094515 0.010455 0.0014637 0.98593 0.99104 3.1665e-006 1.2666e-005 0.16524 0.78317 0.84513 0.0014375 0.91068 0.40098 0.001935 0.41899 1.8521 1.8499 16.0226 144.9032 0.00027326 -85.3263 0.36094
8.465 0.98814 5.4649e-005 3.8183 0.01192 0.00011003 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5808 0.57944 0.17714 0.020355 17.4428 0.12612 0.00016486 0.76404 0.0094519 0.010455 0.0014631 0.98594 0.99105 3.1651e-006 1.2661e-005 0.16524 0.78379 0.84548 0.0014371 0.91123 0.40119 0.0019346 0.419 1.8535 1.8513 16.0227 144.9033 0.00027272 -85.3287 0.36194
8.466 0.98814 5.4649e-005 3.8183 0.01192 0.00011004 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5809 0.57948 0.17715 0.020356 17.4459 0.12613 0.00016487 0.76404 0.0094523 0.010455 0.0014625 0.98595 0.99105 3.1638e-006 1.2655e-005 0.16524 0.78441 0.84583 0.0014368 0.91177 0.40139 0.0019342 0.41902 1.8549 1.8527 16.0227 144.9033 0.00027219 -85.3311 0.36294
8.467 0.98814 5.4649e-005 3.8183 0.01192 0.00011005 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.581 0.57953 0.17716 0.020357 17.449 0.12613 0.00016487 0.76403 0.0094526 0.010456 0.0014619 0.98596 0.99106 3.1624e-006 1.265e-005 0.16524 0.78503 0.84617 0.0014365 0.9123 0.4016 0.0019338 0.41903 1.8562 1.8541 16.0227 144.9033 0.00027165 -85.3336 0.36394
8.468 0.98814 5.4649e-005 3.8183 0.01192 0.00011007 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5811 0.57957 0.17718 0.020358 17.4521 0.12614 0.00016488 0.76402 0.009453 0.010456 0.0014613 0.98597 0.99106 3.1611e-006 1.2644e-005 0.16525 0.78565 0.84652 0.0014362 0.91284 0.40181 0.0019334 0.41904 1.8576 1.8555 16.0227 144.9033 0.00027112 -85.3359 0.36494
8.469 0.98814 5.4649e-005 3.8183 0.01192 0.00011008 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5812 0.57962 0.17719 0.020359 17.4551 0.12615 0.00016489 0.76402 0.0094534 0.010456 0.0014607 0.98597 0.99107 3.1597e-006 1.2639e-005 0.16525 0.78627 0.84686 0.0014359 0.91337 0.40201 0.0019331 0.41906 1.859 1.8569 16.0227 144.9033 0.00027059 -85.3383 0.36594
8.47 0.98814 5.4649e-005 3.8183 0.01192 0.00011009 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5812 0.57966 0.1772 0.02036 17.4582 0.12615 0.0001649 0.76401 0.0094537 0.010457 0.0014601 0.98598 0.99107 3.1584e-006 1.2634e-005 0.16525 0.78688 0.8472 0.0014356 0.9139 0.40222 0.0019327 0.41907 1.8604 1.8583 16.0227 144.9033 0.00027006 -85.3407 0.36694
8.471 0.98814 5.4649e-005 3.8183 0.01192 0.00011011 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5813 0.57971 0.17722 0.020361 17.4613 0.12616 0.00016491 0.76401 0.0094541 0.010457 0.0014596 0.98599 0.99108 3.1571e-006 1.2628e-005 0.16525 0.7875 0.84754 0.0014353 0.91442 0.40242 0.0019323 0.41908 1.8618 1.8597 16.0227 144.9034 0.00026953 -85.343 0.36794
8.472 0.98814 5.4649e-005 3.8183 0.01192 0.00011012 0.0011743 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5814 0.57975 0.17723 0.020362 17.4644 0.12617 0.00016492 0.764 0.0094545 0.010458 0.001459 0.986 0.99108 3.1558e-006 1.2623e-005 0.16526 0.78811 0.84788 0.0014351 0.91494 0.40263 0.0019319 0.4191 1.8632 1.861 16.0227 144.9034 0.00026901 -85.3454 0.36894
8.473 0.98814 5.4649e-005 3.8183 0.01192 0.00011013 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5815 0.5798 0.17724 0.020363 17.4675 0.12617 0.00016493 0.76399 0.0094548 0.010458 0.0014584 0.986 0.99109 3.1545e-006 1.2618e-005 0.16526 0.78872 0.84822 0.0014348 0.91546 0.40284 0.0019315 0.41911 1.8645 1.8624 16.0227 144.9034 0.00026849 -85.3477 0.36994
8.474 0.98814 5.4649e-005 3.8183 0.011919 0.00011014 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5816 0.57984 0.17726 0.020364 17.4706 0.12618 0.00016494 0.76399 0.0094552 0.010458 0.0014579 0.98601 0.99109 3.1532e-006 1.2613e-005 0.16526 0.78932 0.84855 0.0014345 0.91598 0.40304 0.0019311 0.41912 1.8659 1.8638 16.0227 144.9034 0.00026797 -85.35 0.37094
8.475 0.98814 5.4649e-005 3.8183 0.011919 0.00011016 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5817 0.57989 0.17727 0.020365 17.4737 0.12619 0.00016495 0.76398 0.0094556 0.010459 0.0014573 0.98602 0.9911 3.152e-006 1.2608e-005 0.16527 0.78993 0.84889 0.0014342 0.91649 0.40325 0.0019308 0.41914 1.8673 1.8652 16.0228 144.9034 0.00026746 -85.3522 0.37194
8.476 0.98814 5.4649e-005 3.8183 0.011919 0.00011017 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5818 0.57993 0.17728 0.020366 17.4768 0.12619 0.00016496 0.76397 0.0094559 0.010459 0.0014568 0.98603 0.9911 3.1507e-006 1.2603e-005 0.16527 0.79053 0.84922 0.0014339 0.917 0.40345 0.0019304 0.41915 1.8686 1.8665 16.0228 144.9035 0.00026694 -85.3545 0.37294
8.477 0.98814 5.4648e-005 3.8183 0.011919 0.00011018 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5818 0.57997 0.1773 0.020367 17.48 0.1262 0.00016497 0.76397 0.0094563 0.01046 0.0014562 0.98603 0.99111 3.1495e-006 1.2598e-005 0.16527 0.79113 0.84955 0.0014336 0.9175 0.40366 0.00193 0.41917 1.87 1.8679 16.0228 144.9035 0.00026643 -85.3567 0.37394
8.478 0.98814 5.4648e-005 3.8183 0.011919 0.0001102 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5819 0.58002 0.17731 0.020369 17.4831 0.1262 0.00016498 0.76396 0.0094567 0.01046 0.0014557 0.98604 0.99111 3.1482e-006 1.2593e-005 0.16527 0.79173 0.84988 0.0014333 0.91801 0.40387 0.0019297 0.41918 1.8713 1.8692 16.0228 144.9035 0.00026592 -85.359 0.37494
8.479 0.98814 5.4648e-005 3.8183 0.011919 0.00011021 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.582 0.58006 0.17732 0.02037 17.4862 0.12621 0.00016499 0.76395 0.009457 0.01046 0.0014551 0.98605 0.99112 3.147e-006 1.2588e-005 0.16528 0.79233 0.85021 0.0014331 0.91851 0.40407 0.0019293 0.41919 1.8727 1.8706 16.0228 144.9035 0.00026541 -85.3612 0.37594
8.48 0.98814 5.4648e-005 3.8183 0.011919 0.00011022 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5821 0.58011 0.17734 0.020371 17.4893 0.12622 0.000165 0.76395 0.0094574 0.010461 0.0014546 0.98605 0.99112 3.1458e-006 1.2583e-005 0.16528 0.79293 0.85054 0.0014328 0.919 0.40428 0.0019289 0.41921 1.874 1.8719 16.0228 144.9035 0.00026491 -85.3634 0.37694
8.481 0.98814 5.4648e-005 3.8183 0.011919 0.00011023 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5822 0.58015 0.17735 0.020372 17.4924 0.12622 0.00016501 0.76394 0.0094577 0.010461 0.0014541 0.98606 0.99113 3.1446e-006 1.2578e-005 0.16528 0.79352 0.85086 0.0014325 0.9195 0.40448 0.0019286 0.41922 1.8754 1.8733 16.0228 144.9035 0.00026441 -85.3655 0.37794
8.482 0.98814 5.4648e-005 3.8183 0.011919 0.00011025 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5823 0.5802 0.17736 0.020373 17.4955 0.12623 0.00016502 0.76394 0.0094581 0.010461 0.0014536 0.98607 0.99113 3.1434e-006 1.2573e-005 0.16529 0.79412 0.85118 0.0014323 0.91999 0.40469 0.0019282 0.41924 1.8767 1.8746 16.0228 144.9036 0.00026391 -85.3677 0.37894
8.483 0.98814 5.4648e-005 3.8183 0.011919 0.00011026 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5823 0.58024 0.17738 0.020374 17.4986 0.12624 0.00016503 0.76393 0.0094585 0.010462 0.0014531 0.98607 0.99113 3.1422e-006 1.2569e-005 0.16529 0.79471 0.85151 0.001432 0.92048 0.40489 0.0019279 0.41925 1.878 1.876 16.0228 144.9036 0.00026341 -85.3699 0.37994
8.484 0.98814 5.4648e-005 3.8183 0.011919 0.00011027 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5824 0.58029 0.17739 0.020375 17.5017 0.12624 0.00016504 0.76392 0.0094588 0.010462 0.0014525 0.98608 0.99114 3.141e-006 1.2564e-005 0.16529 0.79529 0.85183 0.0014317 0.92096 0.4051 0.0019275 0.41926 1.8794 1.8773 16.0228 144.9036 0.00026291 -85.372 0.38094
8.485 0.98814 5.4648e-005 3.8183 0.011919 0.00011028 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5825 0.58033 0.1774 0.020376 17.5048 0.12625 0.00016505 0.76392 0.0094592 0.010463 0.001452 0.98609 0.99114 3.1398e-006 1.2559e-005 0.16529 0.79588 0.85215 0.0014314 0.92144 0.40531 0.0019272 0.41928 1.8807 1.8786 16.0228 144.9036 0.00026242 -85.3741 0.38194
8.486 0.98814 5.4648e-005 3.8183 0.011919 0.0001103 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5826 0.58038 0.17742 0.020377 17.5079 0.12625 0.00016506 0.76391 0.0094596 0.010463 0.0014515 0.98609 0.99115 3.1386e-006 1.2555e-005 0.1653 0.79647 0.85246 0.0014312 0.92192 0.40551 0.0019268 0.41929 1.882 1.88 16.0228 144.9036 0.00026193 -85.3762 0.38294
8.487 0.98814 5.4648e-005 3.8183 0.011919 0.00011031 0.0011744 0.23369 0.00065931 0.23434 0.21625 0 0.03226 0.0389 0 1.5827 0.58042 0.17743 0.020378 17.511 0.12626 0.00016507 0.7639 0.0094599 0.010463 0.001451 0.9861 0.99115 3.1375e-006 1.255e-005 0.1653 0.79705 0.85278 0.0014309 0.9224 0.40572 0.0019265 0.41931 1.8833 1.8813 16.0228 144.9037 0.00026144 -85.3783 0.38394
8.488 0.98814 5.4648e-005 3.8183 0.011919 0.00011032 0.0011744 0.23369 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5828 0.58047 0.17744 0.020379 17.5141 0.12627 0.00016508 0.7639 0.0094603 0.010464 0.0014505 0.98611 0.99116 3.1363e-006 1.2545e-005 0.1653 0.79763 0.85309 0.0014307 0.92287 0.40592 0.0019262 0.41932 1.8846 1.8826 16.0229 144.9037 0.00026095 -85.3803 0.38494
8.489 0.98814 5.4647e-005 3.8183 0.011919 0.00011034 0.0011744 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5829 0.58051 0.17746 0.02038 17.5172 0.12627 0.00016509 0.76389 0.0094607 0.010464 0.00145 0.98611 0.99116 3.1352e-006 1.2541e-005 0.16531 0.79821 0.85341 0.0014304 0.92334 0.40613 0.0019258 0.41933 1.8859 1.8839 16.0229 144.9037 0.00026047 -85.3824 0.38594
8.49 0.98814 5.4647e-005 3.8183 0.011919 0.00011035 0.0011744 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5829 0.58055 0.17747 0.020381 17.5203 0.12628 0.0001651 0.76389 0.009461 0.010465 0.0014495 0.98612 0.99117 3.1341e-006 1.2536e-005 0.16531 0.79879 0.85372 0.0014301 0.92381 0.40633 0.0019255 0.41935 1.8873 1.8853 16.0229 144.9037 0.00025998 -85.3844 0.38694
8.491 0.98814 5.4647e-005 3.8183 0.011919 0.00011036 0.0011744 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.583 0.5806 0.17748 0.020382 17.5234 0.12629 0.00016511 0.76388 0.0094614 0.010465 0.001449 0.98613 0.99117 3.1329e-006 1.2532e-005 0.16531 0.79936 0.85403 0.0014299 0.92427 0.40654 0.0019252 0.41936 1.8886 1.8866 16.0229 144.9037 0.0002595 -85.3865 0.38794
8.492 0.98814 5.4647e-005 3.8183 0.011919 0.00011037 0.0011744 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5831 0.58064 0.1775 0.020383 17.5265 0.12629 0.00016512 0.76387 0.0094618 0.010465 0.0014486 0.98613 0.99117 3.1318e-006 1.2527e-005 0.16531 0.79994 0.85434 0.0014297 0.92473 0.40674 0.0019248 0.41938 1.8899 1.8879 16.0229 144.9037 0.00025902 -85.3885 0.38894
8.493 0.98814 5.4647e-005 3.8183 0.011919 0.00011039 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5832 0.58069 0.17751 0.020384 17.5296 0.1263 0.00016513 0.76387 0.0094621 0.010466 0.0014481 0.98614 0.99118 3.1307e-006 1.2523e-005 0.16532 0.80051 0.85465 0.0014294 0.92519 0.40695 0.0019245 0.41939 1.8912 1.8892 16.0229 144.9038 0.00025855 -85.3905 0.38994
8.494 0.98814 5.4647e-005 3.8183 0.011919 0.0001104 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5833 0.58073 0.17752 0.020385 17.5327 0.12631 0.00016514 0.76386 0.0094625 0.010466 0.0014476 0.98615 0.99118 3.1296e-006 1.2519e-005 0.16532 0.80108 0.85495 0.0014292 0.92565 0.40715 0.0019242 0.4194 1.8924 1.8905 16.0229 144.9038 0.00025807 -85.3924 0.39094
8.495 0.98814 5.4647e-005 3.8183 0.011919 0.00011041 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5834 0.58078 0.17754 0.020387 17.5358 0.12631 0.00016514 0.76385 0.0094628 0.010467 0.0014471 0.98615 0.99119 3.1285e-006 1.2514e-005 0.16532 0.80165 0.85526 0.0014289 0.9261 0.40736 0.0019239 0.41942 1.8937 1.8918 16.0229 144.9038 0.0002576 -85.3944 0.39194
8.496 0.98814 5.4647e-005 3.8183 0.011919 0.00011043 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5834 0.58082 0.17755 0.020388 17.5389 0.12632 0.00016515 0.76385 0.0094632 0.010467 0.0014466 0.98616 0.99119 3.1275e-006 1.251e-005 0.16532 0.80222 0.85556 0.0014287 0.92655 0.40756 0.0019235 0.41943 1.895 1.8931 16.0229 144.9038 0.00025713 -85.3964 0.39294
8.497 0.98814 5.4647e-005 3.8183 0.011919 0.00011044 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5835 0.58087 0.17756 0.020389 17.542 0.12632 0.00016516 0.76384 0.0094636 0.010467 0.0014462 0.98616 0.99119 3.1264e-006 1.2506e-005 0.16533 0.80278 0.85587 0.0014284 0.927 0.40777 0.0019232 0.41945 1.8963 1.8944 16.0229 144.9038 0.00025666 -85.3983 0.39394
8.498 0.98814 5.4647e-005 3.8183 0.011919 0.00011045 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5836 0.58091 0.17758 0.02039 17.5452 0.12633 0.00016517 0.76383 0.0094639 0.010468 0.0014457 0.98617 0.9912 3.1253e-006 1.2501e-005 0.16533 0.80335 0.85617 0.0014282 0.92744 0.40797 0.0019229 0.41946 1.8976 1.8956 16.0229 144.9039 0.0002562 -85.4002 0.39494
8.499 0.98814 5.4647e-005 3.8183 0.011919 0.00011046 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5837 0.58096 0.17759 0.020391 17.5483 0.12634 0.00016518 0.76383 0.0094643 0.010468 0.0014452 0.98618 0.9912 3.1243e-006 1.2497e-005 0.16533 0.80391 0.85647 0.0014279 0.92788 0.40818 0.0019226 0.41947 1.8989 1.8969 16.0229 144.9039 0.00025573 -85.4021 0.39594
8.5 0.98814 5.4647e-005 3.8183 0.011919 0.00011048 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5838 0.581 0.1776 0.020392 17.5514 0.12634 0.00016519 0.76382 0.0094647 0.010468 0.0014448 0.98618 0.99121 3.1232e-006 1.2493e-005 0.16534 0.80447 0.85677 0.0014277 0.92832 0.40838 0.0019223 0.41949 1.9001 1.8982 16.0229 144.9039 0.00025527 -85.404 0.39694
8.501 0.98814 5.4646e-005 3.8183 0.011919 0.00011049 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5839 0.58105 0.17762 0.020393 17.5545 0.12635 0.0001652 0.76382 0.009465 0.010469 0.0014443 0.98619 0.99121 3.1222e-006 1.2489e-005 0.16534 0.80503 0.85706 0.0014275 0.92876 0.40859 0.001922 0.4195 1.9014 1.8995 16.0229 144.9039 0.00025481 -85.4059 0.39794
8.502 0.98814 5.4646e-005 3.8183 0.011919 0.0001105 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.584 0.58109 0.17763 0.020394 17.5576 0.12636 0.00016521 0.76381 0.0094654 0.010469 0.0014439 0.98619 0.99121 3.1212e-006 1.2485e-005 0.16534 0.80558 0.85736 0.0014272 0.92919 0.40879 0.0019217 0.41952 1.9027 1.9008 16.0229 144.9039 0.00025435 -85.4078 0.39894
8.503 0.98814 5.4646e-005 3.8183 0.011919 0.00011052 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.584 0.58113 0.17764 0.020395 17.5607 0.12636 0.00016522 0.7638 0.0094658 0.01047 0.0014435 0.9862 0.99122 3.1201e-006 1.2481e-005 0.16534 0.80614 0.85765 0.001427 0.92963 0.40899 0.0019214 0.41953 1.9039 1.902 16.0229 144.904 0.0002539 -85.4096 0.39994
8.504 0.98814 5.4646e-005 3.8183 0.011919 0.00011053 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5841 0.58118 0.17766 0.020396 17.5638 0.12637 0.00016523 0.7638 0.0094661 0.01047 0.001443 0.98621 0.99122 3.1191e-006 1.2476e-005 0.16535 0.80669 0.85795 0.0014268 0.93005 0.4092 0.0019211 0.41955 1.9052 1.9033 16.0229 144.904 0.00025344 -85.4114 0.40094
8.505 0.98814 5.4646e-005 3.8183 0.011919 0.00011054 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5842 0.58122 0.17767 0.020397 17.5669 0.12637 0.00016524 0.76379 0.0094665 0.01047 0.0014426 0.98621 0.99123 3.1181e-006 1.2472e-005 0.16535 0.80724 0.85824 0.0014266 0.93048 0.4094 0.0019208 0.41956 1.9064 1.9045 16.0229 144.904 0.00025299 -85.4133 0.40194
8.506 0.98814 5.4646e-005 3.8183 0.011919 0.00011055 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5843 0.58127 0.17768 0.020398 17.57 0.12638 0.00016525 0.76378 0.0094669 0.010471 0.0014422 0.98622 0.99123 3.1171e-006 1.2468e-005 0.16535 0.80779 0.85853 0.0014263 0.9309 0.40961 0.0019205 0.41957 1.9077 1.9058 16.0229 144.904 0.00025254 -85.4151 0.40294
8.507 0.98814 5.4646e-005 3.8183 0.011919 0.00011057 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5844 0.58131 0.1777 0.020399 17.5731 0.12639 0.00016526 0.76378 0.0094672 0.010471 0.0014417 0.98622 0.99123 3.1161e-006 1.2464e-005 0.16536 0.80834 0.85882 0.0014261 0.93133 0.40981 0.0019202 0.41959 1.9089 1.9071 16.0229 144.904 0.00025209 -85.4169 0.40394
8.508 0.98814 5.4646e-005 3.8183 0.011919 0.00011058 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5845 0.58136 0.17771 0.0204 17.5763 0.12639 0.00016527 0.76377 0.0094676 0.010472 0.0014413 0.98623 0.99124 3.1151e-006 1.2461e-005 0.16536 0.80889 0.85911 0.0014259 0.93174 0.41002 0.0019199 0.4196 1.9102 1.9083 16.0229 144.904 0.00025165 -85.4187 0.40494
8.509 0.98814 5.4646e-005 3.8183 0.011919 0.00011059 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5845 0.5814 0.17772 0.020401 17.5794 0.1264 0.00016528 0.76377 0.0094679 0.010472 0.0014409 0.98623 0.99124 3.1142e-006 1.2457e-005 0.16536 0.80943 0.85939 0.0014257 0.93216 0.41022 0.0019196 0.41962 1.9114 1.9096 16.0229 144.9041 0.0002512 -85.4204 0.40594
8.51 0.98814 5.4646e-005 3.8183 0.011919 0.0001106 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5846 0.58145 0.17774 0.020402 17.5825 0.12641 0.00016529 0.76376 0.0094683 0.010472 0.0014404 0.98624 0.99124 3.1132e-006 1.2453e-005 0.16536 0.80998 0.85968 0.0014255 0.93257 0.41042 0.0019193 0.41963 1.9127 1.9108 16.0229 144.9041 0.00025076 -85.4222 0.40694
8.511 0.98814 5.4646e-005 3.8183 0.011919 0.00011062 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5847 0.58149 0.17775 0.020404 17.5856 0.12641 0.0001653 0.76375 0.0094687 0.010473 0.00144 0.98625 0.99125 3.1122e-006 1.2449e-005 0.16537 0.81052 0.85996 0.0014252 0.93298 0.41063 0.001919 0.41965 1.9139 1.912 16.023 144.9041 0.00025032 -85.4239 0.40794
8.512 0.98814 5.4646e-005 3.8183 0.011919 0.00011063 0.0011745 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5848 0.58154 0.17776 0.020405 17.5887 0.12642 0.00016531 0.76375 0.009469 0.010473 0.0014396 0.98625 0.99125 3.1113e-006 1.2445e-005 0.16537 0.81106 0.86024 0.001425 0.93339 0.41083 0.0019188 0.41966 1.9151 1.9133 16.023 144.9041 0.00024988 -85.4257 0.40894
8.513 0.98814 5.4645e-005 3.8183 0.011919 0.00011064 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5849 0.58158 0.17777 0.020406 17.5918 0.12643 0.00016532 0.76374 0.0094694 0.010473 0.0014392 0.98626 0.99125 3.1103e-006 1.2441e-005 0.16537 0.81159 0.86053 0.0014248 0.9338 0.41104 0.0019185 0.41967 1.9164 1.9145 16.023 144.9041 0.00024945 -85.4274 0.40994
8.514 0.98814 5.4645e-005 3.8183 0.011919 0.00011066 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.585 0.58163 0.17779 0.020407 17.5949 0.12643 0.00016533 0.76373 0.0094698 0.010474 0.0014388 0.98626 0.99126 3.1094e-006 1.2438e-005 0.16538 0.81213 0.86081 0.0014246 0.9342 0.41124 0.0019182 0.41969 1.9176 1.9157 16.023 144.9042 0.00024901 -85.4291 0.41094
8.515 0.98814 5.4645e-005 3.8183 0.011919 0.00011067 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5851 0.58167 0.1778 0.020408 17.598 0.12644 0.00016534 0.76373 0.0094701 0.010474 0.0014384 0.98627 0.99126 3.1085e-006 1.2434e-005 0.16538 0.81266 0.86109 0.0014244 0.9346 0.41144 0.0019179 0.4197 1.9188 1.917 16.023 144.9042 0.00024858 -85.4308 0.41194
8.516 0.98814 5.4645e-005 3.8183 0.011919 0.00011068 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5851 0.58171 0.17781 0.020409 17.6012 0.12644 0.00016535 0.76372 0.0094705 0.010475 0.001438 0.98627 0.99127 3.1075e-006 1.243e-005 0.16538 0.8132 0.86136 0.0014242 0.935 0.41165 0.0019176 0.41972 1.92 1.9182 16.023 144.9042 0.00024815 -85.4325 0.41294
8.517 0.98814 5.4645e-005 3.8183 0.011919 0.00011069 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5852 0.58176 0.17783 0.02041 17.6043 0.12645 0.00016536 0.76372 0.0094708 0.010475 0.0014376 0.98628 0.99127 3.1066e-006 1.2426e-005 0.16538 0.81373 0.86164 0.001424 0.93539 0.41185 0.0019174 0.41973 1.9212 1.9194 16.023 144.9042 0.00024772 -85.4341 0.41394
8.518 0.98814 5.4645e-005 3.8183 0.011919 0.00011071 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5853 0.5818 0.17784 0.020411 17.6074 0.12646 0.00016537 0.76371 0.0094712 0.010475 0.0014372 0.98628 0.99127 3.1057e-006 1.2423e-005 0.16539 0.81426 0.86192 0.0014238 0.93579 0.41205 0.0019171 0.41975 1.9224 1.9206 16.023 144.9042 0.0002473 -85.4358 0.41494
8.519 0.98814 5.4645e-005 3.8183 0.011919 0.00011072 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5854 0.58185 0.17785 0.020412 17.6105 0.12646 0.00016538 0.7637 0.0094716 0.010476 0.0014368 0.98629 0.99128 3.1048e-006 1.2419e-005 0.16539 0.81479 0.86219 0.0014236 0.93618 0.41226 0.0019168 0.41976 1.9237 1.9218 16.023 144.9043 0.00024687 -85.4375 0.41594
8.52 0.98814 5.4645e-005 3.8183 0.011919 0.00011073 0.0011746 0.23368 0.00065931 0.23434 0.21624 0 0.03226 0.0389 0 1.5855 0.58189 0.17787 0.020413 17.6136 0.12647 0.00016538 0.7637 0.0094719 0.010476 0.0014364 0.98629 0.99128 3.1039e-006 1.2416e-005 0.16539 0.81531 0.86246 0.0014234 0.93657 0.41246 0.0019166 0.41978 1.9249 1.9231 16.023 144.9043 0.00024645 -85.4391 0.41694
8.521 0.98814 5.4645e-005 3.8183 0.011919 0.00011075 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5856 0.58194 0.17788 0.020414 17.6167 0.12648 0.00016539 0.76369 0.0094723 0.010477 0.001436 0.9863 0.99128 3.103e-006 1.2412e-005 0.16539 0.81584 0.86274 0.0014232 0.93695 0.41266 0.0019163 0.41979 1.9261 1.9243 16.023 144.9043 0.00024603 -85.4407 0.41794
8.522 0.98814 5.4645e-005 3.8183 0.011919 0.00011076 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5856 0.58198 0.17789 0.020415 17.6198 0.12648 0.0001654 0.76368 0.0094727 0.010477 0.0014356 0.9863 0.99129 3.1021e-006 1.2408e-005 0.1654 0.81636 0.86301 0.001423 0.93733 0.41287 0.001916 0.4198 1.9273 1.9255 16.023 144.9043 0.00024561 -85.4423 0.41894
8.523 0.98814 5.4645e-005 3.8183 0.011919 0.00011077 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5857 0.58203 0.17791 0.020416 17.623 0.12649 0.00016541 0.76368 0.009473 0.010477 0.0014352 0.98631 0.99129 3.1012e-006 1.2405e-005 0.1654 0.81688 0.86328 0.0014228 0.93772 0.41307 0.0019158 0.41982 1.9285 1.9267 16.023 144.9043 0.00024519 -85.4439 0.41994
8.524 0.98814 5.4645e-005 3.8183 0.011919 0.00011078 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5858 0.58207 0.17792 0.020417 17.6261 0.12649 0.00016542 0.76367 0.0094734 0.010478 0.0014349 0.98631 0.99129 3.1004e-006 1.2401e-005 0.1654 0.8174 0.86355 0.0014225 0.93809 0.41327 0.0019155 0.41983 1.9296 1.9279 16.023 144.9043 0.00024477 -85.4455 0.42094
8.525 0.98814 5.4644e-005 3.8183 0.011919 0.0001108 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5859 0.58212 0.17793 0.020418 17.6292 0.1265 0.00016543 0.76366 0.0094737 0.010478 0.0014345 0.98632 0.9913 3.0995e-006 1.2398e-005 0.16541 0.81792 0.86381 0.0014223 0.93847 0.41348 0.0019153 0.41985 1.9308 1.9291 16.023 144.9044 0.00024436 -85.4471 0.42194
8.526 0.98814 5.4644e-005 3.8183 0.011919 0.00011081 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.586 0.58216 0.17795 0.020419 17.6323 0.12651 0.00016544 0.76366 0.0094741 0.010478 0.0014341 0.98632 0.9913 3.0987e-006 1.2395e-005 0.16541 0.81844 0.86408 0.0014221 0.93884 0.41368 0.001915 0.41986 1.932 1.9302 16.023 144.9044 0.00024395 -85.4486 0.42294
8.527 0.98814 5.4644e-005 3.8183 0.011919 0.00011082 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5861 0.5822 0.17796 0.02042 17.6354 0.12651 0.00016545 0.76365 0.0094745 0.010479 0.0014337 0.98633 0.9913 3.0978e-006 1.2391e-005 0.16541 0.81895 0.86435 0.001422 0.93922 0.41388 0.0019148 0.41988 1.9332 1.9314 16.023 144.9044 0.00024354 -85.4502 0.42394
8.528 0.98814 5.4644e-005 3.8183 0.011919 0.00011084 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5862 0.58225 0.17797 0.020422 17.6386 0.12652 0.00016546 0.76365 0.0094748 0.010479 0.0014333 0.98633 0.99131 3.097e-006 1.2388e-005 0.16541 0.81947 0.86461 0.0014218 0.93959 0.41409 0.0019145 0.41989 1.9344 1.9326 16.023 144.9044 0.00024313 -85.4517 0.42494
8.529 0.98814 5.4644e-005 3.8183 0.011919 0.00011085 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5862 0.58229 0.17799 0.020423 17.6417 0.12653 0.00016547 0.76364 0.0094752 0.01048 0.001433 0.98634 0.99131 3.0961e-006 1.2384e-005 0.16542 0.81998 0.86487 0.0014216 0.93995 0.41429 0.0019143 0.41991 1.9355 1.9338 16.023 144.9044 0.00024272 -85.4533 0.42594
8.53 0.98814 5.4644e-005 3.8183 0.011918 0.00011086 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5863 0.58234 0.178 0.020424 17.6448 0.12653 0.00016548 0.76363 0.0094756 0.01048 0.0014326 0.98634 0.99131 3.0953e-006 1.2381e-005 0.16542 0.82049 0.86513 0.0014214 0.94032 0.41449 0.001914 0.41992 1.9367 1.935 16.023 144.9045 0.00024232 -85.4548 0.42694
8.531 0.98814 5.4644e-005 3.8183 0.011918 0.00011087 0.0011746 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5864 0.58238 0.17801 0.020425 17.6479 0.12654 0.00016549 0.76363 0.0094759 0.01048 0.0014323 0.98635 0.99131 3.0945e-006 1.2378e-005 0.16542 0.821 0.86539 0.0014212 0.94068 0.41469 0.0019138 0.41993 1.9379 1.9361 16.023 144.9045 0.00024191 -85.4563 0.42794
8.532 0.98814 5.4644e-005 3.8183 0.011918 0.00011089 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5865 0.58243 0.17803 0.020426 17.651 0.12654 0.0001655 0.76362 0.0094763 0.010481 0.0014319 0.98635 0.99132 3.0936e-006 1.2375e-005 0.16543 0.8215 0.86565 0.001421 0.94104 0.4149 0.0019135 0.41995 1.939 1.9373 16.023 144.9045 0.00024151 -85.4578 0.42894
8.533 0.98814 5.4644e-005 3.8183 0.011918 0.0001109 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5866 0.58247 0.17804 0.020427 17.6541 0.12655 0.00016551 0.76361 0.0094766 0.010481 0.0014316 0.98636 0.99132 3.0928e-006 1.2371e-005 0.16543 0.82201 0.86591 0.0014208 0.9414 0.4151 0.0019133 0.41996 1.9402 1.9385 16.023 144.9045 0.00024111 -85.4593 0.42994
8.534 0.98814 5.4644e-005 3.8183 0.011918 0.00011091 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5867 0.58252 0.17805 0.020428 17.6573 0.12656 0.00016552 0.76361 0.009477 0.010482 0.0014312 0.98636 0.99132 3.092e-006 1.2368e-005 0.16543 0.82251 0.86617 0.0014207 0.94175 0.4153 0.001913 0.41998 1.9414 1.9396 16.023 144.9045 0.00024071 -85.4608 0.43094
8.535 0.98814 5.4644e-005 3.8183 0.011918 0.00011092 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5867 0.58256 0.17807 0.020429 17.6604 0.12656 0.00016553 0.7636 0.0094774 0.010482 0.0014309 0.98637 0.99133 3.0912e-006 1.2365e-005 0.16543 0.82301 0.86643 0.0014205 0.94211 0.41551 0.0019128 0.41999 1.9425 1.9408 16.023 144.9046 0.00024032 -85.4622 0.43194
8.536 0.98814 5.4644e-005 3.8183 0.011918 0.00011094 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5868 0.58261 0.17808 0.02043 17.6635 0.12657 0.00016554 0.7636 0.0094777 0.010482 0.0014305 0.98637 0.99133 3.0904e-006 1.2362e-005 0.16544 0.82352 0.86668 0.0014203 0.94246 0.41571 0.0019126 0.42001 1.9437 1.942 16.023 144.9046 0.00023992 -85.4637 0.43294
8.537 0.98814 5.4643e-005 3.8183 0.011918 0.00011095 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5869 0.58265 0.17809 0.020431 17.6666 0.12658 0.00016555 0.76359 0.0094781 0.010483 0.0014302 0.98637 0.99133 3.0896e-006 1.2359e-005 0.16544 0.82401 0.86693 0.0014201 0.94281 0.41591 0.0019123 0.42002 1.9448 1.9431 16.023 144.9046 0.00023953 -85.4651 0.43394
8.538 0.98814 5.4643e-005 3.8183 0.011918 0.00011096 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.587 0.58269 0.17811 0.020432 17.6698 0.12658 0.00016556 0.76358 0.0094785 0.010483 0.0014298 0.98638 0.99134 3.0888e-006 1.2355e-005 0.16544 0.82451 0.86719 0.0014199 0.94316 0.41611 0.0019121 0.42004 1.946 1.9443 16.023 144.9046 0.00023914 -85.4666 0.43494
8.539 0.98814 5.4643e-005 3.8183 0.011918 0.00011098 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5871 0.58274 0.17812 0.020433 17.6729 0.12659 0.00016557 0.76358 0.0094788 0.010483 0.0014295 0.98638 0.99134 3.0881e-006 1.2352e-005 0.16544 0.82501 0.86744 0.0014198 0.9435 0.41631 0.0019119 0.42005 1.9471 1.9454 16.023 144.9046 0.00023875 -85.468 0.43594
8.54 0.98814 5.4643e-005 3.8183 0.011918 0.00011099 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5872 0.58278 0.17813 0.020434 17.676 0.1266 0.00016558 0.76357 0.0094792 0.010484 0.0014292 0.98639 0.99134 3.0873e-006 1.2349e-005 0.16545 0.8255 0.86769 0.0014196 0.94384 0.41652 0.0019116 0.42007 1.9483 1.9466 16.023 144.9047 0.00023836 -85.4694 0.43694
8.541 0.98814 5.4643e-005 3.8183 0.011918 0.000111 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5873 0.58283 0.17815 0.020435 17.6791 0.1266 0.00016559 0.76356 0.0094795 0.010484 0.0014288 0.98639 0.99134 3.0865e-006 1.2346e-005 0.16545 0.826 0.86794 0.0014194 0.94418 0.41672 0.0019114 0.42008 1.9494 1.9477 16.023 144.9047 0.00023797 -85.4708 0.43794
8.542 0.98814 5.4643e-005 3.8183 0.011918 0.00011101 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5873 0.58287 0.17816 0.020436 17.6822 0.12661 0.0001656 0.76356 0.0094799 0.010485 0.0014285 0.9864 0.99135 3.0858e-006 1.2343e-005 0.16545 0.82649 0.86819 0.0014192 0.94452 0.41692 0.0019112 0.4201 1.9505 1.9488 16.023 144.9047 0.00023759 -85.4722 0.43894
8.543 0.98814 5.4643e-005 3.8183 0.011918 0.00011103 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5874 0.58292 0.17817 0.020437 17.6854 0.12661 0.00016561 0.76355 0.0094803 0.010485 0.0014282 0.9864 0.99135 3.085e-006 1.234e-005 0.16546 0.82698 0.86844 0.0014191 0.94486 0.41712 0.001911 0.42011 1.9517 1.95 16.0229 144.9047 0.0002372 -85.4736 0.43994
8.544 0.98814 5.4643e-005 3.8183 0.011918 0.00011104 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5875 0.58296 0.17819 0.020438 17.6885 0.12662 0.00016561 0.76355 0.0094806 0.010485 0.0014278 0.98641 0.99135 3.0843e-006 1.2337e-005 0.16546 0.82747 0.86868 0.0014189 0.94519 0.41733 0.0019107 0.42013 1.9528 1.9511 16.0229 144.9047 0.00023682 -85.4749 0.44094
8.545 0.98814 5.4643e-005 3.8183 0.011918 0.00011105 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5876 0.58301 0.1782 0.020439 17.6916 0.12663 0.00016562 0.76354 0.009481 0.010486 0.0014275 0.98641 0.99136 3.0835e-006 1.2334e-005 0.16546 0.82795 0.86893 0.0014187 0.94553 0.41753 0.0019105 0.42014 1.9539 1.9522 16.0229 144.9047 0.00023644 -85.4763 0.44194
8.546 0.98814 5.4643e-005 3.8183 0.011918 0.00011107 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5877 0.58305 0.17821 0.020441 17.6947 0.12663 0.00016563 0.76353 0.0094813 0.010486 0.0014272 0.98641 0.99136 3.0828e-006 1.2331e-005 0.16546 0.82844 0.86917 0.0014185 0.94586 0.41773 0.0019103 0.42015 1.955 1.9534 16.0229 144.9048 0.00023606 -85.4776 0.44294
8.547 0.98814 5.4643e-005 3.8183 0.011918 0.00011108 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5878 0.5831 0.17823 0.020442 17.6979 0.12664 0.00016564 0.76353 0.0094817 0.010486 0.0014268 0.98642 0.99136 3.0821e-006 1.2328e-005 0.16547 0.82892 0.86941 0.0014184 0.94618 0.41793 0.0019101 0.42017 1.9561 1.9545 16.0229 144.9048 0.00023569 -85.479 0.44394
8.548 0.98814 5.4643e-005 3.8183 0.011918 0.00011109 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5878 0.58314 0.17824 0.020443 17.701 0.12665 0.00016565 0.76352 0.0094821 0.010487 0.0014265 0.98642 0.99136 3.0813e-006 1.2325e-005 0.16547 0.8294 0.86966 0.0014182 0.94651 0.41813 0.0019099 0.42018 1.9573 1.9556 16.0229 144.9048 0.00023531 -85.4803 0.44494
8.549 0.98814 5.4643e-005 3.8183 0.011918 0.0001111 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5879 0.58319 0.17825 0.020444 17.7041 0.12665 0.00016566 0.76351 0.0094824 0.010487 0.0014262 0.98643 0.99137 3.0806e-006 1.2322e-005 0.16547 0.82989 0.8699 0.001418 0.94683 0.41833 0.0019096 0.4202 1.9584 1.9567 16.0229 144.9048 0.00023494 -85.4816 0.44594
8.55 0.98814 5.4642e-005 3.8183 0.011918 0.00011112 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.588 0.58323 0.17826 0.020445 17.7072 0.12666 0.00016567 0.76351 0.0094828 0.010488 0.0014259 0.98643 0.99137 3.0799e-006 1.232e-005 0.16548 0.83036 0.87014 0.0014179 0.94716 0.41854 0.0019094 0.42021 1.9595 1.9578 16.0229 144.9048 0.00023457 -85.483 0.44694
8.551 0.98814 5.4642e-005 3.8183 0.011918 0.00011113 0.0011747 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5881 0.58327 0.17828 0.020446 17.7104 0.12666 0.00016568 0.7635 0.0094832 0.010488 0.0014256 0.98643 0.99137 3.0792e-006 1.2317e-005 0.16548 0.83084 0.87038 0.0014177 0.94748 0.41874 0.0019092 0.42023 1.9606 1.959 16.0229 144.9049 0.0002342 -85.4843 0.44794
8.552 0.98814 5.4642e-005 3.8183 0.011918 0.00011114 0.0011748 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5882 0.58332 0.17829 0.020447 17.7135 0.12667 0.00016569 0.7635 0.0094835 0.010488 0.0014253 0.98644 0.99137 3.0785e-006 1.2314e-005 0.16548 0.83132 0.87062 0.0014176 0.94779 0.41894 0.001909 0.42024 1.9617 1.9601 16.0229 144.9049 0.00023383 -85.4856 0.44894
8.553 0.98814 5.4642e-005 3.8183 0.011918 0.00011116 0.0011748 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5883 0.58336 0.1783 0.020448 17.7166 0.12668 0.0001657 0.76349 0.0094839 0.010489 0.001425 0.98644 0.99138 3.0778e-006 1.2311e-005 0.16548 0.83179 0.87085 0.0014174 0.94811 0.41914 0.0019088 0.42026 1.9628 1.9612 16.0229 144.9049 0.00023346 -85.4868 0.44994
8.554 0.98814 5.4642e-005 3.8183 0.011918 0.00011117 0.0011748 0.23368 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5884 0.58341 0.17832 0.020449 17.7197 0.12668 0.00016571 0.76348 0.0094842 0.010489 0.0014247 0.98645 0.99138 3.0771e-006 1.2308e-005 0.16549 0.83227 0.87109 0.0014172 0.94842 0.41934 0.0019086 0.42027 1.9639 1.9623 16.0229 144.9049 0.0002331 -85.4881 0.45094
8.555 0.98814 5.4642e-005 3.8183 0.011918 0.00011118 0.0011748 0.23367 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5884 0.58345 0.17833 0.02045 17.7229 0.12669 0.00016572 0.76348 0.0094846 0.01049 0.0014244 0.98645 0.99138 3.0764e-006 1.2306e-005 0.16549 0.83274 0.87132 0.0014171 0.94873 0.41954 0.0019084 0.42029 1.965 1.9634 16.0229 144.9049 0.00023273 -85.4894 0.45194
8.556 0.98814 5.4642e-005 3.8183 0.011918 0.00011119 0.0011748 0.23367 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5885 0.5835 0.17834 0.020451 17.726 0.1267 0.00016573 0.76347 0.009485 0.01049 0.0014241 0.98645 0.99138 3.0757e-006 1.2303e-005 0.16549 0.83321 0.87156 0.0014169 0.94904 0.41974 0.0019082 0.4203 1.9661 1.9645 16.0229 144.905 0.00023237 -85.4906 0.45294
8.557 0.98814 5.4642e-005 3.8183 0.011918 0.00011121 0.0011748 0.23367 0.00065931 0.23433 0.21624 0 0.03226 0.0389 0 1.5886 0.58354 0.17836 0.020452 17.7291 0.1267 0.00016574 0.76346 0.0094853 0.01049 0.0014238 0.98646 0.99139 3.075e-006 1.23e-005 0.16549 0.83368 0.87179 0.0014168 0.94935 0.41995 0.001908 0.42032 1.9671 1.9656 16.0229 144.905 0.00023201 -85.4919 0.45394
8.558 0.98814 5.4642e-005 3.8183 0.011918 0.00011122 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5887 0.58359 0.17837 0.020453 17.7322 0.12671 0.00016575 0.76346 0.0094857 0.010491 0.0014235 0.98646 0.99139 3.0744e-006 1.2297e-005 0.1655 0.83415 0.87202 0.0014166 0.94966 0.42015 0.0019078 0.42033 1.9682 1.9666 16.0229 144.905 0.00023165 -85.4931 0.45494
8.559 0.98814 5.4642e-005 3.8183 0.011918 0.00011123 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5888 0.58363 0.17838 0.020454 17.7354 0.12671 0.00016576 0.76345 0.009486 0.010491 0.0014232 0.98647 0.99139 3.0737e-006 1.2295e-005 0.1655 0.83461 0.87226 0.0014165 0.94996 0.42035 0.0019076 0.42035 1.9693 1.9677 16.0229 144.905 0.00023129 -85.4944 0.45594
8.56 0.98814 5.4642e-005 3.8183 0.011918 0.00011124 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5889 0.58368 0.1784 0.020455 17.7385 0.12672 0.00016577 0.76345 0.0094864 0.010491 0.0014229 0.98647 0.99139 3.073e-006 1.2292e-005 0.1655 0.83508 0.87249 0.0014163 0.95027 0.42055 0.0019074 0.42036 1.9704 1.9688 16.0229 144.905 0.00023093 -85.4956 0.45694
8.561 0.98814 5.4642e-005 3.8183 0.011918 0.00011126 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5889 0.58372 0.17841 0.020456 17.7416 0.12673 0.00016578 0.76344 0.0094868 0.010492 0.0014226 0.98647 0.9914 3.0724e-006 1.2289e-005 0.16551 0.83554 0.87272 0.0014162 0.95057 0.42075 0.0019072 0.42038 1.9715 1.9699 16.0229 144.9051 0.00023058 -85.4968 0.45794
8.562 0.98814 5.4641e-005 3.8183 0.011918 0.00011127 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.589 0.58376 0.17842 0.020457 17.7448 0.12673 0.00016579 0.76343 0.0094871 0.010492 0.0014223 0.98648 0.9914 3.0717e-006 1.2287e-005 0.16551 0.836 0.87294 0.001416 0.95086 0.42095 0.001907 0.42039 1.9725 1.971 16.0229 144.9051 0.00023023 -85.498 0.45894
8.563 0.98814 5.4641e-005 3.8183 0.011918 0.00011128 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5891 0.58381 0.17844 0.020458 17.7479 0.12674 0.0001658 0.76343 0.0094875 0.010493 0.0014221 0.98648 0.9914 3.0711e-006 1.2284e-005 0.16551 0.83646 0.87317 0.0014159 0.95116 0.42115 0.0019068 0.42041 1.9736 1.972 16.0229 144.9051 0.00022987 -85.4992 0.45994
8.564 0.98814 5.4641e-005 3.8183 0.011918 0.0001113 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5892 0.58385 0.17845 0.020459 17.751 0.12675 0.00016581 0.76342 0.0094878 0.010493 0.0014218 0.98648 0.9914 3.0704e-006 1.2282e-005 0.16551 0.83692 0.8734 0.0014157 0.95146 0.42135 0.0019066 0.42042 1.9747 1.9731 16.0229 144.9051 0.00022952 -85.5004 0.46094
8.565 0.98814 5.4641e-005 3.8183 0.011918 0.00011131 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5893 0.5839 0.17846 0.020461 17.7542 0.12675 0.00016582 0.76341 0.0094882 0.010493 0.0014215 0.98649 0.99141 3.0698e-006 1.2279e-005 0.16552 0.83738 0.87362 0.0014156 0.95175 0.42155 0.0019064 0.42044 1.9757 1.9742 16.0229 144.9051 0.00022918 -85.5015 0.46194
8.566 0.98814 5.4641e-005 3.8183 0.011918 0.00011132 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5894 0.58394 0.17848 0.020462 17.7573 0.12676 0.00016583 0.76341 0.0094886 0.010494 0.0014212 0.98649 0.99141 3.0691e-006 1.2277e-005 0.16552 0.83784 0.87385 0.0014154 0.95204 0.42175 0.0019062 0.42045 1.9768 1.9752 16.0229 144.9052 0.00022883 -85.5027 0.46294
8.567 0.98814 5.4641e-005 3.8183 0.011918 0.00011133 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.03226 0.0389 0 1.5895 0.58399 0.17849 0.020463 17.7604 0.12676 0.00016583 0.7634 0.0094889 0.010494 0.0014209 0.98649 0.99141 3.0685e-006 1.2274e-005 0.16552 0.83829 0.87407 0.0014153 0.95233 0.42195 0.001906 0.42047 1.9779 1.9763 16.0229 144.9052 0.00022848 -85.5039 0.46394
8.568 0.98814 5.4641e-005 3.8183 0.011918 0.00011135 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5895 0.58403 0.1785 0.020464 17.7635 0.12677 0.00016584 0.7634 0.0094893 0.010495 0.0014206 0.9865 0.99141 3.0679e-006 1.2272e-005 0.16553 0.83874 0.87429 0.0014151 0.95262 0.42215 0.0019059 0.42048 1.9789 1.9774 16.0228 144.9052 0.00022814 -85.505 0.46494
8.569 0.98814 5.4641e-005 3.8183 0.011918 0.00011136 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5896 0.58408 0.17852 0.020465 17.7667 0.12678 0.00016585 0.76339 0.0094896 0.010495 0.0014204 0.9865 0.99142 3.0673e-006 1.2269e-005 0.16553 0.8392 0.87452 0.001415 0.9529 0.42236 0.0019057 0.4205 1.98 1.9784 16.0228 144.9052 0.00022779 -85.5062 0.46594
8.57 0.98814 5.4641e-005 3.8183 0.011918 0.00011137 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5897 0.58412 0.17853 0.020466 17.7698 0.12678 0.00016586 0.76338 0.00949 0.010495 0.0014201 0.98651 0.99142 3.0666e-006 1.2267e-005 0.16553 0.83965 0.87474 0.0014149 0.95319 0.42256 0.0019055 0.42051 1.981 1.9795 16.0228 144.9052 0.00022745 -85.5073 0.46694
8.571 0.98814 5.4641e-005 3.8183 0.011918 0.00011139 0.0011748 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5898 0.58417 0.17854 0.020467 17.7729 0.12679 0.00016587 0.76338 0.0094904 0.010496 0.0014198 0.98651 0.99142 3.066e-006 1.2264e-005 0.16553 0.84009 0.87496 0.0014147 0.95347 0.42276 0.0019053 0.42052 1.9821 1.9805 16.0228 144.9053 0.00022711 -85.5084 0.46794
8.572 0.98814 5.4641e-005 3.8183 0.011918 0.0001114 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5899 0.58421 0.17856 0.020468 17.7761 0.1268 0.00016588 0.76337 0.0094907 0.010496 0.0014196 0.98651 0.99142 3.0654e-006 1.2262e-005 0.16554 0.84054 0.87518 0.0014146 0.95375 0.42296 0.0019051 0.42054 1.9831 1.9816 16.0228 144.9053 0.00022677 -85.5096 0.46894
8.573 0.98814 5.4641e-005 3.8183 0.011918 0.00011141 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.59 0.58425 0.17857 0.020469 17.7792 0.1268 0.00016589 0.76336 0.0094911 0.010496 0.0014193 0.98652 0.99143 3.0648e-006 1.2259e-005 0.16554 0.84099 0.8754 0.0014144 0.95403 0.42316 0.0019049 0.42055 1.9841 1.9826 16.0228 144.9053 0.00022644 -85.5107 0.46994
8.574 0.98814 5.464e-005 3.8183 0.011918 0.00011142 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.59 0.5843 0.17858 0.02047 17.7823 0.12681 0.0001659 0.76336 0.0094914 0.010497 0.0014191 0.98652 0.99143 3.0642e-006 1.2257e-005 0.16554 0.84143 0.87561 0.0014143 0.9543 0.42336 0.0019048 0.42057 1.9852 1.9837 16.0228 144.9053 0.0002261 -85.5118 0.47094
8.575 0.98814 5.464e-005 3.8183 0.011918 0.00011144 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5901 0.58434 0.1786 0.020471 17.7855 0.12681 0.00016591 0.76335 0.0094918 0.010497 0.0014188 0.98652 0.99143 3.0636e-006 1.2255e-005 0.16554 0.84188 0.87583 0.0014142 0.95458 0.42356 0.0019046 0.42058 1.9862 1.9847 16.0228 144.9053 0.00022577 -85.5129 0.47194
8.576 0.98814 5.464e-005 3.8183 0.011918 0.00011145 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5902 0.58439 0.17861 0.020472 17.7886 0.12682 0.00016592 0.76335 0.0094922 0.010498 0.0014186 0.98653 0.99143 3.063e-006 1.2252e-005 0.16555 0.84232 0.87604 0.001414 0.95485 0.42376 0.0019044 0.4206 1.9872 1.9857 16.0228 144.9053 0.00022543 -85.514 0.47294
8.577 0.98814 5.464e-005 3.8183 0.011918 0.00011146 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5903 0.58443 0.17862 0.020473 17.7917 0.12683 0.00016593 0.76334 0.0094925 0.010498 0.0014183 0.98653 0.99143 3.0625e-006 1.225e-005 0.16555 0.84276 0.87626 0.0014139 0.95512 0.42396 0.0019042 0.42061 1.9883 1.9868 16.0228 144.9054 0.0002251 -85.515 0.47394
8.578 0.98814 5.464e-005 3.8183 0.011918 0.00011148 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5904 0.58448 0.17864 0.020474 17.7949 0.12683 0.00016594 0.76333 0.0094929 0.010498 0.0014181 0.98653 0.99144 3.0619e-006 1.2247e-005 0.16555 0.8432 0.87647 0.0014138 0.95539 0.42416 0.0019041 0.42063 1.9893 1.9878 16.0228 144.9054 0.00022477 -85.5161 0.47494
8.579 0.98814 5.464e-005 3.8183 0.011918 0.00011149 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5905 0.58452 0.17865 0.020475 17.798 0.12684 0.00016595 0.76333 0.0094932 0.010499 0.0014178 0.98654 0.99144 3.0613e-006 1.2245e-005 0.16556 0.84364 0.87669 0.0014137 0.95566 0.42436 0.0019039 0.42064 1.9903 1.9888 16.0228 144.9054 0.00022444 -85.5172 0.47594
8.58 0.98814 5.464e-005 3.8183 0.011918 0.0001115 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5906 0.58457 0.17866 0.020476 17.8011 0.12685 0.00016596 0.76332 0.0094936 0.010499 0.0014175 0.98654 0.99144 3.0607e-006 1.2243e-005 0.16556 0.84407 0.8769 0.0014135 0.95593 0.42456 0.0019037 0.42066 1.9913 1.9899 16.0228 144.9054 0.00022411 -85.5182 0.47694
8.581 0.98814 5.464e-005 3.8183 0.011918 0.00011151 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5906 0.58461 0.17867 0.020477 17.8043 0.12685 0.00016597 0.76331 0.009494 0.010499 0.0014173 0.98654 0.99144 3.0602e-006 1.2241e-005 0.16556 0.84451 0.87711 0.0014134 0.95619 0.42476 0.0019036 0.42067 1.9924 1.9909 16.0228 144.9054 0.00022379 -85.5193 0.47794
8.582 0.98814 5.464e-005 3.8183 0.011918 0.00011153 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5907 0.58466 0.17869 0.020478 17.8074 0.12686 0.00016598 0.76331 0.0094943 0.0105 0.001417 0.98655 0.99144 3.0596e-006 1.2238e-005 0.16556 0.84494 0.87732 0.0014133 0.95646 0.42496 0.0019034 0.42069 1.9934 1.9919 16.0228 144.9055 0.00022346 -85.5203 0.47894
8.583 0.98814 5.464e-005 3.8183 0.011918 0.00011154 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5908 0.5847 0.1787 0.020479 17.8106 0.12686 0.00016599 0.7633 0.0094947 0.0105 0.0014168 0.98655 0.99145 3.059e-006 1.2236e-005 0.16557 0.84538 0.87753 0.0014131 0.95672 0.42516 0.0019032 0.4207 1.9944 1.9929 16.0227 144.9055 0.00022314 -85.5214 0.47994
8.584 0.98814 5.464e-005 3.8183 0.011918 0.00011155 0.0011749 0.23367 0.00065931 0.23433 0.21623 0 0.032261 0.0389 0 1.5909 0.58474 0.17871 0.020481 17.8137 0.12687 0.000166 0.7633 0.009495 0.010501 0.0014166 0.98655 0.99145 3.0585e-006 1.2234e-005 0.16557 0.84581 0.87774 0.001413 0.95698 0.42535 0.001903 0.42072 1.9954 1.9939 16.0227 144.9055 0.00022282 -85.5224 0.48094
8.585 0.98814 5.464e-005 3.8183 0.011918 0.00011156 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.591 0.58479 0.17873 0.020482 17.8168 0.12688 0.00016601 0.76329 0.0094954 0.010501 0.0014163 0.98655 0.99145 3.0579e-006 1.2232e-005 0.16557 0.84624 0.87794 0.0014129 0.95724 0.42555 0.0019029 0.42073 1.9964 1.995 16.0227 144.9055 0.0002225 -85.5234 0.48194
8.586 0.98814 5.4639e-005 3.8183 0.011917 0.00011158 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5911 0.58483 0.17874 0.020483 17.82 0.12688 0.00016602 0.76328 0.0094958 0.010501 0.0014161 0.98656 0.99145 3.0574e-006 1.2229e-005 0.16557 0.84667 0.87815 0.0014128 0.95749 0.42575 0.0019027 0.42075 1.9974 1.996 16.0227 144.9055 0.00022218 -85.5244 0.48294
8.587 0.98814 5.4639e-005 3.8183 0.011917 0.00011159 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5911 0.58488 0.17875 0.020484 17.8231 0.12689 0.00016603 0.76328 0.0094961 0.010502 0.0014159 0.98656 0.99146 3.0568e-006 1.2227e-005 0.16558 0.84709 0.87836 0.0014126 0.95775 0.42595 0.0019026 0.42076 1.9984 1.997 16.0227 144.9056 0.00022186 -85.5254 0.48394
8.588 0.98814 5.4639e-005 3.8183 0.011917 0.0001116 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5912 0.58492 0.17877 0.020485 17.8262 0.1269 0.00016604 0.76327 0.0094965 0.010502 0.0014156 0.98656 0.99146 3.0563e-006 1.2225e-005 0.16558 0.84752 0.87856 0.0014125 0.958 0.42615 0.0019024 0.42078 1.9994 1.998 16.0227 144.9056 0.00022154 -85.5264 0.48494
8.589 0.98814 5.4639e-005 3.8183 0.011917 0.00011162 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5913 0.58497 0.17878 0.020486 17.8294 0.1269 0.00016604 0.76326 0.0094968 0.010502 0.0014154 0.98657 0.99146 3.0558e-006 1.2223e-005 0.16558 0.84794 0.87877 0.0014124 0.95825 0.42635 0.0019022 0.42079 2.0004 1.999 16.0227 144.9056 0.00022122 -85.5274 0.48594
8.59 0.98814 5.4639e-005 3.8183 0.011917 0.00011163 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5914 0.58501 0.17879 0.020487 17.8325 0.12691 0.00016605 0.76326 0.0094972 0.010503 0.0014151 0.98657 0.99146 3.0552e-006 1.2221e-005 0.16559 0.84837 0.87897 0.0014123 0.9585 0.42655 0.0019021 0.42081 2.0014 2 16.0227 144.9056 0.00022091 -85.5284 0.48694
8.591 0.98814 5.4639e-005 3.8183 0.011917 0.00011164 0.0011749 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5915 0.58506 0.17881 0.020488 17.8357 0.12691 0.00016606 0.76325 0.0094976 0.010503 0.0014149 0.98657 0.99146 3.0547e-006 1.2219e-005 0.16559 0.84879 0.87917 0.0014121 0.95875 0.42675 0.0019019 0.42082 2.0024 2.001 16.0227 144.9056 0.0002206 -85.5294 0.48794
8.592 0.98814 5.4639e-005 3.8183 0.011917 0.00011165 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5916 0.5851 0.17882 0.020489 17.8388 0.12692 0.00016607 0.76325 0.0094979 0.010504 0.0014147 0.98658 0.99147 3.0542e-006 1.2217e-005 0.16559 0.84921 0.87937 0.001412 0.959 0.42695 0.0019018 0.42084 2.0034 2.002 16.0227 144.9057 0.00022029 -85.5303 0.48894
8.593 0.98814 5.4639e-005 3.8183 0.011917 0.00011167 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5917 0.58515 0.17883 0.02049 17.8419 0.12693 0.00016608 0.76324 0.0094983 0.010504 0.0014144 0.98658 0.99147 3.0537e-006 1.2215e-005 0.16559 0.84963 0.87957 0.0014119 0.95924 0.42715 0.0019016 0.42085 2.0044 2.0029 16.0227 144.9057 0.00021998 -85.5313 0.48994
8.594 0.98814 5.4639e-005 3.8183 0.011917 0.00011168 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5917 0.58519 0.17885 0.020491 17.8451 0.12693 0.00016609 0.76323 0.0094986 0.010504 0.0014142 0.98658 0.99147 3.0531e-006 1.2213e-005 0.1656 0.85005 0.87978 0.0014118 0.95949 0.42735 0.0019015 0.42087 2.0054 2.0039 16.0227 144.9057 0.00021967 -85.5322 0.49094
8.595 0.98814 5.4639e-005 3.8183 0.011917 0.00011169 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5918 0.58523 0.17886 0.020492 17.8482 0.12694 0.0001661 0.76323 0.009499 0.010505 0.001414 0.98658 0.99147 3.0526e-006 1.221e-005 0.1656 0.85046 0.87997 0.0014117 0.95973 0.42755 0.0019013 0.42088 2.0063 2.0049 16.0226 144.9057 0.00021936 -85.5332 0.49194
8.596 0.98814 5.4639e-005 3.8183 0.011917 0.00011171 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5919 0.58528 0.17887 0.020493 17.8514 0.12695 0.00016611 0.76322 0.0094993 0.010505 0.0014138 0.98659 0.99147 3.0521e-006 1.2208e-005 0.1656 0.85088 0.88017 0.0014116 0.95997 0.42774 0.0019011 0.4209 2.0073 2.0059 16.0226 144.9057 0.00021905 -85.5341 0.49294
8.597 0.98814 5.4639e-005 3.8183 0.011917 0.00011172 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.592 0.58532 0.17889 0.020494 17.8545 0.12695 0.00016612 0.76321 0.0094997 0.010506 0.0014136 0.98659 0.99147 3.0516e-006 1.2206e-005 0.16561 0.85129 0.88037 0.0014115 0.96021 0.42794 0.001901 0.42091 2.0083 2.0069 16.0226 144.9058 0.00021875 -85.5351 0.49394
8.598 0.98814 5.4638e-005 3.8183 0.011917 0.00011173 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5921 0.58537 0.1789 0.020495 17.8576 0.12696 0.00016613 0.76321 0.0095001 0.010506 0.0014134 0.98659 0.99148 3.0511e-006 1.2204e-005 0.16561 0.8517 0.88057 0.0014113 0.96045 0.42814 0.0019008 0.42093 2.0093 2.0079 16.0226 144.9058 0.00021844 -85.536 0.49494
8.599 0.98814 5.4638e-005 3.8183 0.011917 0.00011174 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5922 0.58541 0.17891 0.020496 17.8608 0.12696 0.00016614 0.7632 0.0095004 0.010506 0.0014131 0.9866 0.99148 3.0506e-006 1.2202e-005 0.16561 0.85212 0.88076 0.0014112 0.96068 0.42834 0.0019007 0.42094 2.0102 2.0088 16.0226 144.9058 0.00021814 -85.5369 0.49594
8.6 0.98814 5.4638e-005 3.8183 0.011917 0.00011176 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5922 0.58546 0.17893 0.020497 17.8639 0.12697 0.00016615 0.7632 0.0095008 0.010507 0.0014129 0.9866 0.99148 3.0501e-006 1.22e-005 0.16561 0.85253 0.88096 0.0014111 0.96092 0.42854 0.0019006 0.42096 2.0112 2.0098 16.0226 144.9058 0.00021784 -85.5378 0.49694
8.601 0.98814 5.4638e-005 3.8183 0.011917 0.00011177 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5923 0.5855 0.17894 0.020498 17.8671 0.12698 0.00016616 0.76319 0.0095011 0.010507 0.0014127 0.9866 0.99148 3.0496e-006 1.2198e-005 0.16562 0.85294 0.88115 0.001411 0.96115 0.42874 0.0019004 0.42097 2.0122 2.0108 16.0226 144.9058 0.00021754 -85.5387 0.49794
8.602 0.98814 5.4638e-005 3.8183 0.011917 0.00011178 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5924 0.58555 0.17895 0.020499 17.8702 0.12698 0.00016617 0.76318 0.0095015 0.010507 0.0014124 0.9866 0.99148 3.0491e-006 1.2197e-005 0.16562 0.85334 0.88135 0.0014108 0.96138 0.42894 0.0019003 0.42099 2.0131 2.0117 16.0226 144.9059 0.00021724 -85.5396 0.49894
8.603 0.98814 5.4638e-005 3.8183 0.011917 0.0001118 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5925 0.58559 0.17897 0.0205 17.8734 0.12699 0.00016618 0.76318 0.0095019 0.010508 0.0014122 0.98661 0.99149 3.0487e-006 1.2195e-005 0.16562 0.85375 0.88154 0.0014107 0.96161 0.42913 0.0019001 0.421 2.0141 2.0127 16.0226 144.9059 0.00021694 -85.5405 0.49994
8.604 0.98814 5.4638e-005 3.8183 0.011917 0.00011181 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5926 0.58563 0.17898 0.020502 17.8765 0.127 0.00016619 0.76317 0.0095022 0.010508 0.0014121 0.98661 0.99149 3.0482e-006 1.2193e-005 0.16562 0.85415 0.88173 0.0014106 0.96184 0.42933 0.0019 0.42102 2.015 2.0137 16.0226 144.9059 0.00021664 -85.5414 0.50094
8.605 0.98814 5.4638e-005 3.8183 0.011917 0.00011182 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5927 0.58568 0.17899 0.020503 17.8796 0.127 0.0001662 0.76316 0.0095026 0.010509 0.0014119 0.98661 0.99149 3.0477e-006 1.2191e-005 0.16563 0.85456 0.88192 0.0014106 0.96207 0.42953 0.0018998 0.42103 2.016 2.0146 16.0225 144.9059 0.00021635 -85.5423 0.50194
8.606 0.98814 5.4638e-005 3.8183 0.011917 0.00011183 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5927 0.58572 0.17901 0.020504 17.8828 0.12701 0.00016621 0.76316 0.0095029 0.010509 0.0014117 0.98662 0.99149 3.0473e-006 1.2189e-005 0.16563 0.85496 0.88211 0.0014105 0.9623 0.42973 0.0018997 0.42105 2.0169 2.0156 16.0225 144.9059 0.00021605 -85.5432 0.50294
8.607 0.98814 5.4638e-005 3.8183 0.011917 0.00011185 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5928 0.58577 0.17902 0.020505 17.8859 0.12701 0.00016622 0.76315 0.0095033 0.010509 0.0014115 0.98662 0.99149 3.0468e-006 1.2187e-005 0.16563 0.85536 0.8823 0.0014104 0.96252 0.42993 0.0018995 0.42106 2.0179 2.0165 16.0225 144.906 0.00021576 -85.544 0.50394
8.608 0.98814 5.4638e-005 3.8183 0.011917 0.00011186 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5929 0.58581 0.17903 0.020506 17.8891 0.12702 0.00016623 0.76315 0.0095036 0.01051 0.0014113 0.98662 0.99149 3.0463e-006 1.2185e-005 0.16564 0.85576 0.88249 0.0014103 0.96274 0.43012 0.0018994 0.42108 2.0188 2.0175 16.0225 144.906 0.00021547 -85.5449 0.50494
8.609 0.98814 5.4638e-005 3.8183 0.011917 0.00011187 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.593 0.58586 0.17904 0.020507 17.8922 0.12703 0.00016624 0.76314 0.009504 0.01051 0.0014111 0.98662 0.9915 3.0459e-006 1.2183e-005 0.16564 0.85616 0.88268 0.0014102 0.96297 0.43032 0.0018993 0.42109 2.0198 2.0184 16.0225 144.906 0.00021518 -85.5458 0.50594
8.61 0.98814 5.4637e-005 3.8183 0.011917 0.00011188 0.001175 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5931 0.5859 0.17906 0.020508 17.8954 0.12703 0.00016624 0.76313 0.0095044 0.01051 0.0014109 0.98663 0.9915 3.0454e-006 1.2182e-005 0.16564 0.85656 0.88287 0.0014101 0.96319 0.43052 0.0018991 0.42111 2.0207 2.0194 16.0225 144.906 0.00021489 -85.5466 0.50694
8.611 0.98814 5.4637e-005 3.8183 0.011917 0.0001119 0.0011751 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5932 0.58595 0.17907 0.020509 17.8985 0.12704 0.00016625 0.76313 0.0095047 0.010511 0.0014107 0.98663 0.9915 3.0449e-006 1.218e-005 0.16564 0.85696 0.88306 0.00141 0.96341 0.43072 0.001899 0.42112 2.0217 2.0203 16.0225 144.906 0.0002146 -85.5475 0.50794
8.612 0.98814 5.4637e-005 3.8183 0.011917 0.00011191 0.0011751 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5933 0.58599 0.17908 0.02051 17.9017 0.12705 0.00016626 0.76312 0.0095051 0.010511 0.0014105 0.98663 0.9915 3.0445e-006 1.2178e-005 0.16565 0.85735 0.88324 0.0014099 0.96362 0.43092 0.0018989 0.42114 2.0226 2.0212 16.0225 144.9061 0.00021431 -85.5483 0.50894
8.613 0.98814 5.4637e-005 3.8183 0.011917 0.00011192 0.0011751 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5933 0.58604 0.1791 0.020511 17.9048 0.12705 0.00016627 0.76311 0.0095054 0.010512 0.0014103 0.98663 0.9915 3.044e-006 1.2176e-005 0.16565 0.85774 0.88343 0.0014097 0.96384 0.43111 0.0018987 0.42115 2.0235 2.0222 16.0225 144.9061 0.00021403 -85.5491 0.50994
8.614 0.98814 5.4637e-005 3.8183 0.011917 0.00011194 0.0011751 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5934 0.58608 0.17911 0.020512 17.9079 0.12706 0.00016628 0.76311 0.0095058 0.010512 0.0014101 0.98664 0.9915 3.0436e-006 1.2174e-005 0.16565 0.85814 0.88361 0.0014096 0.96405 0.43131 0.0018986 0.42117 2.0245 2.0231 16.0225 144.9061 0.00021374 -85.55 0.51094
8.615 0.98814 5.4637e-005 3.8183 0.011917 0.00011195 0.0011751 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5935 0.58612 0.17912 0.020513 17.9111 0.12706 0.00016629 0.7631 0.0095061 0.010512 0.0014099 0.98664 0.99151 3.0432e-006 1.2173e-005 0.16565 0.85853 0.88379 0.0014095 0.96427 0.43151 0.0018985 0.42118 2.0254 2.0241 16.0224 144.9061 0.00021346 -85.5508 0.51194
8.616 0.98814 5.4637e-005 3.8183 0.011917 0.00011196 0.0011751 0.23367 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5936 0.58617 0.17914 0.020514 17.9142 0.12707 0.0001663 0.7631 0.0095065 0.010513 0.0014097 0.98664 0.99151 3.0427e-006 1.2171e-005 0.16566 0.85892 0.88398 0.0014094 0.96448 0.43171 0.0018983 0.4212 2.0263 2.025 16.0224 144.9061 0.00021318 -85.5516 0.51294
8.617 0.98814 5.4637e-005 3.8183 0.011917 0.00011197 0.0011751 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5937 0.58621 0.17915 0.020515 17.9174 0.12708 0.00016631 0.76309 0.0095069 0.010513 0.0014095 0.98664 0.99151 3.0423e-006 1.2169e-005 0.16566 0.85931 0.88416 0.0014093 0.96469 0.4319 0.0018982 0.42121 2.0272 2.0259 16.0224 144.9062 0.0002129 -85.5524 0.51394
8.618 0.98814 5.4637e-005 3.8183 0.011917 0.00011199 0.0011751 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5938 0.58626 0.17916 0.020516 17.9205 0.12708 0.00016632 0.76308 0.0095072 0.010513 0.0014093 0.98665 0.99151 3.0418e-006 1.2167e-005 0.16566 0.8597 0.88434 0.0014092 0.9649 0.4321 0.0018981 0.42123 2.0282 2.0268 16.0224 144.9062 0.00021262 -85.5532 0.51494
8.619 0.98814 5.4637e-005 3.8183 0.011917 0.000112 0.0011751 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5938 0.5863 0.17918 0.020517 17.9237 0.12709 0.00016633 0.76308 0.0095076 0.010514 0.0014091 0.98665 0.99151 3.0414e-006 1.2166e-005 0.16567 0.86008 0.88452 0.0014091 0.96511 0.4323 0.0018979 0.42125 2.0291 2.0278 16.0224 144.9062 0.00021234 -85.554 0.51594
8.62 0.98814 5.4637e-005 3.8183 0.011917 0.00011201 0.0011751 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5939 0.58635 0.17919 0.020518 17.9268 0.1271 0.00016634 0.76307 0.0095079 0.010514 0.0014089 0.98665 0.99151 3.041e-006 1.2164e-005 0.16567 0.86047 0.8847 0.001409 0.96531 0.4325 0.0018978 0.42126 2.03 2.0287 16.0224 144.9062 0.00021206 -85.5548 0.51694
8.621 0.98814 5.4637e-005 3.8183 0.011917 0.00011203 0.0011751 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.594 0.58639 0.1792 0.020519 17.93 0.1271 0.00016635 0.76306 0.0095083 0.010515 0.0014087 0.98665 0.99152 3.0406e-006 1.2162e-005 0.16567 0.86085 0.88488 0.0014089 0.96552 0.43269 0.0018977 0.42128 2.0309 2.0296 16.0224 144.9062 0.00021178 -85.5556 0.51794
8.622 0.98814 5.4636e-005 3.8183 0.011917 0.00011204 0.0011751 0.23366 0.00065931 0.23432 0.21623 0 0.032261 0.0389 0 1.5941 0.58644 0.17922 0.02052 17.9331 0.12711 0.00016636 0.76306 0.0095087 0.010515 0.0014086 0.98666 0.99152 3.0401e-006 1.2161e-005 0.16567 0.86124 0.88506 0.0014088 0.96572 0.43289 0.0018976 0.42129 2.0318 2.0305 16.0224 144.9063 0.00021151 -85.5564 0.51894
8.623 0.98814 5.4636e-005 3.8183 0.011917 0.00011205 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5942 0.58648 0.17923 0.020521 17.9363 0.12711 0.00016637 0.76305 0.009509 0.010515 0.0014084 0.98666 0.99152 3.0397e-006 1.2159e-005 0.16568 0.86162 0.88524 0.0014087 0.96593 0.43309 0.0018974 0.42131 2.0327 2.0314 16.0223 144.9063 0.00021123 -85.5571 0.51994
8.624 0.98814 5.4636e-005 3.8183 0.011917 0.00011206 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5943 0.58653 0.17924 0.020522 17.9394 0.12712 0.00016638 0.76305 0.0095094 0.010516 0.0014082 0.98666 0.99152 3.0393e-006 1.2157e-005 0.16568 0.862 0.88542 0.0014086 0.96613 0.43328 0.0018973 0.42132 2.0336 2.0323 16.0223 144.9063 0.00021096 -85.5579 0.52094
8.625 0.98814 5.4636e-005 3.8183 0.011917 0.00011208 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5944 0.58657 0.17926 0.020524 17.9426 0.12713 0.00016639 0.76304 0.0095097 0.010516 0.001408 0.98666 0.99152 3.0389e-006 1.2156e-005 0.16568 0.86238 0.88559 0.0014085 0.96633 0.43348 0.0018972 0.42134 2.0345 2.0332 16.0223 144.9063 0.00021069 -85.5587 0.52194
8.626 0.98814 5.4636e-005 3.8183 0.011917 0.00011209 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5944 0.58661 0.17927 0.020525 17.9457 0.12713 0.0001664 0.76303 0.0095101 0.010517 0.0014078 0.98667 0.99152 3.0385e-006 1.2154e-005 0.16568 0.86276 0.88577 0.0014084 0.96653 0.43368 0.0018971 0.42135 2.0354 2.0341 16.0223 144.9063 0.00021041 -85.5594 0.52294
8.627 0.98814 5.4636e-005 3.8183 0.011917 0.0001121 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5945 0.58666 0.17928 0.020526 17.9489 0.12714 0.00016641 0.76303 0.0095104 0.010517 0.0014077 0.98667 0.99152 3.0381e-006 1.2152e-005 0.16569 0.86313 0.88594 0.0014083 0.96672 0.43387 0.0018969 0.42137 2.0363 2.035 16.0223 144.9064 0.00021014 -85.5602 0.52394
8.628 0.98814 5.4636e-005 3.8183 0.011917 0.00011212 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5946 0.5867 0.1793 0.020527 17.952 0.12715 0.00016642 0.76302 0.0095108 0.010517 0.0014075 0.98667 0.99153 3.0377e-006 1.2151e-005 0.16569 0.86351 0.88612 0.0014083 0.96692 0.43407 0.0018968 0.42138 2.0372 2.0359 16.0223 144.9064 0.00020987 -85.5609 0.52494
8.629 0.98814 5.4636e-005 3.8183 0.011917 0.00011213 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5947 0.58675 0.17931 0.020528 17.9552 0.12715 0.00016643 0.76301 0.0095111 0.010518 0.0014073 0.98667 0.99153 3.0373e-006 1.2149e-005 0.16569 0.86388 0.88629 0.0014082 0.96712 0.43427 0.0018967 0.4214 2.0381 2.0368 16.0223 144.9064 0.00020961 -85.5617 0.52594
8.63 0.98814 5.4636e-005 3.8183 0.011917 0.00011214 0.0011751 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5948 0.58679 0.17932 0.020529 17.9583 0.12716 0.00016644 0.76301 0.0095115 0.010518 0.0014071 0.98667 0.99153 3.0369e-006 1.2148e-005 0.1657 0.86426 0.88646 0.0014081 0.96731 0.43446 0.0018966 0.42141 2.039 2.0377 16.0223 144.9064 0.00020934 -85.5624 0.52694
8.631 0.98814 5.4636e-005 3.8183 0.011917 0.00011215 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5949 0.58684 0.17933 0.02053 17.9615 0.12716 0.00016644 0.763 0.0095119 0.010518 0.001407 0.98668 0.99153 3.0365e-006 1.2146e-005 0.1657 0.86463 0.88664 0.001408 0.9675 0.43466 0.0018965 0.42143 2.0399 2.0386 16.0222 144.9064 0.00020907 -85.5631 0.52794
8.632 0.98814 5.4636e-005 3.8183 0.011917 0.00011217 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5949 0.58688 0.17935 0.020531 17.9646 0.12717 0.00016645 0.763 0.0095122 0.010519 0.0014068 0.98668 0.99153 3.0361e-006 1.2144e-005 0.1657 0.865 0.88681 0.0014079 0.96769 0.43486 0.0018964 0.42144 2.0408 2.0395 16.0222 144.9065 0.00020881 -85.5639 0.52894
8.633 0.98814 5.4636e-005 3.8183 0.011917 0.00011218 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.595 0.58693 0.17936 0.020532 17.9678 0.12718 0.00016646 0.76299 0.0095126 0.010519 0.0014066 0.98668 0.99153 3.0357e-006 1.2143e-005 0.1657 0.86537 0.88698 0.0014078 0.96788 0.43505 0.0018962 0.42146 2.0417 2.0404 16.0222 144.9065 0.00020855 -85.5646 0.52994
8.634 0.98814 5.4635e-005 3.8183 0.011917 0.00011219 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5951 0.58697 0.17937 0.020533 17.9709 0.12718 0.00016647 0.76298 0.0095129 0.01052 0.0014064 0.98668 0.99153 3.0353e-006 1.2141e-005 0.16571 0.86574 0.88715 0.0014077 0.96807 0.43525 0.0018961 0.42147 2.0426 2.0413 16.0222 144.9065 0.00020828 -85.5653 0.53094
8.635 0.98814 5.4635e-005 3.8183 0.011917 0.0001122 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5952 0.58701 0.17939 0.020534 17.9741 0.12719 0.00016648 0.76298 0.0095133 0.01052 0.0014063 0.98669 0.99154 3.035e-006 1.214e-005 0.16571 0.86611 0.88732 0.0014076 0.96826 0.43545 0.001896 0.42149 2.0434 2.0422 16.0222 144.9065 0.00020802 -85.566 0.53194
8.636 0.98814 5.4635e-005 3.8183 0.011917 0.00011222 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5953 0.58706 0.1794 0.020535 17.9772 0.1272 0.00016649 0.76297 0.0095136 0.01052 0.0014061 0.98669 0.99154 3.0346e-006 1.2138e-005 0.16571 0.86647 0.88749 0.0014075 0.96845 0.43564 0.0018959 0.4215 2.0443 2.0431 16.0222 144.9065 0.00020776 -85.5667 0.53294
8.637 0.98814 5.4635e-005 3.8183 0.011917 0.00011223 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5954 0.5871 0.17941 0.020536 17.9804 0.1272 0.0001665 0.76297 0.009514 0.010521 0.001406 0.98669 0.99154 3.0342e-006 1.2137e-005 0.16571 0.86684 0.88766 0.0014074 0.96863 0.43584 0.0018958 0.42152 2.0452 2.0439 16.0222 144.9066 0.0002075 -85.5674 0.53394
8.638 0.98814 5.4635e-005 3.8183 0.011917 0.00011224 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5954 0.58715 0.17943 0.020537 17.9836 0.12721 0.00016651 0.76296 0.0095144 0.010521 0.0014058 0.98669 0.99154 3.0338e-006 1.2135e-005 0.16572 0.8672 0.88782 0.0014073 0.96882 0.43604 0.0018957 0.42153 2.0461 2.0448 16.0222 144.9066 0.00020724 -85.5681 0.53494
8.639 0.98814 5.4635e-005 3.8183 0.011917 0.00011226 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5955 0.58719 0.17944 0.020538 17.9867 0.12721 0.00016652 0.76295 0.0095147 0.010521 0.0014056 0.98669 0.99154 3.0335e-006 1.2134e-005 0.16572 0.86757 0.88799 0.0014073 0.969 0.43623 0.0018956 0.42155 2.0469 2.0457 16.0221 144.9066 0.00020699 -85.5688 0.53594
8.64 0.98814 5.4635e-005 3.8183 0.011917 0.00011227 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5956 0.58724 0.17945 0.020539 17.9899 0.12722 0.00016653 0.76295 0.0095151 0.010522 0.0014055 0.9867 0.99154 3.0331e-006 1.2132e-005 0.16572 0.86793 0.88816 0.0014072 0.96918 0.43643 0.0018954 0.42156 2.0478 2.0466 16.0221 144.9066 0.00020673 -85.5695 0.53694
8.641 0.98814 5.4635e-005 3.8183 0.011917 0.00011228 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5957 0.58728 0.17947 0.02054 17.993 0.12723 0.00016654 0.76294 0.0095154 0.010522 0.0014053 0.9867 0.99154 3.0327e-006 1.2131e-005 0.16573 0.86829 0.88832 0.0014071 0.96936 0.43662 0.0018953 0.42158 2.0487 2.0474 16.0221 144.9066 0.00020647 -85.5702 0.53794
8.642 0.98814 5.4635e-005 3.8183 0.011916 0.00011229 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5958 0.58733 0.17948 0.020541 17.9962 0.12723 0.00016655 0.76293 0.0095158 0.010523 0.0014051 0.9867 0.99155 3.0324e-006 1.2129e-005 0.16573 0.86865 0.88849 0.001407 0.96954 0.43682 0.0018952 0.42159 2.0495 2.0483 16.0221 144.9067 0.00020622 -85.5708 0.53894
8.643 0.98814 5.4635e-005 3.8183 0.011916 0.00011231 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.5959 0.58737 0.17949 0.020542 17.9993 0.12724 0.00016656 0.76293 0.0095161 0.010523 0.001405 0.9867 0.99155 3.032e-006 1.2128e-005 0.16573 0.86901 0.88865 0.0014069 0.96972 0.43702 0.0018951 0.42161 2.0504 2.0492 16.0221 144.9067 0.00020597 -85.5715 0.53994
8.644 0.98814 5.4635e-005 3.8183 0.011916 0.00011232 0.0011752 0.23366 0.00065931 0.23432 0.21622 0 0.032261 0.0389 0 1.596 0.58742 0.17951 0.020543 18.0025 0.12724 0.00016657 0.76292 0.0095165 0.010523 0.0014048 0.9867 0.99155 3.0317e-006 1.2127e-005 0.16573 0.86937 0.88882 0.0014069 0.9699 0.43721 0.001895 0.42162 2.0513 2.05 16.0221 144.9067 0.00020571 -85.5722 0.54094
8.645 0.98814 5.4635e-005 3.8183 0.011916 0.00011233 0.0011752 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.596 0.58746 0.17952 0.020544 18.0056 0.12725 0.00016658 0.76292 0.0095169 0.010524 0.0014047 0.98671 0.99155 3.0313e-006 1.2125e-005 0.16574 0.86972 0.88898 0.0014068 0.97007 0.43741 0.0018949 0.42164 2.0521 2.0509 16.0221 144.9067 0.00020546 -85.5728 0.54194
8.646 0.98814 5.4634e-005 3.8183 0.011916 0.00011235 0.0011752 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5961 0.5875 0.17953 0.020545 18.0088 0.12726 0.00016659 0.76291 0.0095172 0.010524 0.0014046 0.98671 0.99155 3.0309e-006 1.2124e-005 0.16574 0.87008 0.88914 0.0014067 0.97025 0.4376 0.0018948 0.42165 2.053 2.0518 16.022 144.9067 0.00020521 -85.5735 0.54294
8.647 0.98814 5.4634e-005 3.8183 0.011916 0.00011236 0.0011752 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5962 0.58755 0.17955 0.020547 18.012 0.12726 0.0001666 0.7629 0.0095176 0.010524 0.0014044 0.98671 0.99155 3.0306e-006 1.2122e-005 0.16574 0.87043 0.8893 0.0014066 0.97042 0.4378 0.0018947 0.42167 2.0538 2.0526 16.022 144.9068 0.00020496 -85.5741 0.54394
8.648 0.98814 5.4634e-005 3.8183 0.011916 0.00011237 0.0011752 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5963 0.58759 0.17956 0.020548 18.0151 0.12727 0.00016661 0.7629 0.0095179 0.010525 0.0014043 0.98671 0.99155 3.0303e-006 1.2121e-005 0.16574 0.87079 0.88946 0.0014066 0.9706 0.43799 0.0018946 0.42168 2.0547 2.0535 16.022 144.9068 0.00020472 -85.5748 0.54494
8.649 0.98814 5.4634e-005 3.8183 0.011916 0.00011238 0.0011752 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5964 0.58764 0.17957 0.020549 18.0183 0.12728 0.00016662 0.76289 0.0095183 0.010525 0.0014041 0.98671 0.99155 3.0299e-006 1.212e-005 0.16575 0.87114 0.88962 0.0014065 0.97077 0.43819 0.0018945 0.4217 2.0555 2.0543 16.022 144.9068 0.00020447 -85.5754 0.54594
8.65 0.98814 5.4634e-005 3.8183 0.011916 0.0001124 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5965 0.58768 0.17959 0.02055 18.0214 0.12728 0.00016662 0.76288 0.0095186 0.010526 0.001404 0.98672 0.99156 3.0296e-006 1.2118e-005 0.16575 0.87149 0.88978 0.0014064 0.97094 0.43838 0.0018944 0.42171 2.0564 2.0552 16.022 144.9068 0.00020422 -85.5761 0.54694
8.651 0.98814 5.4634e-005 3.8183 0.011916 0.00011241 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5965 0.58773 0.1796 0.020551 18.0246 0.12729 0.00016663 0.76288 0.009519 0.010526 0.0014038 0.98672 0.99156 3.0292e-006 1.2117e-005 0.16575 0.87184 0.88994 0.0014063 0.97111 0.43858 0.0018943 0.42173 2.0572 2.056 16.022 144.9068 0.00020398 -85.5767 0.54794
8.652 0.98814 5.4634e-005 3.8183 0.011916 0.00011242 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5966 0.58777 0.17961 0.020552 18.0278 0.12729 0.00016664 0.76287 0.0095193 0.010526 0.0014037 0.98672 0.99156 3.0289e-006 1.2115e-005 0.16576 0.87219 0.8901 0.0014062 0.97128 0.43877 0.0018942 0.42174 2.058 2.0569 16.022 144.9069 0.00020373 -85.5773 0.54894
8.653 0.98814 5.4634e-005 3.8183 0.011916 0.00011243 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5967 0.58782 0.17962 0.020553 18.0309 0.1273 0.00016665 0.76287 0.0095197 0.010527 0.0014035 0.98672 0.99156 3.0286e-006 1.2114e-005 0.16576 0.87254 0.89026 0.0014062 0.97144 0.43897 0.0018941 0.42176 2.0589 2.0577 16.0219 144.9069 0.00020349 -85.5779 0.54994
8.654 0.98814 5.4634e-005 3.8183 0.011916 0.00011245 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5968 0.58786 0.17964 0.020554 18.0341 0.12731 0.00016666 0.76286 0.0095201 0.010527 0.0014034 0.98672 0.99156 3.0282e-006 1.2113e-005 0.16576 0.87288 0.89042 0.0014061 0.97161 0.43916 0.001894 0.42177 2.0597 2.0585 16.0219 144.9069 0.00020325 -85.5786 0.55094
8.655 0.98814 5.4634e-005 3.8183 0.011916 0.00011246 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5969 0.5879 0.17965 0.020555 18.0372 0.12731 0.00016667 0.76285 0.0095204 0.010527 0.0014032 0.98673 0.99156 3.0279e-006 1.2111e-005 0.16576 0.87323 0.89057 0.001406 0.97177 0.43936 0.0018939 0.42179 2.0606 2.0594 16.0219 144.9069 0.00020301 -85.5792 0.55194
8.656 0.98814 5.4634e-005 3.8183 0.011916 0.00011247 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.597 0.58795 0.17966 0.020556 18.0404 0.12732 0.00016668 0.76285 0.0095208 0.010528 0.0014031 0.98673 0.99156 3.0276e-006 1.211e-005 0.16577 0.87357 0.89073 0.0014059 0.97194 0.43955 0.0018938 0.4218 2.0614 2.0602 16.0219 144.9069 0.00020277 -85.5798 0.55294
8.657 0.98814 5.4634e-005 3.8183 0.011916 0.00011249 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.597 0.58799 0.17968 0.020557 18.0436 0.12733 0.00016669 0.76284 0.0095211 0.010528 0.0014029 0.98673 0.99156 3.0272e-006 1.2109e-005 0.16577 0.87392 0.89088 0.0014058 0.9721 0.43975 0.0018937 0.42182 2.0622 2.061 16.0219 144.907 0.00020253 -85.5804 0.55394
8.658 0.98814 5.4633e-005 3.8183 0.011916 0.0001125 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5971 0.58804 0.17969 0.020558 18.0467 0.12733 0.0001667 0.76283 0.0095215 0.010529 0.0014028 0.98673 0.99157 3.0269e-006 1.2108e-005 0.16577 0.87426 0.89104 0.0014058 0.97226 0.43994 0.0018936 0.42183 2.063 2.0619 16.0219 144.907 0.00020229 -85.581 0.55494
8.659 0.98814 5.4633e-005 3.8183 0.011916 0.00011251 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5972 0.58808 0.1797 0.020559 18.0499 0.12734 0.00016671 0.76283 0.0095218 0.010529 0.0014026 0.98673 0.99157 3.0266e-006 1.2106e-005 0.16577 0.8746 0.89119 0.0014057 0.97242 0.44014 0.0018935 0.42185 2.0639 2.0627 16.0219 144.907 0.00020205 -85.5816 0.55594
8.66 0.98814 5.4633e-005 3.8183 0.011916 0.00011252 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5973 0.58813 0.17972 0.02056 18.053 0.12734 0.00016672 0.76282 0.0095222 0.010529 0.0014025 0.98673 0.99157 3.0263e-006 1.2105e-005 0.16578 0.87494 0.89135 0.0014056 0.97258 0.44033 0.0018934 0.42186 2.0647 2.0635 16.0218 144.907 0.00020181 -85.5822 0.55694
8.661 0.98814 5.4633e-005 3.8183 0.011916 0.00011254 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5974 0.58817 0.17973 0.020561 18.0562 0.12735 0.00016673 0.76282 0.0095225 0.01053 0.0014024 0.98674 0.99157 3.026e-006 1.2104e-005 0.16578 0.87528 0.8915 0.0014055 0.97274 0.44053 0.0018933 0.42188 2.0655 2.0644 16.0218 144.907 0.00020158 -85.5828 0.55794
8.662 0.98814 5.4633e-005 3.8183 0.011916 0.00011255 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5975 0.58822 0.17974 0.020562 18.0594 0.12736 0.00016674 0.76281 0.0095229 0.01053 0.0014022 0.98674 0.99157 3.0256e-006 1.2103e-005 0.16578 0.87562 0.89165 0.0014055 0.9729 0.44072 0.0018932 0.42189 2.0663 2.0652 16.0218 144.9071 0.00020134 -85.5834 0.55894
8.663 0.98814 5.4633e-005 3.8183 0.011916 0.00011256 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5976 0.58826 0.17976 0.020563 18.0625 0.12736 0.00016675 0.7628 0.0095232 0.01053 0.0014021 0.98674 0.99157 3.0253e-006 1.2101e-005 0.16579 0.87595 0.8918 0.0014054 0.97306 0.44092 0.0018931 0.42191 2.0671 2.066 16.0218 144.9071 0.00020111 -85.5839 0.55994
8.664 0.98814 5.4633e-005 3.8183 0.011916 0.00011258 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5976 0.5883 0.17977 0.020564 18.0657 0.12737 0.00016676 0.7628 0.0095236 0.010531 0.0014019 0.98674 0.99157 3.025e-006 1.21e-005 0.16579 0.87629 0.89196 0.0014053 0.97321 0.44111 0.001893 0.42192 2.068 2.0668 16.0218 144.9071 0.00020088 -85.5845 0.56094
8.665 0.98814 5.4633e-005 3.8183 0.011916 0.00011259 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5977 0.58835 0.17978 0.020565 18.0688 0.12738 0.00016677 0.76279 0.009524 0.010531 0.0014018 0.98674 0.99157 3.0247e-006 1.2099e-005 0.16579 0.87662 0.89211 0.0014053 0.97337 0.44131 0.0018929 0.42194 2.0688 2.0676 16.0218 144.9071 0.00020064 -85.5851 0.56194
8.666 0.98814 5.4633e-005 3.8183 0.011916 0.0001126 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5978 0.58839 0.1798 0.020566 18.072 0.12738 0.00016678 0.76279 0.0095243 0.010532 0.0014017 0.98674 0.99158 3.0244e-006 1.2098e-005 0.16579 0.87696 0.89226 0.0014052 0.97352 0.4415 0.0018928 0.42195 2.0696 2.0684 16.0217 144.9071 0.00020041 -85.5857 0.56294
8.667 0.98814 5.4633e-005 3.8183 0.011916 0.00011261 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5979 0.58844 0.17981 0.020567 18.0752 0.12739 0.00016679 0.76278 0.0095247 0.010532 0.0014015 0.98675 0.99158 3.0241e-006 1.2096e-005 0.1658 0.87729 0.89241 0.0014051 0.97368 0.4417 0.0018928 0.42197 2.0704 2.0693 16.0217 144.9072 0.00020018 -85.5862 0.56394
8.668 0.98814 5.4633e-005 3.8183 0.011916 0.00011263 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.598 0.58848 0.17982 0.020568 18.0783 0.12739 0.0001668 0.76277 0.009525 0.010532 0.0014014 0.98675 0.99158 3.0238e-006 1.2095e-005 0.1658 0.87762 0.89256 0.0014051 0.97383 0.44189 0.0018927 0.42199 2.0712 2.0701 16.0217 144.9072 0.00019995 -85.5868 0.56494
8.669 0.98814 5.4633e-005 3.8183 0.011916 0.00011264 0.0011753 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5981 0.58853 0.17984 0.020569 18.0815 0.1274 0.0001668 0.76277 0.0095254 0.010533 0.0014013 0.98675 0.99158 3.0235e-006 1.2094e-005 0.1658 0.87795 0.8927 0.001405 0.97398 0.44208 0.0018926 0.422 2.072 2.0709 16.0217 144.9072 0.00019972 -85.5874 0.56594
8.67 0.98814 5.4632e-005 3.8183 0.011916 0.00011265 0.0011754 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5981 0.58857 0.17985 0.020571 18.0847 0.12741 0.00016681 0.76276 0.0095257 0.010533 0.0014012 0.98675 0.99158 3.0232e-006 1.2093e-005 0.1658 0.87828 0.89285 0.0014049 0.97413 0.44228 0.0018925 0.42202 2.0728 2.0717 16.0217 144.9072 0.0001995 -85.5879 0.56694
8.671 0.98814 5.4632e-005 3.8183 0.011916 0.00011267 0.0011754 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5982 0.58862 0.17986 0.020572 18.0878 0.12741 0.00016682 0.76275 0.0095261 0.010533 0.001401 0.98675 0.99158 3.0229e-006 1.2092e-005 0.16581 0.87861 0.893 0.0014049 0.97428 0.44247 0.0018924 0.42203 2.0736 2.0725 16.0217 144.9072 0.00019927 -85.5885 0.56794
8.672 0.98814 5.4632e-005 3.8183 0.011916 0.00011268 0.0011754 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5983 0.58866 0.17987 0.020573 18.091 0.12742 0.00016683 0.76275 0.0095264 0.010534 0.0014009 0.98675 0.99158 3.0226e-006 1.209e-005 0.16581 0.87894 0.89314 0.0014048 0.97443 0.44267 0.0018923 0.42205 2.0744 2.0733 16.0216 144.9073 0.00019904 -85.589 0.56894
8.673 0.98815 5.4632e-005 3.8183 0.011916 0.00011269 0.0011754 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5984 0.5887 0.17989 0.020574 18.0942 0.12742 0.00016684 0.76274 0.0095268 0.010534 0.0014008 0.98676 0.99158 3.0224e-006 1.2089e-005 0.16581 0.87927 0.89329 0.0014047 0.97457 0.44286 0.0018922 0.42206 2.0752 2.0741 16.0216 144.9073 0.00019882 -85.5895 0.56994
8.674 0.98815 5.4632e-005 3.8183 0.011916 0.0001127 0.0011754 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5985 0.58875 0.1799 0.020575 18.0973 0.12743 0.00016685 0.76274 0.0095272 0.010535 0.0014007 0.98676 0.99158 3.0221e-006 1.2088e-005 0.16582 0.87959 0.89344 0.0014047 0.97472 0.44305 0.0018921 0.42208 2.076 2.0749 16.0216 144.9073 0.0001986 -85.5901 0.57094
8.675 0.98815 5.4632e-005 3.8183 0.011916 0.00011272 0.0011754 0.23366 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5986 0.58879 0.17991 0.020576 18.1005 0.12744 0.00016686 0.76273 0.0095275 0.010535 0.0014005 0.98676 0.99158 3.0218e-006 1.2087e-005 0.16582 0.87992 0.89358 0.0014046 0.97486 0.44325 0.001892 0.42209 2.0768 2.0757 16.0216 144.9073 0.00019837 -85.5906 0.57194
8.676 0.98815 5.4632e-005 3.8183 0.011916 0.00011273 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5986 0.58884 0.17993 0.020577 18.1037 0.12744 0.00016687 0.76272 0.0095279 0.010535 0.0014004 0.98676 0.99159 3.0215e-006 1.2086e-005 0.16582 0.88024 0.89373 0.0014045 0.97501 0.44344 0.001892 0.42211 2.0776 2.0765 16.0216 144.9073 0.00019815 -85.5911 0.57294
8.677 0.98815 5.4632e-005 3.8183 0.011916 0.00011274 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5987 0.58888 0.17994 0.020578 18.1068 0.12745 0.00016688 0.76272 0.0095282 0.010536 0.0014003 0.98676 0.99159 3.0212e-006 1.2085e-005 0.16582 0.88056 0.89387 0.0014045 0.97515 0.44363 0.0018919 0.42212 2.0784 2.0773 16.0216 144.9074 0.00019793 -85.5917 0.57394
8.678 0.98815 5.4632e-005 3.8183 0.011916 0.00011275 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5988 0.58893 0.17995 0.020579 18.11 0.12746 0.00016689 0.76271 0.0095286 0.010536 0.0014001 0.98676 0.99159 3.0209e-006 1.2084e-005 0.16583 0.88088 0.89401 0.0014044 0.97529 0.44383 0.0018918 0.42214 2.0792 2.0781 16.0215 144.9074 0.00019771 -85.5922 0.57494
8.679 0.98815 5.4632e-005 3.8183 0.011916 0.00011277 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5989 0.58897 0.17997 0.02058 18.1132 0.12746 0.0001669 0.7627 0.0095289 0.010536 0.0014 0.98677 0.99159 3.0206e-006 1.2083e-005 0.16583 0.8812 0.89416 0.0014043 0.97544 0.44402 0.0018917 0.42215 2.0799 2.0788 16.0215 144.9074 0.00019749 -85.5927 0.57594
8.68 0.98815 5.4632e-005 3.8183 0.011916 0.00011278 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.599 0.58902 0.17998 0.020581 18.1163 0.12747 0.00016691 0.7627 0.0095293 0.010537 0.0013999 0.98677 0.99159 3.0204e-006 1.2081e-005 0.16583 0.88152 0.8943 0.0014043 0.97558 0.44421 0.0018916 0.42217 2.0807 2.0796 16.0215 144.9074 0.00019727 -85.5932 0.57694
8.681 0.98815 5.4632e-005 3.8183 0.011916 0.00011279 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5991 0.58906 0.17999 0.020582 18.1195 0.12747 0.00016692 0.76269 0.0095296 0.010537 0.0013998 0.98677 0.99159 3.0201e-006 1.208e-005 0.16583 0.88184 0.89444 0.0014042 0.97572 0.44441 0.0018915 0.42218 2.0815 2.0804 16.0215 144.9074 0.00019705 -85.5937 0.57794
8.682 0.98815 5.4631e-005 3.8183 0.011916 0.00011281 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5992 0.58911 0.18001 0.020583 18.1227 0.12748 0.00016693 0.76269 0.00953 0.010538 0.0013997 0.98677 0.99159 3.0198e-006 1.2079e-005 0.16584 0.88216 0.89458 0.0014041 0.97586 0.4446 0.0018915 0.4222 2.0823 2.0812 16.0215 144.9075 0.00019684 -85.5942 0.57894
8.683 0.98815 5.4631e-005 3.8183 0.011916 0.00011282 0.0011754 0.23365 0.00065931 0.23431 0.21622 0 0.032261 0.0389 0 1.5992 0.58915 0.18002 0.020584 18.1258 0.12749 0.00016694 0.76268 0.0095303 0.010538 0.0013996 0.98677 0.99159 3.0196e-006 1.2078e-005 0.16584 0.88248 0.89472 0.0014041 0.97599 0.44479 0.0018914 0.42221 2.0831 2.082 16.0215 144.9075 0.00019662 -85.5947 0.57994
8.684 0.98815 5.4631e-005 3.8183 0.011916 0.00011283 0.0011754 0.23365 0.00065931 0.23431 0.21621 0 0.032261 0.0389 0 1.5993 0.58919 0.18003 0.020585 18.129 0.12749 0.00016695 0.76267 0.0095307 0.010538 0.0013994 0.98677 0.99159 3.0193e-006 1.2077e-005 0.16584 0.88279 0.89486 0.001404 0.97613 0.44499 0.0018913 0.42223 2.0838 2.0827 16.0214 144.9075 0.0001964 -85.5952 0.58094
8.685 0.98815 5.4631e-005 3.8183 0.011916 0.00011284 0.0011754 0.23365 0.00065931 0.23431 0.21621 0 0.032261 0.0389 0 1.5994 0.58924 0.18005 0.020586 18.1322 0.1275 0.00016696 0.76267 0.009531 0.010539 0.0013993 0.98678 0.99159 3.019e-006 1.2076e-005 0.16585 0.88311 0.895 0.001404 0.97627 0.44518 0.0018912 0.42224 2.0846 2.0835 16.0214 144.9075 0.00019619 -85.5957 0.58194
8.686 0.98815 5.4631e-005 3.8183 0.011916 0.00011286 0.0011754 0.23365 0.00065931 0.23431 0.21621 0 0.032261 0.0389 0 1.5995 0.58928 0.18006 0.020587 18.1354 0.12751 0.00016697 0.76266 0.0095314 0.010539 0.0013992 0.98678 0.9916 3.0188e-006 1.2075e-005 0.16585 0.88342 0.89514 0.0014039 0.9764 0.44537 0.0018911 0.42226 2.0854 2.0843 16.0214 144.9075 0.00019598 -85.5962 0.58294
8.687 0.98815 5.4631e-005 3.8183 0.011916 0.00011287 0.0011754 0.23365 0.00065931 0.23431 0.21621 0 0.032261 0.0389 0 1.5996 0.58933 0.18007 0.020588 18.1385 0.12751 0.00016698 0.76266 0.0095318 0.010539 0.0013991 0.98678 0.9916 3.0185e-006 1.2074e-005 0.16585 0.88373 0.89528 0.0014038 0.97654 0.44557 0.0018911 0.42227 2.0861 2.0851 16.0214 144.9076 0.00019576 -85.5967 0.58394
8.688 0.98815 5.4631e-005 3.8183 0.011916 0.00011288 0.0011754 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.5997 0.58937 0.18009 0.020589 18.1417 0.12752 0.00016698 0.76265 0.0095321 0.01054 0.001399 0.98678 0.9916 3.0182e-006 1.2073e-005 0.16585 0.88405 0.89541 0.0014038 0.97667 0.44576 0.001891 0.42229 2.0869 2.0858 16.0214 144.9076 0.00019555 -85.5972 0.58494
8.689 0.98815 5.4631e-005 3.8183 0.011916 0.0001129 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.5997 0.58942 0.1801 0.02059 18.1449 0.12752 0.00016699 0.76264 0.0095325 0.01054 0.0013989 0.98678 0.9916 3.018e-006 1.2072e-005 0.16586 0.88436 0.89555 0.0014037 0.9768 0.44595 0.0018909 0.4223 2.0877 2.0866 16.0213 144.9076 0.00019534 -85.5977 0.58594
8.69 0.98815 5.4631e-005 3.8183 0.011916 0.00011291 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.5998 0.58946 0.18011 0.020591 18.148 0.12753 0.000167 0.76264 0.0095328 0.010541 0.0013988 0.98678 0.9916 3.0177e-006 1.2071e-005 0.16586 0.88467 0.89569 0.0014037 0.97694 0.44615 0.0018908 0.42232 2.0884 2.0874 16.0213 144.9076 0.00019513 -85.5982 0.58694
8.691 0.98815 5.4631e-005 3.8183 0.011916 0.00011292 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.5999 0.58951 0.18012 0.020592 18.1512 0.12754 0.00016701 0.76263 0.0095332 0.010541 0.0013987 0.98678 0.9916 3.0175e-006 1.207e-005 0.16586 0.88497 0.89582 0.0014036 0.97707 0.44634 0.0018908 0.42233 2.0892 2.0881 16.0213 144.9076 0.00019492 -85.5986 0.58794
8.692 0.98815 5.4631e-005 3.8183 0.011916 0.00011293 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6 0.58955 0.18014 0.020593 18.1544 0.12754 0.00016702 0.76262 0.0095335 0.010541 0.0013986 0.98679 0.9916 3.0172e-006 1.2069e-005 0.16586 0.88528 0.89596 0.0014036 0.9772 0.44653 0.0018907 0.42235 2.0899 2.0889 16.0213 144.9077 0.00019471 -85.5991 0.58894
8.693 0.98815 5.4631e-005 3.8183 0.011916 0.00011295 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6001 0.58959 0.18015 0.020594 18.1576 0.12755 0.00016703 0.76262 0.0095339 0.010542 0.0013984 0.98679 0.9916 3.017e-006 1.2068e-005 0.16587 0.88559 0.8961 0.0014035 0.97733 0.44672 0.0018906 0.42236 2.0907 2.0897 16.0213 144.9077 0.0001945 -85.5996 0.58994
8.694 0.98815 5.463e-005 3.8183 0.011916 0.00011296 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6002 0.58964 0.18016 0.020596 18.1607 0.12755 0.00016704 0.76261 0.0095342 0.010542 0.0013983 0.98679 0.9916 3.0167e-006 1.2067e-005 0.16587 0.8859 0.89623 0.0014034 0.97745 0.44692 0.0018905 0.42238 2.0915 2.0904 16.0213 144.9077 0.0001943 -85.6 0.59094
8.695 0.98815 5.463e-005 3.8183 0.011916 0.00011297 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6002 0.58968 0.18018 0.020597 18.1639 0.12756 0.00016705 0.76261 0.0095346 0.010542 0.0013982 0.98679 0.9916 3.0165e-006 1.2066e-005 0.16587 0.8862 0.89636 0.0014034 0.97758 0.44711 0.0018905 0.42239 2.0922 2.0912 16.0212 144.9077 0.00019409 -85.6005 0.59194
8.696 0.98815 5.463e-005 3.8183 0.011916 0.00011298 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6003 0.58973 0.18019 0.020598 18.1671 0.12757 0.00016706 0.7626 0.0095349 0.010543 0.0013981 0.98679 0.99161 3.0162e-006 1.2065e-005 0.16588 0.8865 0.8965 0.0014033 0.97771 0.4473 0.0018904 0.42241 2.093 2.0919 16.0212 144.9077 0.00019388 -85.601 0.59294
8.697 0.98815 5.463e-005 3.8183 0.011916 0.000113 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6004 0.58977 0.1802 0.020599 18.1702 0.12757 0.00016707 0.76259 0.0095353 0.010543 0.001398 0.98679 0.99161 3.016e-006 1.2064e-005 0.16588 0.88681 0.89663 0.0014033 0.97784 0.44749 0.0018903 0.42242 2.0937 2.0927 16.0212 144.9078 0.00019368 -85.6014 0.59394
8.698 0.98815 5.463e-005 3.8183 0.011915 0.00011301 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6005 0.58982 0.18022 0.0206 18.1734 0.12758 0.00016708 0.76259 0.0095356 0.010544 0.0013979 0.98679 0.99161 3.0158e-006 1.2063e-005 0.16588 0.88711 0.89676 0.0014032 0.97796 0.44769 0.0018902 0.42244 2.0945 2.0934 16.0212 144.9078 0.00019348 -85.6019 0.59494
8.699 0.98815 5.463e-005 3.8183 0.011915 0.00011302 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6006 0.58986 0.18023 0.020601 18.1766 0.12759 0.00016709 0.76258 0.009536 0.010544 0.0013978 0.9868 0.99161 3.0155e-006 1.2062e-005 0.16588 0.88741 0.8969 0.0014032 0.97808 0.44788 0.0018902 0.42245 2.0952 2.0942 16.0212 144.9078 0.00019327 -85.6023 0.59594
8.7 0.98815 5.463e-005 3.8183 0.011915 0.00011304 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6007 0.58991 0.18024 0.020602 18.1798 0.12759 0.0001671 0.76258 0.0095363 0.010544 0.0013977 0.9868 0.99161 3.0153e-006 1.2061e-005 0.16589 0.88771 0.89703 0.0014031 0.97821 0.44807 0.0018901 0.42247 2.0959 2.0949 16.0211 144.9078 0.00019307 -85.6028 0.59694
8.701 0.98815 5.463e-005 3.8183 0.011915 0.00011305 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6007 0.58995 0.18026 0.020603 18.1829 0.1276 0.00016711 0.76257 0.0095367 0.010545 0.0013976 0.9868 0.99161 3.0151e-006 1.206e-005 0.16589 0.88801 0.89716 0.0014031 0.97833 0.44826 0.00189 0.42248 2.0967 2.0957 16.0211 144.9078 0.00019287 -85.6032 0.59794
8.702 0.98815 5.463e-005 3.8183 0.011915 0.00011306 0.0011755 0.23365 0.00065931 0.23431 0.21621 0 0.032262 0.0389 0 1.6008 0.58999 0.18027 0.020604 18.1861 0.1276 0.00016712 0.76256 0.0095371 0.010545 0.0013975 0.9868 0.99161 3.0148e-006 1.2059e-005 0.16589 0.88831 0.89729 0.001403 0.97845 0.44845 0.00189 0.4225 2.0974 2.0964 16.0211 144.9079 0.00019267 -85.6036 0.59894
8.703 0.98815 5.463e-005 3.8183 0.011915 0.00011307 0.0011755 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6009 0.59004 0.18028 0.020605 18.1893 0.12761 0.00016713 0.76256 0.0095374 0.010545 0.0013974 0.9868 0.99161 3.0146e-006 1.2058e-005 0.16589 0.88861 0.89742 0.001403 0.97857 0.44865 0.0018899 0.42251 2.0982 2.0971 16.0211 144.9079 0.00019247 -85.6041 0.59994
8.704 0.98815 5.463e-005 3.8183 0.011915 0.00011309 0.0011755 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.601 0.59008 0.1803 0.020606 18.1925 0.12762 0.00016714 0.76255 0.0095378 0.010546 0.0013973 0.9868 0.99161 3.0144e-006 1.2057e-005 0.1659 0.8889 0.89755 0.0014029 0.9787 0.44884 0.0018898 0.42253 2.0989 2.0979 16.0211 144.9079 0.00019227 -85.6045 0.60094
8.705 0.98815 5.463e-005 3.8183 0.011915 0.0001131 0.0011755 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6011 0.59013 0.18031 0.020607 18.1956 0.12762 0.00016714 0.76254 0.0095381 0.010546 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.1659 0.8892 0.89768 0.0014028 0.97882 0.44903 0.0018897 0.42254 2.0996 2.0986 16.0211 144.9079 0.00019207 -85.6049 0.60194
8.706 0.98815 5.4629e-005 3.8183 0.011915 0.00011311 0.0011755 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6012 0.59017 0.18032 0.020608 18.1988 0.12763 0.00016715 0.76254 0.0095385 0.010547 0.0013971 0.9868 0.99161 3.0139e-006 1.2056e-005 0.1659 0.88949 0.89781 0.0014028 0.97893 0.44922 0.0018897 0.42256 2.1004 2.0993 16.021 144.9079 0.00019187 -85.6054 0.60294
8.707 0.98815 5.4629e-005 3.8183 0.011915 0.00011313 0.0011755 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6013 0.59022 0.18033 0.020609 18.202 0.12763 0.00016716 0.76253 0.0095388 0.010547 0.001397 0.98681 0.99161 3.0137e-006 1.2055e-005 0.16591 0.88979 0.89793 0.0014027 0.97905 0.44941 0.0018896 0.42257 2.1011 2.1001 16.021 144.908 0.00019168 -85.6058 0.60394
8.708 0.98815 5.4629e-005 3.8183 0.011915 0.00011314 0.0011755 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6013 0.59026 0.18035 0.02061 18.2052 0.12764 0.00016717 0.76253 0.0095392 0.010547 0.0013969 0.98681 0.99162 3.0134e-006 1.2054e-005 0.16591 0.89008 0.89806 0.0014027 0.97917 0.4496 0.0018895 0.42259 2.1018 2.1008 16.021 144.908 0.00019148 -85.6062 0.60494
8.709 0.98815 5.4629e-005 3.8183 0.011915 0.00011315 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6014 0.59031 0.18036 0.020611 18.2084 0.12765 0.00016718 0.76252 0.0095395 0.010548 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.16591 0.89037 0.89819 0.0014026 0.97929 0.4498 0.0018895 0.4226 2.1025 2.1015 16.021 144.908 0.00019128 -85.6066 0.60594
8.71 0.98815 5.4629e-005 3.8183 0.011915 0.00011316 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6015 0.59035 0.18037 0.020612 18.2115 0.12765 0.00016719 0.76251 0.0095399 0.010548 0.0013967 0.98681 0.99162 3.013e-006 1.2052e-005 0.16591 0.89066 0.89831 0.0014026 0.9794 0.44999 0.0018894 0.42262 2.1033 2.1023 16.021 144.908 0.00019109 -85.607 0.60694
8.711 0.98815 5.4629e-005 3.8183 0.011915 0.00011318 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6016 0.59039 0.18039 0.020613 18.2147 0.12766 0.0001672 0.76251 0.0095402 0.010548 0.0013966 0.98681 0.99162 3.0128e-006 1.2051e-005 0.16592 0.89095 0.89844 0.0014025 0.97952 0.45018 0.0018893 0.42263 2.104 2.103 16.0209 144.908 0.0001909 -85.6075 0.60794
8.712 0.98815 5.4629e-005 3.8183 0.011915 0.00011319 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6017 0.59044 0.1804 0.020614 18.2179 0.12767 0.00016721 0.7625 0.0095406 0.010549 0.0013965 0.98681 0.99162 3.0126e-006 1.205e-005 0.16592 0.89124 0.89857 0.0014025 0.97963 0.45037 0.0018893 0.42265 2.1047 2.1037 16.0209 144.9081 0.0001907 -85.6079 0.60894
8.713 0.98815 5.4629e-005 3.8183 0.011915 0.0001132 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6018 0.59048 0.18041 0.020615 18.2211 0.12767 0.00016722 0.7625 0.0095409 0.010549 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.16592 0.89153 0.89869 0.0014024 0.97975 0.45056 0.0018892 0.42266 2.1054 2.1044 16.0209 144.9081 0.00019051 -85.6083 0.60994
8.714 0.98815 5.4629e-005 3.8183 0.011915 0.00011322 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6018 0.59053 0.18043 0.020616 18.2243 0.12768 0.00016723 0.76249 0.0095413 0.01055 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.16592 0.89182 0.89882 0.0014024 0.97986 0.45075 0.0018891 0.42268 2.1061 2.1052 16.0209 144.9081 0.00019032 -85.6087 0.61094
8.715 0.98815 5.4629e-005 3.8183 0.011915 0.00011323 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6019 0.59057 0.18044 0.020617 18.2274 0.12768 0.00016724 0.76248 0.0095416 0.01055 0.0013962 0.98682 0.99162 3.0119e-006 1.2048e-005 0.16593 0.8921 0.89894 0.0014023 0.97997 0.45094 0.0018891 0.42269 2.1069 2.1059 16.0209 144.9081 0.00019013 -85.6091 0.61194
8.716 0.98815 5.4629e-005 3.8183 0.011915 0.00011324 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.602 0.59062 0.18045 0.020618 18.2306 0.12769 0.00016725 0.76248 0.009542 0.01055 0.0013961 0.98682 0.99162 3.0117e-006 1.2047e-005 0.16593 0.89239 0.89906 0.0014023 0.98008 0.45114 0.001889 0.42271 2.1076 2.1066 16.0208 144.9081 0.00018994 -85.6095 0.61294
8.717 0.98815 5.4629e-005 3.8183 0.011915 0.00011325 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6021 0.59066 0.18047 0.020619 18.2338 0.1277 0.00016726 0.76247 0.0095423 0.010551 0.001396 0.98682 0.99162 3.0115e-006 1.2046e-005 0.16593 0.89267 0.89919 0.0014022 0.98019 0.45133 0.001889 0.42272 2.1083 2.1073 16.0208 144.9082 0.00018975 -85.6099 0.61394
8.718 0.98815 5.4628e-005 3.8183 0.011915 0.00011327 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6022 0.59071 0.18048 0.02062 18.237 0.1277 0.00016727 0.76246 0.0095427 0.010551 0.0013959 0.98682 0.99162 3.0113e-006 1.2045e-005 0.16593 0.89296 0.89931 0.0014022 0.9803 0.45152 0.0018889 0.42274 2.109 2.108 16.0208 144.9082 0.00018956 -85.6103 0.61494
8.719 0.98815 5.4628e-005 3.8183 0.011915 0.00011328 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6023 0.59075 0.18049 0.020621 18.2402 0.12771 0.00016728 0.76246 0.009543 0.010551 0.0013959 0.98682 0.99162 3.0111e-006 1.2044e-005 0.16594 0.89324 0.89943 0.0014021 0.98041 0.45171 0.0018888 0.42275 2.1097 2.1087 16.0208 144.9082 0.00018937 -85.6107 0.61594
8.72 0.98815 5.4628e-005 3.8183 0.011915 0.00011329 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6023 0.59079 0.18051 0.020623 18.2433 0.12772 0.00016729 0.76245 0.0095434 0.010552 0.0013958 0.98682 0.99163 3.0109e-006 1.2043e-005 0.16594 0.89352 0.89955 0.0014021 0.98052 0.4519 0.0018888 0.42277 2.1104 2.1094 16.0208 144.9082 0.00018918 -85.611 0.61694
8.721 0.98815 5.4628e-005 3.8183 0.011915 0.0001133 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6024 0.59084 0.18052 0.020624 18.2465 0.12772 0.0001673 0.76245 0.0095437 0.010552 0.0013957 0.98682 0.99163 3.0107e-006 1.2043e-005 0.16594 0.8938 0.89968 0.001402 0.98063 0.45209 0.0018887 0.42278 2.1111 2.1101 16.0207 144.9082 0.000189 -85.6114 0.61794
8.722 0.98815 5.4628e-005 3.8183 0.011915 0.00011332 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6025 0.59088 0.18053 0.020625 18.2497 0.12773 0.00016731 0.76244 0.0095441 0.010553 0.0013956 0.98682 0.99163 3.0105e-006 1.2042e-005 0.16595 0.89408 0.8998 0.001402 0.98074 0.45228 0.0018886 0.4228 2.1118 2.1108 16.0207 144.9083 0.00018881 -85.6118 0.61894
8.723 0.98815 5.4628e-005 3.8183 0.011915 0.00011333 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6026 0.59093 0.18054 0.020626 18.2529 0.12773 0.00016731 0.76243 0.0095445 0.010553 0.0013955 0.98682 0.99163 3.0103e-006 1.2041e-005 0.16595 0.89436 0.89992 0.001402 0.98084 0.45247 0.0018886 0.42281 2.1125 2.1116 16.0207 144.9083 0.00018863 -85.6122 0.61994
8.724 0.98815 5.4628e-005 3.8183 0.011915 0.00011334 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6027 0.59097 0.18056 0.020627 18.2561 0.12774 0.00016732 0.76243 0.0095448 0.010553 0.0013954 0.98683 0.99163 3.0101e-006 1.204e-005 0.16595 0.89464 0.90004 0.0014019 0.98095 0.45266 0.0018885 0.42283 2.1132 2.1123 16.0207 144.9083 0.00018844 -85.6126 0.62094
8.725 0.98815 5.4628e-005 3.8183 0.011915 0.00011336 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6028 0.59102 0.18057 0.020628 18.2592 0.12775 0.00016733 0.76242 0.0095452 0.010554 0.0013953 0.98683 0.99163 3.0099e-006 1.2039e-005 0.16595 0.89492 0.90016 0.0014019 0.98105 0.45285 0.0018885 0.42284 2.1139 2.113 16.0207 144.9083 0.00018826 -85.6129 0.62194
8.726 0.98815 5.4628e-005 3.8183 0.011915 0.00011337 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6029 0.59106 0.18058 0.020629 18.2624 0.12775 0.00016734 0.76242 0.0095455 0.010554 0.0013953 0.98683 0.99163 3.0097e-006 1.2039e-005 0.16596 0.8952 0.90028 0.0014018 0.98116 0.45304 0.0018884 0.42286 2.1146 2.1137 16.0206 144.9083 0.00018807 -85.6133 0.62294
8.727 0.98815 5.4628e-005 3.8183 0.011915 0.00011338 0.0011756 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6029 0.59111 0.1806 0.02063 18.2656 0.12776 0.00016735 0.76241 0.0095459 0.010554 0.0013952 0.98683 0.99163 3.0095e-006 1.2038e-005 0.16596 0.89547 0.90039 0.0014018 0.98126 0.45323 0.0018883 0.42287 2.1153 2.1143 16.0206 144.9084 0.00018789 -85.6137 0.62394
8.728 0.98815 5.4628e-005 3.8183 0.011915 0.00011339 0.0011757 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.603 0.59115 0.18061 0.020631 18.2688 0.12776 0.00016736 0.7624 0.0095462 0.010555 0.0013951 0.98683 0.99163 3.0093e-006 1.2037e-005 0.16596 0.89575 0.90051 0.0014017 0.98137 0.45342 0.0018883 0.42289 2.116 2.115 16.0206 144.9084 0.00018771 -85.614 0.62494
8.729 0.98815 5.4628e-005 3.8183 0.011915 0.00011341 0.0011757 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6031 0.59119 0.18062 0.020632 18.272 0.12777 0.00016737 0.7624 0.0095466 0.010555 0.001395 0.98683 0.99163 3.0091e-006 1.2036e-005 0.16596 0.89602 0.90063 0.0014017 0.98147 0.45361 0.0018882 0.4229 2.1167 2.1157 16.0206 144.9084 0.00018753 -85.6144 0.62594
8.73 0.98815 5.4627e-005 3.8183 0.011915 0.00011342 0.0011757 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6032 0.59124 0.18064 0.020633 18.2752 0.12778 0.00016738 0.76239 0.0095469 0.010555 0.0013949 0.98683 0.99163 3.0089e-006 1.2035e-005 0.16597 0.8963 0.90075 0.0014016 0.98157 0.4538 0.0018882 0.42292 2.1174 2.1164 16.0205 144.9084 0.00018735 -85.6147 0.62694
8.731 0.98815 5.4627e-005 3.8183 0.011915 0.00011343 0.0011757 0.23365 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6033 0.59128 0.18065 0.020634 18.2784 0.12778 0.00016739 0.76238 0.0095473 0.010556 0.0013948 0.98683 0.99163 3.0087e-006 1.2035e-005 0.16597 0.89657 0.90086 0.0014016 0.98167 0.45399 0.0018881 0.42293 2.1181 2.1171 16.0205 144.9084 0.00018717 -85.6151 0.62794
8.732 0.98815 5.4627e-005 3.8183 0.011915 0.00011345 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6034 0.59133 0.18066 0.020635 18.2815 0.12779 0.0001674 0.76238 0.0095476 0.010556 0.0013947 0.98683 0.99163 3.0085e-006 1.2034e-005 0.16597 0.89684 0.90098 0.0014015 0.98177 0.45418 0.0018881 0.42295 2.1188 2.1178 16.0205 144.9085 0.00018699 -85.6155 0.62894
8.733 0.98815 5.4627e-005 3.8183 0.011915 0.00011346 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6034 0.59137 0.18068 0.020636 18.2847 0.1278 0.00016741 0.76237 0.009548 0.010557 0.0013947 0.98684 0.99163 3.0083e-006 1.2033e-005 0.16598 0.89711 0.9011 0.0014015 0.98187 0.45437 0.001888 0.42296 2.1194 2.1185 16.0205 144.9085 0.00018681 -85.6158 0.62994
8.734 0.98815 5.4627e-005 3.8183 0.011915 0.00011347 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6035 0.59142 0.18069 0.020637 18.2879 0.1278 0.00016742 0.76237 0.0095483 0.010557 0.0013946 0.98684 0.99164 3.0081e-006 1.2032e-005 0.16598 0.89738 0.90121 0.0014015 0.98197 0.45456 0.0018879 0.42298 2.1201 2.1192 16.0205 144.9085 0.00018663 -85.6162 0.63094
8.735 0.98815 5.4627e-005 3.8183 0.011915 0.00011348 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6036 0.59146 0.1807 0.020638 18.2911 0.12781 0.00016743 0.76236 0.0095487 0.010557 0.0013945 0.98684 0.99164 3.008e-006 1.2032e-005 0.16598 0.89765 0.90133 0.0014014 0.98207 0.45475 0.0018879 0.42299 2.1208 2.1199 16.0204 144.9085 0.00018646 -85.6165 0.63194
8.736 0.98815 5.4627e-005 3.8183 0.011915 0.0001135 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6037 0.59151 0.18072 0.020639 18.2943 0.12781 0.00016744 0.76235 0.009549 0.010558 0.0013944 0.98684 0.99164 3.0078e-006 1.2031e-005 0.16598 0.89792 0.90144 0.0014014 0.98217 0.45494 0.0018878 0.42301 2.1215 2.1205 16.0204 144.9085 0.00018628 -85.6168 0.63294
8.737 0.98815 5.4627e-005 3.8183 0.011915 0.00011351 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6038 0.59155 0.18073 0.02064 18.2975 0.12782 0.00016745 0.76235 0.0095494 0.010558 0.0013943 0.98684 0.99164 3.0076e-006 1.203e-005 0.16599 0.89819 0.90156 0.0014013 0.98227 0.45513 0.0018878 0.42302 2.1222 2.1212 16.0204 144.9086 0.00018611 -85.6172 0.63394
8.738 0.98815 5.4627e-005 3.8183 0.011915 0.00011352 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6039 0.59159 0.18074 0.020641 18.3007 0.12783 0.00016746 0.76234 0.0095497 0.010558 0.0013943 0.98684 0.99164 3.0074e-006 1.203e-005 0.16599 0.89845 0.90167 0.0014013 0.98236 0.45532 0.0018877 0.42304 2.1228 2.1219 16.0204 144.9086 0.00018593 -85.6175 0.63494
8.739 0.98815 5.4627e-005 3.8183 0.011915 0.00011353 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6039 0.59164 0.18075 0.020642 18.3038 0.12783 0.00016747 0.76234 0.0095501 0.010559 0.0013942 0.98684 0.99164 3.0072e-006 1.2029e-005 0.16599 0.89872 0.90178 0.0014013 0.98246 0.45551 0.0018877 0.42305 2.1235 2.1226 16.0204 144.9086 0.00018576 -85.6179 0.63594
8.74 0.98815 5.4627e-005 3.8183 0.011915 0.00011355 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.604 0.59168 0.18077 0.020643 18.307 0.12784 0.00016747 0.76233 0.0095504 0.010559 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.16599 0.89898 0.9019 0.0014012 0.98255 0.4557 0.0018876 0.42307 2.1242 2.1233 16.0203 144.9086 0.00018558 -85.6182 0.63694
8.741 0.98815 5.4627e-005 3.8183 0.011915 0.00011356 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6041 0.59173 0.18078 0.020644 18.3102 0.12784 0.00016748 0.76232 0.0095508 0.01056 0.001394 0.98684 0.99164 3.0069e-006 1.2027e-005 0.166 0.89925 0.90201 0.0014012 0.98265 0.45589 0.0018876 0.42308 2.1248 2.1239 16.0203 144.9086 0.00018541 -85.6185 0.63794
8.742 0.98815 5.4626e-005 3.8183 0.011915 0.00011357 0.0011757 0.23364 0.00065931 0.2343 0.21621 0 0.032262 0.0389 0 1.6042 0.59177 0.18079 0.020645 18.3134 0.12785 0.00016749 0.76232 0.0095511 0.01056 0.001394 0.98684 0.99164 3.0067e-006 1.2027e-005 0.166 0.89951 0.90212 0.0014011 0.98274 0.45608 0.0018875 0.4231 2.1255 2.1246 16.0203 144.9087 0.00018524 -85.6189 0.63894
8.743 0.98815 5.4626e-005 3.8183 0.011915 0.00011359 0.0011757 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6043 0.59182 0.18081 0.020646 18.3166 0.12786 0.0001675 0.76231 0.0095515 0.01056 0.0013939 0.98685 0.99164 3.0065e-006 1.2026e-005 0.166 0.89977 0.90223 0.0014011 0.98284 0.45627 0.0018875 0.42311 2.1262 2.1253 16.0203 144.9087 0.00018507 -85.6192 0.63994
8.744 0.98815 5.4626e-005 3.8183 0.011915 0.0001136 0.0011757 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6044 0.59186 0.18082 0.020647 18.3198 0.12786 0.00016751 0.7623 0.0095518 0.010561 0.0013938 0.98685 0.99164 3.0064e-006 1.2025e-005 0.166 0.90004 0.90234 0.001401 0.98293 0.45646 0.0018874 0.42313 2.1268 2.1259 16.0202 144.9087 0.00018489 -85.6195 0.64094
8.745 0.98815 5.4626e-005 3.8183 0.011915 0.00011361 0.0011757 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6044 0.5919 0.18083 0.020648 18.323 0.12787 0.00016752 0.7623 0.0095522 0.010561 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.16601 0.9003 0.90246 0.001401 0.98302 0.45665 0.0018874 0.42314 2.1275 2.1266 16.0202 144.9087 0.00018472 -85.6198 0.64194
8.746 0.98815 5.4626e-005 3.8183 0.011915 0.00011362 0.0011757 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6045 0.59195 0.18085 0.020649 18.3262 0.12788 0.00016753 0.76229 0.0095525 0.010561 0.0013936 0.98685 0.99164 3.006e-006 1.2024e-005 0.16601 0.90056 0.90257 0.001401 0.98311 0.45684 0.0018873 0.42316 2.1282 2.1273 16.0202 144.9087 0.00018455 -85.6202 0.64294
8.747 0.98815 5.4626e-005 3.8183 0.011915 0.00011364 0.0011757 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6046 0.59199 0.18086 0.02065 18.3294 0.12788 0.00016754 0.76229 0.0095529 0.010562 0.0013935 0.98685 0.99164 3.0058e-006 1.2023e-005 0.16601 0.90082 0.90268 0.0014009 0.9832 0.45703 0.0018873 0.42317 2.1288 2.1279 16.0202 144.9088 0.00018439 -85.6205 0.64394
8.748 0.98815 5.4626e-005 3.8183 0.011915 0.00011365 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6047 0.59204 0.18087 0.020651 18.3325 0.12789 0.00016755 0.76228 0.0095532 0.010562 0.0013935 0.98685 0.99164 3.0057e-006 1.2023e-005 0.16602 0.90107 0.90279 0.0014009 0.9833 0.45722 0.0018872 0.42319 2.1295 2.1286 16.0202 144.9088 0.00018422 -85.6208 0.64494
8.749 0.98815 5.4626e-005 3.8183 0.011915 0.00011366 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6048 0.59208 0.18089 0.020653 18.3357 0.12789 0.00016756 0.76227 0.0095536 0.010563 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.16602 0.90133 0.90289 0.0014009 0.98339 0.45741 0.0018872 0.4232 2.1301 2.1292 16.0201 144.9088 0.00018405 -85.6211 0.64594
8.75 0.98815 5.4626e-005 3.8183 0.011915 0.00011368 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6049 0.59213 0.1809 0.020654 18.3389 0.1279 0.00016757 0.76227 0.0095539 0.010563 0.0013933 0.98685 0.99165 3.0053e-006 1.2021e-005 0.16602 0.90159 0.903 0.0014008 0.98347 0.4576 0.0018871 0.42322 2.1308 2.1299 16.0201 144.9088 0.00018388 -85.6214 0.64694
8.751 0.98815 5.4626e-005 3.8183 0.011915 0.00011369 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6049 0.59217 0.18091 0.020655 18.3421 0.12791 0.00016758 0.76226 0.0095543 0.010563 0.0013933 0.98685 0.99165 3.0052e-006 1.2021e-005 0.16602 0.90184 0.90311 0.0014008 0.98356 0.45778 0.0018871 0.42323 2.1315 2.1306 16.0201 144.9089 0.00018372 -85.6217 0.64794
8.752 0.98815 5.4626e-005 3.8183 0.011915 0.0001137 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.605 0.59222 0.18092 0.020656 18.3453 0.12791 0.00016759 0.76226 0.0095546 0.010564 0.0013932 0.98685 0.99165 3.005e-006 1.202e-005 0.16603 0.9021 0.90322 0.0014007 0.98365 0.45797 0.001887 0.42325 2.1321 2.1312 16.0201 144.9089 0.00018355 -85.622 0.64894
8.753 0.98815 5.4625e-005 3.8183 0.011915 0.00011371 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6051 0.59226 0.18094 0.020657 18.3485 0.12792 0.0001676 0.76225 0.009555 0.010564 0.0013931 0.98686 0.99165 3.0049e-006 1.2019e-005 0.16603 0.90235 0.90333 0.0014007 0.98374 0.45816 0.001887 0.42326 2.1328 2.1319 16.02 144.9089 0.00018338 -85.6223 0.64994
8.754 0.98815 5.4625e-005 3.8183 0.011914 0.00011373 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6052 0.5923 0.18095 0.020658 18.3517 0.12792 0.00016761 0.76224 0.0095553 0.010564 0.0013931 0.98686 0.99165 3.0047e-006 1.2019e-005 0.16603 0.90261 0.90343 0.0014007 0.98383 0.45835 0.0018869 0.42328 2.1334 2.1325 16.02 144.9089 0.00018322 -85.6226 0.65094
8.755 0.98815 5.4625e-005 3.8183 0.011914 0.00011374 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6053 0.59235 0.18096 0.020659 18.3549 0.12793 0.00016762 0.76224 0.0095557 0.010565 0.001393 0.98686 0.99165 3.0045e-006 1.2018e-005 0.16603 0.90286 0.90354 0.0014006 0.98391 0.45854 0.0018869 0.42329 2.1341 2.1332 16.02 144.9089 0.00018306 -85.6229 0.65194
8.756 0.98815 5.4625e-005 3.8183 0.011914 0.00011375 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6054 0.59239 0.18098 0.02066 18.3581 0.12794 0.00016762 0.76223 0.009556 0.010565 0.0013929 0.98686 0.99165 3.0044e-006 1.2017e-005 0.16604 0.90311 0.90365 0.0014006 0.984 0.45873 0.0018868 0.42331 2.1347 2.1338 16.02 144.909 0.00018289 -85.6232 0.65294
8.757 0.98815 5.4625e-005 3.8183 0.011914 0.00011377 0.0011758 0.23364 0.00065931 0.2343 0.2162 0 0.032262 0.0389 0 1.6055 0.59244 0.18099 0.020661 18.3613 0.12794 0.00016763 0.76222 0.0095564 0.010566 0.0013928 0.98686 0.99165 3.0042e-006 1.2017e-005 0.16604 0.90336 0.90375 0.0014006 0.98409 0.45892 0.0018868 0.42332 2.1354 2.1345 16.02 144.909 0.00018273 -85.6235 0.65394
8.758 0.98815 5.4625e-005 3.8183 0.011914 0.00011378 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6055 0.59248 0.181 0.020662 18.3645 0.12795 0.00016764 0.76222 0.0095567 0.010566 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.16604 0.90361 0.90386 0.0014005 0.98417 0.4591 0.0018867 0.42334 2.136 2.1351 16.0199 144.909 0.00018257 -85.6238 0.65494
8.759 0.98815 5.4625e-005 3.8183 0.011914 0.00011379 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6056 0.59253 0.18102 0.020663 18.3677 0.12795 0.00016765 0.76221 0.0095571 0.010566 0.0013927 0.98686 0.99165 3.0039e-006 1.2016e-005 0.16605 0.90386 0.90396 0.0014005 0.98425 0.45929 0.0018867 0.42335 2.1366 2.1358 16.0199 144.909 0.00018241 -85.6241 0.65594
8.76 0.98815 5.4625e-005 3.8183 0.011914 0.0001138 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6057 0.59257 0.18103 0.020664 18.3709 0.12796 0.00016766 0.76221 0.0095574 0.010567 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.16605 0.90411 0.90407 0.0014004 0.98434 0.45948 0.0018866 0.42337 2.1373 2.1364 16.0199 144.909 0.00018224 -85.6244 0.65694
8.761 0.98815 5.4625e-005 3.8183 0.011914 0.00011382 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6058 0.59262 0.18104 0.020665 18.3741 0.12797 0.00016767 0.7622 0.0095578 0.010567 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.16605 0.90436 0.90417 0.0014004 0.98442 0.45967 0.0018866 0.42338 2.1379 2.137 16.0199 144.9091 0.00018208 -85.6247 0.65794
8.762 0.98815 5.4625e-005 3.8183 0.011914 0.00011383 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6059 0.59266 0.18106 0.020666 18.3772 0.12797 0.00016768 0.76219 0.0095581 0.010567 0.0013925 0.98686 0.99165 3.0035e-006 1.2014e-005 0.16605 0.90461 0.90428 0.0014004 0.9845 0.45986 0.0018865 0.4234 2.1386 2.1377 16.0198 144.9091 0.00018192 -85.625 0.65894
8.763 0.98815 5.4625e-005 3.8183 0.011914 0.00011384 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.606 0.5927 0.18107 0.020667 18.3804 0.12798 0.00016769 0.76219 0.0095585 0.010568 0.0013925 0.98686 0.99165 3.0033e-006 1.2013e-005 0.16606 0.90485 0.90438 0.0014003 0.98459 0.46005 0.0018865 0.42341 2.1392 2.1383 16.0198 144.9091 0.00018176 -85.6253 0.65994
8.764 0.98815 5.4625e-005 3.8183 0.011914 0.00011385 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.606 0.59275 0.18108 0.020668 18.3836 0.12799 0.0001677 0.76218 0.0095588 0.010568 0.0013924 0.98686 0.99165 3.0032e-006 1.2013e-005 0.16606 0.9051 0.90448 0.0014003 0.98467 0.46023 0.0018864 0.42343 2.1398 2.139 16.0198 144.9091 0.00018161 -85.6255 0.66094
8.765 0.98815 5.4624e-005 3.8183 0.011914 0.00011387 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6061 0.59279 0.1811 0.020669 18.3868 0.12799 0.00016771 0.76218 0.0095592 0.010568 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.16606 0.90535 0.90459 0.0014003 0.98475 0.46042 0.0018864 0.42344 2.1405 2.1396 16.0198 144.9091 0.00018145 -85.6258 0.66194
8.766 0.98815 5.4624e-005 3.8183 0.011914 0.00011388 0.0011758 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6062 0.59284 0.18111 0.02067 18.39 0.128 0.00016772 0.76217 0.0095595 0.010569 0.0013922 0.98687 0.99165 3.0029e-006 1.2011e-005 0.16606 0.90559 0.90469 0.0014002 0.98483 0.46061 0.0018863 0.42346 2.1411 2.1402 16.0197 144.9092 0.00018129 -85.6261 0.66294
8.767 0.98815 5.4624e-005 3.8183 0.011914 0.00011389 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6063 0.59288 0.18112 0.020671 18.3932 0.128 0.00016773 0.76216 0.0095599 0.010569 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.16607 0.90583 0.90479 0.0014002 0.98491 0.4608 0.0018863 0.42347 2.1417 2.1409 16.0197 144.9092 0.00018113 -85.6264 0.66394
8.768 0.98815 5.4624e-005 3.8183 0.011914 0.00011391 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6064 0.59293 0.18113 0.020672 18.3964 0.12801 0.00016774 0.76216 0.0095602 0.01057 0.0013921 0.98687 0.99166 3.0026e-006 1.201e-005 0.16607 0.90608 0.90489 0.0014002 0.98499 0.46098 0.0018863 0.42348 2.1423 2.1415 16.0197 144.9092 0.00018098 -85.6266 0.66494
8.769 0.98815 5.4624e-005 3.8183 0.011914 0.00011392 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6065 0.59297 0.18115 0.020673 18.3996 0.12802 0.00016775 0.76215 0.0095606 0.01057 0.001392 0.98687 0.99166 3.0024e-006 1.201e-005 0.16607 0.90632 0.90499 0.0014001 0.98507 0.46117 0.0018862 0.4235 2.143 2.1421 16.0197 144.9092 0.00018082 -85.6269 0.66594
8.77 0.98815 5.4624e-005 3.8183 0.011914 0.00011393 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6065 0.59302 0.18116 0.020674 18.4028 0.12802 0.00016776 0.76215 0.0095609 0.01057 0.001392 0.98687 0.99166 3.0023e-006 1.2009e-005 0.16607 0.90656 0.9051 0.0014001 0.98515 0.46136 0.0018862 0.42351 2.1436 2.1427 16.0197 144.9092 0.00018067 -85.6272 0.66694
8.771 0.98815 5.4624e-005 3.8183 0.011914 0.00011394 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6066 0.59306 0.18117 0.020675 18.406 0.12803 0.00016777 0.76214 0.0095613 0.010571 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.16608 0.9068 0.9052 0.0014001 0.98523 0.46155 0.0018861 0.42353 2.1442 2.1434 16.0196 144.9093 0.00018051 -85.6275 0.66794
8.772 0.98815 5.4624e-005 3.8183 0.011914 0.00011396 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6067 0.5931 0.18119 0.020676 18.4092 0.12803 0.00016777 0.76213 0.0095616 0.010571 0.0013919 0.98687 0.99166 3.002e-006 1.2008e-005 0.16608 0.90704 0.9053 0.0014 0.9853 0.46174 0.0018861 0.42354 2.1448 2.144 16.0196 144.9093 0.00018036 -85.6277 0.66894
8.773 0.98815 5.4624e-005 3.8183 0.011914 0.00011397 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6068 0.59315 0.1812 0.020677 18.4124 0.12804 0.00016778 0.76213 0.009562 0.010571 0.0013918 0.98687 0.99166 3.0019e-006 1.2007e-005 0.16608 0.90728 0.9054 0.0014 0.98538 0.46192 0.001886 0.42356 2.1455 2.1446 16.0196 144.9093 0.00018021 -85.628 0.66994
8.774 0.98815 5.4624e-005 3.8183 0.011914 0.00011398 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6069 0.59319 0.18121 0.020678 18.4156 0.12805 0.00016779 0.76212 0.0095623 0.010572 0.0013918 0.98687 0.99166 3.0017e-006 1.2007e-005 0.16609 0.90752 0.9055 0.0014 0.98546 0.46211 0.001886 0.42357 2.1461 2.1452 16.0196 144.9093 0.00018005 -85.6282 0.67094
8.775 0.98815 5.4624e-005 3.8183 0.011914 0.000114 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.607 0.59324 0.18123 0.020679 18.4188 0.12805 0.0001678 0.76211 0.0095627 0.010572 0.0013917 0.98687 0.99166 3.0016e-006 1.2006e-005 0.16609 0.90775 0.90559 0.0013999 0.98553 0.4623 0.001886 0.42359 2.1467 2.1459 16.0195 144.9093 0.0001799 -85.6285 0.67194
8.776 0.98815 5.4624e-005 3.8183 0.011914 0.00011401 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.607 0.59328 0.18124 0.02068 18.422 0.12806 0.00016781 0.76211 0.009563 0.010573 0.0013916 0.98687 0.99166 3.0014e-006 1.2006e-005 0.16609 0.90799 0.90569 0.0013999 0.98561 0.46248 0.0018859 0.4236 2.1473 2.1465 16.0195 144.9094 0.00017975 -85.6288 0.67294
8.777 0.98815 5.4623e-005 3.8183 0.011914 0.00011402 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6071 0.59333 0.18125 0.020681 18.4252 0.12807 0.00016782 0.7621 0.0095634 0.010573 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.16609 0.90823 0.90579 0.0013999 0.98568 0.46267 0.0018859 0.42362 2.1479 2.1471 16.0195 144.9094 0.0001796 -85.629 0.67394
8.778 0.98815 5.4623e-005 3.8183 0.011914 0.00011403 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6072 0.59337 0.18127 0.020682 18.4284 0.12807 0.00016783 0.7621 0.0095637 0.010573 0.0013915 0.98688 0.99166 3.0012e-006 1.2005e-005 0.1661 0.90846 0.90589 0.0013999 0.98576 0.46286 0.0018858 0.42363 2.1485 2.1477 16.0195 144.9094 0.00017945 -85.6293 0.67494
8.779 0.98815 5.4623e-005 3.8183 0.011914 0.00011405 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6073 0.59341 0.18128 0.020683 18.4316 0.12808 0.00016784 0.76209 0.0095641 0.010574 0.0013915 0.98688 0.99166 3.001e-006 1.2004e-005 0.1661 0.9087 0.90599 0.0013998 0.98583 0.46305 0.0018858 0.42365 2.1492 2.1483 16.0194 144.9094 0.0001793 -85.6295 0.67594
8.78 0.98815 5.4623e-005 3.8183 0.011914 0.00011406 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6074 0.59346 0.18129 0.020685 18.4348 0.12808 0.00016785 0.76208 0.0095644 0.010574 0.0013914 0.98688 0.99166 3.0009e-006 1.2004e-005 0.1661 0.90893 0.90608 0.0013998 0.98591 0.46323 0.0018858 0.42366 2.1498 2.1489 16.0194 144.9094 0.00017915 -85.6298 0.67694
8.781 0.98815 5.4623e-005 3.8183 0.011914 0.00011407 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6075 0.5935 0.1813 0.020686 18.438 0.12809 0.00016786 0.76208 0.0095648 0.010574 0.0013914 0.98688 0.99166 3.0008e-006 1.2003e-005 0.1661 0.90916 0.90618 0.0013998 0.98598 0.46342 0.0018857 0.42368 2.1504 2.1495 16.0194 144.9095 0.000179 -85.63 0.67794
8.782 0.98815 5.4623e-005 3.8183 0.011914 0.00011408 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6075 0.59355 0.18132 0.020687 18.4412 0.1281 0.00016787 0.76207 0.0095651 0.010575 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.16611 0.9094 0.90628 0.0013997 0.98605 0.46361 0.0018857 0.42369 2.151 2.1502 16.0194 144.9095 0.00017885 -85.6303 0.67894
8.783 0.98815 5.4623e-005 3.8183 0.011914 0.0001141 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6076 0.59359 0.18133 0.020688 18.4444 0.1281 0.00016788 0.76207 0.0095655 0.010575 0.0013912 0.98688 0.99166 3.0005e-006 1.2002e-005 0.16611 0.90963 0.90637 0.0013997 0.98613 0.46379 0.0018856 0.42371 2.1516 2.1508 16.0193 144.9095 0.0001787 -85.6305 0.67994
8.784 0.98815 5.4623e-005 3.8183 0.011914 0.00011411 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6077 0.59364 0.18134 0.020689 18.4476 0.12811 0.00016789 0.76206 0.0095658 0.010575 0.0013912 0.98688 0.99166 3.0004e-006 1.2001e-005 0.16611 0.90986 0.90647 0.0013997 0.9862 0.46398 0.0018856 0.42372 2.1522 2.1514 16.0193 144.9095 0.00017856 -85.6308 0.68094
8.785 0.98815 5.4623e-005 3.8183 0.011914 0.00011412 0.0011759 0.23364 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6078 0.59368 0.18136 0.02069 18.4508 0.12811 0.0001679 0.76205 0.0095662 0.010576 0.0013911 0.98688 0.99166 3.0003e-006 1.2001e-005 0.16611 0.91009 0.90657 0.0013996 0.98627 0.46417 0.0018856 0.42374 2.1528 2.152 16.0193 144.9095 0.00017841 -85.631 0.68194
8.786 0.98815 5.4623e-005 3.8183 0.011914 0.00011414 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6079 0.59373 0.18137 0.020691 18.454 0.12812 0.00016791 0.76205 0.0095665 0.010576 0.0013911 0.98688 0.99166 3.0001e-006 1.2e-005 0.16612 0.91032 0.90666 0.0013996 0.98634 0.46435 0.0018855 0.42375 2.1534 2.1526 16.0193 144.9096 0.00017826 -85.6312 0.68294
8.787 0.98815 5.4623e-005 3.8183 0.011914 0.00011415 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.608 0.59377 0.18138 0.020692 18.4572 0.12813 0.00016792 0.76204 0.0095669 0.010577 0.001391 0.98688 0.99166 3e-006 1.2e-005 0.16612 0.91055 0.90676 0.0013996 0.98641 0.46454 0.0018855 0.42377 2.154 2.1532 16.0192 144.9096 0.00017812 -85.6315 0.68394
8.788 0.98815 5.4623e-005 3.8183 0.011914 0.00011416 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6081 0.59381 0.1814 0.020693 18.4604 0.12813 0.00016792 0.76204 0.0095672 0.010577 0.0013909 0.98688 0.99167 2.9999e-006 1.1999e-005 0.16612 0.91078 0.90685 0.0013996 0.98648 0.46473 0.0018854 0.42378 2.1546 2.1538 16.0192 144.9096 0.00017797 -85.6317 0.68494
8.789 0.98815 5.4622e-005 3.8183 0.011914 0.00011417 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6081 0.59386 0.18141 0.020694 18.4636 0.12814 0.00016793 0.76203 0.0095676 0.010577 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.16613 0.911 0.90694 0.0013995 0.98655 0.46491 0.0018854 0.4238 2.1552 2.1544 16.0192 144.9096 0.00017783 -85.632 0.68594
8.79 0.98815 5.4622e-005 3.8183 0.011914 0.00011419 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6082 0.5939 0.18142 0.020695 18.4668 0.12814 0.00016794 0.76202 0.0095679 0.010578 0.0013908 0.98688 0.99167 2.9996e-006 1.1998e-005 0.16613 0.91123 0.90704 0.0013995 0.98662 0.4651 0.0018854 0.42381 2.1558 2.155 16.0192 144.9096 0.00017768 -85.6322 0.68694
8.791 0.98815 5.4622e-005 3.8183 0.011914 0.0001142 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6083 0.59395 0.18144 0.020696 18.47 0.12815 0.00016795 0.76202 0.0095682 0.010578 0.0013908 0.98689 0.99167 2.9995e-006 1.1998e-005 0.16613 0.91146 0.90713 0.0013995 0.98669 0.46529 0.0018853 0.42383 2.1564 2.1556 16.0191 144.9097 0.00017754 -85.6324 0.68794
8.792 0.98815 5.4622e-005 3.8183 0.011914 0.00011421 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6084 0.59399 0.18145 0.020697 18.4732 0.12816 0.00016796 0.76201 0.0095686 0.010578 0.0013907 0.98689 0.99167 2.9994e-006 1.1997e-005 0.16613 0.91168 0.90722 0.0013994 0.98675 0.46547 0.0018853 0.42384 2.157 2.1562 16.0191 144.9097 0.0001774 -85.6326 0.68894
8.793 0.98815 5.4622e-005 3.8183 0.011914 0.00011423 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6085 0.59404 0.18146 0.020698 18.4765 0.12816 0.00016797 0.762 0.0095689 0.010579 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.16614 0.91191 0.90732 0.0013994 0.98682 0.46566 0.0018853 0.42385 2.1576 2.1568 16.0191 144.9097 0.00017725 -85.6329 0.68994
8.794 0.98815 5.4622e-005 3.8183 0.011914 0.00011424 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6086 0.59408 0.18147 0.020699 18.4797 0.12817 0.00016798 0.762 0.0095693 0.010579 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.16614 0.91213 0.90741 0.0013994 0.98689 0.46584 0.0018852 0.42387 2.1582 2.1574 16.0191 144.9097 0.00017711 -85.6331 0.69094
8.795 0.98815 5.4622e-005 3.8183 0.011914 0.00011425 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6086 0.59412 0.18149 0.0207 18.4829 0.12818 0.00016799 0.76199 0.0095696 0.01058 0.0013906 0.98689 0.99167 2.999e-006 1.1996e-005 0.16614 0.91235 0.9075 0.0013994 0.98696 0.46603 0.0018852 0.42388 2.1587 2.1579 16.019 144.9097 0.00017697 -85.6333 0.69194
8.796 0.98815 5.4622e-005 3.8183 0.011914 0.00011426 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032262 0.0389 0 1.6087 0.59417 0.1815 0.020701 18.4861 0.12818 0.000168 0.76199 0.00957 0.01058 0.0013905 0.98689 0.99167 2.9989e-006 1.1995e-005 0.16614 0.91257 0.90759 0.0013993 0.98702 0.46622 0.0018852 0.4239 2.1593 2.1585 16.019 144.9098 0.00017683 -85.6335 0.69294
8.797 0.98815 5.4622e-005 3.8183 0.011914 0.00011428 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032263 0.0389 0 1.6088 0.59421 0.18151 0.020702 18.4893 0.12819 0.00016801 0.76198 0.0095703 0.01058 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.16615 0.9128 0.90768 0.0013993 0.98709 0.4664 0.0018851 0.42391 2.1599 2.1591 16.019 144.9098 0.00017669 -85.6338 0.69394
8.798 0.98815 5.4622e-005 3.8183 0.011914 0.00011429 0.001176 0.23363 0.00065931 0.23429 0.2162 0 0.032263 0.0389 0 1.6089 0.59426 0.18153 0.020703 18.4925 0.12819 0.00016802 0.76197 0.0095707 0.010581 0.0013904 0.98689 0.99167 2.9987e-006 1.1995e-005 0.16615 0.91302 0.90777 0.0013993 0.98715 0.46659 0.0018851 0.42393 2.1605 2.1597 16.019 144.9098 0.00017655 -85.634 0.69494
8.799 0.98815 5.4622e-005 3.8183 0.011914 0.0001143 0.001176 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.609 0.5943 0.18154 0.020704 18.4957 0.1282 0.00016803 0.76197 0.009571 0.010581 0.0013904 0.98689 0.99167 2.9985e-006 1.1994e-005 0.16615 0.91324 0.90787 0.0013992 0.98722 0.46677 0.0018851 0.42394 2.1611 2.1603 16.0189 144.9098 0.00017641 -85.6342 0.69594
8.8 0.98815 5.4622e-005 3.8183 0.011914 0.00011432 0.001176 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6091 0.59435 0.18155 0.020705 18.4989 0.12821 0.00016804 0.76196 0.0095714 0.010581 0.0013903 0.98689 0.99167 2.9984e-006 1.1994e-005 0.16615 0.91346 0.90796 0.0013992 0.98728 0.46696 0.001885 0.42396 2.1617 2.1609 16.0189 144.9099 0.00017627 -85.6344 0.69694
8.801 0.98815 5.4621e-005 3.8183 0.011914 0.00011433 0.001176 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6091 0.59439 0.18157 0.020706 18.5021 0.12821 0.00016805 0.76196 0.0095717 0.010582 0.0013903 0.98689 0.99167 2.9983e-006 1.1993e-005 0.16616 0.91368 0.90805 0.0013992 0.98735 0.46715 0.001885 0.42397 2.1623 2.1615 16.0189 144.9099 0.00017613 -85.6346 0.69794
8.802 0.98815 5.4621e-005 3.8183 0.011914 0.00011434 0.001176 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6092 0.59444 0.18158 0.020707 18.5053 0.12822 0.00016806 0.76195 0.0095721 0.010582 0.0013902 0.98689 0.99167 2.9982e-006 1.1993e-005 0.16616 0.91389 0.90814 0.0013992 0.98741 0.46733 0.0018849 0.42399 2.1628 2.1621 16.0189 144.9099 0.000176 -85.6349 0.69894
8.803 0.98815 5.4621e-005 3.8183 0.011914 0.00011435 0.001176 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6093 0.59448 0.18159 0.020708 18.5085 0.12822 0.00016807 0.76194 0.0095724 0.010582 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.16616 0.91411 0.90822 0.0013991 0.98748 0.46752 0.0018849 0.424 2.1634 2.1626 16.0188 144.9099 0.00017586 -85.6351 0.69994
8.804 0.98815 5.4621e-005 3.8183 0.011914 0.00011437 0.001176 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6094 0.59452 0.18161 0.020709 18.5117 0.12823 0.00016807 0.76194 0.0095728 0.010583 0.0013901 0.98689 0.99167 2.998e-006 1.1992e-005 0.16617 0.91433 0.90831 0.0013991 0.98754 0.4677 0.0018849 0.42402 2.164 2.1632 16.0188 144.9099 0.00017572 -85.6353 0.70094
8.805 0.98815 5.4621e-005 3.8183 0.011914 0.00011438 0.0011761 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6095 0.59457 0.18162 0.02071 18.5149 0.12824 0.00016808 0.76193 0.0095731 0.010583 0.0013901 0.98689 0.99167 2.9979e-006 1.1991e-005 0.16617 0.91455 0.9084 0.0013991 0.9876 0.46789 0.0018848 0.42403 2.1646 2.1638 16.0188 144.91 0.00017559 -85.6355 0.70194
8.806 0.98815 5.4621e-005 3.8183 0.011914 0.00011439 0.0011761 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6096 0.59461 0.18163 0.020711 18.5182 0.12824 0.00016809 0.76193 0.0095735 0.010584 0.00139 0.9869 0.99167 2.9978e-006 1.1991e-005 0.16617 0.91476 0.90849 0.0013991 0.98766 0.46807 0.0018848 0.42405 2.1651 2.1644 16.0188 144.91 0.00017545 -85.6357 0.70294
8.807 0.98815 5.4621e-005 3.8183 0.011914 0.0001144 0.0011761 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6096 0.59466 0.18164 0.020712 18.5214 0.12825 0.0001681 0.76192 0.0095738 0.010584 0.00139 0.9869 0.99167 2.9976e-006 1.1991e-005 0.16617 0.91498 0.90858 0.001399 0.98773 0.46826 0.0018848 0.42406 2.1657 2.1649 16.0187 144.91 0.00017531 -85.6359 0.70394
8.808 0.98815 5.4621e-005 3.8183 0.011914 0.00011442 0.0011761 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6097 0.5947 0.18166 0.020713 18.5246 0.12825 0.00016811 0.76191 0.0095742 0.010584 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.16618 0.91519 0.90867 0.001399 0.98779 0.46844 0.0018847 0.42408 2.1663 2.1655 16.0187 144.91 0.00017518 -85.6361 0.70494
8.809 0.98815 5.4621e-005 3.8183 0.011913 0.00011443 0.0011761 0.23363 0.00065931 0.23429 0.21619 0 0.032263 0.0389 0 1.6098 0.59475 0.18167 0.020714 18.5278 0.12826 0.00016812 0.76191 0.0095745 0.010585 0.0013899 0.9869 0.99167 2.9974e-006 1.199e-005 0.16618 0.9154 0.90875 0.001399 0.98785 0.46863 0.0018847 0.42409 2.1669 2.1661 16.0187 144.91 0.00017505 -85.6363 0.70594
8.81 0.98815 5.4621e-005 3.8183 0.011913 0.00011444 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6099 0.59479 0.18168 0.020715 18.531 0.12827 0.00016813 0.7619 0.0095749 0.010585 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.16618 0.91562 0.90884 0.001399 0.98791 0.46881 0.0018847 0.4241 2.1674 2.1667 16.0187 144.9101 0.00017491 -85.6365 0.70694
8.811 0.98815 5.4621e-005 3.8183 0.011913 0.00011446 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.61 0.59483 0.1817 0.020716 18.5342 0.12827 0.00016814 0.7619 0.0095752 0.010585 0.0013898 0.9869 0.99168 2.9972e-006 1.1989e-005 0.16618 0.91583 0.90893 0.0013989 0.98797 0.469 0.0018847 0.42412 2.168 2.1672 16.0186 144.9101 0.00017478 -85.6367 0.70794
8.812 0.98815 5.4621e-005 3.8183 0.011913 0.00011447 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6101 0.59488 0.18171 0.020717 18.5374 0.12828 0.00016815 0.76189 0.0095755 0.010586 0.0013897 0.9869 0.99168 2.9971e-006 1.1988e-005 0.16619 0.91604 0.90901 0.0013989 0.98803 0.46918 0.0018846 0.42413 2.1686 2.1678 16.0186 144.9101 0.00017465 -85.6369 0.70894
8.813 0.98815 5.462e-005 3.8183 0.011913 0.00011448 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6101 0.59492 0.18172 0.020718 18.5406 0.12829 0.00016816 0.76188 0.0095759 0.010586 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.16619 0.91625 0.9091 0.0013989 0.98809 0.46937 0.0018846 0.42415 2.1691 2.1684 16.0186 144.9101 0.00017451 -85.6371 0.70994
8.814 0.98815 5.462e-005 3.8183 0.011913 0.00011449 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6102 0.59497 0.18174 0.020719 18.5438 0.12829 0.00016817 0.76188 0.0095762 0.010587 0.0013897 0.9869 0.99168 2.9969e-006 1.1988e-005 0.16619 0.91646 0.90919 0.0013989 0.98815 0.46955 0.0018846 0.42416 2.1697 2.1689 16.0186 144.9101 0.00017438 -85.6373 0.71094
8.815 0.98815 5.462e-005 3.8183 0.011913 0.00011451 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6103 0.59501 0.18175 0.020721 18.5471 0.1283 0.00016818 0.76187 0.0095766 0.010587 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.16619 0.91667 0.90927 0.0013988 0.98821 0.46974 0.0018845 0.42418 2.1703 2.1695 16.0185 144.9102 0.00017425 -85.6375 0.71194
8.816 0.98815 5.462e-005 3.8183 0.011913 0.00011452 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6104 0.59506 0.18176 0.020722 18.5503 0.1283 0.00016819 0.76186 0.0095769 0.010587 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.1662 0.91688 0.90936 0.0013988 0.98826 0.46992 0.0018845 0.42419 2.1708 2.1701 16.0185 144.9102 0.00017412 -85.6377 0.71294
8.817 0.98815 5.462e-005 3.8183 0.011913 0.00011453 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6105 0.5951 0.18178 0.020723 18.5535 0.12831 0.0001682 0.76186 0.0095773 0.010588 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.1662 0.91709 0.90944 0.0013988 0.98832 0.47011 0.0018845 0.42421 2.1714 2.1706 16.0185 144.9102 0.00017399 -85.6379 0.71394
8.818 0.98815 5.462e-005 3.8183 0.011913 0.00011455 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6106 0.59515 0.18179 0.020724 18.5567 0.12832 0.00016821 0.76185 0.0095776 0.010588 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.1662 0.9173 0.90953 0.0013988 0.98838 0.47029 0.0018844 0.42422 2.1719 2.1712 16.0185 144.9102 0.00017386 -85.6381 0.71494
8.819 0.98815 5.462e-005 3.8183 0.011913 0.00011456 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6106 0.59519 0.1818 0.020725 18.5599 0.12832 0.00016821 0.76185 0.009578 0.010588 0.0013894 0.9869 0.99168 2.9964e-006 1.1986e-005 0.16621 0.9175 0.90961 0.0013988 0.98844 0.47048 0.0018844 0.42424 2.1725 2.1717 16.0184 144.9102 0.00017373 -85.6383 0.71594
8.82 0.98815 5.462e-005 3.8183 0.011913 0.00011457 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6107 0.59523 0.18181 0.020726 18.5631 0.12833 0.00016822 0.76184 0.0095783 0.010589 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.16621 0.91771 0.90969 0.0013987 0.98849 0.47066 0.0018844 0.42425 2.173 2.1723 16.0184 144.9103 0.0001736 -85.6384 0.71694
8.821 0.98815 5.462e-005 3.8183 0.011913 0.00011458 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6108 0.59528 0.18183 0.020727 18.5663 0.12833 0.00016823 0.76183 0.0095787 0.010589 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.16621 0.91792 0.90978 0.0013987 0.98855 0.47085 0.0018843 0.42427 2.1736 2.1729 16.0184 144.9103 0.00017347 -85.6386 0.71794
8.822 0.98815 5.462e-005 3.8183 0.011913 0.0001146 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6109 0.59532 0.18184 0.020728 18.5695 0.12834 0.00016824 0.76183 0.009579 0.010589 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.16621 0.91812 0.90986 0.0013987 0.98861 0.47103 0.0018843 0.42428 2.1742 2.1734 16.0184 144.9103 0.00017334 -85.6388 0.71894
8.823 0.98815 5.462e-005 3.8183 0.011913 0.00011461 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.611 0.59537 0.18185 0.020729 18.5728 0.12835 0.00016825 0.76182 0.0095794 0.01059 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.16622 0.91832 0.90994 0.0013987 0.98866 0.47121 0.0018843 0.42429 2.1747 2.174 16.0183 144.9103 0.00017322 -85.639 0.71994
8.824 0.98815 5.462e-005 3.8183 0.011913 0.00011462 0.0011761 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6111 0.59541 0.18187 0.02073 18.576 0.12835 0.00016826 0.76182 0.0095797 0.01059 0.0013892 0.98691 0.99168 2.9959e-006 1.1984e-005 0.16622 0.91853 0.91003 0.0013986 0.98872 0.4714 0.0018843 0.42431 2.1753 2.1745 16.0183 144.9103 0.00017309 -85.6392 0.72094
8.825 0.98815 5.4619e-005 3.8183 0.011913 0.00011463 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6112 0.59546 0.18188 0.020731 18.5792 0.12836 0.00016827 0.76181 0.0095801 0.010591 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.16622 0.91873 0.91011 0.0013986 0.98877 0.47158 0.0018842 0.42432 2.1758 2.1751 16.0183 144.9104 0.00017296 -85.6394 0.72194
8.826 0.98815 5.4619e-005 3.8183 0.011913 0.00011465 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6112 0.5955 0.18189 0.020732 18.5824 0.12836 0.00016828 0.7618 0.0095804 0.010591 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.16622 0.91893 0.91019 0.0013986 0.98883 0.47177 0.0018842 0.42434 2.1764 2.1756 16.0183 144.9104 0.00017284 -85.6395 0.72294
8.827 0.98815 5.4619e-005 3.8183 0.011913 0.00011466 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6113 0.59554 0.18191 0.020733 18.5856 0.12837 0.00016829 0.7618 0.0095807 0.010591 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.16623 0.91914 0.91027 0.0013986 0.98888 0.47195 0.0018842 0.42435 2.1769 2.1762 16.0182 144.9104 0.00017271 -85.6397 0.72394
8.828 0.98815 5.4619e-005 3.8183 0.011913 0.00011467 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6114 0.59559 0.18192 0.020734 18.5888 0.12838 0.0001683 0.76179 0.0095811 0.010592 0.0013891 0.98691 0.99168 2.9955e-006 1.1982e-005 0.16623 0.91934 0.91036 0.0013986 0.98893 0.47214 0.0018841 0.42437 2.1775 2.1767 16.0182 144.9104 0.00017259 -85.6399 0.72494
8.829 0.98815 5.4619e-005 3.8183 0.011913 0.00011469 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6115 0.59563 0.18193 0.020735 18.5921 0.12838 0.00016831 0.76179 0.0095814 0.010592 0.001389 0.98691 0.99168 2.9954e-006 1.1982e-005 0.16623 0.91954 0.91044 0.0013985 0.98899 0.47232 0.0018841 0.42438 2.178 2.1773 16.0182 144.9104 0.00017246 -85.6401 0.72594
8.83 0.98815 5.4619e-005 3.8183 0.011913 0.0001147 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6116 0.59568 0.18194 0.020736 18.5953 0.12839 0.00016832 0.76178 0.0095818 0.010592 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.16623 0.91974 0.91052 0.0013985 0.98904 0.4725 0.0018841 0.4244 2.1785 2.1778 16.0181 144.9105 0.00017234 -85.6402 0.72694
8.831 0.98815 5.4619e-005 3.8183 0.011913 0.00011471 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6117 0.59572 0.18196 0.020737 18.5985 0.12839 0.00016833 0.76177 0.0095821 0.010593 0.001389 0.98691 0.99168 2.9953e-006 1.1981e-005 0.16624 0.91994 0.9106 0.0013985 0.98909 0.47269 0.0018841 0.42441 2.1791 2.1784 16.0181 144.9105 0.00017221 -85.6404 0.72794
8.832 0.98815 5.4619e-005 3.8183 0.011913 0.00011472 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6117 0.59577 0.18197 0.020738 18.6017 0.1284 0.00016834 0.76177 0.0095825 0.010593 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.16624 0.92014 0.91068 0.0013985 0.98915 0.47287 0.001884 0.42443 2.1796 2.1789 16.0181 144.9105 0.00017209 -85.6406 0.72894
8.833 0.98815 5.4619e-005 3.8183 0.011913 0.00011474 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6118 0.59581 0.18198 0.020739 18.6049 0.12841 0.00016835 0.76176 0.0095828 0.010593 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.16624 0.92033 0.91076 0.0013984 0.9892 0.47305 0.001884 0.42444 2.1802 2.1794 16.0181 144.9105 0.00017197 -85.6408 0.72994
8.834 0.98815 5.4619e-005 3.8183 0.011913 0.00011475 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6119 0.59586 0.182 0.02074 18.6082 0.12841 0.00016835 0.76176 0.0095832 0.010594 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.16625 0.92053 0.91084 0.0013984 0.98925 0.47324 0.001884 0.42445 2.1807 2.18 16.018 144.9105 0.00017184 -85.6409 0.73094
8.835 0.98815 5.4619e-005 3.8183 0.011913 0.00011476 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.612 0.5959 0.18201 0.020741 18.6114 0.12842 0.00016836 0.76175 0.0095835 0.010594 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.16625 0.92073 0.91092 0.0013984 0.9893 0.47342 0.0018839 0.42447 2.1812 2.1805 16.018 144.9106 0.00017172 -85.6411 0.73194
8.836 0.98815 5.4619e-005 3.8183 0.011913 0.00011478 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6121 0.59594 0.18202 0.020742 18.6146 0.12843 0.00016837 0.76174 0.0095839 0.010595 0.0013888 0.98691 0.99168 2.9948e-006 1.1979e-005 0.16625 0.92092 0.911 0.0013984 0.98935 0.4736 0.0018839 0.42448 2.1818 2.1811 16.018 144.9106 0.0001716 -85.6413 0.73294
8.837 0.98815 5.4618e-005 3.8183 0.011913 0.00011479 0.0011762 0.23363 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6122 0.59599 0.18204 0.020743 18.6178 0.12843 0.00016838 0.76174 0.0095842 0.010595 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.16625 0.92112 0.91108 0.0013984 0.9894 0.47379 0.0018839 0.4245 2.1823 2.1816 16.018 144.9106 0.00017148 -85.6414 0.73394
8.838 0.98815 5.4618e-005 3.8183 0.011913 0.0001148 0.0011762 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6122 0.59603 0.18205 0.020744 18.621 0.12844 0.00016839 0.76173 0.0095846 0.010595 0.0013887 0.98691 0.99168 2.9946e-006 1.1978e-005 0.16626 0.92132 0.91115 0.0013983 0.98945 0.47397 0.0018839 0.42451 2.1829 2.1821 16.0179 144.9106 0.00017136 -85.6416 0.73494
8.839 0.98815 5.4618e-005 3.8183 0.011913 0.00011481 0.0011762 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6123 0.59608 0.18206 0.020745 18.6242 0.12844 0.0001684 0.76172 0.0095849 0.010596 0.0013886 0.98691 0.99168 2.9946e-006 1.1978e-005 0.16626 0.92151 0.91123 0.0013983 0.98951 0.47415 0.0018838 0.42453 2.1834 2.1827 16.0179 144.9106 0.00017124 -85.6417 0.73594
8.84 0.98815 5.4618e-005 3.8183 0.011913 0.00011483 0.0011762 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6124 0.59612 0.18208 0.020746 18.6275 0.12845 0.00016841 0.76172 0.0095852 0.010596 0.0013886 0.98691 0.99169 2.9945e-006 1.1978e-005 0.16626 0.9217 0.91131 0.0013983 0.98955 0.47434 0.0018838 0.42454 2.1839 2.1832 16.0179 144.9107 0.00017112 -85.6419 0.73694
8.841 0.98815 5.4618e-005 3.8183 0.011913 0.00011484 0.0011762 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6125 0.59617 0.18209 0.020747 18.6307 0.12846 0.00016842 0.76171 0.0095856 0.010596 0.0013886 0.98691 0.99169 2.9944e-006 1.1977e-005 0.16626 0.9219 0.91139 0.0013983 0.9896 0.47452 0.0018838 0.42456 2.1844 2.1837 16.0179 144.9107 0.000171 -85.6421 0.73794
8.842 0.98815 5.4618e-005 3.8183 0.011913 0.00011485 0.0011762 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6126 0.59621 0.1821 0.020748 18.6339 0.12846 0.00016843 0.76171 0.0095859 0.010597 0.0013885 0.98691 0.99169 2.9943e-006 1.1977e-005 0.16627 0.92209 0.91147 0.0013983 0.98965 0.4747 0.0018838 0.42457 2.185 2.1843 16.0178 144.9107 0.00017088 -85.6422 0.73894
8.843 0.98815 5.4618e-005 3.8183 0.011913 0.00011486 0.0011762 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6127 0.59625 0.18211 0.020749 18.6371 0.12847 0.00016844 0.7617 0.0095863 0.010597 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.16627 0.92228 0.91154 0.0013982 0.9897 0.47489 0.0018837 0.42459 2.1855 2.1848 16.0178 144.9107 0.00017076 -85.6424 0.73994
8.844 0.98815 5.4618e-005 3.8183 0.011913 0.00011488 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6127 0.5963 0.18213 0.02075 18.6404 0.12847 0.00016845 0.76169 0.0095866 0.010597 0.0013885 0.98692 0.99169 2.9941e-006 1.1976e-005 0.16627 0.92247 0.91162 0.0013982 0.98975 0.47507 0.0018837 0.4246 2.186 2.1853 16.0178 144.9108 0.00017064 -85.6425 0.74094
8.845 0.98815 5.4618e-005 3.8183 0.011913 0.00011489 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6128 0.59634 0.18214 0.020751 18.6436 0.12848 0.00016846 0.76169 0.009587 0.010598 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.16627 0.92266 0.9117 0.0013982 0.9898 0.47525 0.0018837 0.42461 2.1866 2.1859 16.0177 144.9108 0.00017052 -85.6427 0.74194
8.846 0.98815 5.4618e-005 3.8183 0.011913 0.0001149 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6129 0.59639 0.18215 0.020752 18.6468 0.12849 0.00016847 0.76168 0.0095873 0.010598 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.16628 0.92285 0.91177 0.0013982 0.98985 0.47544 0.0018837 0.42463 2.1871 2.1864 16.0177 144.9108 0.00017041 -85.6429 0.74294
8.847 0.98815 5.4618e-005 3.8183 0.011913 0.00011492 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.613 0.59643 0.18217 0.020753 18.65 0.12849 0.00016848 0.76168 0.0095877 0.010599 0.0013883 0.98692 0.99169 2.9939e-006 1.1975e-005 0.16628 0.92304 0.91185 0.0013982 0.9899 0.47562 0.0018836 0.42464 2.1876 2.1869 16.0177 144.9108 0.00017029 -85.643 0.74394
8.848 0.98815 5.4618e-005 3.8183 0.011913 0.00011493 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6131 0.59648 0.18218 0.020754 18.6532 0.1285 0.00016848 0.76167 0.009588 0.010599 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.16628 0.92323 0.91193 0.0013982 0.98994 0.4758 0.0018836 0.42466 2.1881 2.1874 16.0177 144.9108 0.00017017 -85.6432 0.74494
8.849 0.98815 5.4617e-005 3.8183 0.011913 0.00011494 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6132 0.59652 0.18219 0.020755 18.6565 0.1285 0.00016849 0.76166 0.0095884 0.010599 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.16628 0.92342 0.912 0.0013981 0.98999 0.47598 0.0018836 0.42467 2.1887 2.188 16.0176 144.9109 0.00017006 -85.6433 0.74594
8.85 0.98815 5.4617e-005 3.8183 0.011913 0.00011495 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6132 0.59656 0.18221 0.020756 18.6597 0.12851 0.0001685 0.76166 0.0095887 0.0106 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16629 0.92361 0.91208 0.0013981 0.99004 0.47617 0.0018836 0.42469 2.1892 2.1885 16.0176 144.9109 0.00016994 -85.6435 0.74694
8.851 0.98815 5.4617e-005 3.8183 0.011913 0.00011497 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6133 0.59661 0.18222 0.020757 18.6629 0.12852 0.00016851 0.76165 0.009589 0.0106 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16629 0.9238 0.91215 0.0013981 0.99008 0.47635 0.0018835 0.4247 2.1897 2.189 16.0176 144.9109 0.00016983 -85.6436 0.74794
8.852 0.98815 5.4617e-005 3.8183 0.011913 0.00011498 0.0011763 0.23362 0.00065931 0.23428 0.21619 0 0.032263 0.0389 0 1.6134 0.59665 0.18223 0.020758 18.6661 0.12852 0.00016852 0.76165 0.0095894 0.0106 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.16629 0.92398 0.91223 0.0013981 0.99013 0.47653 0.0018835 0.42472 2.1902 2.1895 16.0175 144.9109 0.00016971 -85.6438 0.74894
8.853 0.98815 5.4617e-005 3.8183 0.011913 0.00011499 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6135 0.5967 0.18224 0.020759 18.6694 0.12853 0.00016853 0.76164 0.0095897 0.010601 0.0013882 0.98692 0.99169 2.9934e-006 1.1974e-005 0.1663 0.92417 0.9123 0.0013981 0.99017 0.47671 0.0018835 0.42473 2.1907 2.19 16.0175 144.9109 0.0001696 -85.6439 0.74994
8.854 0.98815 5.4617e-005 3.8183 0.011913 0.00011501 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6136 0.59674 0.18226 0.02076 18.6726 0.12853 0.00016854 0.76163 0.0095901 0.010601 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.1663 0.92435 0.91237 0.001398 0.99022 0.4769 0.0018835 0.42474 2.1912 2.1906 16.0175 144.911 0.00016948 -85.644 0.75094
8.855 0.98815 5.4617e-005 3.8183 0.011913 0.00011502 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6137 0.59679 0.18227 0.020762 18.6758 0.12854 0.00016855 0.76163 0.0095904 0.010601 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.1663 0.92454 0.91245 0.001398 0.99027 0.47708 0.0018835 0.42476 2.1918 2.1911 16.0175 144.911 0.00016937 -85.6442 0.75194
8.856 0.98815 5.4617e-005 3.8183 0.011913 0.00011503 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6137 0.59683 0.18228 0.020763 18.679 0.12855 0.00016856 0.76162 0.0095908 0.010602 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.1663 0.92472 0.91252 0.001398 0.99031 0.47726 0.0018834 0.42477 2.1923 2.1916 16.0174 144.911 0.00016926 -85.6443 0.75294
8.857 0.98815 5.4617e-005 3.8183 0.011913 0.00011504 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6138 0.59688 0.1823 0.020764 18.6823 0.12855 0.00016857 0.76162 0.0095911 0.010602 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.16631 0.92491 0.9126 0.001398 0.99035 0.47744 0.0018834 0.42479 2.1928 2.1921 16.0174 144.911 0.00016914 -85.6445 0.75394
8.858 0.98815 5.4617e-005 3.8183 0.011913 0.00011506 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6139 0.59692 0.18231 0.020765 18.6855 0.12856 0.00016858 0.76161 0.0095915 0.010603 0.001388 0.98692 0.99169 2.993e-006 1.1972e-005 0.16631 0.92509 0.91267 0.001398 0.9904 0.47762 0.0018834 0.4248 2.1933 2.1926 16.0174 144.911 0.00016903 -85.6446 0.75494
8.859 0.98815 5.4617e-005 3.8183 0.011913 0.00011507 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.614 0.59696 0.18232 0.020766 18.6887 0.12857 0.00016859 0.7616 0.0095918 0.010603 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.16631 0.92527 0.91274 0.001398 0.99044 0.47781 0.0018834 0.42482 2.1938 2.1931 16.0174 144.9111 0.00016892 -85.6448 0.75594
8.86 0.98815 5.4617e-005 3.8183 0.011913 0.00011508 0.0011763 0.23362 0.00065931 0.23428 0.21618 0 0.032263 0.0389 0 1.6141 0.59701 0.18234 0.020767 18.6919 0.12857 0.0001686 0.7616 0.0095921 0.010603 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.16631 0.92546 0.91281 0.0013979 0.99049 0.47799 0.0018833 0.42483 2.1943 2.1936 16.0173 144.9111 0.00016881 -85.6449 0.75694
8.861 0.98815 5.4616e-005 3.8183 0.011913 0.00011509 0.0011763 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6142 0.59705 0.18235 0.020768 18.6952 0.12858 0.00016861 0.76159 0.0095925 0.010604 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.16632 0.92564 0.91289 0.0013979 0.99053 0.47817 0.0018833 0.42485 2.1948 2.1941 16.0173 144.9111 0.0001687 -85.645 0.75794
8.862 0.98815 5.4616e-005 3.8183 0.011913 0.00011511 0.0011763 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6142 0.5971 0.18236 0.020769 18.6984 0.12858 0.00016861 0.76159 0.0095928 0.010604 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.16632 0.92582 0.91296 0.0013979 0.99057 0.47835 0.0018833 0.42486 2.1953 2.1947 16.0173 144.9111 0.00016858 -85.6452 0.75894
8.863 0.98815 5.4616e-005 3.8183 0.011913 0.00011512 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6143 0.59714 0.18238 0.02077 18.7016 0.12859 0.00016862 0.76158 0.0095932 0.010604 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.16632 0.926 0.91303 0.0013979 0.99062 0.47853 0.0018833 0.42487 2.1958 2.1952 16.0172 144.9111 0.00016847 -85.6453 0.75994
8.864 0.98815 5.4616e-005 3.8183 0.011913 0.00011513 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6144 0.59719 0.18239 0.020771 18.7049 0.1286 0.00016863 0.76157 0.0095935 0.010605 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.16632 0.92618 0.9131 0.0013979 0.99066 0.47872 0.0018833 0.42489 2.1963 2.1957 16.0172 144.9112 0.00016836 -85.6454 0.76094
8.865 0.98815 5.4616e-005 3.8183 0.011912 0.00011515 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6145 0.59723 0.1824 0.020772 18.7081 0.1286 0.00016864 0.76157 0.0095939 0.010605 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.16633 0.92636 0.91317 0.0013979 0.9907 0.4789 0.0018832 0.4249 2.1968 2.1962 16.0172 144.9112 0.00016825 -85.6456 0.76194
8.866 0.98815 5.4616e-005 3.8183 0.011912 0.00011516 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6146 0.59727 0.18241 0.020773 18.7113 0.12861 0.00016865 0.76156 0.0095942 0.010605 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.16633 0.92654 0.91324 0.0013978 0.99074 0.47908 0.0018832 0.42492 2.1973 2.1967 16.0172 144.9112 0.00016815 -85.6457 0.76294
8.867 0.98815 5.4616e-005 3.8183 0.011912 0.00011517 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6147 0.59732 0.18243 0.020774 18.7145 0.12861 0.00016866 0.76156 0.0095946 0.010606 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.16633 0.92671 0.91332 0.0013978 0.99079 0.47926 0.0018832 0.42493 2.1979 2.1972 16.0171 144.9112 0.00016804 -85.6458 0.76394
8.868 0.98815 5.4616e-005 3.8183 0.011912 0.00011518 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6147 0.59736 0.18244 0.020775 18.7178 0.12862 0.00016867 0.76155 0.0095949 0.010606 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.16634 0.92689 0.91339 0.0013978 0.99083 0.47944 0.0018832 0.42495 2.1984 2.1977 16.0171 144.9112 0.00016793 -85.646 0.76494
8.869 0.98815 5.4616e-005 3.8183 0.011912 0.0001152 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6148 0.59741 0.18245 0.020776 18.721 0.12863 0.00016868 0.76154 0.0095952 0.010607 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.16634 0.92707 0.91346 0.0013978 0.99087 0.47962 0.0018831 0.42496 2.1989 2.1982 16.0171 144.9113 0.00016782 -85.6461 0.76594
8.87 0.98815 5.4616e-005 3.8183 0.011912 0.00011521 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6149 0.59745 0.18247 0.020777 18.7242 0.12863 0.00016869 0.76154 0.0095956 0.010607 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.16634 0.92725 0.91353 0.0013978 0.99091 0.4798 0.0018831 0.42498 2.1993 2.1987 16.017 144.9113 0.00016771 -85.6462 0.76694
8.871 0.98815 5.4616e-005 3.8183 0.011912 0.00011522 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.615 0.5975 0.18248 0.020778 18.7275 0.12864 0.0001687 0.76153 0.0095959 0.010607 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.16634 0.92742 0.9136 0.0013978 0.99095 0.47999 0.0018831 0.42499 2.1998 2.1992 16.017 144.9113 0.0001676 -85.6464 0.76794
8.872 0.98815 5.4616e-005 3.8183 0.011912 0.00011524 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6151 0.59754 0.18249 0.020779 18.7307 0.12864 0.00016871 0.76152 0.0095963 0.010608 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16635 0.9276 0.91367 0.0013977 0.99099 0.48017 0.0018831 0.425 2.2003 2.1997 16.017 144.9113 0.0001675 -85.6465 0.76894
8.873 0.98815 5.4615e-005 3.8183 0.011912 0.00011525 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6152 0.59758 0.18251 0.02078 18.7339 0.12865 0.00016872 0.76152 0.0095966 0.010608 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16635 0.92777 0.91374 0.0013977 0.99103 0.48035 0.0018831 0.42502 2.2008 2.2002 16.017 144.9113 0.00016739 -85.6466 0.76994
8.874 0.98815 5.4615e-005 3.8183 0.011912 0.00011526 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6152 0.59763 0.18252 0.020781 18.7372 0.12866 0.00016873 0.76151 0.009597 0.010608 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.16635 0.92795 0.9138 0.0013977 0.99107 0.48053 0.001883 0.42503 2.2013 2.2007 16.0169 144.9114 0.00016729 -85.6467 0.77094
8.875 0.98815 5.4615e-005 3.8183 0.011912 0.00011527 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6153 0.59767 0.18253 0.020782 18.7404 0.12866 0.00016874 0.76151 0.0095973 0.010609 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.16635 0.92812 0.91387 0.0013977 0.99111 0.48071 0.001883 0.42505 2.2018 2.2012 16.0169 144.9114 0.00016718 -85.6469 0.77194
8.876 0.98815 5.4615e-005 3.8183 0.011912 0.00011529 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6154 0.59772 0.18254 0.020783 18.7436 0.12867 0.00016874 0.7615 0.0095977 0.010609 0.0013874 0.98693 0.9917 2.9918e-006 1.1967e-005 0.16636 0.92829 0.91394 0.0013977 0.99115 0.48089 0.001883 0.42506 2.2023 2.2017 16.0169 144.9114 0.00016707 -85.647 0.77294
8.877 0.98815 5.4615e-005 3.8183 0.011912 0.0001153 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6155 0.59776 0.18256 0.020784 18.7469 0.12867 0.00016875 0.76149 0.009598 0.010609 0.0013874 0.98693 0.9917 2.9917e-006 1.1967e-005 0.16636 0.92847 0.91401 0.0013977 0.99119 0.48107 0.001883 0.42508 2.2028 2.2022 16.0168 144.9114 0.00016697 -85.6471 0.77394
8.878 0.98815 5.4615e-005 3.8183 0.011912 0.00011531 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6156 0.59781 0.18257 0.020785 18.7501 0.12868 0.00016876 0.76149 0.0095983 0.01061 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.16636 0.92864 0.91408 0.0013977 0.99123 0.48125 0.001883 0.42509 2.2033 2.2026 16.0168 144.9115 0.00016686 -85.6472 0.77494
8.879 0.98815 5.4615e-005 3.8183 0.011912 0.00011533 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6157 0.59785 0.18258 0.020786 18.7533 0.12869 0.00016877 0.76148 0.0095987 0.01061 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.16636 0.92881 0.91415 0.0013976 0.99127 0.48143 0.0018829 0.4251 2.2038 2.2031 16.0168 144.9115 0.00016676 -85.6474 0.77594
8.88 0.98815 5.4615e-005 3.8183 0.011912 0.00011534 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6157 0.59789 0.1826 0.020787 18.7566 0.12869 0.00016878 0.76148 0.009599 0.010611 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.16637 0.92898 0.91421 0.0013976 0.99131 0.48161 0.0018829 0.42512 2.2043 2.2036 16.0168 144.9115 0.00016666 -85.6475 0.77694
8.881 0.98815 5.4615e-005 3.8183 0.011912 0.00011535 0.0011764 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6158 0.59794 0.18261 0.020788 18.7598 0.1287 0.00016879 0.76147 0.0095994 0.010611 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.16637 0.92915 0.91428 0.0013976 0.99134 0.48179 0.0018829 0.42513 2.2048 2.2041 16.0167 144.9115 0.00016655 -85.6476 0.77794
8.882 0.98815 5.4615e-005 3.8183 0.011912 0.00011536 0.0011765 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6159 0.59798 0.18262 0.020789 18.763 0.1287 0.0001688 0.76146 0.0095997 0.010611 0.0013872 0.98693 0.9917 2.9914e-006 1.1965e-005 0.16637 0.92932 0.91435 0.0013976 0.99138 0.48198 0.0018829 0.42515 2.2053 2.2046 16.0167 144.9115 0.00016645 -85.6477 0.77894
8.883 0.98815 5.4615e-005 3.8183 0.011912 0.00011538 0.0011765 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.616 0.59803 0.18264 0.02079 18.7663 0.12871 0.00016881 0.76146 0.0096001 0.010612 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16637 0.92949 0.91441 0.0013976 0.99142 0.48216 0.0018829 0.42516 2.2057 2.2051 16.0167 144.9116 0.00016635 -85.6478 0.77994
8.884 0.98815 5.4615e-005 3.8183 0.011912 0.00011539 0.0011765 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6161 0.59807 0.18265 0.020791 18.7695 0.12872 0.00016882 0.76145 0.0096004 0.010612 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16638 0.92966 0.91448 0.0013976 0.99146 0.48234 0.0018829 0.42518 2.2062 2.2056 16.0166 144.9116 0.00016624 -85.6479 0.78094
8.885 0.98815 5.4614e-005 3.8183 0.011912 0.0001154 0.0011765 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6162 0.59812 0.18266 0.020792 18.7727 0.12872 0.00016883 0.76145 0.0096007 0.010612 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.16638 0.92983 0.91455 0.0013976 0.99149 0.48252 0.0018828 0.42519 2.2067 2.2061 16.0166 144.9116 0.00016614 -85.6481 0.78194
8.886 0.98815 5.4614e-005 3.8183 0.011912 0.00011541 0.0011765 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6162 0.59816 0.18267 0.020793 18.776 0.12873 0.00016884 0.76144 0.0096011 0.010613 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.16638 0.93 0.91461 0.0013975 0.99153 0.4827 0.0018828 0.4252 2.2072 2.2065 16.0166 144.9116 0.00016604 -85.6482 0.78294
8.887 0.98815 5.4614e-005 3.8183 0.011912 0.00011543 0.0011765 0.23362 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6163 0.5982 0.18269 0.020794 18.7792 0.12873 0.00016885 0.76143 0.0096014 0.010613 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.16639 0.93016 0.91468 0.0013975 0.99157 0.48288 0.0018828 0.42522 2.2077 2.207 16.0166 144.9116 0.00016594 -85.6483 0.78394
8.888 0.98815 5.4614e-005 3.8183 0.011912 0.00011544 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6164 0.59825 0.1827 0.020795 18.7824 0.12874 0.00016886 0.76143 0.0096018 0.010613 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16639 0.93033 0.91475 0.0013975 0.9916 0.48306 0.0018828 0.42523 2.2081 2.2075 16.0165 144.9117 0.00016584 -85.6484 0.78494
8.889 0.98815 5.4614e-005 3.8183 0.011912 0.00011545 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6165 0.59829 0.18271 0.020796 18.7857 0.12875 0.00016887 0.76142 0.0096021 0.010614 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16639 0.9305 0.91481 0.0013975 0.99164 0.48324 0.0018828 0.42525 2.2086 2.208 16.0165 144.9117 0.00016574 -85.6485 0.78594
8.89 0.98815 5.4614e-005 3.8183 0.011912 0.00011547 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6166 0.59834 0.18273 0.020797 18.7889 0.12875 0.00016887 0.76142 0.0096025 0.010614 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.16639 0.93066 0.91488 0.0013975 0.99168 0.48342 0.0018827 0.42526 2.2091 2.2085 16.0165 144.9117 0.00016564 -85.6486 0.78694
8.891 0.98815 5.4614e-005 3.8183 0.011912 0.00011548 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6167 0.59838 0.18274 0.020798 18.7922 0.12876 0.00016888 0.76141 0.0096028 0.010615 0.001387 0.98693 0.9917 2.9909e-006 1.1963e-005 0.1664 0.93083 0.91494 0.0013975 0.99171 0.4836 0.0018827 0.42528 2.2096 2.2089 16.0164 144.9117 0.00016554 -85.6487 0.78794
8.892 0.98815 5.4614e-005 3.8183 0.011912 0.00011549 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6168 0.59843 0.18275 0.020799 18.7954 0.12876 0.00016889 0.7614 0.0096032 0.010615 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.1664 0.93099 0.91501 0.0013975 0.99175 0.48378 0.0018827 0.42529 2.2101 2.2094 16.0164 144.9117 0.00016544 -85.6488 0.78894
8.893 0.98815 5.4614e-005 3.8183 0.011912 0.0001155 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6168 0.59847 0.18277 0.0208 18.7986 0.12877 0.0001689 0.7614 0.0096035 0.010615 0.001387 0.98694 0.9917 2.9907e-006 1.1963e-005 0.1664 0.93116 0.91507 0.0013974 0.99178 0.48396 0.0018827 0.4253 2.2105 2.2099 16.0164 144.9118 0.00016534 -85.649 0.78994
8.894 0.98815 5.4614e-005 3.8183 0.011912 0.00011552 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6169 0.59851 0.18278 0.020801 18.8019 0.12878 0.00016891 0.76139 0.0096038 0.010616 0.0013869 0.98694 0.9917 2.9907e-006 1.1963e-005 0.1664 0.93132 0.91513 0.0013974 0.99182 0.48414 0.0018827 0.42532 2.211 2.2104 16.0164 144.9118 0.00016524 -85.6491 0.79094
8.895 0.98815 5.4614e-005 3.8183 0.011912 0.00011553 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.617 0.59856 0.18279 0.020802 18.8051 0.12878 0.00016892 0.76139 0.0096042 0.010616 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16641 0.93148 0.9152 0.0013974 0.99185 0.48432 0.0018827 0.42533 2.2115 2.2108 16.0163 144.9118 0.00016514 -85.6492 0.79194
8.896 0.98815 5.4614e-005 3.8183 0.011912 0.00011554 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6171 0.5986 0.1828 0.020803 18.8083 0.12879 0.00016893 0.76138 0.0096045 0.010616 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16641 0.93165 0.91526 0.0013974 0.99189 0.4845 0.0018826 0.42535 2.2119 2.2113 16.0163 144.9118 0.00016504 -85.6493 0.79294
8.897 0.98815 5.4613e-005 3.8183 0.011912 0.00011556 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6172 0.59865 0.18282 0.020804 18.8116 0.1288 0.00016894 0.76137 0.0096049 0.010617 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16641 0.93181 0.91533 0.0013974 0.99192 0.48468 0.0018826 0.42536 2.2124 2.2118 16.0163 144.9118 0.00016494 -85.6494 0.79394
8.898 0.98815 5.4613e-005 3.8183 0.011912 0.00011557 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032263 0.0389 0 1.6173 0.59869 0.18283 0.020805 18.8148 0.1288 0.00016895 0.76137 0.0096052 0.010617 0.0013868 0.98694 0.9917 2.9904e-006 1.1962e-005 0.16641 0.93197 0.91539 0.0013974 0.99196 0.48486 0.0018826 0.42538 2.2129 2.2123 16.0162 144.9119 0.00016485 -85.6495 0.79494
8.899 0.98815 5.4613e-005 3.8183 0.011912 0.00011558 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.6173 0.59874 0.18284 0.020806 18.8181 0.12881 0.00016896 0.76136 0.0096055 0.010617 0.0013868 0.98694 0.9917 2.9904e-006 1.1961e-005 0.16642 0.93213 0.91545 0.0013974 0.99199 0.48504 0.0018826 0.42539 2.2134 2.2127 16.0162 144.9119 0.00016475 -85.6496 0.79594
8.9 0.98815 5.4613e-005 3.8183 0.011912 0.00011559 0.0011765 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.6174 0.59878 0.18286 0.020807 18.8213 0.12881 0.00016897 0.76136 0.0096059 0.010618 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16642 0.93229 0.91552 0.0013974 0.99202 0.48521 0.0018826 0.4254 2.2138 2.2132 16.0162 144.9119 0.00016465 -85.6497 0.79694
8.901 0.98815 5.4613e-005 3.8183 0.011912 0.00011561 0.0011766 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.6175 0.59883 0.18287 0.020808 18.8245 0.12882 0.00016898 0.76135 0.0096062 0.010618 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16642 0.93245 0.91558 0.0013973 0.99206 0.48539 0.0018826 0.42542 2.2143 2.2137 16.0161 144.9119 0.00016456 -85.6498 0.79794
8.902 0.98815 5.4613e-005 3.8183 0.011912 0.00011562 0.0011766 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.6176 0.59887 0.18288 0.020809 18.8278 0.12883 0.00016899 0.76134 0.0096066 0.010619 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16642 0.93261 0.91564 0.0013973 0.99209 0.48557 0.0018825 0.42543 2.2148 2.2141 16.0161 144.9119 0.00016446 -85.6499 0.79894
8.903 0.98815 5.4613e-005 3.8183 0.011912 0.00011563 0.0011766 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.6177 0.59891 0.1829 0.02081 18.831 0.12883 0.000169 0.76134 0.0096069 0.010619 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16643 0.93277 0.9157 0.0013973 0.99212 0.48575 0.0018825 0.42545 2.2152 2.2146 16.0161 144.912 0.00016436 -85.65 0.79994
8.904 0.98815 5.4613e-005 3.8183 0.011912 0.00011564 0.0011766 0.23361 0.00065931 0.23427 0.21618 0 0.032264 0.0389 0 1.6178 0.59896 0.18291 0.020811 18.8343 0.12884 0.000169 0.76133 0.0096073 0.010619 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.16643 0.93293 0.91577 0.0013973 0.99216 0.48593 0.0018825 0.42546 2.2157 2.2151 16.0161 144.912 0.00016427 -85.6501 0.80094
8.905 0.98815 5.4613e-005 3.8183 0.011912 0.00011566 0.0011766 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.6178 0.599 0.18292 0.020813 18.8375 0.12884 0.00016901 0.76133 0.0096076 0.01062 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.16643 0.93309 0.91583 0.0013973 0.99219 0.48611 0.0018825 0.42547 2.2162 2.2155 16.016 144.912 0.00016417 -85.6502 0.80194
8.906 0.98815 5.4613e-005 3.8183 0.011912 0.00011567 0.0011766 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.6179 0.59905 0.18293 0.020814 18.8407 0.12885 0.00016902 0.76132 0.0096079 0.01062 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.16644 0.93324 0.91589 0.0013973 0.99222 0.48629 0.0018825 0.42549 2.2166 2.216 16.016 144.912 0.00016408 -85.6503 0.80294
8.907 0.98815 5.4613e-005 3.8183 0.011912 0.00011568 0.0011766 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.618 0.59909 0.18295 0.020815 18.844 0.12886 0.00016903 0.76131 0.0096083 0.01062 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.16644 0.9334 0.91595 0.0013973 0.99225 0.48647 0.0018825 0.4255 2.2171 2.2165 16.016 144.912 0.00016399 -85.6504 0.80394
8.908 0.98815 5.4613e-005 3.8183 0.011912 0.0001157 0.0011766 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.6181 0.59914 0.18296 0.020816 18.8472 0.12886 0.00016904 0.76131 0.0096086 0.010621 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.16644 0.93356 0.91601 0.0013973 0.99229 0.48665 0.0018824 0.42552 2.2175 2.2169 16.0159 144.9121 0.00016389 -85.6505 0.80494
8.909 0.98815 5.4612e-005 3.8183 0.011912 0.00011571 0.0011766 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.6182 0.59918 0.18297 0.020817 18.8505 0.12887 0.00016905 0.7613 0.009609 0.010621 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.16644 0.93371 0.91607 0.0013972 0.99232 0.48683 0.0018824 0.42553 2.218 2.2174 16.0159 144.9121 0.0001638 -85.6506 0.80594
8.91 0.98815 5.4612e-005 3.8183 0.011912 0.00011572 0.0011766 0.23361 0.00065931 0.23427 0.21617 0 0.032264 0.0389 0 1.6183 0.59922 0.18299 0.020818 18.8537 0.12887 0.00016906 0.7613 0.0096093 0.010621 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.16645 0.93387 0.91613 0.0013972 0.99235 0.48701 0.0018824 0.42555 2.2185 2.2178 16.0159 144.9121 0.0001637 -85.6507 0.80694
8.911 0.98815 5.4612e-005 3.8183 0.011912 0.00011573 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6183 0.59927 0.183 0.020819 18.857 0.12888 0.00016907 0.76129 0.0096097 0.010622 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.16645 0.93403 0.91619 0.0013972 0.99238 0.48718 0.0018824 0.42556 2.2189 2.2183 16.0158 144.9121 0.00016361 -85.6508 0.80794
8.912 0.98815 5.4612e-005 3.8183 0.011912 0.00011575 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6184 0.59931 0.18301 0.02082 18.8602 0.12889 0.00016908 0.76128 0.00961 0.010622 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.16645 0.93418 0.91625 0.0013972 0.99241 0.48736 0.0018824 0.42557 2.2194 2.2188 16.0158 144.9121 0.00016352 -85.6509 0.80894
8.913 0.98815 5.4612e-005 3.8183 0.011912 0.00011576 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6185 0.59936 0.18303 0.020821 18.8635 0.12889 0.00016909 0.76128 0.0096103 0.010623 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.16645 0.93433 0.91631 0.0013972 0.99244 0.48754 0.0018824 0.42559 2.2198 2.2192 16.0158 144.9122 0.00016343 -85.651 0.80994
8.914 0.98815 5.4612e-005 3.8183 0.011912 0.00011577 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6186 0.5994 0.18304 0.020822 18.8667 0.1289 0.0001691 0.76127 0.0096107 0.010623 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16646 0.93449 0.91637 0.0013972 0.99247 0.48772 0.0018824 0.4256 2.2203 2.2197 16.0158 144.9122 0.00016333 -85.6511 0.81094
8.915 0.98815 5.4612e-005 3.8183 0.011912 0.00011579 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6187 0.59945 0.18305 0.020823 18.8699 0.1289 0.00016911 0.76127 0.009611 0.010623 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16646 0.93464 0.91643 0.0013972 0.9925 0.4879 0.0018823 0.42562 2.2207 2.2201 16.0157 144.9122 0.00016324 -85.6511 0.81194
8.916 0.98815 5.4612e-005 3.8183 0.011912 0.0001158 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6188 0.59949 0.18306 0.020824 18.8732 0.12891 0.00016912 0.76126 0.0096114 0.010624 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16646 0.93479 0.91649 0.0013972 0.99253 0.48808 0.0018823 0.42563 2.2212 2.2206 16.0157 144.9122 0.00016315 -85.6512 0.81294
8.917 0.98815 5.4612e-005 3.8183 0.011912 0.00011581 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6188 0.59953 0.18308 0.020825 18.8764 0.12892 0.00016912 0.76125 0.0096117 0.010624 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16646 0.93495 0.91655 0.0013972 0.99256 0.48826 0.0018823 0.42564 2.2216 2.221 16.0157 144.9123 0.00016306 -85.6513 0.81394
8.918 0.98815 5.4612e-005 3.8183 0.011912 0.00011582 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6189 0.59958 0.18309 0.020826 18.8797 0.12892 0.00016913 0.76125 0.009612 0.010624 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.16647 0.9351 0.91661 0.0013971 0.99259 0.48843 0.0018823 0.42566 2.2221 2.2215 16.0156 144.9123 0.00016297 -85.6514 0.81494
8.919 0.98815 5.4612e-005 3.8183 0.011912 0.00011584 0.0011766 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.619 0.59962 0.1831 0.020827 18.8829 0.12893 0.00016914 0.76124 0.0096124 0.010625 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.16647 0.93525 0.91667 0.0013971 0.99262 0.48861 0.0018823 0.42567 2.2225 2.2219 16.0156 144.9123 0.00016288 -85.6515 0.81594
8.92 0.98815 5.4612e-005 3.8183 0.011911 0.00011585 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6191 0.59967 0.18312 0.020828 18.8862 0.12893 0.00016915 0.76124 0.0096127 0.010625 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16647 0.9354 0.91673 0.0013971 0.99265 0.48879 0.0018823 0.42569 2.223 2.2224 16.0156 144.9123 0.00016279 -85.6516 0.81694
8.921 0.98815 5.4611e-005 3.8183 0.011911 0.00011586 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6192 0.59971 0.18313 0.020829 18.8894 0.12894 0.00016916 0.76123 0.0096131 0.010625 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.16647 0.93555 0.91679 0.0013971 0.99268 0.48897 0.0018823 0.4257 2.2234 2.2228 16.0155 144.9123 0.0001627 -85.6517 0.81794
8.922 0.98815 5.4611e-005 3.8183 0.011911 0.00011587 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6193 0.59976 0.18314 0.02083 18.8927 0.12895 0.00016917 0.76122 0.0096134 0.010626 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16648 0.9357 0.91685 0.0013971 0.99271 0.48915 0.0018822 0.42571 2.2239 2.2233 16.0155 144.9124 0.00016261 -85.6518 0.81894
8.923 0.98815 5.4611e-005 3.8183 0.011911 0.00011589 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6193 0.5998 0.18316 0.020831 18.8959 0.12895 0.00016918 0.76122 0.0096138 0.010626 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16648 0.93585 0.9169 0.0013971 0.99274 0.48932 0.0018822 0.42573 2.2243 2.2237 16.0155 144.9124 0.00016252 -85.6519 0.81994
8.924 0.98815 5.4611e-005 3.8183 0.011911 0.0001159 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6194 0.59984 0.18317 0.020832 18.8992 0.12896 0.00016919 0.76121 0.0096141 0.010626 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.16648 0.936 0.91696 0.0013971 0.99277 0.4895 0.0018822 0.42574 2.2248 2.2242 16.0155 144.9124 0.00016243 -85.6519 0.82094
8.925 0.98815 5.4611e-005 3.8183 0.011911 0.00011591 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6195 0.59989 0.18318 0.020833 18.9024 0.12896 0.0001692 0.76121 0.0096144 0.010627 0.0013862 0.98694 0.9917 2.9891e-006 1.1956e-005 0.16648 0.93615 0.91702 0.0013971 0.9928 0.48968 0.0018822 0.42576 2.2252 2.2246 16.0154 144.9124 0.00016234 -85.652 0.82194
8.926 0.98815 5.4611e-005 3.8183 0.011911 0.00011593 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6196 0.59993 0.18319 0.020834 18.9057 0.12897 0.00016921 0.7612 0.0096148 0.010627 0.0013862 0.98694 0.99171 2.9891e-006 1.1956e-005 0.16649 0.9363 0.91708 0.0013971 0.99283 0.48986 0.0018822 0.42577 2.2257 2.2251 16.0154 144.9124 0.00016225 -85.6521 0.82294
8.927 0.98815 5.4611e-005 3.8183 0.011911 0.00011594 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6197 0.59998 0.18321 0.020835 18.9089 0.12898 0.00016922 0.76119 0.0096151 0.010628 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16649 0.93644 0.91713 0.001397 0.99286 0.49004 0.0018822 0.42578 2.2261 2.2255 16.0154 144.9125 0.00016216 -85.6522 0.82394
8.928 0.98815 5.4611e-005 3.8183 0.011911 0.00011595 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6198 0.60002 0.18322 0.020836 18.9122 0.12898 0.00016923 0.76119 0.0096155 0.010628 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16649 0.93659 0.91719 0.001397 0.99288 0.49021 0.0018822 0.4258 2.2266 2.226 16.0153 144.9125 0.00016208 -85.6523 0.82494
8.929 0.98815 5.4611e-005 3.8183 0.011911 0.00011596 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6198 0.60007 0.18323 0.020837 18.9154 0.12899 0.00016924 0.76118 0.0096158 0.010628 0.0013862 0.98695 0.99171 2.9889e-006 1.1956e-005 0.1665 0.93674 0.91725 0.001397 0.99291 0.49039 0.0018821 0.42581 2.227 2.2264 16.0153 144.9125 0.00016199 -85.6524 0.82594
8.93 0.98815 5.4611e-005 3.8183 0.011911 0.00011598 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6199 0.60011 0.18325 0.020838 18.9187 0.12899 0.00016924 0.76117 0.0096161 0.010629 0.0013862 0.98695 0.99171 2.9889e-006 1.1955e-005 0.1665 0.93688 0.9173 0.001397 0.99294 0.49057 0.0018821 0.42583 2.2274 2.2269 16.0153 144.9125 0.0001619 -85.6524 0.82694
8.931 0.98815 5.4611e-005 3.8183 0.011911 0.00011599 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.62 0.60015 0.18326 0.020839 18.9219 0.129 0.00016925 0.76117 0.0096165 0.010629 0.0013861 0.98695 0.99171 2.9889e-006 1.1955e-005 0.1665 0.93703 0.91736 0.001397 0.99297 0.49075 0.0018821 0.42584 2.2279 2.2273 16.0152 144.9125 0.00016182 -85.6525 0.82794
8.932 0.98815 5.4611e-005 3.8183 0.011911 0.000116 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6201 0.6002 0.18327 0.02084 18.9252 0.12901 0.00016926 0.76116 0.0096168 0.010629 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.1665 0.93718 0.91742 0.001397 0.99299 0.49092 0.0018821 0.42585 2.2283 2.2277 16.0152 144.9126 0.00016173 -85.6526 0.82894
8.933 0.98815 5.461e-005 3.8183 0.011911 0.00011602 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6202 0.60024 0.18329 0.020841 18.9284 0.12901 0.00016927 0.76116 0.0096172 0.01063 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16651 0.93732 0.91747 0.001397 0.99302 0.4911 0.0018821 0.42587 2.2288 2.2282 16.0152 144.9126 0.00016164 -85.6527 0.82994
8.934 0.98815 5.461e-005 3.8183 0.011911 0.00011603 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6203 0.60029 0.1833 0.020842 18.9317 0.12902 0.00016928 0.76115 0.0096175 0.01063 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16651 0.93746 0.91753 0.001397 0.99305 0.49128 0.0018821 0.42588 2.2292 2.2286 16.0152 144.9126 0.00016156 -85.6528 0.83094
8.935 0.98815 5.461e-005 3.8183 0.011911 0.00011604 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6203 0.60033 0.18331 0.020843 18.9349 0.12902 0.00016929 0.76114 0.0096178 0.01063 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16651 0.93761 0.91758 0.001397 0.99308 0.49146 0.0018821 0.4259 2.2296 2.2291 16.0151 144.9126 0.00016147 -85.6528 0.83194
8.936 0.98815 5.461e-005 3.8183 0.011911 0.00011605 0.0011767 0.23361 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6204 0.60038 0.18332 0.020844 18.9382 0.12903 0.0001693 0.76114 0.0096182 0.010631 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16651 0.93775 0.91764 0.001397 0.9931 0.49163 0.0018821 0.42591 2.2301 2.2295 16.0151 144.9126 0.00016139 -85.6529 0.83294
8.937 0.98815 5.461e-005 3.8183 0.011911 0.00011607 0.0011767 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6205 0.60042 0.18334 0.020845 18.9414 0.12904 0.00016931 0.76113 0.0096185 0.010631 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16652 0.9379 0.9177 0.001397 0.99313 0.49181 0.001882 0.42592 2.2305 2.2299 16.0151 144.9127 0.0001613 -85.653 0.83394
8.938 0.98815 5.461e-005 3.8183 0.011911 0.00011608 0.0011767 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6206 0.60046 0.18335 0.020846 18.9447 0.12904 0.00016932 0.76113 0.0096189 0.010632 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16652 0.93804 0.91775 0.0013969 0.99315 0.49199 0.001882 0.42594 2.2309 2.2304 16.015 144.9127 0.00016122 -85.6531 0.83494
8.939 0.98815 5.461e-005 3.8183 0.011911 0.00011609 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6207 0.60051 0.18336 0.020847 18.9479 0.12905 0.00016933 0.76112 0.0096192 0.010632 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16652 0.93818 0.91781 0.0013969 0.99318 0.49216 0.001882 0.42595 2.2314 2.2308 16.015 144.9127 0.00016113 -85.6531 0.83594
8.94 0.98815 5.461e-005 3.8183 0.011911 0.0001161 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6208 0.60055 0.18338 0.020848 18.9512 0.12905 0.00016934 0.76111 0.0096196 0.010632 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16652 0.93832 0.91786 0.0013969 0.99321 0.49234 0.001882 0.42597 2.2318 2.2312 16.015 144.9127 0.00016105 -85.6532 0.83694
8.941 0.98815 5.461e-005 3.8183 0.011911 0.00011612 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6208 0.6006 0.18339 0.020849 18.9544 0.12906 0.00016935 0.76111 0.0096199 0.010633 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.16653 0.93846 0.91791 0.0013969 0.99323 0.49252 0.001882 0.42598 2.2322 2.2317 16.0149 144.9127 0.00016096 -85.6533 0.83794
8.942 0.98815 5.461e-005 3.8183 0.011911 0.00011613 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6209 0.60064 0.1834 0.02085 18.9577 0.12907 0.00016936 0.7611 0.0096202 0.010633 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.16653 0.9386 0.91797 0.0013969 0.99326 0.4927 0.001882 0.42599 2.2327 2.2321 16.0149 144.9128 0.00016088 -85.6534 0.83894
8.943 0.98815 5.461e-005 3.8183 0.011911 0.00011614 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.621 0.60069 0.18342 0.020851 18.9609 0.12907 0.00016936 0.7611 0.0096206 0.010633 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.16653 0.93874 0.91802 0.0013969 0.99328 0.49287 0.001882 0.42601 2.2331 2.2325 16.0149 144.9128 0.0001608 -85.6534 0.83994
8.944 0.98815 5.4609e-005 3.8183 0.011911 0.00011616 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6211 0.60073 0.18343 0.020852 18.9642 0.12908 0.00016937 0.76109 0.0096209 0.010634 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16653 0.93888 0.91808 0.0013969 0.99331 0.49305 0.001882 0.42602 2.2335 2.233 16.0148 144.9128 0.00016071 -85.6535 0.84094
8.945 0.98815 5.4609e-005 3.8183 0.011911 0.00011617 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6212 0.60077 0.18344 0.020853 18.9674 0.12908 0.00016938 0.76108 0.0096213 0.010634 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16654 0.93902 0.91813 0.0013969 0.99333 0.49323 0.0018819 0.42604 2.2339 2.2334 16.0148 144.9128 0.00016063 -85.6536 0.84194
8.946 0.98815 5.4609e-005 3.8183 0.011911 0.00011618 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6213 0.60082 0.18345 0.020854 18.9707 0.12909 0.00016939 0.76108 0.0096216 0.010634 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16654 0.93916 0.91818 0.0013969 0.99336 0.4934 0.0018819 0.42605 2.2344 2.2338 16.0148 144.9128 0.00016055 -85.6537 0.84294
8.947 0.98815 5.4609e-005 3.8183 0.011911 0.00011619 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6213 0.60086 0.18347 0.020855 18.974 0.1291 0.0001694 0.76107 0.0096219 0.010635 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16654 0.9393 0.91824 0.0013969 0.99338 0.49358 0.0018819 0.42606 2.2348 2.2342 16.0147 144.9129 0.00016047 -85.6537 0.84394
8.948 0.98815 5.4609e-005 3.8183 0.011911 0.00011621 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6214 0.60091 0.18348 0.020856 18.9772 0.1291 0.00016941 0.76107 0.0096223 0.010635 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16654 0.93944 0.91829 0.0013969 0.99341 0.49376 0.0018819 0.42608 2.2352 2.2347 16.0147 144.9129 0.00016038 -85.6538 0.84494
8.949 0.98815 5.4609e-005 3.8183 0.011911 0.00011622 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6215 0.60095 0.18349 0.020857 18.9805 0.12911 0.00016942 0.76106 0.0096226 0.010635 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16655 0.93958 0.91834 0.0013968 0.99343 0.49393 0.0018819 0.42609 2.2357 2.2351 16.0147 144.9129 0.0001603 -85.6539 0.84594
8.95 0.98815 5.4609e-005 3.8183 0.011911 0.00011623 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6216 0.601 0.18351 0.020858 18.9837 0.12911 0.00016943 0.76105 0.009623 0.010636 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16655 0.93972 0.9184 0.0013968 0.99346 0.49411 0.0018819 0.42611 2.2361 2.2355 16.0147 144.9129 0.00016022 -85.6539 0.84694
8.951 0.98815 5.4609e-005 3.8183 0.011911 0.00011625 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6217 0.60104 0.18352 0.020859 18.987 0.12912 0.00016944 0.76105 0.0096233 0.010636 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16655 0.93985 0.91845 0.0013968 0.99348 0.49428 0.0018819 0.42612 2.2365 2.2359 16.0146 144.913 0.00016014 -85.654 0.84794
8.952 0.98815 5.4609e-005 3.8183 0.011911 0.00011626 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6218 0.60108 0.18353 0.02086 18.9902 0.12913 0.00016945 0.76104 0.0096236 0.010637 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16656 0.93999 0.9185 0.0013968 0.99351 0.49446 0.0018819 0.42613 2.2369 2.2364 16.0146 144.913 0.00016006 -85.6541 0.84894
8.953 0.98815 5.4609e-005 3.8183 0.011911 0.00011627 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6218 0.60113 0.18354 0.020861 18.9935 0.12913 0.00016946 0.76104 0.009624 0.010637 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16656 0.94012 0.91855 0.0013968 0.99353 0.49464 0.0018819 0.42615 2.2373 2.2368 16.0146 144.913 0.00015998 -85.6541 0.84994
8.954 0.98815 5.4609e-005 3.8183 0.011911 0.00011628 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.6219 0.60117 0.18356 0.020862 18.9968 0.12914 0.00016947 0.76103 0.0096243 0.010637 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16656 0.94026 0.91861 0.0013968 0.99355 0.49481 0.0018818 0.42616 2.2378 2.2372 16.0145 144.913 0.0001599 -85.6542 0.85094
8.955 0.98815 5.4609e-005 3.8183 0.011911 0.0001163 0.0011768 0.2336 0.00065931 0.23426 0.21617 0 0.032264 0.0389 0 1.622 0.60122 0.18357 0.020863 19 0.12914 0.00016948 0.76102 0.0096247 0.010638 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.16656 0.9404 0.91866 0.0013968 0.99358 0.49499 0.0018818 0.42618 2.2382 2.2376 16.0145 144.913 0.00015982 -85.6543 0.85194
8.956 0.98815 5.4608e-005 3.8183 0.011911 0.00011631 0.0011768 0.2336 0.00065931 0.23426 0.21616 0 0.032264 0.0389 0 1.6221 0.60126 0.18358 0.020864 19.0033 0.12915 0.00016948 0.76102 0.009625 0.010638 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.16657 0.94053 0.91871 0.0013968 0.9936 0.49516 0.0018818 0.42619 2.2386 2.2381 16.0145 144.9131 0.00015974 -85.6543 0.85294
8.957 0.98815 5.4608e-005 3.8183 0.011911 0.00011632 0.0011768 0.2336 0.00065931 0.23426 0.21616 0 0.032264 0.0389 0 1.6222 0.6013 0.1836 0.020865 19.0065 0.12916 0.00016949 0.76101 0.0096253 0.010638 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16657 0.94066 0.91876 0.0013968 0.99362 0.49534 0.0018818 0.4262 2.239 2.2385 16.0144 144.9131 0.00015966 -85.6544 0.85394
8.958 0.98815 5.4608e-005 3.8183 0.011911 0.00011633 0.0011769 0.2336 0.00065931 0.23426 0.21616 0 0.032264 0.0389 0 1.6223 0.60135 0.18361 0.020866 19.0098 0.12916 0.0001695 0.76101 0.0096257 0.010639 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16657 0.9408 0.91881 0.0013968 0.99365 0.49552 0.0018818 0.42622 2.2394 2.2389 16.0144 144.9131 0.00015958 -85.6545 0.85494
8.959 0.98815 5.4608e-005 3.8183 0.011911 0.00011635 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6223 0.60139 0.18362 0.020867 19.013 0.12917 0.00016951 0.761 0.009626 0.010639 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16657 0.94093 0.91886 0.0013968 0.99367 0.49569 0.0018818 0.42623 2.2399 2.2393 16.0144 144.9131 0.0001595 -85.6545 0.85594
8.96 0.98815 5.4608e-005 3.8183 0.011911 0.00011636 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6224 0.60144 0.18364 0.020868 19.0163 0.12917 0.00016952 0.76099 0.0096264 0.010639 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16658 0.94107 0.91891 0.0013968 0.99369 0.49587 0.0018818 0.42624 2.2403 2.2397 16.0143 144.9131 0.00015942 -85.6546 0.85694
8.961 0.98815 5.4608e-005 3.8183 0.011911 0.00011637 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6225 0.60148 0.18365 0.020869 19.0196 0.12918 0.00016953 0.76099 0.0096267 0.01064 0.0013857 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16658 0.9412 0.91896 0.0013967 0.99371 0.49604 0.0018818 0.42626 2.2407 2.2401 16.0143 144.9132 0.00015935 -85.6547 0.85794
8.962 0.98815 5.4608e-005 3.8183 0.011911 0.00011639 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6226 0.60153 0.18366 0.02087 19.0228 0.12919 0.00016954 0.76098 0.009627 0.01064 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16658 0.94133 0.91902 0.0013967 0.99374 0.49622 0.0018818 0.42627 2.2411 2.2406 16.0143 144.9132 0.00015927 -85.6547 0.85894
8.963 0.98815 5.4608e-005 3.8183 0.011911 0.0001164 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6227 0.60157 0.18367 0.020871 19.0261 0.12919 0.00016955 0.76098 0.0096274 0.010641 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16658 0.94146 0.91907 0.0013967 0.99376 0.49639 0.0018818 0.42629 2.2415 2.241 16.0142 144.9132 0.00015919 -85.6548 0.85994
8.964 0.98815 5.4608e-005 3.8183 0.011911 0.00011641 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6228 0.60161 0.18369 0.020872 19.0293 0.1292 0.00016956 0.76097 0.0096277 0.010641 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16659 0.94159 0.91912 0.0013967 0.99378 0.49657 0.0018817 0.4263 2.2419 2.2414 16.0142 144.9132 0.00015911 -85.6549 0.86094
8.965 0.98815 5.4608e-005 3.8183 0.011911 0.00011642 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6228 0.60166 0.1837 0.020873 19.0326 0.1292 0.00016957 0.76096 0.009628 0.010641 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16659 0.94173 0.91917 0.0013967 0.9938 0.49675 0.0018817 0.42631 2.2423 2.2418 16.0142 144.9132 0.00015904 -85.6549 0.86194
8.966 0.98815 5.4608e-005 3.8183 0.011911 0.00011644 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6229 0.6017 0.18371 0.020874 19.0359 0.12921 0.00016958 0.76096 0.0096284 0.010642 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.16659 0.94186 0.91922 0.0013967 0.99383 0.49692 0.0018817 0.42633 2.2428 2.2422 16.0142 144.9133 0.00015896 -85.655 0.86294
8.967 0.98815 5.4608e-005 3.8183 0.011911 0.00011645 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.623 0.60175 0.18373 0.020875 19.0391 0.12922 0.00016959 0.76095 0.0096287 0.010642 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.16659 0.94199 0.91927 0.0013967 0.99385 0.4971 0.0018817 0.42634 2.2432 2.2426 16.0141 144.9133 0.00015888 -85.655 0.86394
8.968 0.98815 5.4607e-005 3.8183 0.011911 0.00011646 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6231 0.60179 0.18374 0.020876 19.0424 0.12922 0.0001696 0.76095 0.0096291 0.010642 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.1666 0.94212 0.91932 0.0013967 0.99387 0.49727 0.0018817 0.42636 2.2436 2.243 16.0141 144.9133 0.00015881 -85.6551 0.86494
8.969 0.98815 5.4607e-005 3.8183 0.011911 0.00011648 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6232 0.60184 0.18375 0.020877 19.0457 0.12923 0.0001696 0.76094 0.0096294 0.010643 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.1666 0.94225 0.91936 0.0013967 0.99389 0.49745 0.0018817 0.42637 2.244 2.2434 16.0141 144.9133 0.00015873 -85.6552 0.86594
8.97 0.98815 5.4607e-005 3.8183 0.011911 0.00011649 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6233 0.60188 0.18377 0.020878 19.0489 0.12923 0.00016961 0.76094 0.0096297 0.010643 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.1666 0.94237 0.91941 0.0013967 0.99391 0.49762 0.0018817 0.42638 2.2444 2.2439 16.014 144.9133 0.00015865 -85.6552 0.86694
8.971 0.98815 5.4607e-005 3.8183 0.011911 0.0001165 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6233 0.60192 0.18378 0.020879 19.0522 0.12924 0.00016962 0.76093 0.0096301 0.010643 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.1666 0.9425 0.91946 0.0013967 0.99393 0.4978 0.0018817 0.4264 2.2448 2.2443 16.014 144.9134 0.00015858 -85.6553 0.86794
8.972 0.98815 5.4607e-005 3.8183 0.011911 0.00011651 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6234 0.60197 0.18379 0.02088 19.0554 0.12925 0.00016963 0.76092 0.0096304 0.010644 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.16661 0.94263 0.91951 0.0013967 0.99395 0.49797 0.0018817 0.42641 2.2452 2.2447 16.014 144.9134 0.0001585 -85.6553 0.86894
8.973 0.98815 5.4607e-005 3.8183 0.011911 0.00011653 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6235 0.60201 0.1838 0.020881 19.0587 0.12925 0.00016964 0.76092 0.0096308 0.010644 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16661 0.94276 0.91956 0.0013967 0.99398 0.49815 0.0018817 0.42642 2.2456 2.2451 16.0139 144.9134 0.00015843 -85.6554 0.86994
8.974 0.98815 5.4607e-005 3.8183 0.011911 0.00011654 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6236 0.60206 0.18382 0.020882 19.062 0.12926 0.00016965 0.76091 0.0096311 0.010644 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16661 0.94289 0.91961 0.0013967 0.994 0.49832 0.0018817 0.42644 2.246 2.2455 16.0139 144.9134 0.00015835 -85.6554 0.87094
8.975 0.98815 5.4607e-005 3.8183 0.011911 0.00011655 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6237 0.6021 0.18383 0.020883 19.0652 0.12926 0.00016966 0.76091 0.0096314 0.010645 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16661 0.94301 0.91966 0.0013966 0.99402 0.4985 0.0018816 0.42645 2.2464 2.2459 16.0139 144.9134 0.00015828 -85.6555 0.87194
8.976 0.98815 5.4607e-005 3.8183 0.01191 0.00011656 0.0011769 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6238 0.60215 0.18384 0.020885 19.0685 0.12927 0.00016967 0.7609 0.0096318 0.010645 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16662 0.94314 0.91971 0.0013966 0.99404 0.49867 0.0018816 0.42647 2.2468 2.2463 16.0138 144.9135 0.00015821 -85.6556 0.87294
8.977 0.98815 5.4607e-005 3.8183 0.01191 0.00011658 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6238 0.60219 0.18386 0.020886 19.0718 0.12928 0.00016968 0.76089 0.0096321 0.010646 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16662 0.94327 0.91975 0.0013966 0.99406 0.49885 0.0018816 0.42648 2.2472 2.2467 16.0138 144.9135 0.00015813 -85.6556 0.87394
8.978 0.98815 5.4607e-005 3.8183 0.01191 0.00011659 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6239 0.60223 0.18387 0.020887 19.075 0.12928 0.00016969 0.76089 0.0096325 0.010646 0.0013854 0.98696 0.99171 2.9872e-006 1.1949e-005 0.16662 0.94339 0.9198 0.0013966 0.99408 0.49902 0.0018816 0.42649 2.2476 2.2471 16.0138 144.9135 0.00015806 -85.6557 0.87494
8.979 0.98815 5.4607e-005 3.8183 0.01191 0.0001166 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.624 0.60228 0.18388 0.020888 19.0783 0.12929 0.0001697 0.76088 0.0096328 0.010646 0.0013854 0.98696 0.99171 2.9872e-006 1.1949e-005 0.16663 0.94352 0.91985 0.0013966 0.9941 0.4992 0.0018816 0.42651 2.248 2.2475 16.0137 144.9135 0.00015798 -85.6557 0.87594
8.98 0.98815 5.4606e-005 3.8183 0.01191 0.00011662 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6241 0.60232 0.18389 0.020889 19.0816 0.12929 0.00016971 0.76088 0.0096331 0.010647 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16663 0.94364 0.9199 0.0013966 0.99412 0.49937 0.0018816 0.42652 2.2484 2.2479 16.0137 144.9136 0.00015791 -85.6558 0.87694
8.981 0.98815 5.4606e-005 3.8183 0.01191 0.00011663 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6242 0.60237 0.18391 0.02089 19.0848 0.1293 0.00016971 0.76087 0.0096335 0.010647 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16663 0.94377 0.91994 0.0013966 0.99414 0.49954 0.0018816 0.42653 2.2488 2.2483 16.0137 144.9136 0.00015784 -85.6558 0.87794
8.982 0.98815 5.4606e-005 3.8183 0.01191 0.00011664 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6242 0.60241 0.18392 0.020891 19.0881 0.12931 0.00016972 0.76086 0.0096338 0.010647 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16663 0.94389 0.91999 0.0013966 0.99416 0.49972 0.0018816 0.42655 2.2492 2.2487 16.0136 144.9136 0.00015777 -85.6559 0.87894
8.983 0.98815 5.4606e-005 3.8183 0.01191 0.00011665 0.001177 0.2336 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6243 0.60246 0.18393 0.020892 19.0914 0.12931 0.00016973 0.76086 0.0096341 0.010648 0.0013854 0.98696 0.99171 2.987e-006 1.1948e-005 0.16664 0.94402 0.92004 0.0013966 0.99418 0.49989 0.0018816 0.42656 2.2496 2.2491 16.0136 144.9136 0.00015769 -85.6559 0.87994
8.984 0.98815 5.4606e-005 3.8183 0.01191 0.00011667 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6244 0.6025 0.18395 0.020893 19.0946 0.12932 0.00016974 0.76085 0.0096345 0.010648 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16664 0.94414 0.92009 0.0013966 0.9942 0.50007 0.0018816 0.42658 2.25 2.2495 16.0136 144.9136 0.00015762 -85.656 0.88094
8.985 0.98815 5.4606e-005 3.8183 0.01191 0.00011668 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6245 0.60254 0.18396 0.020894 19.0979 0.12932 0.00016975 0.76085 0.0096348 0.010648 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16664 0.94426 0.92013 0.0013966 0.99422 0.50024 0.0018816 0.42659 2.2504 2.2499 16.0135 144.9137 0.00015755 -85.656 0.88194
8.986 0.98815 5.4606e-005 3.8183 0.01191 0.00011669 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6246 0.60259 0.18397 0.020895 19.1012 0.12933 0.00016976 0.76084 0.0096352 0.010649 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16664 0.94439 0.92018 0.0013966 0.99424 0.50042 0.0018815 0.4266 2.2508 2.2503 16.0135 144.9137 0.00015748 -85.6561 0.88294
8.987 0.98815 5.4606e-005 3.8183 0.01191 0.00011671 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6247 0.60263 0.18399 0.020896 19.1044 0.12934 0.00016977 0.76083 0.0096355 0.010649 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16665 0.94451 0.92022 0.0013966 0.99425 0.50059 0.0018815 0.42662 2.2512 2.2507 16.0135 144.9137 0.00015741 -85.6562 0.88394
8.988 0.98815 5.4606e-005 3.8183 0.01191 0.00011672 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6247 0.60268 0.184 0.020897 19.1077 0.12934 0.00016978 0.76083 0.0096358 0.010649 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16665 0.94463 0.92027 0.0013966 0.99427 0.50076 0.0018815 0.42663 2.2516 2.2511 16.0134 144.9137 0.00015733 -85.6562 0.88494
8.989 0.98815 5.4606e-005 3.8183 0.01191 0.00011673 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6248 0.60272 0.18401 0.020898 19.111 0.12935 0.00016979 0.76082 0.0096362 0.01065 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16665 0.94475 0.92032 0.0013966 0.99429 0.50094 0.0018815 0.42664 2.252 2.2515 16.0134 144.9137 0.00015726 -85.6563 0.88594
8.99 0.98815 5.4606e-005 3.8183 0.01191 0.00011674 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6249 0.60277 0.18402 0.020899 19.1142 0.12935 0.0001698 0.76082 0.0096365 0.01065 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16665 0.94487 0.92036 0.0013965 0.99431 0.50111 0.0018815 0.42666 2.2524 2.2519 16.0134 144.9138 0.00015719 -85.6563 0.88694
8.991 0.98815 5.4606e-005 3.8183 0.01191 0.00011676 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.625 0.60281 0.18404 0.0209 19.1175 0.12936 0.00016981 0.76081 0.0096369 0.010651 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16666 0.94499 0.92041 0.0013965 0.99433 0.50129 0.0018815 0.42667 2.2528 2.2523 16.0134 144.9138 0.00015712 -85.6564 0.88794
8.992 0.98815 5.4605e-005 3.8183 0.01191 0.00011677 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6251 0.60285 0.18405 0.020901 19.1208 0.12937 0.00016982 0.7608 0.0096372 0.010651 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16666 0.94511 0.92045 0.0013965 0.99435 0.50146 0.0018815 0.42669 2.2532 2.2527 16.0133 144.9138 0.00015705 -85.6564 0.88894
8.993 0.98815 5.4605e-005 3.8183 0.01191 0.00011678 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6252 0.6029 0.18406 0.020902 19.1241 0.12937 0.00016983 0.7608 0.0096375 0.010651 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16666 0.94523 0.9205 0.0013965 0.99437 0.50163 0.0018815 0.4267 2.2536 2.2531 16.0133 144.9138 0.00015698 -85.6564 0.88994
8.994 0.98815 5.4605e-005 3.8183 0.01191 0.00011679 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032264 0.0389 0 1.6252 0.60294 0.18408 0.020903 19.1273 0.12938 0.00016983 0.76079 0.0096379 0.010652 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16666 0.94535 0.92055 0.0013965 0.99438 0.50181 0.0018815 0.42671 2.254 2.2535 16.0133 144.9138 0.00015691 -85.6565 0.89094
8.995 0.98815 5.4605e-005 3.8183 0.01191 0.00011681 0.001177 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6253 0.60299 0.18409 0.020904 19.1306 0.12938 0.00016984 0.76079 0.0096382 0.010652 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16667 0.94547 0.92059 0.0013965 0.9944 0.50198 0.0018815 0.42673 2.2544 2.2538 16.0132 144.9139 0.00015684 -85.6565 0.89194
8.996 0.98815 5.4605e-005 3.8183 0.01191 0.00011682 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6254 0.60303 0.1841 0.020905 19.1339 0.12939 0.00016985 0.76078 0.0096385 0.010652 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16667 0.94559 0.92064 0.0013965 0.99442 0.50215 0.0018815 0.42674 2.2547 2.2542 16.0132 144.9139 0.00015677 -85.6566 0.89294
8.997 0.98815 5.4605e-005 3.8183 0.01191 0.00011683 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6255 0.60307 0.18411 0.020906 19.1371 0.1294 0.00016986 0.76077 0.0096389 0.010653 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16667 0.94571 0.92068 0.0013965 0.99444 0.50233 0.0018815 0.42675 2.2551 2.2546 16.0132 144.9139 0.0001567 -85.6566 0.89394
8.998 0.98815 5.4605e-005 3.8183 0.01191 0.00011685 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6256 0.60312 0.18413 0.020907 19.1404 0.1294 0.00016987 0.76077 0.0096392 0.010653 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16667 0.94583 0.92072 0.0013965 0.99446 0.5025 0.0018815 0.42677 2.2555 2.255 16.0131 144.9139 0.00015663 -85.6567 0.89494
8.999 0.98815 5.4605e-005 3.8183 0.01191 0.00011686 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6257 0.60316 0.18414 0.020908 19.1437 0.12941 0.00016988 0.76076 0.0096396 0.010653 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16668 0.94595 0.92077 0.0013965 0.99447 0.50267 0.0018814 0.42678 2.2559 2.2554 16.0131 144.9139 0.00015657 -85.6567 0.89594
9 0.98815 5.4605e-005 3.8183 0.01191 0.00011687 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6257 0.60321 0.18415 0.020909 19.147 0.12941 0.00016989 0.76076 0.0096399 0.010654 0.0013852 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16668 0.94606 0.92081 0.0013965 0.99449 0.50285 0.0018814 0.42679 2.2563 2.2558 16.0131 144.914 0.0001565 -85.6568 0.89694
9.001 0.98815 5.4605e-005 3.8183 0.01191 0.00011688 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6258 0.60325 0.18417 0.02091 19.1502 0.12942 0.0001699 0.76075 0.0096402 0.010654 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16668 0.94618 0.92086 0.0013965 0.99451 0.50302 0.0018814 0.42681 2.2567 2.2562 16.013 144.914 0.00015643 -85.6568 0.89794
9.002 0.98815 5.4605e-005 3.8183 0.01191 0.0001169 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6259 0.6033 0.18418 0.020911 19.1535 0.12943 0.00016991 0.76074 0.0096406 0.010654 0.0013851 0.98696 0.99171 2.9866e-006 1.1946e-005 0.16668 0.9463 0.9209 0.0013965 0.99453 0.50319 0.0018814 0.42682 2.2571 2.2566 16.013 144.914 0.00015636 -85.6569 0.89894
9.003 0.98815 5.4605e-005 3.8183 0.01191 0.00011691 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.626 0.60334 0.18419 0.020912 19.1568 0.12943 0.00016992 0.76074 0.0096409 0.010655 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16669 0.94641 0.92095 0.0013965 0.99454 0.50337 0.0018814 0.42683 2.2574 2.2569 16.013 144.914 0.00015629 -85.6569 0.89994
9.004 0.98815 5.4604e-005 3.8183 0.01191 0.00011692 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6261 0.60338 0.18421 0.020913 19.1601 0.12944 0.00016993 0.76073 0.0096412 0.010655 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16669 0.94653 0.92099 0.0013965 0.99456 0.50354 0.0018814 0.42685 2.2578 2.2573 16.0129 144.914 0.00015623 -85.657 0.90094
9.005 0.98815 5.4604e-005 3.8183 0.01191 0.00011694 0.0011771 0.23359 0.00065931 0.23425 0.21616 0 0.032265 0.0389 0 1.6262 0.60343 0.18422 0.020914 19.1633 0.12944 0.00016994 0.76073 0.0096416 0.010656 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.16669 0.94665 0.92103 0.0013965 0.99458 0.50371 0.0018814 0.42686 2.2582 2.2577 16.0129 144.9141 0.00015616 -85.657 0.90194
9.006 0.98815 5.4604e-005 3.8183 0.01191 0.00011695 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6262 0.60347 0.18423 0.020915 19.1666 0.12945 0.00016994 0.76072 0.0096419 0.010656 0.0013851 0.98696 0.99171 2.9865e-006 1.1946e-005 0.1667 0.94676 0.92108 0.0013965 0.99459 0.50389 0.0018814 0.42688 2.2586 2.2581 16.0129 144.9141 0.00015609 -85.657 0.90294
9.007 0.98815 5.4604e-005 3.8183 0.01191 0.00011696 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6263 0.60352 0.18424 0.020916 19.1699 0.12946 0.00016995 0.76071 0.0096423 0.010656 0.0013851 0.98696 0.99171 2.9864e-006 1.1946e-005 0.1667 0.94688 0.92112 0.0013965 0.99461 0.50406 0.0018814 0.42689 2.259 2.2585 16.0128 144.9141 0.00015603 -85.6571 0.90394
9.008 0.98815 5.4604e-005 3.8183 0.01191 0.00011697 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6264 0.60356 0.18426 0.020917 19.1731 0.12946 0.00016996 0.76071 0.0096426 0.010657 0.001385 0.98696 0.99171 2.9864e-006 1.1946e-005 0.1667 0.94699 0.92116 0.0013964 0.99463 0.50423 0.0018814 0.4269 2.2594 2.2589 16.0128 144.9141 0.00015596 -85.6571 0.90494
9.009 0.98815 5.4604e-005 3.8183 0.01191 0.00011699 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6265 0.60361 0.18427 0.020918 19.1764 0.12947 0.00016997 0.7607 0.0096429 0.010657 0.001385 0.98696 0.99172 2.9864e-006 1.1945e-005 0.1667 0.9471 0.92121 0.0013964 0.99464 0.5044 0.0018814 0.42692 2.2597 2.2592 16.0128 144.9141 0.00015589 -85.6572 0.90594
9.01 0.98815 5.4604e-005 3.8183 0.01191 0.000117 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6266 0.60365 0.18428 0.020919 19.1797 0.12947 0.00016998 0.7607 0.0096433 0.010657 0.001385 0.98696 0.99172 2.9864e-006 1.1945e-005 0.16671 0.94722 0.92125 0.0013964 0.99466 0.50458 0.0018814 0.42693 2.2601 2.2596 16.0127 144.9142 0.00015583 -85.6572 0.90694
9.011 0.98815 5.4604e-005 3.8183 0.01191 0.00011701 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6267 0.60369 0.1843 0.02092 19.183 0.12948 0.00016999 0.76069 0.0096436 0.010658 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16671 0.94733 0.92129 0.0013964 0.99468 0.50475 0.0018814 0.42694 2.2605 2.26 16.0127 144.9142 0.00015576 -85.6573 0.90794
9.012 0.98815 5.4604e-005 3.8183 0.01191 0.00011702 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6267 0.60374 0.18431 0.020921 19.1863 0.12949 0.00017 0.76068 0.0096439 0.010658 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16671 0.94745 0.92133 0.0013964 0.99469 0.50492 0.0018814 0.42696 2.2609 2.2604 16.0127 144.9142 0.0001557 -85.6573 0.90894
9.013 0.98815 5.4604e-005 3.8183 0.01191 0.00011704 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6268 0.60378 0.18432 0.020922 19.1895 0.12949 0.00017001 0.76068 0.0096443 0.010658 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16671 0.94756 0.92138 0.0013964 0.99471 0.50509 0.0018813 0.42697 2.2613 2.2608 16.0126 144.9142 0.00015563 -85.6573 0.90994
9.014 0.98815 5.4604e-005 3.8183 0.01191 0.00011705 0.0011771 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6269 0.60383 0.18433 0.020923 19.1928 0.1295 0.00017002 0.76067 0.0096446 0.010659 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16672 0.94767 0.92142 0.0013964 0.99473 0.50527 0.0018813 0.42698 2.2616 2.2611 16.0126 144.9143 0.00015556 -85.6574 0.91094
9.015 0.98815 5.4604e-005 3.8183 0.01191 0.00011706 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.627 0.60387 0.18435 0.020924 19.1961 0.1295 0.00017003 0.76067 0.0096449 0.010659 0.001385 0.98696 0.99172 2.9863e-006 1.1945e-005 0.16672 0.94778 0.92146 0.0013964 0.99474 0.50544 0.0018813 0.427 2.262 2.2615 16.0126 144.9143 0.0001555 -85.6574 0.91194
9.016 0.98815 5.4603e-005 3.8183 0.01191 0.00011708 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6271 0.60392 0.18436 0.020925 19.1994 0.12951 0.00017004 0.76066 0.0096453 0.010659 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16672 0.94789 0.9215 0.0013964 0.99476 0.50561 0.0018813 0.42701 2.2624 2.2619 16.0125 144.9143 0.00015544 -85.6575 0.91294
9.017 0.98815 5.4603e-005 3.8183 0.01191 0.00011709 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6272 0.60396 0.18437 0.020926 19.2026 0.12952 0.00017005 0.76065 0.0096456 0.01066 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16672 0.94801 0.92155 0.0013964 0.99477 0.50578 0.0018813 0.42702 2.2628 2.2623 16.0125 144.9143 0.00015537 -85.6575 0.91394
9.018 0.98815 5.4603e-005 3.8183 0.01191 0.0001171 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6272 0.604 0.18439 0.020927 19.2059 0.12952 0.00017005 0.76065 0.009646 0.01066 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16673 0.94812 0.92159 0.0013964 0.99479 0.50596 0.0018813 0.42704 2.2631 2.2626 16.0125 144.9143 0.00015531 -85.6575 0.91494
9.019 0.98815 5.4603e-005 3.8183 0.01191 0.00011711 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6273 0.60405 0.1844 0.020928 19.2092 0.12953 0.00017006 0.76064 0.0096463 0.01066 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16673 0.94823 0.92163 0.0013964 0.9948 0.50613 0.0018813 0.42705 2.2635 2.263 16.0124 144.9144 0.00015524 -85.6576 0.91594
9.02 0.98815 5.4603e-005 3.8183 0.01191 0.00011713 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6274 0.60409 0.18441 0.020929 19.2125 0.12953 0.00017007 0.76064 0.0096466 0.010661 0.001385 0.98696 0.99172 2.9862e-006 1.1945e-005 0.16673 0.94834 0.92167 0.0013964 0.99482 0.5063 0.0018813 0.42707 2.2639 2.2634 16.0124 144.9144 0.00015518 -85.6576 0.91694
9.021 0.98815 5.4603e-005 3.8183 0.01191 0.00011714 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6275 0.60414 0.18443 0.02093 19.2158 0.12954 0.00017008 0.76063 0.009647 0.010661 0.001385 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16673 0.94845 0.92171 0.0013964 0.99484 0.50647 0.0018813 0.42708 2.2643 2.2638 16.0124 144.9144 0.00015511 -85.6577 0.91794
9.022 0.98815 5.4603e-005 3.8183 0.01191 0.00011715 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6276 0.60418 0.18444 0.020931 19.219 0.12955 0.00017009 0.76062 0.0096473 0.010662 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16674 0.94856 0.92175 0.0013964 0.99485 0.50664 0.0018813 0.42709 2.2646 2.2641 16.0123 144.9144 0.00015505 -85.6577 0.91894
9.023 0.98815 5.4603e-005 3.8183 0.01191 0.00011717 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6277 0.60422 0.18445 0.020932 19.2223 0.12955 0.0001701 0.76062 0.0096476 0.010662 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16674 0.94867 0.92179 0.0013964 0.99487 0.50682 0.0018813 0.42711 2.265 2.2645 16.0123 144.9144 0.00015499 -85.6577 0.91994
9.024 0.98815 5.4603e-005 3.8183 0.01191 0.00011718 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6277 0.60427 0.18446 0.020933 19.2256 0.12956 0.00017011 0.76061 0.009648 0.010662 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16674 0.94878 0.92183 0.0013964 0.99488 0.50699 0.0018813 0.42712 2.2654 2.2649 16.0123 144.9145 0.00015493 -85.6578 0.92094
9.025 0.98815 5.4603e-005 3.8183 0.01191 0.00011719 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6278 0.60431 0.18448 0.020934 19.2289 0.12956 0.00017012 0.76061 0.0096483 0.010663 0.0013849 0.98696 0.99172 2.9861e-006 1.1944e-005 0.16674 0.94888 0.92187 0.0013964 0.9949 0.50716 0.0018813 0.42713 2.2657 2.2653 16.0122 144.9145 0.00015486 -85.6578 0.92194
9.026 0.98815 5.4603e-005 3.8183 0.01191 0.0001172 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6279 0.60436 0.18449 0.020935 19.2322 0.12957 0.00017013 0.7606 0.0096486 0.010663 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16675 0.94899 0.92192 0.0013964 0.99491 0.50733 0.0018813 0.42715 2.2661 2.2656 16.0122 144.9145 0.0001548 -85.6578 0.92294
9.027 0.98815 5.4603e-005 3.8183 0.01191 0.00011722 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.628 0.6044 0.1845 0.020936 19.2354 0.12958 0.00017014 0.76059 0.009649 0.010663 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16675 0.9491 0.92196 0.0013964 0.99492 0.5075 0.0018813 0.42716 2.2665 2.266 16.0122 144.9145 0.00015474 -85.6579 0.92394
9.028 0.98815 5.4602e-005 3.8183 0.01191 0.00011723 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6281 0.60445 0.18452 0.020937 19.2387 0.12958 0.00017015 0.76059 0.0096493 0.010664 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16675 0.94921 0.922 0.0013963 0.99494 0.50768 0.0018813 0.42717 2.2668 2.2664 16.0121 144.9145 0.00015468 -85.6579 0.92494
9.029 0.98815 5.4602e-005 3.8183 0.01191 0.00011724 0.0011772 0.23359 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6282 0.60449 0.18453 0.020938 19.242 0.12959 0.00017016 0.76058 0.0096497 0.010664 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16675 0.94932 0.92204 0.0013963 0.99495 0.50785 0.0018813 0.42719 2.2672 2.2667 16.0121 144.9146 0.00015461 -85.6579 0.92594
9.03 0.98815 5.4602e-005 3.8183 0.01191 0.00011725 0.0011772 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6282 0.60453 0.18454 0.020939 19.2453 0.12959 0.00017016 0.76058 0.00965 0.010664 0.0013849 0.98696 0.99172 2.986e-006 1.1944e-005 0.16676 0.94942 0.92208 0.0013963 0.99497 0.50802 0.0018812 0.4272 2.2676 2.2671 16.0121 144.9146 0.00015455 -85.658 0.92694
9.031 0.98815 5.4602e-005 3.8183 0.011909 0.00011727 0.0011772 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6283 0.60458 0.18455 0.02094 19.2486 0.1296 0.00017017 0.76057 0.0096503 0.010665 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16676 0.94953 0.92212 0.0013963 0.99498 0.50819 0.0018812 0.42721 2.2679 2.2675 16.012 144.9146 0.00015449 -85.658 0.92794
9.032 0.98815 5.4602e-005 3.8183 0.011909 0.00011728 0.0011772 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6284 0.60462 0.18457 0.020941 19.2519 0.12961 0.00017018 0.76057 0.0096507 0.010665 0.0013849 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16676 0.94964 0.92216 0.0013963 0.995 0.50836 0.0018812 0.42723 2.2683 2.2678 16.012 144.9146 0.00015443 -85.658 0.92894
9.033 0.98815 5.4602e-005 3.8183 0.011909 0.00011729 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6285 0.60467 0.18458 0.020942 19.2551 0.12961 0.00017019 0.76056 0.009651 0.010665 0.0013848 0.98696 0.99172 2.9859e-006 1.1944e-005 0.16676 0.94974 0.9222 0.0013963 0.99501 0.50853 0.0018812 0.42724 2.2687 2.2682 16.012 144.9146 0.00015437 -85.6581 0.92994
9.034 0.98815 5.4602e-005 3.8183 0.011909 0.00011731 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6286 0.60471 0.18459 0.020943 19.2584 0.12962 0.0001702 0.76055 0.0096513 0.010666 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16677 0.94985 0.92223 0.0013963 0.99503 0.5087 0.0018812 0.42725 2.269 2.2686 16.0119 144.9147 0.00015431 -85.6581 0.93094
9.035 0.98815 5.4602e-005 3.8183 0.011909 0.00011732 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6287 0.60476 0.18461 0.020944 19.2617 0.12962 0.00017021 0.76055 0.0096517 0.010666 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16677 0.94995 0.92227 0.0013963 0.99504 0.50888 0.0018812 0.42727 2.2694 2.2689 16.0119 144.9147 0.00015425 -85.6582 0.93194
9.036 0.98815 5.4602e-005 3.8183 0.011909 0.00011733 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6287 0.6048 0.18462 0.020945 19.265 0.12963 0.00017022 0.76054 0.009652 0.010667 0.0013848 0.98696 0.99172 2.9859e-006 1.1943e-005 0.16677 0.95006 0.92231 0.0013963 0.99505 0.50905 0.0018812 0.42728 2.2698 2.2693 16.0119 144.9147 0.00015419 -85.6582 0.93294
9.037 0.98815 5.4602e-005 3.8183 0.011909 0.00011734 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6288 0.60484 0.18463 0.020946 19.2683 0.12963 0.00017023 0.76054 0.0096523 0.010667 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16677 0.95016 0.92235 0.0013963 0.99507 0.50922 0.0018812 0.42729 2.2701 2.2697 16.0118 144.9147 0.00015413 -85.6582 0.93394
9.038 0.98815 5.4602e-005 3.8183 0.011909 0.00011736 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6289 0.60489 0.18464 0.020947 19.2716 0.12964 0.00017024 0.76053 0.0096527 0.010667 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16678 0.95027 0.92239 0.0013963 0.99508 0.50939 0.0018812 0.42731 2.2705 2.27 16.0118 144.9147 0.00015407 -85.6582 0.93494
9.039 0.98815 5.4602e-005 3.8183 0.011909 0.00011737 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.629 0.60493 0.18466 0.020948 19.2748 0.12965 0.00017025 0.76052 0.009653 0.010668 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16678 0.95037 0.92243 0.0013963 0.99509 0.50956 0.0018812 0.42732 2.2708 2.2704 16.0118 144.9148 0.00015401 -85.6583 0.93594
9.04 0.98815 5.4601e-005 3.8183 0.011909 0.00011738 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6291 0.60498 0.18467 0.020949 19.2781 0.12965 0.00017026 0.76052 0.0096533 0.010668 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16678 0.95047 0.92247 0.0013963 0.99511 0.50973 0.0018812 0.42733 2.2712 2.2707 16.0117 144.9148 0.00015395 -85.6583 0.93694
9.041 0.98815 5.4601e-005 3.8183 0.011909 0.0001174 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6292 0.60502 0.18468 0.02095 19.2814 0.12966 0.00017026 0.76051 0.0096537 0.010668 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16679 0.95058 0.92251 0.0013963 0.99512 0.5099 0.0018812 0.42735 2.2716 2.2711 16.0117 144.9148 0.00015389 -85.6583 0.93794
9.042 0.98815 5.4601e-005 3.8183 0.011909 0.00011741 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6292 0.60506 0.1847 0.020951 19.2847 0.12966 0.00017027 0.76051 0.009654 0.010669 0.0013848 0.98696 0.99172 2.9858e-006 1.1943e-005 0.16679 0.95068 0.92255 0.0013963 0.99513 0.51007 0.0018812 0.42736 2.2719 2.2715 16.0117 144.9148 0.00015383 -85.6584 0.93894
9.043 0.98815 5.4601e-005 3.8183 0.011909 0.00011742 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6293 0.60511 0.18471 0.020952 19.288 0.12967 0.00017028 0.7605 0.0096544 0.010669 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16679 0.95078 0.92258 0.0013963 0.99515 0.51024 0.0018812 0.42737 2.2723 2.2718 16.0116 144.9148 0.00015377 -85.6584 0.93994
9.044 0.98815 5.4601e-005 3.8183 0.011909 0.00011743 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6294 0.60515 0.18472 0.020953 19.2913 0.12968 0.00017029 0.76049 0.0096547 0.010669 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.16679 0.95089 0.92262 0.0013963 0.99516 0.51041 0.0018812 0.42739 2.2726 2.2722 16.0116 144.9149 0.00015371 -85.6584 0.94094
9.045 0.98815 5.4601e-005 3.8183 0.011909 0.00011745 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6295 0.6052 0.18474 0.020954 19.2946 0.12968 0.0001703 0.76049 0.009655 0.01067 0.0013848 0.98696 0.99172 2.9857e-006 1.1943e-005 0.1668 0.95099 0.92266 0.0013963 0.99517 0.51058 0.0018812 0.4274 2.273 2.2725 16.0116 144.9149 0.00015365 -85.6585 0.94194
9.046 0.98815 5.4601e-005 3.8183 0.011909 0.00011746 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6296 0.60524 0.18475 0.020955 19.2978 0.12969 0.00017031 0.76048 0.0096554 0.01067 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.1668 0.95109 0.9227 0.0013963 0.99519 0.51075 0.0018812 0.42741 2.2734 2.2729 16.0115 144.9149 0.00015359 -85.6585 0.94294
9.047 0.98815 5.4601e-005 3.8183 0.011909 0.00011747 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6296 0.60529 0.18476 0.020956 19.3011 0.12969 0.00017032 0.76048 0.0096557 0.01067 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.1668 0.95119 0.92274 0.0013963 0.9952 0.51092 0.0018812 0.42743 2.2737 2.2733 16.0115 144.9149 0.00015353 -85.6585 0.94394
9.048 0.98815 5.4601e-005 3.8183 0.011909 0.00011748 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6297 0.60533 0.18477 0.020957 19.3044 0.1297 0.00017033 0.76047 0.009656 0.010671 0.0013847 0.98696 0.99172 2.9857e-006 1.1943e-005 0.1668 0.95129 0.92277 0.0013963 0.99521 0.5111 0.0018812 0.42744 2.2741 2.2736 16.0115 144.915 0.00015348 -85.6586 0.94494
9.049 0.98815 5.4601e-005 3.8183 0.011909 0.0001175 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6298 0.60537 0.18479 0.020958 19.3077 0.12971 0.00017034 0.76046 0.0096564 0.010671 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16681 0.95139 0.92281 0.0013963 0.99523 0.51127 0.0018811 0.42745 2.2744 2.274 16.0114 144.915 0.00015342 -85.6586 0.94594
9.05 0.98815 5.4601e-005 3.8183 0.011909 0.00011751 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.6299 0.60542 0.1848 0.020959 19.311 0.12971 0.00017035 0.76046 0.0096567 0.010671 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16681 0.95149 0.92285 0.0013963 0.99524 0.51144 0.0018811 0.42747 2.2748 2.2743 16.0114 144.915 0.00015336 -85.6586 0.94694
9.051 0.98815 5.46e-005 3.8183 0.011909 0.00011752 0.0011773 0.23358 0.00065931 0.23424 0.21615 0 0.032265 0.0389 0 1.63 0.60546 0.18481 0.02096 19.3143 0.12972 0.00017036 0.76045 0.009657 0.010672 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16681 0.95159 0.92289 0.0013963 0.99525 0.51161 0.0018811 0.42748 2.2751 2.2747 16.0114 144.915 0.0001533 -85.6586 0.94794
9.052 0.98815 5.46e-005 3.8183 0.011909 0.00011754 0.0011774 0.23358 0.00065931 0.23423 0.21615 0 0.032265 0.0389 0 1.6301 0.60551 0.18483 0.020961 19.3176 0.12972 0.00017037 0.76045 0.0096574 0.010672 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16681 0.95169 0.92292 0.0013963 0.99526 0.51178 0.0018811 0.42749 2.2755 2.275 16.0113 144.915 0.00015325 -85.6587 0.94894
9.053 0.98815 5.46e-005 3.8183 0.011909 0.00011755 0.0011774 0.23358 0.00065931 0.23423 0.21615 0 0.032265 0.0389 0 1.6301 0.60555 0.18484 0.020962 19.3209 0.12973 0.00017037 0.76044 0.0096577 0.010673 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16682 0.95179 0.92296 0.0013963 0.99528 0.51195 0.0018811 0.42751 2.2758 2.2754 16.0113 144.9151 0.00015319 -85.6587 0.94994
9.054 0.98815 5.46e-005 3.8183 0.011909 0.00011756 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6302 0.60559 0.18485 0.020963 19.3242 0.12974 0.00017038 0.76043 0.009658 0.010673 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16682 0.95189 0.923 0.0013963 0.99529 0.51212 0.0018811 0.42752 2.2762 2.2757 16.0113 144.9151 0.00015313 -85.6587 0.95094
9.055 0.98815 5.46e-005 3.8183 0.011909 0.00011757 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6303 0.60564 0.18486 0.020964 19.3275 0.12974 0.00017039 0.76043 0.0096584 0.010673 0.0013847 0.98696 0.99172 2.9856e-006 1.1942e-005 0.16682 0.95199 0.92303 0.0013962 0.9953 0.51229 0.0018811 0.42753 2.2765 2.2761 16.0112 144.9151 0.00015308 -85.6588 0.95194
9.056 0.98815 5.46e-005 3.8183 0.011909 0.00011759 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6304 0.60568 0.18488 0.020965 19.3307 0.12975 0.0001704 0.76042 0.0096587 0.010674 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16682 0.95209 0.92307 0.0013962 0.99531 0.51246 0.0018811 0.42755 2.2769 2.2764 16.0112 144.9151 0.00015302 -85.6588 0.95294
9.057 0.98815 5.46e-005 3.8183 0.011909 0.0001176 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6305 0.60573 0.18489 0.020966 19.334 0.12975 0.00017041 0.76042 0.009659 0.010674 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16683 0.95219 0.92311 0.0013962 0.99532 0.51263 0.0018811 0.42756 2.2772 2.2768 16.0112 144.9151 0.00015296 -85.6588 0.95394
9.058 0.98815 5.46e-005 3.8183 0.011909 0.00011761 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6306 0.60577 0.1849 0.020967 19.3373 0.12976 0.00017042 0.76041 0.0096594 0.010674 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16683 0.95229 0.92314 0.0013962 0.99534 0.5128 0.0018811 0.42757 2.2776 2.2771 16.0111 144.9152 0.00015291 -85.6588 0.95494
9.059 0.98815 5.46e-005 3.8183 0.011909 0.00011763 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6306 0.60582 0.18492 0.020968 19.3406 0.12977 0.00017043 0.7604 0.0096597 0.010675 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16683 0.95238 0.92318 0.0013962 0.99535 0.51297 0.0018811 0.42759 2.2779 2.2775 16.0111 144.9152 0.00015285 -85.6589 0.95594
9.06 0.98815 5.46e-005 3.8183 0.011909 0.00011764 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6307 0.60586 0.18493 0.020969 19.3439 0.12977 0.00017044 0.7604 0.00966 0.010675 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16683 0.95248 0.92322 0.0013962 0.99536 0.51314 0.0018811 0.4276 2.2783 2.2778 16.0111 144.9152 0.00015279 -85.6589 0.95694
9.061 0.98815 5.46e-005 3.8183 0.011909 0.00011765 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6308 0.6059 0.18494 0.02097 19.3472 0.12978 0.00017045 0.76039 0.0096604 0.010675 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16684 0.95258 0.92325 0.0013962 0.99537 0.51331 0.0018811 0.42761 2.2786 2.2782 16.011 144.9152 0.00015274 -85.6589 0.95794
9.062 0.98815 5.46e-005 3.8183 0.011909 0.00011766 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6309 0.60595 0.18495 0.020971 19.3505 0.12978 0.00017046 0.76039 0.0096607 0.010676 0.0013847 0.98696 0.99172 2.9855e-006 1.1942e-005 0.16684 0.95267 0.92329 0.0013962 0.99538 0.51347 0.0018811 0.42763 2.279 2.2785 16.011 144.9152 0.00015268 -85.6589 0.95894
9.063 0.98815 5.4599e-005 3.8183 0.011909 0.00011768 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.631 0.60599 0.18497 0.020972 19.3538 0.12979 0.00017047 0.76038 0.0096611 0.010676 0.0013847 0.98696 0.99172 2.9854e-006 1.1942e-005 0.16684 0.95277 0.92332 0.0013962 0.9954 0.51364 0.0018811 0.42764 2.2793 2.2789 16.011 144.9153 0.00015263 -85.659 0.95994
9.064 0.98815 5.4599e-005 3.8183 0.011909 0.00011769 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6311 0.60604 0.18498 0.020973 19.3571 0.1298 0.00017047 0.76038 0.0096614 0.010676 0.0013846 0.98697 0.99172 2.9854e-006 1.1942e-005 0.16684 0.95287 0.92336 0.0013962 0.99541 0.51381 0.0018811 0.42765 2.2797 2.2792 16.0109 144.9153 0.00015257 -85.659 0.96094
9.065 0.98815 5.4599e-005 3.8183 0.011909 0.0001177 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6311 0.60608 0.18499 0.020974 19.3604 0.1298 0.00017048 0.76037 0.0096617 0.010677 0.0013846 0.98697 0.99172 2.9854e-006 1.1942e-005 0.16685 0.95296 0.92339 0.0013962 0.99542 0.51398 0.0018811 0.42767 2.28 2.2796 16.0109 144.9153 0.00015252 -85.659 0.96194
9.066 0.98815 5.4599e-005 3.8183 0.011909 0.00011771 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6312 0.60613 0.18501 0.020975 19.3637 0.12981 0.00017049 0.76036 0.0096621 0.010677 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16685 0.95306 0.92343 0.0013962 0.99543 0.51415 0.0018811 0.42768 2.2804 2.2799 16.0109 144.9153 0.00015246 -85.659 0.96294
9.067 0.98815 5.4599e-005 3.8183 0.011909 0.00011773 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6313 0.60617 0.18502 0.020976 19.367 0.12981 0.0001705 0.76036 0.0096624 0.010677 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16685 0.95315 0.92346 0.0013962 0.99544 0.51432 0.0018811 0.42769 2.2807 2.2803 16.0108 144.9153 0.00015241 -85.6591 0.96394
9.068 0.98815 5.4599e-005 3.8183 0.011909 0.00011774 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6314 0.60621 0.18503 0.020977 19.3703 0.12982 0.00017051 0.76035 0.0096627 0.010678 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16685 0.95325 0.9235 0.0013962 0.99545 0.51449 0.0018811 0.42771 2.2811 2.2806 16.0108 144.9154 0.00015236 -85.6591 0.96494
9.069 0.98815 5.4599e-005 3.8183 0.011909 0.00011775 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6315 0.60626 0.18504 0.020978 19.3736 0.12982 0.00017052 0.76035 0.0096631 0.010678 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16686 0.95334 0.92353 0.0013962 0.99546 0.51466 0.0018811 0.42772 2.2814 2.281 16.0108 144.9154 0.0001523 -85.6591 0.96594
9.07 0.98815 5.4599e-005 3.8183 0.011909 0.00011777 0.0011774 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6316 0.6063 0.18506 0.020979 19.3768 0.12983 0.00017053 0.76034 0.0096634 0.010679 0.0013846 0.98697 0.99172 2.9854e-006 1.1941e-005 0.16686 0.95344 0.92357 0.0013962 0.99547 0.51483 0.0018811 0.42773 2.2818 2.2813 16.0107 144.9154 0.00015225 -85.6591 0.96694
9.071 0.98815 5.4599e-005 3.8183 0.011909 0.00011778 0.0011775 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6316 0.60635 0.18507 0.02098 19.3801 0.12984 0.00017054 0.76033 0.0096637 0.010679 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16686 0.95353 0.9236 0.0013962 0.99549 0.515 0.0018811 0.42775 2.2821 2.2817 16.0107 144.9154 0.00015219 -85.6592 0.96794
9.072 0.98815 5.4599e-005 3.8183 0.011909 0.00011779 0.0011775 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6317 0.60639 0.18508 0.020981 19.3834 0.12984 0.00017055 0.76033 0.0096641 0.010679 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16686 0.95362 0.92364 0.0013962 0.9955 0.51517 0.0018811 0.42776 2.2824 2.282 16.0106 144.9154 0.00015214 -85.6592 0.96894
9.073 0.98815 5.4599e-005 3.8183 0.011909 0.0001178 0.0011775 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6318 0.60643 0.1851 0.020982 19.3867 0.12985 0.00017056 0.76032 0.0096644 0.01068 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16687 0.95372 0.92367 0.0013962 0.99551 0.51534 0.001881 0.42777 2.2828 2.2823 16.0106 144.9155 0.00015209 -85.6592 0.96994
9.074 0.98815 5.4599e-005 3.8183 0.011909 0.00011782 0.0011775 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6319 0.60648 0.18511 0.020983 19.39 0.12985 0.00017057 0.76032 0.0096647 0.01068 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16687 0.95381 0.92371 0.0013962 0.99552 0.51551 0.001881 0.42779 2.2831 2.2827 16.0106 144.9155 0.00015203 -85.6592 0.97094
9.075 0.98815 5.4598e-005 3.8183 0.011909 0.00011783 0.0011775 0.23358 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.632 0.60652 0.18512 0.020984 19.3933 0.12986 0.00017058 0.76031 0.0096651 0.01068 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16687 0.9539 0.92374 0.0013962 0.99553 0.51567 0.001881 0.4278 2.2835 2.283 16.0105 144.9155 0.00015198 -85.6593 0.97194
9.076 0.98815 5.4598e-005 3.8183 0.011909 0.00011784 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6321 0.60657 0.18514 0.020985 19.3966 0.12987 0.00017058 0.7603 0.0096654 0.010681 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16687 0.954 0.92378 0.0013962 0.99554 0.51584 0.001881 0.42781 2.2838 2.2834 16.0105 144.9155 0.00015193 -85.6593 0.97294
9.077 0.98815 5.4598e-005 3.8183 0.011909 0.00011786 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6321 0.60661 0.18515 0.020986 19.3999 0.12987 0.00017059 0.7603 0.0096657 0.010681 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16688 0.95409 0.92381 0.0013962 0.99555 0.51601 0.001881 0.42782 2.2841 2.2837 16.0105 144.9156 0.00015188 -85.6593 0.97394
9.078 0.98815 5.4598e-005 3.8183 0.011909 0.00011787 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6322 0.60666 0.18516 0.020987 19.4032 0.12988 0.0001706 0.76029 0.0096661 0.010681 0.0013846 0.98697 0.99172 2.9853e-006 1.1941e-005 0.16688 0.95418 0.92384 0.0013962 0.99556 0.51618 0.001881 0.42784 2.2845 2.284 16.0104 144.9156 0.00015182 -85.6593 0.97494
9.079 0.98815 5.4598e-005 3.8183 0.011909 0.00011788 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6323 0.6067 0.18517 0.020988 19.4065 0.12988 0.00017061 0.76029 0.0096664 0.010682 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16688 0.95427 0.92388 0.0013962 0.99557 0.51635 0.001881 0.42785 2.2848 2.2844 16.0104 144.9156 0.00015177 -85.6593 0.97594
9.08 0.98815 5.4598e-005 3.8183 0.011909 0.00011789 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6324 0.60674 0.18519 0.020989 19.4098 0.12989 0.00017062 0.76028 0.0096667 0.010682 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16689 0.95436 0.92391 0.0013962 0.99558 0.51652 0.001881 0.42786 2.2852 2.2847 16.0104 144.9156 0.00015172 -85.6594 0.97694
9.081 0.98815 5.4598e-005 3.8183 0.011909 0.00011791 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6325 0.60679 0.1852 0.02099 19.4131 0.1299 0.00017063 0.76027 0.0096671 0.010682 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16689 0.95446 0.92395 0.0013962 0.99559 0.51669 0.001881 0.42788 2.2855 2.2851 16.0103 144.9156 0.00015167 -85.6594 0.97794
9.082 0.98815 5.4598e-005 3.8183 0.011909 0.00011792 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6326 0.60683 0.18521 0.020991 19.4164 0.1299 0.00017064 0.76027 0.0096674 0.010683 0.0013846 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16689 0.95455 0.92398 0.0013962 0.9956 0.51685 0.001881 0.42789 2.2858 2.2854 16.0103 144.9157 0.00015162 -85.6594 0.97894
9.083 0.98815 5.4598e-005 3.8183 0.011909 0.00011793 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6326 0.60688 0.18523 0.020992 19.4197 0.12991 0.00017065 0.76026 0.0096677 0.010683 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.16689 0.95464 0.92401 0.0013962 0.99561 0.51702 0.001881 0.4279 2.2862 2.2857 16.0103 144.9157 0.00015156 -85.6594 0.97994
9.084 0.98815 5.4598e-005 3.8183 0.011909 0.00011794 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6327 0.60692 0.18524 0.020993 19.423 0.12991 0.00017066 0.76026 0.0096681 0.010683 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1669 0.95473 0.92405 0.0013962 0.99562 0.51719 0.001881 0.42792 2.2865 2.2861 16.0102 144.9157 0.00015151 -85.6594 0.98094
9.085 0.98815 5.4598e-005 3.8183 0.011909 0.00011796 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6328 0.60696 0.18525 0.020994 19.4263 0.12992 0.00017067 0.76025 0.0096684 0.010684 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1669 0.95482 0.92408 0.0013962 0.99563 0.51736 0.001881 0.42793 2.2868 2.2864 16.0102 144.9157 0.00015146 -85.6595 0.98194
9.086 0.98815 5.4598e-005 3.8183 0.011908 0.00011797 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032265 0.0389 0 1.6329 0.60701 0.18526 0.020995 19.4296 0.12993 0.00017068 0.76024 0.0096687 0.010684 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1669 0.95491 0.92411 0.0013962 0.99564 0.51753 0.001881 0.42794 2.2872 2.2867 16.0102 144.9157 0.00015141 -85.6595 0.98294
9.087 0.98815 5.4597e-005 3.8183 0.011908 0.00011798 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.633 0.60705 0.18528 0.020996 19.4329 0.12993 0.00017068 0.76024 0.0096691 0.010685 0.0013845 0.98697 0.99172 2.9852e-006 1.1941e-005 0.1669 0.955 0.92415 0.0013962 0.99565 0.5177 0.001881 0.42796 2.2875 2.2871 16.0101 144.9158 0.00015136 -85.6595 0.98394
9.088 0.98815 5.4597e-005 3.8183 0.011908 0.000118 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.633 0.6071 0.18529 0.020997 19.4362 0.12994 0.00017069 0.76023 0.0096694 0.010685 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16691 0.95509 0.92418 0.0013962 0.99566 0.51786 0.001881 0.42797 2.2878 2.2874 16.0101 144.9158 0.00015131 -85.6595 0.98494
9.089 0.98815 5.4597e-005 3.8183 0.011908 0.00011801 0.0011775 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6331 0.60714 0.1853 0.020998 19.4395 0.12994 0.0001707 0.76023 0.0096697 0.010685 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16691 0.95517 0.92421 0.0013962 0.99567 0.51803 0.001881 0.42798 2.2882 2.2877 16.0101 144.9158 0.00015126 -85.6595 0.98594
9.09 0.98815 5.4597e-005 3.8183 0.011908 0.00011802 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6332 0.60719 0.18532 0.020999 19.4428 0.12995 0.00017071 0.76022 0.0096701 0.010686 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16691 0.95526 0.92424 0.0013961 0.99568 0.5182 0.001881 0.428 2.2885 2.2881 16.01 144.9158 0.00015121 -85.6596 0.98694
9.091 0.98815 5.4597e-005 3.8183 0.011908 0.00011803 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6333 0.60723 0.18533 0.021 19.4461 0.12996 0.00017072 0.76022 0.0096704 0.010686 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16691 0.95535 0.92428 0.0013961 0.99569 0.51837 0.001881 0.42801 2.2888 2.2884 16.01 144.9158 0.00015116 -85.6596 0.98794
9.092 0.98815 5.4597e-005 3.8183 0.011908 0.00011805 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6334 0.60727 0.18534 0.021001 19.4494 0.12996 0.00017073 0.76021 0.0096707 0.010686 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16692 0.95544 0.92431 0.0013961 0.9957 0.51854 0.001881 0.42802 2.2892 2.2887 16.01 144.9159 0.00015111 -85.6596 0.98894
9.093 0.98815 5.4597e-005 3.8183 0.011908 0.00011806 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6335 0.60732 0.18535 0.021002 19.4527 0.12997 0.00017074 0.7602 0.0096711 0.010687 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16692 0.95553 0.92434 0.0013961 0.99571 0.5187 0.001881 0.42803 2.2895 2.2891 16.0099 144.9159 0.00015106 -85.6596 0.98994
9.094 0.98815 5.4597e-005 3.8183 0.011908 0.00011807 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6335 0.60736 0.18537 0.021003 19.456 0.12997 0.00017075 0.7602 0.0096714 0.010687 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16692 0.95562 0.92437 0.0013961 0.99572 0.51887 0.001881 0.42805 2.2898 2.2894 16.0099 144.9159 0.00015101 -85.6596 0.99094
9.095 0.98815 5.4597e-005 3.8183 0.011908 0.00011808 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6336 0.60741 0.18538 0.021004 19.4593 0.12998 0.00017076 0.76019 0.0096717 0.010687 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16692 0.9557 0.92441 0.0013961 0.99573 0.51904 0.001881 0.42806 2.2902 2.2897 16.0099 144.9159 0.00015096 -85.6597 0.99194
9.096 0.98815 5.4597e-005 3.8183 0.011908 0.0001181 0.0011776 0.23357 0.00065931 0.23423 0.21614 0 0.032266 0.0389 0 1.6337 0.60745 0.18539 0.021005 19.4626 0.12998 0.00017077 0.76019 0.0096721 0.010688 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16693 0.95579 0.92444 0.0013961 0.99574 0.51921 0.001881 0.42807 2.2905 2.2901 16.0098 144.9159 0.00015091 -85.6597 0.99294
9.097 0.98815 5.4597e-005 3.8183 0.011908 0.00011811 0.0011776 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.6338 0.60749 0.18541 0.021006 19.4659 0.12999 0.00017078 0.76018 0.0096724 0.010688 0.0013845 0.98697 0.99172 2.9851e-006 1.194e-005 0.16693 0.95588 0.92447 0.0013961 0.99575 0.51937 0.001881 0.42809 2.2908 2.2904 16.0098 144.916 0.00015086 -85.6597 0.99394
9.098 0.98815 5.4597e-005 3.8183 0.011908 0.00011812 0.0011776 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.6339 0.60754 0.18542 0.021007 19.4692 0.13 0.00017078 0.76017 0.0096727 0.010688 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16693 0.95596 0.9245 0.0013961 0.99576 0.51954 0.001881 0.4281 2.2911 2.2907 16.0098 144.916 0.00015081 -85.6597 0.99494
9.099 0.98815 5.4596e-005 3.8183 0.011908 0.00011814 0.0011776 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.634 0.60758 0.18543 0.021008 19.4726 0.13 0.00017079 0.76017 0.0096731 0.010689 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16693 0.95605 0.92453 0.0013961 0.99577 0.51971 0.001881 0.42811 2.2915 2.2911 16.0097 144.916 0.00015076 -85.6597 0.99594
9.1 0.98815 5.4596e-005 3.8183 0.011908 0.00011815 0.0011776 0.23357 0.00065931 0.23422 0.21614 0 0.032266 0.0389 0 1.634 0.60763 0.18544 0.021009 19.4759 0.13001 0.0001708 0.76016 0.0096734 0.010689 0.0013845 0.98697 0.99172 2.985e-006 1.194e-005 0.16694 0.95613 0.92456 0.0013961 0.99578 0.51988 0.001881 0.42813 2.2918 2.2914 16.0097 144.916 0.00015071 -85.6587 0.99694
9.101 0.98815 5.4596e-005 3.8183 0.011908 0.00011816 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6341 0.60767 0.18546 0.02101 19.4792 0.13001 0.00017081 0.76016 0.0096737 0.010689 0.0064781 0.98322 0.99099 1.453e-005 5.3377e-005 0.16694 0.95617 0.9246 0.0027742 0.99577 0.52002 0.0023962 0.42809 2.2921 2.2917 16.0096 144.916 0.00015067 -76.1561 0.99794
9.102 0.98815 5.4596e-005 3.8183 0.011908 0.00011817 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6342 0.60772 0.18547 0.021011 19.4825 0.13002 0.00017082 0.76015 0.0096741 0.01069 0.026238 0.97169 0.98766 6.6022e-005 0.00022964 0.16694 0.95598 0.92463 0.0053023 0.99572 0.52015 0.003337 0.42797 2.2925 2.292 16.0096 144.916 0.00015066 -67.1424 0.99894
9.103 0.98815 5.4596e-005 3.8183 0.011908 0.00011819 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6343 0.60776 0.18548 0.021012 19.4858 0.13003 0.00017083 0.76014 0.0096744 0.01069 0.094933 0.94719 0.97731 0.0002846 0.00091374 0.16694 0.95525 0.92466 0.0092499 0.99546 0.52026 0.0044258 0.4278 2.2928 2.2924 16.0095 144.916 0.00015066 -58.0105 0.99994
9.104 0.98815 5.4596e-005 3.8183 0.011908 0.0001182 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6344 0.6078 0.1855 0.021013 19.4891 0.13003 0.00017084 0.76014 0.0096747 0.01069 0.48872 0.85607 0.93868 0.0021841 0.005486 0.16695 0.95326 0.92468 0.015758 0.99134 0.52031 0.0056249 0.42762 2.2931 2.2927 16.0102 144.916 0.00015069 -37.1797 0.15534
9.105 0.98815 5.4596e-005 3.8183 0.011908 0.00011821 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6345 0.60785 0.18551 0.021014 19.4924 0.13004 0.00017085 0.76013 0.009675 0.010691 0.99964 0.0021546 0.712 0.94446 0.99675 0.16695 0.91998 0.9216 0.3364 0.96393 0.50888 0.044611 0.42741 2.2318 0.98885 16.0141 144.9156 0.00025144 25.3853 0.0019369
9.106 0.98815 5.4596e-005 3.8183 0.011908 0.00011823 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6345 0.60789 0.18552 0.021015 19.4957 0.13004 0.00017086 0.76013 0.0096754 0.010691 0.99956 1.2714e-006 0.52802 0.9985 0.99965 0.16695 0.88011 0.90292 0.6333 0.93678 0.49462 0.10213 0.42721 2.0065 0.63489 16.0137 144.9142 0.00037358 22.8929 0.0029369
9.107 0.98815 5.4596e-005 3.8183 0.011908 0.00011824 0.0011776 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6346 0.60794 0.18553 0.021016 19.499 0.13005 0.00017087 0.76012 0.0096757 0.010692 0.99928 4.2151e-010 0.39179 0.99714 0.99921 0.16695 0.84227 0.87857 0.76383 0.91039 0.48086 0.14776 0.42701 1.7981 0.62469 16.0133 144.9124 0.00045468 18.129 0.0039369
9.108 0.98815 5.4596e-005 3.8183 0.011908 0.00011825 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6347 0.60798 0.18555 0.021017 19.5023 0.13006 0.00017088 0.76012 0.009676 0.010692 0.99896 -6.315e-011 0.29093 0.9948 0.99856 0.16696 0.80668 0.85106 0.82103 0.88475 0.46767 0.18401 0.4268 1.626 0.67806 16.013 144.9105 0.00051737 14.7797 0.0049369
9.109 0.98815 5.4596e-005 3.8183 0.011908 0.00011826 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6348 0.60802 0.18556 0.021018 19.5056 0.13006 0.00017088 0.76011 0.0096764 0.010692 0.99868 1.7443e-011 0.2162 0.99215 0.99784 0.16696 0.77336 0.82169 0.84634 0.85984 0.45506 0.21454 0.4266 1.4904 0.75137 16.0127 144.9086 0.00056668 12.56 0.0059369
9.11 0.98815 5.4596e-005 3.8183 0.011908 0.00011828 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6349 0.60807 0.18557 0.021019 19.5089 0.13007 0.00017089 0.7601 0.0096767 0.010693 0.99842 -2.4766e-010 0.16077 0.98936 0.99709 0.16696 0.74211 0.79137 0.85607 0.83563 0.44301 0.24121 0.4264 1.3871 0.82835 16.0123 144.9067 0.00060509 10.9002 0.0069369
9.111 0.98815 5.4595e-005 3.8183 0.011908 0.00011829 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.635 0.60811 0.18559 0.02102 19.5122 0.13007 0.0001709 0.7601 0.009677 0.010693 0.99816 -2.5756e-011 0.11962 0.98636 0.99627 0.16696 0.71277 0.76084 0.85738 0.8121 0.43149 0.26495 0.42619 1.311 0.90027 16.012 144.9049 0.0006347 9.5027 0.0079369
9.112 0.98815 5.4595e-005 3.8183 0.011908 0.0001183 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.635 0.60816 0.1856 0.021021 19.5155 0.13008 0.00017091 0.76009 0.0096774 0.010693 0.99789 -4.0083e-011 0.089057 0.98305 0.99535 0.16697 0.68523 0.73062 0.85373 0.78923 0.42049 0.28624 0.42599 1.2568 0.96237 16.0117 144.9032 0.00065751 8.2304 0.0089369
9.113 0.98815 5.4595e-005 3.8183 0.011908 0.00011831 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6351 0.6082 0.18561 0.021022 19.5189 0.13009 0.00017092 0.76009 0.0096777 0.010694 0.9976 2.1143e-011 0.066345 0.97928 0.99429 0.16697 0.65937 0.70109 0.84691 0.76702 0.41001 0.3054 0.42579 1.2194 1.0128 16.0114 144.9016 0.00067526 7.0172 0.0099369
9.114 0.98815 5.4595e-005 3.8183 0.011908 0.00011833 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6352 0.60825 0.18562 0.021023 19.5222 0.13009 0.00017093 0.76008 0.009678 0.010694 0.99726 -9.583e-011 0.049461 0.9749 0.99301 0.16697 0.63513 0.6725 0.8379 0.74543 0.40006 0.32265 0.42558 1.1946 1.052 16.0111 144.9001 0.00068934 5.828 0.010937
9.115 0.98815 5.4595e-005 3.8183 0.011908 0.00011834 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6353 0.60829 0.18564 0.021024 19.5255 0.1301 0.00017094 0.76007 0.0096784 0.010694 0.99689 9.346e-011 0.036902 0.96976 0.99152 0.16697 0.61244 0.64505 0.82722 0.72445 0.39063 0.33816 0.42538 1.1787 1.0813 16.0108 144.8986 0.00070082 4.6414 0.011937
9.116 0.98815 5.4595e-005 3.8183 0.011908 0.00011835 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6354 0.60833 0.18565 0.021025 19.5288 0.1301 0.00017095 0.76007 0.0096787 0.010695 0.99645 -5.6312e-011 0.027556 0.96366 0.98966 0.16698 0.59125 0.61886 0.81515 0.70406 0.38175 0.35206 0.42518 1.1691 1.1027 16.0105 144.8972 0.00071043 3.442 0.012937
9.117 0.98815 5.4595e-005 3.8183 0.011908 0.00011837 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6354 0.60838 0.18566 0.021026 19.5321 0.13011 0.00017096 0.76006 0.009679 0.010695 0.99594 3.2188e-011 0.020597 0.95637 0.98741 0.16698 0.5715 0.59401 0.80182 0.68426 0.37342 0.36445 0.42498 1.1637 1.1183 16.0103 144.8959 0.00071868 2.2164 0.013937
9.118 0.98815 5.4595e-005 3.8183 0.011908 0.00011838 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6355 0.60842 0.18568 0.021027 19.5354 0.13011 0.00017097 0.76006 0.0096794 0.010695 0.99533 -1.3534e-011 0.015413 0.94761 0.98463 0.16698 0.55315 0.57059 0.78726 0.66502 0.36565 0.37544 0.42478 1.1612 1.1297 16.01 144.8946 0.0007259 0.95059 0.014937
9.119 0.98815 5.4595e-005 3.8183 0.011908 0.00011839 0.0011777 0.23357 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6356 0.60847 0.18569 0.021028 19.5387 0.13012 0.00017098 0.76005 0.0096797 0.010696 0.9946 4.2255e-012 0.011549 0.937 0.98115 0.16698 0.53619 0.54865 0.77143 0.64632 0.35848 0.38507 0.42457 1.1606 1.1381 16.0097 144.8935 0.00073228 -0.37247 0.015937
9.12 0.98815 5.4595e-005 3.8183 0.011908 0.0001184 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6357 0.60851 0.1857 0.021029 19.542 0.13013 0.00017098 0.76004 0.00968 0.010696 0.9937 4.6821e-012 0.0086681 0.92405 0.97674 0.16699 0.52057 0.52826 0.75421 0.62816 0.35191 0.39342 0.42437 1.1612 1.1446 16.0095 144.8924 0.00073795 -1.7744 0.016937
9.121 0.98815 5.4595e-005 3.8183 0.011908 0.00011842 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6358 0.60855 0.18571 0.02103 19.5453 0.13013 0.00017099 0.76004 0.0096804 0.010696 0.99256 -6.1171e-012 0.0065182 0.90807 0.97108 0.16699 0.50629 0.5095 0.73546 0.61053 0.34598 0.40052 0.42417 1.1625 1.1497 16.0092 144.8914 0.00074297 -3.2847 0.017937
9.122 0.98815 5.4595e-005 3.8183 0.011908 0.00011843 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6359 0.6086 0.18573 0.021031 19.5486 0.13014 0.000171 0.76003 0.0096807 0.010697 0.99106 2.9285e-012 0.0049134 0.88811 0.96364 0.16699 0.49335 0.49244 0.71493 0.5934 0.34071 0.4064 0.42397 1.1644 1.154 16.009 144.8904 0.00074737 -4.9441 0.018937
9.123 0.98815 5.4594e-005 3.8183 0.011908 0.00011844 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6359 0.60864 0.18574 0.021032 19.552 0.13014 0.00017101 0.76003 0.009681 0.010697 0.989 -5.8955e-012 0.0037152 0.86283 0.95367 0.16699 0.48178 0.47718 0.69231 0.57678 0.33614 0.41105 0.42377 1.1666 1.1577 16.0087 144.8896 0.00075114 -6.8105 0.019937
9.124 0.98815 5.4594e-005 3.8183 0.011908 0.00011846 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.636 0.60869 0.18575 0.021033 19.5553 0.13015 0.00017102 0.76002 0.0096814 0.010697 0.98602 7.2152e-012 0.002821 0.83024 0.93993 0.167 0.4716 0.46387 0.66721 0.56065 0.33228 0.41446 0.42356 1.169 1.161 16.0085 144.8888 0.00075424 -8.9663 0.020937
9.125 0.98815 5.4594e-005 3.8183 0.011908 0.00011847 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6361 0.60873 0.18577 0.021034 19.5586 0.13016 0.00017103 0.76001 0.0096817 0.010698 0.9814 -4.6544e-012 0.0021547 0.78746 0.92042 0.167 0.46287 0.45263 0.63919 0.54503 0.32918 0.41663 0.42336 1.1716 1.1642 16.0083 144.888 0.00075659 -11.5266 0.021937
9.126 0.98815 5.4594e-005 3.8183 0.011908 0.00011848 0.0011777 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6362 0.60877 0.18578 0.021035 19.5619 0.13016 0.00017104 0.76001 0.009682 0.010698 0.97367 -1.461e-012 0.0016601 0.73032 0.89191 0.167 0.45565 0.44362 0.60783 0.52994 0.32682 0.41754 0.42316 1.1742 1.1672 16.0081 144.8874 0.00075811 -14.643 0.022937
9.127 0.98815 5.4594e-005 3.8183 0.011908 0.00011849 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6363 0.60882 0.18579 0.021036 19.5652 0.13017 0.00017105 0.76 0.0096823 0.010699 0.95959 -5.2198e-013 0.0012964 0.65314 0.84918 0.167 0.44993 0.43693 0.57291 0.51544 0.32516 0.41721 0.42296 1.1768 1.1701 16.0079 144.8868 0.00075867 -18.4832 0.023937
9.128 0.98815 5.4594e-005 3.8183 0.011908 0.00011851 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6364 0.60886 0.1858 0.021037 19.5685 0.13017 0.00017106 0.76 0.0096827 0.010699 0.93212 1.8206e-012 0.0010339 0.54974 0.78444 0.16701 0.44563 0.43251 0.53458 0.50172 0.32411 0.41572 0.42276 1.1795 1.1729 16.0078 144.8864 0.00075819 -23.1398 0.024937
9.129 0.98815 5.4594e-005 3.8183 0.011908 0.00011852 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6364 0.60891 0.18582 0.021038 19.5718 0.13018 0.00017107 0.75999 0.009683 0.010699 0.87835 -5.7788e-013 0.0008506 0.41813 0.68853 0.16701 0.44252 0.42999 0.49298 0.4892 0.32351 0.41321 0.42256 1.1823 1.1758 16.0076 144.886 0.00075675 -28.441 0.025937
9.13 0.98815 5.4594e-005 3.8183 0.011908 0.00011853 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6365 0.60895 0.18583 0.021039 19.5752 0.13019 0.00017107 0.75999 0.0096833 0.0107 0.78483 -6.3224e-014 0.00072753 0.27119 0.55736 0.16701 0.44027 0.42872 0.44732 0.47882 0.32322 0.4097 0.42236 1.185 1.1785 16.0075 144.8856 0.00075467 -33.8259 0.026937
9.131 0.98815 5.4594e-005 3.8183 0.011908 0.00011854 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6366 0.609 0.18584 0.02104 19.5785 0.13019 0.00017108 0.75998 0.0096837 0.0107 0.65637 -6.1804e-014 0.00064636 0.14122 0.40304 0.16701 0.4386 0.42816 0.39575 0.47185 0.32311 0.40499 0.42216 1.1877 1.1813 16.0074 144.8854 0.0007523 -38.6762 0.027937
9.132 0.98815 5.4594e-005 3.8183 0.011908 0.00011856 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6367 0.60904 0.18586 0.021041 19.5818 0.1302 0.00017109 0.75997 0.009684 0.0107 0.51947 0.00029421 0.00069002 0.0569 0.25405 0.16702 0.43736 0.42831 0.33747 0.46884 0.32312 0.39868 0.42197 1.1905 1.1841 16.0074 144.8852 0.00074982 -42.7692 0.028937
9.133 0.98815 5.4594e-005 3.8183 0.011908 0.00011857 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6368 0.60908 0.18587 0.021042 19.5851 0.1302 0.0001711 0.75997 0.0096843 0.010701 0.39952 0.00094179 0.00096905 0.018085 0.13787 0.16702 0.43646 0.42953 0.2745 0.46885 0.3232 0.3904 0.42177 1.1932 1.1868 16.0073 144.885 0.0007473 -46.1575 0.029937
9.134 0.98815 5.4593e-005 3.8183 0.011908 0.00011858 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6369 0.60913 0.18588 0.021043 19.5884 0.13021 0.00017111 0.75996 0.0096847 0.010701 0.30699 0.0019574 0.0014995 0.0052935 0.064766 0.16702 0.43588 0.4319 0.21161 0.47037 0.32332 0.37991 0.42158 1.1959 1.1896 16.0073 144.8849 0.00074473 -48.9426 0.030937
9.135 0.98815 5.4593e-005 3.8183 0.011908 0.0001186 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6369 0.60917 0.18589 0.021044 19.5917 0.13022 0.00017112 0.75996 0.009685 0.010701 0.24007 0.0034304 0.0023034 0.0020001 0.027285 0.16702 0.43555 0.43509 0.15449 0.47242 0.32347 0.36717 0.42139 1.1987 1.1924 16.0073 144.8848 0.00074214 -51.2304 0.031937
9.136 0.98815 5.4593e-005 3.8183 0.011908 0.00011861 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.637 0.60922 0.18591 0.021045 19.5951 0.13022 0.00017113 0.75995 0.0096853 0.010702 0.19235 0.0054272 0.0033905 0.0011316 0.011241 0.16703 0.43546 0.4387 0.10753 0.47455 0.32362 0.35232 0.42121 1.2014 1.1951 16.0073 144.8847 0.00073952 -53.129 0.032937
9.137 0.98815 5.4593e-005 3.8183 0.011908 0.00011862 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6371 0.60926 0.18592 0.021046 19.5984 0.13023 0.00017114 0.75994 0.0096857 0.010702 0.15768 0.0079986 0.0047637 0.00079241 0.0052141 0.16703 0.43556 0.44246 0.072398 0.47662 0.32378 0.33559 0.42103 1.2041 1.1979 16.0073 144.8847 0.00073689 -54.7402 0.033937
9.138 0.98815 5.4593e-005 3.8183 0.011908 0.00011863 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6372 0.6093 0.18593 0.021047 19.6017 0.13023 0.00017115 0.75994 0.009686 0.010702 0.13158 0.011191 0.0064255 0.00060012 0.0030209 0.16703 0.43582 0.44625 0.048255 0.47858 0.32395 0.3173 0.42085 1.2069 1.2006 16.0073 144.8846 0.00073424 -56.1501 0.034937
9.139 0.98815 5.4593e-005 3.8183 0.011908 0.00011865 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6373 0.60935 0.18595 0.021048 19.605 0.13024 0.00017116 0.75993 0.0096863 0.010703 0.11117 0.015057 0.0083818 0.00047123 0.002113 0.16703 0.43623 0.45002 0.032819 0.48042 0.32412 0.29773 0.42067 1.2096 1.2033 16.0073 144.8846 0.00073159 -57.4241 0.035937
9.14 0.98815 5.4593e-005 3.8183 0.011908 0.00011866 0.0011778 0.23356 0.00065931 0.23422 0.21613 0 0.032266 0.0389 0 1.6374 0.60939 0.18596 0.021049 19.6083 0.13024 0.00017117 0.75993 0.0096866 0.010703 0.094696 0.019664 0.010644 0.00037846 0.0016264 0.16704 0.43677 0.45375 0.023478 0.48216 0.32429 0.27716 0.42049 1.2123 1.2061 16.0074 144.8845 0.00072893 -58.6071 0.036937
9.141 0.98815 5.4593e-005 3.8183 0.011907 0.00011867 0.0011778 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.6374 0.60944 0.18597 0.02105 19.6116 0.13025 0.00017117 0.75992 0.009687 0.010703 0.081089 0.025094 0.013229 0.00030806 0.0013022 0.16704 0.43741 0.45745 0.017985 0.48381 0.32446 0.25589 0.42032 1.215 1.2088 16.0074 144.8845 0.00072626 -59.7277 0.037937
9.142 0.98815 5.4593e-005 3.8183 0.011907 0.00011869 0.0011778 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.6375 0.60948 0.18598 0.021051 19.615 0.13026 0.00017118 0.75991 0.0096873 0.010704 0.069689 0.031444 0.016158 0.00025296 0.0010611 0.16704 0.43816 0.46111 0.014719 0.48537 0.32463 0.23417 0.42015 1.2178 1.2116 16.0074 144.8845 0.00072359 -60.8025 0.038937
9.143 0.98815 5.4593e-005 3.8183 0.011907 0.0001187 0.0011778 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.6376 0.60953 0.186 0.021052 19.6183 0.13026 0.00017119 0.75991 0.0096876 0.010704 0.060061 0.038823 0.019456 0.00020967 0.00087354 0.16705 0.439 0.46473 0.012656 0.48686 0.3248 0.21228 0.41999 1.2205 1.2143 16.0075 144.8845 0.00072092 -61.8407 0.039937
9.144 0.98815 5.4593e-005 3.8183 0.011907 0.00011871 0.0011778 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.6377 0.60957 0.18601 0.021053 19.6216 0.13027 0.0001712 0.7599 0.009688 0.010704 0.051892 0.04735 0.02315 0.00017476 0.00072466 0.16705 0.43993 0.46831 0.011219 0.48829 0.32497 0.19053 0.41983 1.2232 1.217 16.0075 144.8844 0.00071825 -62.8475 0.040937
9.145 0.98815 5.4593e-005 3.8183 0.011907 0.00011872 0.0011778 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.6378 0.60961 0.18602 0.021054 19.6249 0.13027 0.00017121 0.7599 0.0096883 0.010705 0.044943 0.05715 0.027268 0.00014644 0.00060502 0.16705 0.44093 0.47185 0.010114 0.48966 0.32514 0.16919 0.41967 1.2259 1.2198 16.0076 144.8844 0.00071557 -63.8256 0.041937
9.146 0.98815 5.4592e-005 3.8183 0.011907 0.00011874 0.0011779 0.23356 0.00065931 0.23421 0.21613 0 0.032266 0.0389 0 1.6378 0.60966 0.18604 0.021055 19.6282 0.13028 0.00017122 0.75989 0.0096886 0.010705 0.039018 0.068352 0.031842 0.00012343 0.00050807 0.16705 0.442 0.47534 0.0092021 0.49099 0.32531 0.14857 0.41951 1.2286 1.2225 16.0076 144.8844 0.0007129 -64.7768 0.042937
9.147 0.98815 5.4592e-005 3.8183 0.011907 0.00011875 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6379 0.6097 0.18605 0.021056 19.6316 0.13029 0.00017123 0.75989 0.009689 0.010706 0.033959 0.081085 0.036904 0.00010451 0.00042896 0.16706 0.44314 0.4788 0.0084183 0.49229 0.32548 0.12893 0.41936 1.2313 1.2252 16.0077 144.8844 0.00071022 -65.7021 0.043937
9.148 0.98815 5.4592e-005 3.8183 0.011907 0.00011876 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.638 0.60975 0.18606 0.021057 19.6349 0.13029 0.00017124 0.75988 0.0096893 0.010706 0.029633 0.095475 0.042489 8.8908e-005 0.00036402 0.16706 0.44432 0.48223 0.0077313 0.49356 0.32565 0.11051 0.41922 1.2341 1.228 16.0078 144.8843 0.00070755 -66.6023 0.044937
9.149 0.98815 5.4592e-005 3.8183 0.011907 0.00011877 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6381 0.60979 0.18607 0.021058 19.6382 0.1303 0.00017125 0.75987 0.0096896 0.010706 0.025927 0.11164 0.048637 7.5989e-005 0.00031043 0.16706 0.44556 0.48561 0.0071233 0.49481 0.32582 0.093537 0.41907 1.2368 1.2307 16.0078 144.8843 0.00070487 -67.4779 0.045937
9.15 0.98815 5.4592e-005 3.8183 0.011907 0.00011879 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6382 0.60983 0.18609 0.021059 19.6415 0.1303 0.00017126 0.75987 0.00969 0.010707 0.022747 0.12969 0.055388 6.5246e-005 0.000266 0.16706 0.44683 0.48895 0.0065823 0.49605 0.32599 0.078155 0.41894 1.2395 1.2334 16.0079 144.8843 0.0007022 -68.3293 0.046937
9.151 0.98815 5.4592e-005 3.8183 0.011907 0.0001188 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6383 0.60988 0.1861 0.02106 19.6448 0.13031 0.00017127 0.75986 0.0096903 0.010707 0.020016 0.14972 0.062786 5.6268e-005 0.000229 0.16707 0.44815 0.49226 0.006099 0.49728 0.32616 0.064468 0.4188 1.2422 1.2361 16.008 144.8842 0.00069953 -69.1565 0.047937
9.152 0.98815 5.4592e-005 3.8183 0.011907 0.00011881 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6383 0.60992 0.18611 0.021061 19.6482 0.13032 0.00017127 0.75986 0.0096906 0.010707 0.017666 0.17179 0.070879 4.8749e-005 0.00019807 0.16707 0.4495 0.49553 0.0056662 0.49851 0.32634 0.052517 0.41868 1.2449 1.2389 16.0081 144.8842 0.00069686 -69.9592 0.048937
9.153 0.98815 5.4592e-005 3.8183 0.011907 0.00011883 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6384 0.60997 0.18613 0.021062 19.6515 0.13032 0.00017128 0.75985 0.0096909 0.010708 0.015642 0.19593 0.07972 4.242e-005 0.00017212 0.16707 0.45088 0.49876 0.0052777 0.49975 0.32651 0.042285 0.41855 1.2476 1.2416 16.0082 144.8842 0.0006942 -70.7372 0.049937
9.154 0.98815 5.4592e-005 3.8183 0.011907 0.00011884 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6385 0.61001 0.18614 0.021063 19.6548 0.13033 0.00017129 0.75984 0.0096913 0.010708 0.013897 0.22216 0.089361 3.7087e-005 0.00015028 0.16707 0.45228 0.50195 0.0049284 0.50099 0.32669 0.0337 0.41843 1.2503 1.2443 16.0082 144.8842 0.00069154 -71.49 0.050937
9.155 0.98815 5.4592e-005 3.8183 0.011907 0.00011885 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6386 0.61005 0.18615 0.021064 19.6581 0.13033 0.0001713 0.75984 0.0096916 0.010708 0.012391 0.25041 0.099856 3.2576e-005 0.00013184 0.16708 0.45371 0.50511 0.0046142 0.50225 0.32686 0.026644 0.41832 1.253 1.247 16.0083 144.8841 0.00068888 -72.2168 0.051937
9.156 0.98815 5.4592e-005 3.8183 0.011907 0.00011886 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6387 0.6101 0.18616 0.021065 19.6615 0.13034 0.00017131 0.75983 0.0096919 0.010709 0.011089 0.28061 0.11126 2.8748e-005 0.00011623 0.16708 0.45516 0.50824 0.0043311 0.50353 0.32704 0.020963 0.41821 1.2557 1.2497 16.0084 144.8841 0.00068623 -72.917 0.052937
9.157 0.98815 5.4592e-005 3.8183 0.011907 0.00011888 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6388 0.61014 0.18618 0.021066 19.6648 0.13034 0.00017132 0.75983 0.0096923 0.010709 0.0099635 0.3126 0.12361 2.5499e-005 0.00010299 0.16708 0.45662 0.51133 0.0040761 0.50483 0.32722 0.016483 0.41811 1.2584 1.2524 16.0085 144.8841 0.00068358 -73.5898 0.053937
9.158 0.98815 5.4591e-005 3.8183 0.011907 0.00011889 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6388 0.61019 0.18619 0.021067 19.6681 0.13035 0.00017133 0.75982 0.0096926 0.010709 0.008989 0.34619 0.13697 2.2731e-005 9.1733e-005 0.16708 0.4581 0.51438 0.0038463 0.50615 0.32739 0.013022 0.41801 1.2611 1.2551 16.0086 144.884 0.00068094 -74.2343 0.054937
9.159 0.98815 5.4591e-005 3.8183 0.011907 0.0001189 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6389 0.61023 0.1862 0.021068 19.6714 0.13036 0.00017134 0.75982 0.0096929 0.01071 0.008145 0.38112 0.15134 2.0369e-005 8.2133e-005 0.16709 0.45958 0.5174 0.0036393 0.5075 0.32757 0.010398 0.41792 1.2637 1.2578 16.0087 144.884 0.00067831 -74.85 0.055937
9.16 0.98815 5.4591e-005 3.8183 0.011907 0.00011892 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.639 0.61028 0.18622 0.021069 19.6747 0.13036 0.00017135 0.75981 0.0096932 0.01071 0.0074131 0.4171 0.16675 1.8349e-005 7.3933e-005 0.16709 0.46108 0.52039 0.0034528 0.50889 0.32776 0.0084423 0.41783 1.2664 1.2605 16.0088 144.884 0.00067568 -75.4362 0.056937
9.161 0.98815 5.4591e-005 3.8183 0.011907 0.00011893 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6391 0.61032 0.18623 0.02107 19.6781 0.13037 0.00017136 0.7598 0.0096936 0.01071 0.0067774 0.45378 0.18318 1.6618e-005 6.6912e-005 0.16709 0.46259 0.52334 0.0032849 0.5103 0.32794 0.0070057 0.41774 1.2691 1.2632 16.009 144.884 0.00067306 -75.9925 0.057937
9.162 0.98815 5.4591e-005 3.8183 0.011907 0.00011894 0.0011779 0.23356 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6392 0.61036 0.18624 0.021071 19.6814 0.13037 0.00017136 0.7598 0.0096939 0.010711 0.0062253 0.4908 0.2006 1.5131e-005 6.0887e-005 0.16709 0.46411 0.52627 0.0031338 0.51176 0.32812 0.0059609 0.41766 1.2718 1.2659 16.0091 144.8839 0.00067045 -76.5189 0.058937
9.163 0.98815 5.4591e-005 3.8183 0.011907 0.00011895 0.0011779 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6393 0.61041 0.18625 0.021072 19.6847 0.13038 0.00017137 0.75979 0.0096942 0.010711 0.0057452 0.52777 0.21897 1.3852e-005 5.5706e-005 0.1671 0.46563 0.52916 0.0029978 0.51325 0.32831 0.0052047 0.41759 1.2745 1.2686 16.0092 144.8839 0.00066784 -77.0151 0.059937
9.164 0.98815 5.4591e-005 3.8183 0.011907 0.00011897 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6393 0.61045 0.18627 0.021073 19.688 0.13039 0.00017138 0.75979 0.0096946 0.010711 0.0053264 0.56431 0.23821 1.2748e-005 5.1241e-005 0.1671 0.46715 0.53201 0.0028755 0.51477 0.3285 0.0046563 0.41752 1.2771 1.2713 16.0093 144.8839 0.00066525 -77.4816 0.060937
9.165 0.98815 5.4591e-005 3.8183 0.011907 0.00011898 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6394 0.6105 0.18628 0.021074 19.6914 0.13039 0.00017139 0.75978 0.0096949 0.010712 0.0049611 0.60006 0.25822 1.1793e-005 4.7383e-005 0.1671 0.46868 0.53484 0.0027655 0.51634 0.32869 0.0042547 0.41745 1.2798 1.274 16.0094 144.8839 0.00066266 -77.9188 0.061937
9.166 0.98815 5.4591e-005 3.8183 0.011907 0.00011899 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6395 0.61054 0.18629 0.021075 19.6947 0.1304 0.0001714 0.75977 0.0096952 0.010712 0.0046421 0.63466 0.27892 1.0967e-005 4.4042e-005 0.1671 0.47021 0.53764 0.0026666 0.51794 0.32888 0.0039553 0.41739 1.2825 1.2767 16.0095 144.8838 0.00066009 -78.3272 0.062937
9.167 0.98815 5.4591e-005 3.8183 0.011907 0.000119 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6396 0.61058 0.18631 0.021076 19.698 0.1304 0.00017141 0.75977 0.0096956 0.010712 0.0043629 0.66781 0.30016 1.0249e-005 4.1142e-005 0.16711 0.47174 0.54041 0.0025778 0.51958 0.32907 0.0037268 0.41733 1.2852 1.2794 16.0097 144.8838 0.00065752 -78.7079 0.063937
9.168 0.98815 5.4591e-005 3.8183 0.011907 0.00011902 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6397 0.61063 0.18632 0.021077 19.7014 0.13041 0.00017142 0.75976 0.0096959 0.010713 0.004118 0.69927 0.32185 9.6233e-006 3.8619e-005 0.16711 0.47327 0.54314 0.0024978 0.52126 0.32926 0.0035475 0.41728 1.2878 1.2821 16.0098 144.8838 0.00065496 -79.0617 0.064937
9.169 0.98815 5.4591e-005 3.8183 0.011907 0.00011903 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6397 0.61067 0.18633 0.021078 19.7047 0.13041 0.00017143 0.75976 0.0096962 0.010713 0.0039029 0.72884 0.34384 9.0777e-006 3.6418e-005 0.16711 0.4748 0.54585 0.002426 0.52297 0.32946 0.0034029 0.41723 1.2905 1.2847 16.0099 144.8838 0.00065242 -79.3898 0.065937
9.17 0.98815 5.459e-005 3.8183 0.011907 0.00011904 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6398 0.61072 0.18634 0.021079 19.708 0.13042 0.00017144 0.75975 0.0096965 0.010713 0.0037137 0.75636 0.36602 8.6005e-006 3.4493e-005 0.16711 0.47634 0.54853 0.0023614 0.52472 0.32966 0.0032831 0.41718 1.2931 1.2874 16.01 144.8838 0.00064988 -79.6935 0.066937
9.171 0.98815 5.459e-005 3.8183 0.011907 0.00011906 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6399 0.61076 0.18636 0.02108 19.7113 0.13043 0.00017145 0.75974 0.0096969 0.010714 0.0035469 0.78177 0.38826 8.1819e-006 3.2806e-005 0.16712 0.47787 0.55118 0.0023032 0.5265 0.32985 0.0031816 0.41713 1.2958 1.2901 16.0101 144.8838 0.00064736 -79.974 0.067937
9.172 0.98815 5.459e-005 3.8183 0.011907 0.00011907 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.64 0.6108 0.18637 0.021081 19.7147 0.13043 0.00017145 0.75974 0.0096972 0.010714 0.0033995 0.80502 0.41047 7.814e-006 3.1324e-005 0.16712 0.4794 0.5538 0.0022509 0.52831 0.33005 0.0030941 0.41709 1.2985 1.2928 16.0103 144.8837 0.00064485 -80.2327 0.068937
9.173 0.98815 5.459e-005 3.8183 0.011907 0.00011908 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6401 0.61085 0.18638 0.021082 19.718 0.13044 0.00017146 0.75973 0.0096975 0.010715 0.0032692 0.82613 0.43253 7.4899e-006 3.0018e-005 0.16712 0.48093 0.5564 0.0022038 0.53016 0.33025 0.0030176 0.41705 1.3011 1.2954 16.0104 144.8837 0.00064235 -80.471 0.069937
9.174 0.98815 5.459e-005 3.8183 0.011907 0.00011909 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032266 0.0389 0 1.6402 0.61089 0.18639 0.021083 19.7213 0.13044 0.00017147 0.75973 0.0096979 0.010715 0.0031536 0.84515 0.45436 7.2037e-006 2.8865e-005 0.16712 0.48245 0.55897 0.0021614 0.53202 0.33045 0.0029504 0.41701 1.3038 1.2981 16.0105 144.8837 0.00063986 -80.6902 0.070937
9.175 0.98815 5.459e-005 3.8183 0.011907 0.00011911 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6402 0.61094 0.18641 0.021084 19.7247 0.13045 0.00017148 0.75972 0.0096982 0.010715 0.0030508 0.86218 0.47587 6.9502e-006 2.7845e-005 0.16713 0.48398 0.56151 0.0021231 0.53392 0.33066 0.0028908 0.41698 1.3064 1.3008 16.0106 144.8837 0.00063739 -80.8917 0.071937
9.176 0.98815 5.459e-005 3.8183 0.011907 0.00011912 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6403 0.61098 0.18642 0.021085 19.728 0.13046 0.00017149 0.75972 0.0096985 0.010716 0.0029592 0.87732 0.497 6.7252e-006 2.694e-005 0.16713 0.4855 0.56402 0.0020885 0.53583 0.33086 0.0028376 0.41694 1.309 1.3034 16.0108 144.8837 0.00063493 -81.0768 0.072937
9.177 0.98815 5.459e-005 3.8183 0.011907 0.00011913 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6404 0.61102 0.18643 0.021086 19.7313 0.13046 0.0001715 0.75971 0.0096988 0.010716 0.0028776 0.8907 0.51768 6.5252e-006 2.6135e-005 0.16713 0.48702 0.56651 0.0020573 0.53777 0.33106 0.0027901 0.41691 1.3117 1.3061 16.0109 144.8837 0.00063248 -81.2468 0.073937
9.178 0.98815 5.459e-005 3.8183 0.011907 0.00011914 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6405 0.61107 0.18645 0.021087 19.7346 0.13047 0.00017151 0.7597 0.0096992 0.010716 0.0028047 0.90247 0.53787 6.3468e-006 2.5417e-005 0.16713 0.48854 0.56898 0.0020291 0.53973 0.33127 0.0027474 0.41688 1.3143 1.3087 16.011 144.8837 0.00063004 -81.4028 0.074937
9.179 0.98815 5.459e-005 3.8183 0.011907 0.00011916 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6406 0.61111 0.18646 0.021088 19.738 0.13047 0.00017152 0.7597 0.0096995 0.010717 0.0027393 0.91276 0.55753 6.1874e-006 2.4776e-005 0.16714 0.49005 0.57141 0.0020035 0.54171 0.33147 0.002709 0.41685 1.317 1.3114 16.0111 144.8837 0.00062762 -81.546 0.075937
9.18 0.98815 5.459e-005 3.8183 0.011907 0.00011917 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6407 0.61116 0.18647 0.021089 19.7413 0.13048 0.00017153 0.75969 0.0096998 0.010717 0.0026804 0.92172 0.57662 6.0444e-006 2.4201e-005 0.16714 0.49156 0.57383 0.0019803 0.5437 0.33168 0.0026745 0.41683 1.3196 1.314 16.0113 144.8837 0.00062521 -81.6775 0.076937
9.181 0.98815 5.459e-005 3.8183 0.011907 0.00011918 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6407 0.6112 0.18648 0.021089 19.7446 0.13049 0.00017154 0.75969 0.0097002 0.010717 0.0026277 0.9295 0.59512 5.9161e-006 2.3685e-005 0.16714 0.49307 0.57621 0.0019593 0.5457 0.33188 0.0026433 0.4168 1.3222 1.3167 16.0114 144.8837 0.00062281 -81.7983 0.077937
9.182 0.98815 5.4589e-005 3.8183 0.011907 0.0001192 0.001178 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6408 0.61125 0.1865 0.02109 19.748 0.13049 0.00017155 0.75968 0.0097005 0.010718 0.0025801 0.93623 0.61302 5.8006e-006 2.3221e-005 0.16714 0.49457 0.57858 0.0019401 0.54772 0.33209 0.0026151 0.41678 1.3248 1.3193 16.0115 144.8837 0.00062042 -81.9093 0.078937
9.183 0.98815 5.4589e-005 3.8183 0.011907 0.00011921 0.0011781 0.23355 0.00065931 0.23421 0.21612 0 0.032267 0.0389 0 1.6409 0.61129 0.18651 0.021091 19.7513 0.1305 0.00017155 0.75967 0.0097008 0.010718 0.0025367 0.94202 0.6303 5.6963e-006 2.2802e-005 0.16715 0.49607 0.58092 0.0019227 0.54974 0.3323 0.0025895 0.41676 1.3275 1.322 16.0117 144.8837 0.00061805 -82.0114 0.079937
9.184 0.98815 5.4589e-005 3.8183 0.011907 0.00011922 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.641 0.61133 0.18652 0.021092 19.7546 0.1305 0.00017156 0.75967 0.0097011 0.010718 0.0024977 0.94701 0.64696 5.6019e-006 2.2423e-005 0.16715 0.49757 0.58323 0.0019068 0.55178 0.33251 0.0025663 0.41673 1.3301 1.3246 16.0118 144.8837 0.0006157 -82.1055 0.080937
9.185 0.98815 5.4589e-005 3.8183 0.011907 0.00011923 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6411 0.61138 0.18654 0.021093 19.758 0.13051 0.00017157 0.75966 0.0097015 0.010719 0.0024621 0.95128 0.66299 5.5163e-006 2.2079e-005 0.16715 0.49906 0.58553 0.0018922 0.55382 0.33272 0.0025451 0.41671 1.3327 1.3272 16.0119 144.8836 0.00061335 -82.1922 0.081937
9.186 0.98815 5.4589e-005 3.8183 0.011907 0.00011925 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6412 0.61142 0.18655 0.021094 19.7613 0.13051 0.00017158 0.75966 0.0097018 0.010719 0.0024297 0.95494 0.67841 5.4384e-006 2.1766e-005 0.16715 0.50055 0.5878 0.0018789 0.55587 0.33293 0.0025258 0.41669 1.3353 1.3299 16.012 144.8836 0.00061102 -82.2723 0.082937
9.187 0.98815 5.4589e-005 3.8183 0.011907 0.00011926 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6412 0.61147 0.18656 0.021095 19.7646 0.13052 0.00017159 0.75965 0.0097021 0.010719 0.0024003 0.95807 0.69322 5.3674e-006 2.148e-005 0.16716 0.50203 0.59004 0.0018666 0.55792 0.33314 0.0025082 0.41667 1.3379 1.3325 16.0121 144.8836 0.0006087 -82.3464 0.083937
9.188 0.98815 5.4589e-005 3.8183 0.011907 0.00011927 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6413 0.61151 0.18657 0.021096 19.768 0.13053 0.0001716 0.75965 0.0097025 0.01072 0.0023732 0.96075 0.70742 5.3024e-006 2.1219e-005 0.16716 0.50351 0.59227 0.0018553 0.55998 0.33334 0.0024921 0.41666 1.3405 1.3351 16.0123 144.8836 0.00060639 -82.415 0.084937
9.189 0.98815 5.4589e-005 3.8183 0.011907 0.00011929 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6414 0.61155 0.18659 0.021097 19.7713 0.13053 0.00017161 0.75964 0.0097028 0.01072 0.0023482 0.96304 0.72102 5.2428e-006 2.098e-005 0.16716 0.50499 0.59447 0.0018449 0.56204 0.33356 0.0024772 0.41664 1.3432 1.3377 16.0124 144.8836 0.0006041 -82.4787 0.085937
9.19 0.98815 5.4589e-005 3.8183 0.011907 0.0001193 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6415 0.6116 0.1866 0.021098 19.7746 0.13054 0.00017162 0.75963 0.0097031 0.01072 0.0023254 0.96499 0.73405 5.1879e-006 2.076e-005 0.16716 0.50646 0.59665 0.0018353 0.56411 0.33377 0.0024635 0.41662 1.3458 1.3404 16.0125 144.8836 0.00060182 -82.538 0.086937
9.191 0.98815 5.4589e-005 3.8183 0.011907 0.00011931 0.0011781 0.23355 0.00065931 0.2342 0.21612 0 0.032267 0.0389 0 1.6416 0.61164 0.18661 0.021099 19.778 0.13054 0.00017163 0.75963 0.0097034 0.010721 0.0023043 0.96666 0.74652 5.1373e-006 2.0557e-005 0.16717 0.50793 0.59881 0.0018264 0.56617 0.33398 0.0024509 0.4166 1.3484 1.343 16.0126 144.8836 0.00059956 -82.5932 0.087937
9.192 0.98815 5.4589e-005 3.8183 0.011907 0.00011932 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6416 0.61169 0.18663 0.0211 19.7813 0.13055 0.00017164 0.75962 0.0097038 0.010721 0.0022847 0.96809 0.75843 5.0905e-006 2.0369e-005 0.16717 0.50939 0.60095 0.0018181 0.56823 0.33419 0.0024392 0.41659 1.3509 1.3456 16.0128 144.8836 0.0005973 -82.6448 0.088937
9.193 0.98815 5.4589e-005 3.8183 0.011907 0.00011934 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6417 0.61173 0.18664 0.021101 19.7846 0.13056 0.00017164 0.75962 0.0097041 0.010721 0.0022665 0.96932 0.76981 5.047e-006 2.0195e-005 0.16717 0.51085 0.60307 0.0018104 0.5703 0.3344 0.0024284 0.41657 1.3535 1.3482 16.0129 144.8836 0.00059506 -82.6932 0.089937
9.194 0.98815 5.4588e-005 3.8183 0.011907 0.00011935 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6418 0.61177 0.18665 0.021102 19.788 0.13056 0.00017165 0.75961 0.0097044 0.010722 0.0022495 0.97037 0.78068 5.0066e-006 2.0032e-005 0.16717 0.51231 0.60517 0.0018032 0.57236 0.33461 0.0024183 0.41656 1.3561 1.3508 16.013 144.8836 0.00059284 -82.7385 0.090937
9.195 0.98815 5.4588e-005 3.8183 0.011907 0.00011936 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6419 0.61182 0.18666 0.021103 19.7913 0.13057 0.00017166 0.7596 0.0097048 0.010722 0.0022337 0.97128 0.79105 4.9688e-006 1.9881e-005 0.16718 0.51376 0.60724 0.0017964 0.57443 0.33482 0.0024088 0.41655 1.3587 1.3534 16.0131 144.8836 0.00059062 -82.7812 0.091937
9.196 0.98815 5.4588e-005 3.8183 0.011907 0.00011937 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.642 0.61186 0.18668 0.021104 19.7946 0.13057 0.00017167 0.7596 0.0097051 0.010723 0.0022188 0.97206 0.80093 4.9334e-006 1.9739e-005 0.16718 0.51521 0.6093 0.00179 0.57649 0.33503 0.0024 0.41653 1.3613 1.356 16.0132 144.8836 0.00058842 -82.8215 0.092937
9.197 0.98815 5.4588e-005 3.8183 0.011906 0.00011939 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6421 0.61191 0.18669 0.021105 19.798 0.13058 0.00017168 0.75959 0.0097054 0.010723 0.0022049 0.97274 0.81036 4.9002e-006 1.9606e-005 0.16718 0.51665 0.61134 0.001784 0.57855 0.33525 0.0023917 0.41652 1.3639 1.3586 16.0134 144.8836 0.00058623 -82.8597 0.093937
9.198 0.98815 5.4588e-005 3.8183 0.011906 0.0001194 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6421 0.61195 0.1867 0.021106 19.8013 0.13058 0.00017169 0.75959 0.0097057 0.010723 0.0021917 0.97333 0.81934 4.8689e-006 1.948e-005 0.16718 0.51809 0.61335 0.0017784 0.5806 0.33546 0.0023839 0.41651 1.3665 1.3612 16.0135 144.8836 0.00058405 -82.8958 0.094937
9.199 0.98815 5.4588e-005 3.8183 0.011906 0.00011941 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6422 0.61199 0.18672 0.021107 19.8046 0.13059 0.0001717 0.75958 0.0097061 0.010724 0.0021793 0.97385 0.8279 4.8393e-006 1.9361e-005 0.16719 0.51952 0.61535 0.001773 0.58265 0.33567 0.0023765 0.41649 1.369 1.3638 16.0136 144.8836 0.00058189 -82.9302 0.095937
9.2 0.98815 5.4588e-005 3.8183 0.011906 0.00011943 0.0011781 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6423 0.61204 0.18673 0.021108 19.808 0.1306 0.00017171 0.75958 0.0097064 0.010724 0.0021675 0.9743 0.83604 4.8112e-006 1.9249e-005 0.16719 0.52095 0.61733 0.0017679 0.5847 0.33588 0.0023695 0.41648 1.3716 1.3664 16.0137 144.8836 0.00057974 -82.963 0.096937
9.201 0.98815 5.4588e-005 3.8183 0.011906 0.00011944 0.0011782 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6424 0.61208 0.18674 0.021109 19.8113 0.1306 0.00017172 0.75957 0.0097067 0.010724 0.0021563 0.9747 0.8438 4.7846e-006 1.9142e-005 0.16719 0.52238 0.61929 0.001763 0.58675 0.3361 0.0023629 0.41647 1.3742 1.3689 16.0138 144.8836 0.0005776 -82.9943 0.097937
9.202 0.98815 5.4588e-005 3.8183 0.011906 0.00011945 0.0011782 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6425 0.61213 0.18675 0.02111 19.8147 0.13061 0.00017173 0.75956 0.009707 0.010725 0.0021456 0.97506 0.85117 4.7592e-006 1.9041e-005 0.16719 0.5238 0.62124 0.0017584 0.58879 0.33631 0.0023566 0.41646 1.3767 1.3715 16.0139 144.8836 0.00057547 -83.0243 0.098937
9.203 0.98815 5.4588e-005 3.8183 0.011906 0.00011946 0.0011782 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6426 0.61217 0.18677 0.021111 19.818 0.13061 0.00017173 0.75956 0.0097074 0.010725 0.0021354 0.97537 0.85819 4.735e-006 1.8944e-005 0.1672 0.52522 0.62316 0.001754 0.59082 0.33652 0.0023506 0.41645 1.3793 1.3741 16.014 144.8836 0.00057336 -83.0531 0.099937
9.204 0.98815 5.4588e-005 3.8183 0.011906 0.00011948 0.0011782 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6426 0.61222 0.18678 0.021112 19.8213 0.13062 0.00017174 0.75955 0.0097077 0.010725 0.0021256 0.97565 0.86486 4.7118e-006 1.8851e-005 0.1672 0.52664 0.62506 0.0017497 0.59285 0.33673 0.0023448 0.41644 1.3819 1.3767 16.0142 144.8836 0.00057125 -83.0808 0.10094
9.205 0.98815 5.4587e-005 3.8183 0.011906 0.00011949 0.0011782 0.23355 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6427 0.61226 0.18679 0.021113 19.8247 0.13063 0.00017175 0.75955 0.009708 0.010726 0.0021162 0.97591 0.87121 4.6895e-006 1.8761e-005 0.1672 0.52805 0.62695 0.0017456 0.59488 0.33695 0.0023392 0.41643 1.3844 1.3792 16.0143 144.8836 0.00056916 -83.1075 0.10194
9.206 0.98815 5.4587e-005 3.8183 0.011906 0.0001195 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6428 0.6123 0.18681 0.021114 19.828 0.13063 0.00017176 0.75954 0.0097084 0.010726 0.0021072 0.97614 0.87724 4.6681e-006 1.8676e-005 0.1672 0.52945 0.62882 0.0017416 0.5969 0.33716 0.0023339 0.41642 1.387 1.3818 16.0144 144.8837 0.00056708 -83.1334 0.10294
9.207 0.98815 5.4587e-005 3.8183 0.011906 0.00011952 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6429 0.61235 0.18682 0.021115 19.8314 0.13064 0.00017177 0.75953 0.0097087 0.010726 0.0020985 0.97636 0.88297 4.6475e-006 1.8593e-005 0.16721 0.53085 0.63068 0.0017378 0.59892 0.33737 0.0023288 0.41641 1.3895 1.3844 16.0145 144.8837 0.00056502 -83.1584 0.10394
9.208 0.98815 5.4587e-005 3.8183 0.011906 0.00011953 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.643 0.61239 0.18683 0.021116 19.8347 0.13064 0.00017178 0.75953 0.009709 0.010727 0.0020901 0.97655 0.88842 4.6275e-006 1.8513e-005 0.16721 0.53225 0.63251 0.0017341 0.60093 0.33759 0.0023238 0.4164 1.3921 1.3869 16.0146 144.8837 0.00056296 -83.1827 0.10494
9.209 0.98815 5.4587e-005 3.8183 0.011906 0.00011954 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.643 0.61244 0.18684 0.021117 19.838 0.13065 0.00017179 0.75952 0.0097093 0.010727 0.0020819 0.97674 0.89359 4.6082e-006 1.8436e-005 0.16721 0.53364 0.63433 0.0017305 0.60294 0.3378 0.002319 0.41639 1.3946 1.3895 16.0147 144.8837 0.00056092 -83.2063 0.10594
9.21 0.98815 5.4587e-005 3.8183 0.011906 0.00011955 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6431 0.61248 0.18686 0.021118 19.8414 0.13065 0.0001718 0.75952 0.0097097 0.010727 0.002074 0.9769 0.8985 4.5895e-006 1.8361e-005 0.16721 0.53503 0.63613 0.0017271 0.60494 0.33801 0.0023144 0.41638 1.3971 1.392 16.0148 144.8837 0.00055889 -83.2292 0.10694
9.211 0.98815 5.4587e-005 3.8183 0.011906 0.00011957 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6432 0.61252 0.18687 0.021119 19.8447 0.13066 0.00017181 0.75951 0.00971 0.010728 0.0020663 0.97706 0.90317 4.5714e-006 1.8288e-005 0.16722 0.53642 0.63792 0.0017237 0.60693 0.33823 0.0023099 0.41637 1.3997 1.3946 16.0149 144.8837 0.00055687 -83.2516 0.10794
9.212 0.98815 5.4587e-005 3.8183 0.011906 0.00011958 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6433 0.61257 0.18688 0.02112 19.8481 0.13067 0.00017182 0.75951 0.0097103 0.010728 0.0020588 0.97721 0.9076 4.5537e-006 1.8217e-005 0.16722 0.5378 0.63969 0.0017204 0.60892 0.33844 0.0023055 0.41636 1.4022 1.3971 16.015 144.8837 0.00055486 -83.2735 0.10894
9.213 0.98815 5.4587e-005 3.8183 0.011906 0.00011959 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6434 0.61261 0.18689 0.021121 19.8514 0.13067 0.00017182 0.7595 0.0097106 0.010728 0.0020516 0.97735 0.9118 4.5365e-006 1.8148e-005 0.16722 0.53917 0.64144 0.0017171 0.6109 0.33865 0.0023012 0.41635 1.4047 1.3997 16.0151 144.8837 0.00055286 -83.2949 0.10994
9.214 0.98815 5.4587e-005 3.8183 0.011906 0.0001196 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6435 0.61266 0.18691 0.021122 19.8547 0.13068 0.00017183 0.75949 0.009711 0.010729 0.0020445 0.97749 0.9158 4.5197e-006 1.8081e-005 0.16722 0.54055 0.64318 0.001714 0.61288 0.33887 0.002297 0.41635 1.4072 1.4022 16.0153 144.8837 0.00055088 -83.3158 0.11094
9.215 0.98815 5.4587e-005 3.8183 0.011906 0.00011962 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6435 0.6127 0.18692 0.021123 19.8581 0.13068 0.00017184 0.75949 0.0097113 0.010729 0.0020375 0.97761 0.91958 4.5033e-006 1.8015e-005 0.16723 0.54192 0.6449 0.0017109 0.61485 0.33908 0.002293 0.41634 1.4098 1.4048 16.0154 144.8837 0.0005489 -83.3364 0.11194
9.216 0.98815 5.4587e-005 3.8183 0.011906 0.00011963 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6436 0.61274 0.18693 0.021124 19.8614 0.13069 0.00017185 0.75948 0.0097116 0.010729 0.0020307 0.97773 0.92318 4.4873e-006 1.7951e-005 0.16723 0.54328 0.64661 0.0017079 0.61681 0.3393 0.002289 0.41633 1.4123 1.4073 16.0155 144.8837 0.00054694 -83.3565 0.11294
9.217 0.98815 5.4586e-005 3.8183 0.011906 0.00011964 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6437 0.61279 0.18695 0.021125 19.8648 0.1307 0.00017186 0.75948 0.009712 0.01073 0.0020241 0.97785 0.92659 4.4716e-006 1.7888e-005 0.16723 0.54464 0.6483 0.0017049 0.61877 0.33951 0.0022851 0.41632 1.4148 1.4098 16.0156 144.8837 0.00054499 -83.3763 0.11394
9.218 0.98815 5.4586e-005 3.8183 0.011906 0.00011966 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6438 0.61283 0.18696 0.021126 19.8681 0.1307 0.00017187 0.75947 0.0097123 0.01073 0.0020176 0.97796 0.92983 4.4562e-006 1.7827e-005 0.16723 0.546 0.64998 0.001702 0.62072 0.33972 0.0022812 0.41632 1.4173 1.4123 16.0157 144.8837 0.00054305 -83.3957 0.11494
9.219 0.98815 5.4586e-005 3.8183 0.011906 0.00011967 0.0011782 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6439 0.61288 0.18697 0.021127 19.8715 0.13071 0.00017188 0.75946 0.0097126 0.01073 0.0020112 0.97807 0.9329 4.4412e-006 1.7767e-005 0.16724 0.54735 0.65164 0.0016992 0.62267 0.33994 0.0022775 0.41631 1.4198 1.4149 16.0158 144.8837 0.00054112 -83.4148 0.11594
9.22 0.98815 5.4586e-005 3.8183 0.011906 0.00011968 0.0011783 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.644 0.61292 0.18698 0.021128 19.8748 0.13071 0.00017189 0.75946 0.0097129 0.010731 0.0020049 0.97818 0.93581 4.4264e-006 1.7708e-005 0.16724 0.5487 0.65329 0.0016964 0.62461 0.34015 0.0022738 0.4163 1.4223 1.4174 16.0159 144.8837 0.0005392 -83.4336 0.11694
9.221 0.98815 5.4586e-005 3.8183 0.011906 0.00011969 0.0011783 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.644 0.61296 0.187 0.021129 19.8781 0.13072 0.0001719 0.75945 0.0097133 0.010731 0.0019988 0.97828 0.93857 4.4119e-006 1.765e-005 0.16724 0.55004 0.65492 0.0016936 0.62654 0.34037 0.0022702 0.4163 1.4248 1.4199 16.016 144.8837 0.00053729 -83.4522 0.11794
9.222 0.98815 5.4586e-005 3.8183 0.011906 0.00011971 0.0011783 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6441 0.61301 0.18701 0.02113 19.8815 0.13072 0.00017191 0.75945 0.0097136 0.010731 0.0019927 0.97838 0.94119 4.3976e-006 1.7592e-005 0.16724 0.55138 0.65654 0.0016909 0.62846 0.34058 0.0022666 0.41629 1.4273 1.4224 16.0161 144.8837 0.00053539 -83.4705 0.11894
9.223 0.98815 5.4586e-005 3.8183 0.011906 0.00011972 0.0011783 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6442 0.61305 0.18702 0.021131 19.8848 0.13073 0.00017191 0.75944 0.0097139 0.010732 0.0019868 0.97847 0.94368 4.3836e-006 1.7536e-005 0.16725 0.55272 0.65814 0.0016883 0.63038 0.34079 0.0022631 0.41628 1.4298 1.4249 16.0162 144.8837 0.00053351 -83.4885 0.11994
9.224 0.98815 5.4586e-005 3.8183 0.011906 0.00011973 0.0011783 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6443 0.6131 0.18704 0.021132 19.8882 0.13074 0.00017192 0.75944 0.0097142 0.010732 0.0019809 0.97857 0.94603 4.3698e-006 1.7481e-005 0.16725 0.55405 0.65973 0.0016856 0.63229 0.34101 0.0022597 0.41628 1.4323 1.4274 16.0163 144.8837 0.00053163 -83.5063 0.12094
9.225 0.98815 5.4586e-005 3.8183 0.011906 0.00011974 0.0011783 0.23354 0.00065931 0.2342 0.21611 0 0.032267 0.0389 0 1.6444 0.61314 0.18705 0.021133 19.8915 0.13074 0.00017193 0.75943 0.0097146 0.010733 0.0019752 0.97866 0.94826 4.3562e-006 1.7427e-005 0.16725 0.55537 0.66131 0.001683 0.6342 0.34122 0.0022563 0.41627 1.4348 1.4299 16.0164 144.8837 0.00052977 -83.5238 0.12194
9.226 0.98815 5.4586e-005 3.8183 0.011906 0.00011976 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6445 0.61318 0.18706 0.021134 19.8949 0.13075 0.00017194 0.75942 0.0097149 0.010733 0.0019695 0.97875 0.95038 4.3429e-006 1.7373e-005 0.16725 0.5567 0.66287 0.0016805 0.6361 0.34144 0.0022529 0.41627 1.4373 1.4324 16.0165 144.8837 0.00052791 -83.5412 0.12294
9.227 0.98815 5.4586e-005 3.8183 0.011906 0.00011977 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6445 0.61323 0.18707 0.021135 19.8982 0.13075 0.00017195 0.75942 0.0097152 0.010733 0.0019639 0.97883 0.95239 4.3297e-006 1.7321e-005 0.16726 0.55802 0.66442 0.001678 0.63799 0.34165 0.0022496 0.41626 1.4397 1.4349 16.0166 144.8837 0.00052607 -83.5584 0.12394
9.228 0.98815 5.4586e-005 3.8183 0.011906 0.00011978 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6446 0.61327 0.18709 0.021136 19.9016 0.13076 0.00017196 0.75941 0.0097155 0.010734 0.0019584 0.97892 0.95429 4.3168e-006 1.7269e-005 0.16726 0.55933 0.66595 0.0016755 0.63988 0.34187 0.0022463 0.41626 1.4422 1.4374 16.0167 144.8837 0.00052423 -83.5753 0.12494
9.229 0.98816 5.4585e-005 3.8183 0.011906 0.0001198 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6447 0.61332 0.1871 0.021137 19.9049 0.13077 0.00017197 0.75941 0.0097159 0.010734 0.0019529 0.97901 0.9561 4.304e-006 1.7218e-005 0.16726 0.56065 0.66748 0.001673 0.64176 0.34208 0.0022431 0.41625 1.4447 1.4399 16.0168 144.8837 0.00052241 -83.5921 0.12594
9.23 0.98816 5.4585e-005 3.8183 0.011906 0.00011981 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6448 0.61336 0.18711 0.021138 19.9083 0.13077 0.00017198 0.7594 0.0097162 0.010734 0.0019476 0.97909 0.95781 4.2914e-006 1.7167e-005 0.16726 0.56195 0.66899 0.0016706 0.64363 0.3423 0.0022399 0.41625 1.4471 1.4424 16.0169 144.8837 0.00052059 -83.6087 0.12694
9.231 0.98816 5.4585e-005 3.8183 0.011906 0.00011982 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6449 0.61341 0.18712 0.021139 19.9116 0.13078 0.00017199 0.75939 0.0097165 0.010735 0.0019423 0.97917 0.95943 4.2789e-006 1.7117e-005 0.16727 0.56326 0.67048 0.0016682 0.64549 0.34251 0.0022368 0.41624 1.4496 1.4448 16.017 144.8838 0.00051879 -83.6251 0.12794
9.232 0.98816 5.4585e-005 3.8183 0.011906 0.00011983 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6449 0.61345 0.18714 0.02114 19.9149 0.13078 0.000172 0.75939 0.0097169 0.010735 0.0019371 0.97925 0.96097 4.2667e-006 1.7068e-005 0.16727 0.56456 0.67197 0.0016658 0.64735 0.34273 0.0022337 0.41624 1.4521 1.4473 16.0171 144.8838 0.000517 -83.6413 0.12894
9.233 0.98816 5.4585e-005 3.8183 0.011906 0.00011985 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.645 0.61349 0.18715 0.021141 19.9183 0.13079 0.000172 0.75938 0.0097172 0.010735 0.0019319 0.97933 0.96242 4.2545e-006 1.702e-005 0.16727 0.56585 0.67344 0.0016635 0.6492 0.34294 0.0022306 0.41623 1.4545 1.4498 16.0172 144.8838 0.00051521 -83.6574 0.12994
9.234 0.98816 5.4585e-005 3.8183 0.011906 0.00011986 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6451 0.61354 0.18716 0.021142 19.9216 0.13079 0.00017201 0.75938 0.0097175 0.010736 0.0019268 0.97941 0.9638 4.2426e-006 1.6972e-005 0.16727 0.56715 0.6749 0.0016612 0.65105 0.34315 0.0022276 0.41623 1.457 1.4522 16.0173 144.8838 0.00051344 -83.6733 0.13094
9.235 0.98816 5.4585e-005 3.8183 0.011906 0.00011987 0.0011783 0.23354 0.00065931 0.23419 0.21611 0 0.032267 0.0389 0 1.6452 0.61358 0.18718 0.021143 19.925 0.1308 0.00017202 0.75937 0.0097178 0.010736 0.0019218 0.97948 0.96511 4.2308e-006 1.6925e-005 0.16728 0.56843 0.67635 0.0016589 0.65289 0.34337 0.0022246 0.41623 1.4594 1.4547 16.0174 144.8838 0.00051167 -83.689 0.13194
9.236 0.98816 5.4585e-005 3.8183 0.011906 0.00011989 0.0011783 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6453 0.61363 0.18719 0.021144 19.9283 0.13081 0.00017203 0.75937 0.0097182 0.010736 0.0019168 0.97956 0.96635 4.2191e-006 1.6878e-005 0.16728 0.56972 0.67778 0.0016566 0.65472 0.34358 0.0022216 0.41622 1.4619 1.4572 16.0175 144.8838 0.00050992 -83.7046 0.13294
9.237 0.98816 5.4585e-005 3.8183 0.011906 0.0001199 0.0011783 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6454 0.61367 0.1872 0.021145 19.9317 0.13081 0.00017204 0.75936 0.0097185 0.010737 0.0019119 0.97963 0.96753 4.2076e-006 1.6832e-005 0.16728 0.571 0.6792 0.0016544 0.65654 0.3438 0.0022187 0.41622 1.4643 1.4596 16.0175 144.8838 0.00050817 -83.7201 0.13394
9.238 0.98816 5.4585e-005 3.8183 0.011906 0.00011991 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6454 0.61371 0.18721 0.021146 19.935 0.13082 0.00017205 0.75935 0.0097188 0.010737 0.0019071 0.9797 0.96864 4.1962e-006 1.6786e-005 0.16728 0.57227 0.68062 0.0016522 0.65836 0.34401 0.0022158 0.41622 1.4667 1.4621 16.0176 144.8838 0.00050644 -83.7354 0.13494
9.239 0.98816 5.4585e-005 3.8183 0.011906 0.00011992 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6455 0.61376 0.18723 0.021147 19.9384 0.13082 0.00017206 0.75935 0.0097191 0.010737 0.0019023 0.97978 0.96969 4.185e-006 1.6741e-005 0.16729 0.57355 0.68202 0.00165 0.66017 0.34423 0.0022129 0.41621 1.4692 1.4645 16.0177 144.8838 0.00050471 -83.7505 0.13594
9.24 0.98816 5.4585e-005 3.8183 0.011906 0.00011994 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6456 0.6138 0.18724 0.021148 19.9417 0.13083 0.00017207 0.75934 0.0097195 0.010738 0.0018975 0.97985 0.97069 4.1738e-006 1.6697e-005 0.16729 0.57482 0.6834 0.0016478 0.66197 0.34444 0.0022101 0.41621 1.4716 1.4669 16.0178 144.8838 0.000503 -83.7655 0.13694
9.241 0.98816 5.4584e-005 3.8183 0.011906 0.00011995 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6457 0.61385 0.18725 0.021149 19.9451 0.13084 0.00017208 0.75934 0.0097198 0.010738 0.0018929 0.97992 0.97164 4.1629e-006 1.6653e-005 0.16729 0.57608 0.68478 0.0016457 0.66377 0.34466 0.0022073 0.41621 1.474 1.4694 16.0179 144.8838 0.00050129 -83.7804 0.13794
9.242 0.98816 5.4584e-005 3.8183 0.011906 0.00011996 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6458 0.61389 0.18727 0.02115 19.9484 0.13084 0.00017208 0.75933 0.0097201 0.010738 0.0018882 0.97998 0.97254 4.152e-006 1.6609e-005 0.16729 0.57734 0.68615 0.0016436 0.66556 0.34487 0.0022045 0.4162 1.4764 1.4718 16.018 144.8838 0.00049959 -83.7952 0.13894
9.243 0.98816 5.4584e-005 3.8183 0.011906 0.00011997 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6459 0.61393 0.18728 0.021151 19.9518 0.13085 0.00017209 0.75932 0.0097204 0.010739 0.0018837 0.98005 0.97339 4.1413e-006 1.6567e-005 0.1673 0.5786 0.6875 0.0016415 0.66734 0.34509 0.0022018 0.4162 1.4788 1.4742 16.0181 144.8838 0.00049791 -83.8098 0.13994
9.244 0.98816 5.4584e-005 3.8183 0.011906 0.00011999 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6459 0.61398 0.18729 0.021152 19.9551 0.13085 0.0001721 0.75932 0.0097208 0.010739 0.0018791 0.98012 0.97419 4.1307e-006 1.6524e-005 0.1673 0.57985 0.68885 0.0016394 0.66911 0.3453 0.002199 0.4162 1.4813 1.4767 16.0182 144.8838 0.00049623 -83.8243 0.14094
9.245 0.98816 5.4584e-005 3.8183 0.011906 0.00012 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.646 0.61402 0.1873 0.021153 19.9585 0.13086 0.00017211 0.75931 0.0097211 0.010739 0.0018747 0.98019 0.97496 4.1202e-006 1.6482e-005 0.1673 0.5811 0.69018 0.0016373 0.67088 0.34552 0.0021964 0.4162 1.4837 1.4791 16.0183 144.8838 0.00049456 -83.8386 0.14194
9.246 0.98816 5.4584e-005 3.8183 0.011906 0.00012001 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6461 0.61407 0.18732 0.021154 19.9618 0.13086 0.00017212 0.75931 0.0097214 0.01074 0.0018702 0.98025 0.97568 4.1098e-006 1.6441e-005 0.1673 0.58235 0.6915 0.0016353 0.67264 0.34573 0.0021937 0.4162 1.4861 1.4815 16.0184 144.8839 0.0004929 -83.8528 0.14294
9.247 0.98816 5.4584e-005 3.8183 0.011906 0.00012003 0.0011784 0.23354 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6462 0.61411 0.18733 0.021155 19.9652 0.13087 0.00017213 0.7593 0.0097217 0.01074 0.0018659 0.98032 0.97637 4.0996e-006 1.64e-005 0.16731 0.58359 0.69281 0.0016333 0.6744 0.34595 0.0021911 0.41619 1.4885 1.4839 16.0184 144.8839 0.00049125 -83.8669 0.14394
9.248 0.98816 5.4584e-005 3.8183 0.011906 0.00012004 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6463 0.61415 0.18734 0.021156 19.9685 0.13088 0.00017214 0.7593 0.0097221 0.01074 0.0018615 0.98038 0.97702 4.0895e-006 1.6359e-005 0.16731 0.58483 0.69411 0.0016313 0.67614 0.34616 0.0021884 0.41619 1.4909 1.4863 16.0185 144.8839 0.0004896 -83.8809 0.14494
9.249 0.98816 5.4584e-005 3.8183 0.011906 0.00012005 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6463 0.6142 0.18735 0.021157 19.9719 0.13088 0.00017215 0.75929 0.0097224 0.010741 0.0018573 0.98044 0.97764 4.0794e-006 1.6319e-005 0.16731 0.58606 0.6954 0.0016293 0.67788 0.34638 0.0021859 0.41619 1.4933 1.4887 16.0186 144.8839 0.00048797 -83.8948 0.14594
9.25 0.98816 5.4584e-005 3.8183 0.011906 0.00012006 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6464 0.61424 0.18737 0.021158 19.9753 0.13089 0.00017216 0.75928 0.0097227 0.010741 0.001853 0.98051 0.97822 4.0695e-006 1.6279e-005 0.16731 0.58729 0.69668 0.0016273 0.67962 0.34659 0.0021833 0.41619 1.4956 1.4911 16.0187 144.8839 0.00048635 -83.9085 0.14694
9.251 0.98816 5.4584e-005 3.8183 0.011905 0.00012008 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6465 0.61429 0.18738 0.021159 19.9786 0.13089 0.00017217 0.75928 0.009723 0.010741 0.0018488 0.98057 0.97877 4.0597e-006 1.624e-005 0.16732 0.58852 0.69795 0.0016254 0.68134 0.34681 0.0021808 0.41619 1.498 1.4935 16.0188 144.8839 0.00048473 -83.9222 0.14794
9.252 0.98816 5.4584e-005 3.8183 0.011905 0.00012009 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6466 0.61433 0.18739 0.02116 19.982 0.1309 0.00017217 0.75927 0.0097234 0.010742 0.0018447 0.98063 0.9793 4.05e-006 1.6201e-005 0.16732 0.58974 0.69921 0.0016235 0.68306 0.34703 0.0021782 0.41619 1.5004 1.4959 16.0189 144.8839 0.00048312 -83.9357 0.14894
9.253 0.98816 5.4583e-005 3.8183 0.011905 0.0001201 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6467 0.61437 0.18741 0.02116 19.9853 0.13091 0.00017218 0.75927 0.0097237 0.010742 0.0018406 0.98069 0.9798 4.0404e-006 1.6163e-005 0.16732 0.59096 0.70046 0.0016216 0.68477 0.34724 0.0021758 0.41619 1.5028 1.4983 16.019 144.8839 0.00048153 -83.9491 0.14994
9.254 0.98816 5.4583e-005 3.8183 0.011905 0.00012012 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6468 0.61442 0.18742 0.021161 19.9887 0.13091 0.00017219 0.75926 0.009724 0.010742 0.0018365 0.98075 0.98027 4.0309e-006 1.6125e-005 0.16732 0.59218 0.70171 0.0016197 0.68648 0.34746 0.0021733 0.41619 1.5052 1.5007 16.019 144.8839 0.00047994 -83.9624 0.15094
9.255 0.98816 5.4583e-005 3.8183 0.011905 0.00012013 0.0011784 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6468 0.61446 0.18743 0.021162 19.992 0.13092 0.0001722 0.75926 0.0097243 0.010743 0.0018325 0.98081 0.98072 4.0215e-006 1.6087e-005 0.16733 0.59339 0.70294 0.0016178 0.68817 0.34767 0.0021709 0.41619 1.5075 1.5031 16.0191 144.8839 0.00047836 -83.9756 0.15194
9.256 0.98816 5.4583e-005 3.8183 0.011905 0.00012014 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6469 0.61451 0.18744 0.021163 19.9954 0.13092 0.00017221 0.75925 0.0097247 0.010743 0.0018286 0.98087 0.98114 4.0123e-006 1.605e-005 0.16733 0.5946 0.70416 0.001616 0.68987 0.34789 0.0021684 0.41619 1.5099 1.5055 16.0192 144.8839 0.00047678 -83.9886 0.15294
9.257 0.98816 5.4583e-005 3.8183 0.011905 0.00012015 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.647 0.61455 0.18746 0.021164 19.9987 0.13093 0.00017222 0.75924 0.009725 0.010743 0.0018246 0.98092 0.98154 4.0031e-006 1.6013e-005 0.16733 0.5958 0.70537 0.0016141 0.69155 0.3481 0.002166 0.41619 1.5123 1.5079 16.0193 144.8839 0.00047522 -84.0016 0.15394
9.258 0.98816 5.4583e-005 3.8183 0.011905 0.00012017 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032267 0.0389 0 1.6471 0.61459 0.18747 0.021165 20.0021 0.13093 0.00017223 0.75924 0.0097253 0.010744 0.0018207 0.98098 0.98193 3.994e-006 1.5977e-005 0.16733 0.597 0.70657 0.0016123 0.69323 0.34832 0.0021637 0.41619 1.5146 1.5102 16.0194 144.8839 0.00047366 -84.0144 0.15494
9.259 0.98816 5.4583e-005 3.8183 0.011905 0.00012018 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6472 0.61464 0.18748 0.021166 20.0054 0.13094 0.00017224 0.75923 0.0097256 0.010744 0.0018169 0.98104 0.98229 3.985e-006 1.5941e-005 0.16734 0.5982 0.70777 0.0016105 0.6949 0.34853 0.0021613 0.41619 1.517 1.5126 16.0195 144.884 0.00047212 -84.0272 0.15594
9.26 0.98816 5.4583e-005 3.8183 0.011905 0.00012019 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6473 0.61468 0.1875 0.021167 20.0088 0.13095 0.00017225 0.75923 0.009726 0.010745 0.0018131 0.98109 0.98263 3.9761e-006 1.5905e-005 0.16734 0.5994 0.70895 0.0016087 0.69656 0.34875 0.002159 0.41619 1.5193 1.5149 16.0195 144.884 0.00047058 -84.0398 0.15694
9.261 0.98816 5.4583e-005 3.8183 0.011905 0.0001202 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6473 0.61473 0.18751 0.021168 20.0122 0.13095 0.00017226 0.75922 0.0097263 0.010745 0.0018093 0.98115 0.98296 3.9673e-006 1.587e-005 0.16734 0.60059 0.71012 0.001607 0.69821 0.34896 0.0021567 0.41619 1.5216 1.5173 16.0196 144.884 0.00046905 -84.0523 0.15794
9.262 0.98816 5.4583e-005 3.8183 0.011905 0.00012022 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6474 0.61477 0.18752 0.021169 20.0155 0.13096 0.00017226 0.75921 0.0097266 0.010745 0.0018056 0.9812 0.98327 3.9586e-006 1.5835e-005 0.16734 0.60177 0.71129 0.0016052 0.69986 0.34918 0.0021544 0.41619 1.524 1.5197 16.0197 144.884 0.00046752 -84.0648 0.15894
9.263 0.98816 5.4583e-005 3.8183 0.011905 0.00012023 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6475 0.61481 0.18753 0.02117 20.0189 0.13096 0.00017227 0.75921 0.0097269 0.010746 0.0018019 0.98125 0.98356 3.9499e-006 1.5801e-005 0.16735 0.60296 0.71245 0.0016035 0.7015 0.34939 0.0021521 0.41619 1.5263 1.522 16.0198 144.884 0.00046601 -84.0771 0.15994
9.264 0.98816 5.4582e-005 3.8183 0.011905 0.00012024 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6476 0.61486 0.18755 0.021171 20.0222 0.13097 0.00017228 0.7592 0.0097273 0.010746 0.0017982 0.98131 0.98384 3.9414e-006 1.5767e-005 0.16735 0.60413 0.7136 0.0016018 0.70314 0.34961 0.0021499 0.41619 1.5287 1.5244 16.0199 144.884 0.0004645 -84.0893 0.16094
9.265 0.98816 5.4582e-005 3.8183 0.011905 0.00012026 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6477 0.6149 0.18756 0.021172 20.0256 0.13098 0.00017229 0.7592 0.0097276 0.010746 0.0017946 0.98136 0.98411 3.9329e-006 1.5733e-005 0.16735 0.60531 0.71474 0.0016001 0.70476 0.34982 0.0021477 0.41619 1.531 1.5267 16.0199 144.884 0.00046301 -84.1014 0.16194
9.266 0.98816 5.4582e-005 3.8183 0.011905 0.00012027 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6477 0.61495 0.18757 0.021173 20.029 0.13098 0.0001723 0.75919 0.0097279 0.010747 0.001791 0.98141 0.98436 3.9246e-006 1.5699e-005 0.16735 0.60648 0.71587 0.0015984 0.70638 0.35004 0.0021455 0.41619 1.5333 1.529 16.02 144.884 0.00046152 -84.1135 0.16294
9.267 0.98816 5.4582e-005 3.8183 0.011905 0.00012028 0.0011785 0.23353 0.00065931 0.23419 0.2161 0 0.032268 0.0389 0 1.6478 0.61499 0.18758 0.021174 20.0323 0.13099 0.00017231 0.75919 0.0097282 0.010747 0.0017875 0.98146 0.9846 3.9163e-006 1.5666e-005 0.16736 0.60765 0.71699 0.0015967 0.708 0.35026 0.0021433 0.41619 1.5356 1.5314 16.0201 144.884 0.00046003 -84.1254 0.16394
9.268 0.98816 5.4582e-005 3.8183 0.011905 0.00012029 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6479 0.61504 0.1876 0.021175 20.0357 0.13099 0.00017232 0.75918 0.0097286 0.010747 0.001784 0.98151 0.98483 3.9081e-006 1.5633e-005 0.16736 0.60882 0.71811 0.0015951 0.7096 0.35047 0.0021411 0.41619 1.5379 1.5337 16.0202 144.884 0.00045856 -84.1372 0.16494
9.269 0.98816 5.4582e-005 3.8183 0.011905 0.00012031 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.648 0.61508 0.18761 0.021176 20.039 0.131 0.00017233 0.75917 0.0097289 0.010748 0.0017805 0.98156 0.98505 3.9e-006 1.5601e-005 0.16736 0.60998 0.71921 0.0015934 0.7112 0.35069 0.002139 0.41619 1.5402 1.536 16.0202 144.884 0.00045709 -84.149 0.16594
9.27 0.98816 5.4582e-005 3.8183 0.011905 0.00012032 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6481 0.61512 0.18762 0.021177 20.0424 0.131 0.00017234 0.75917 0.0097292 0.010748 0.0017771 0.98161 0.98525 3.892e-006 1.5569e-005 0.16736 0.61113 0.72031 0.0015918 0.7128 0.3509 0.0021369 0.4162 1.5426 1.5383 16.0203 144.884 0.00045564 -84.1606 0.16694
9.271 0.98816 5.4582e-005 3.8183 0.011905 0.00012033 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6482 0.61517 0.18764 0.021178 20.0457 0.13101 0.00017234 0.75916 0.0097295 0.010748 0.0017737 0.98166 0.98545 3.884e-006 1.5537e-005 0.16737 0.61229 0.7214 0.0015902 0.71438 0.35112 0.0021348 0.4162 1.5449 1.5407 16.0204 144.8841 0.00045418 -84.1721 0.16794
9.272 0.98816 5.4582e-005 3.8183 0.011905 0.00012034 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6482 0.61521 0.18765 0.021179 20.0491 0.13102 0.00017235 0.75916 0.0097299 0.010749 0.0017703 0.98171 0.98563 3.8762e-006 1.5506e-005 0.16737 0.61344 0.72248 0.0015886 0.71596 0.35133 0.0021327 0.4162 1.5472 1.543 16.0205 144.8841 0.00045274 -84.1836 0.16894
9.273 0.98816 5.4582e-005 3.8183 0.011905 0.00012036 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6483 0.61526 0.18766 0.02118 20.0525 0.13102 0.00017236 0.75915 0.0097302 0.010749 0.001767 0.98176 0.98581 3.8684e-006 1.5475e-005 0.16737 0.61459 0.72356 0.0015871 0.71753 0.35155 0.0021306 0.4162 1.5494 1.5453 16.0205 144.8841 0.00045131 -84.1949 0.16994
9.274 0.98816 5.4582e-005 3.8183 0.011905 0.00012037 0.0011785 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6484 0.6153 0.18767 0.021181 20.0558 0.13103 0.00017237 0.75914 0.0097305 0.010749 0.0017637 0.9818 0.98598 3.8607e-006 1.5444e-005 0.16737 0.61573 0.72462 0.0015855 0.7191 0.35176 0.0021286 0.4162 1.5517 1.5476 16.0206 144.8841 0.00044988 -84.2062 0.17094
9.275 0.98816 5.4582e-005 3.8183 0.011905 0.00012038 0.0011786 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6485 0.61534 0.18769 0.021182 20.0592 0.13103 0.00017238 0.75914 0.0097308 0.01075 0.0017604 0.98185 0.98614 3.8531e-006 1.5413e-005 0.16738 0.61687 0.72568 0.0015839 0.72065 0.35198 0.0021266 0.41621 1.554 1.5499 16.0207 144.8841 0.00044846 -84.2174 0.17194
9.276 0.98816 5.4581e-005 3.8183 0.011905 0.0001204 0.0011786 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6486 0.61539 0.1877 0.021183 20.0626 0.13104 0.00017239 0.75913 0.0097312 0.01075 0.0017571 0.9819 0.98629 3.8455e-006 1.5383e-005 0.16738 0.61801 0.72673 0.0015824 0.7222 0.35219 0.0021246 0.41621 1.5563 1.5522 16.0208 144.8841 0.00044704 -84.2285 0.17294
9.277 0.98816 5.4581e-005 3.8183 0.011905 0.00012041 0.0011786 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6487 0.61543 0.18771 0.021184 20.0659 0.13104 0.0001724 0.75913 0.0097315 0.01075 0.0017539 0.98194 0.98644 3.838e-006 1.5353e-005 0.16738 0.61914 0.72778 0.0015809 0.72375 0.35241 0.0021226 0.41621 1.5586 1.5545 16.0208 144.8841 0.00044564 -84.2395 0.17394
9.278 0.98816 5.4581e-005 3.8183 0.011905 0.00012042 0.0011786 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6487 0.61548 0.18773 0.021185 20.0693 0.13105 0.00017241 0.75912 0.0097318 0.010751 0.0017507 0.98199 0.98658 3.8306e-006 1.5323e-005 0.16738 0.62027 0.72881 0.0015794 0.72528 0.35263 0.0021206 0.41621 1.5609 1.5567 16.0209 144.8841 0.00044424 -84.2504 0.17494
9.279 0.98816 5.4581e-005 3.8183 0.011905 0.00012043 0.0011786 0.23353 0.00065931 0.23418 0.2161 0 0.032268 0.0389 0 1.6488 0.61552 0.18774 0.021186 20.0726 0.13106 0.00017242 0.75912 0.0097321 0.010751 0.0017476 0.98203 0.98671 3.8233e-006 1.5294e-005 0.16739 0.6214 0.72984 0.0015779 0.72681 0.35284 0.0021186 0.41622 1.5631 1.559 16.021 144.8841 0.00044285 -84.2612 0.17594
9.28 0.98816 5.4581e-005 3.8183 0.011905 0.00012045 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6489 0.61556 0.18775 0.021187 20.076 0.13106 0.00017243 0.75911 0.0097324 0.010751 0.0017445 0.98208 0.98684 3.816e-006 1.5265e-005 0.16739 0.62252 0.73086 0.0015764 0.72833 0.35306 0.0021167 0.41622 1.5654 1.5613 16.021 144.8841 0.00044147 -84.2719 0.17694
9.281 0.98816 5.4581e-005 3.8183 0.011905 0.00012046 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.649 0.61561 0.18776 0.021188 20.0794 0.13107 0.00017243 0.7591 0.0097328 0.010752 0.0017414 0.98212 0.98696 3.8089e-006 1.5236e-005 0.16739 0.62364 0.73188 0.0015749 0.72985 0.35327 0.0021148 0.41622 1.5676 1.5636 16.0211 144.8842 0.00044009 -84.2825 0.17794
9.282 0.98816 5.4581e-005 3.8183 0.011905 0.00012047 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6491 0.61565 0.18778 0.021189 20.0827 0.13107 0.00017244 0.7591 0.0097331 0.010752 0.0017384 0.98217 0.98707 3.8018e-006 1.5208e-005 0.16739 0.62476 0.73288 0.0015735 0.73136 0.35349 0.0021129 0.41622 1.5699 1.5658 16.0212 144.8842 0.00043872 -84.2931 0.17894
9.283 0.98816 5.4581e-005 3.8183 0.011905 0.00012049 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6491 0.6157 0.18779 0.02119 20.0861 0.13108 0.00017245 0.75909 0.0097334 0.010752 0.0017354 0.98221 0.98718 3.7948e-006 1.518e-005 0.1674 0.62587 0.73388 0.0015721 0.73286 0.3537 0.002111 0.41623 1.5722 1.5681 16.0212 144.8842 0.00043736 -84.3036 0.17994
9.284 0.98816 5.4581e-005 3.8183 0.011905 0.0001205 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6492 0.61574 0.1878 0.021191 20.0895 0.13109 0.00017246 0.75909 0.0097337 0.010753 0.0017324 0.98225 0.98729 3.7878e-006 1.5152e-005 0.1674 0.62698 0.73488 0.0015706 0.73436 0.35392 0.0021091 0.41623 1.5744 1.5704 16.0213 144.8842 0.00043601 -84.314 0.18094
9.285 0.98816 5.4581e-005 3.8183 0.011905 0.00012051 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6493 0.61578 0.18781 0.021192 20.0928 0.13109 0.00017247 0.75908 0.0097341 0.010753 0.0017294 0.98229 0.98739 3.7809e-006 1.5124e-005 0.1674 0.62808 0.73586 0.0015692 0.73584 0.35413 0.0021073 0.41623 1.5766 1.5726 16.0214 144.8842 0.00043466 -84.3243 0.18194
9.286 0.98816 5.4581e-005 3.8183 0.011905 0.00012052 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6494 0.61583 0.18783 0.021193 20.0962 0.1311 0.00017248 0.75908 0.0097344 0.010753 0.0017264 0.98234 0.98748 3.774e-006 1.5097e-005 0.1674 0.62919 0.73684 0.0015678 0.73733 0.35435 0.0021055 0.41624 1.5789 1.5749 16.0215 144.8842 0.00043332 -84.3345 0.18294
9.287 0.98816 5.4581e-005 3.8183 0.011905 0.00012054 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6495 0.61587 0.18784 0.021194 20.0996 0.1311 0.00017249 0.75907 0.0097347 0.010754 0.0017233 0.98238 0.98758 3.7671e-006 1.5069e-005 0.1674 0.63029 0.73781 0.0015663 0.7388 0.35457 0.0021036 0.41624 1.5811 1.5771 16.0215 144.8842 0.00043199 -84.3446 0.18394
9.288 0.98816 5.458e-005 3.8183 0.011905 0.00012055 0.0011786 0.23353 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6496 0.61592 0.18785 0.021195 20.1029 0.13111 0.0001725 0.75906 0.009735 0.010754 0.0017203 0.98242 0.98766 3.7603e-006 1.5042e-005 0.16741 0.63138 0.73878 0.0015649 0.74027 0.35478 0.0021018 0.41625 1.5833 1.5794 16.0216 144.8842 0.00043066 -84.3547 0.18494
9.289 0.98816 5.458e-005 3.8183 0.011905 0.00012056 0.0011786 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6496 0.61596 0.18787 0.021196 20.1063 0.13111 0.00017251 0.75906 0.0097354 0.010754 0.0017174 0.98246 0.98775 3.7537e-006 1.5015e-005 0.16741 0.63247 0.73973 0.0015635 0.74173 0.355 0.0021 0.41625 1.5856 1.5816 16.0217 144.8842 0.00042934 -84.3647 0.18594
9.29 0.98816 5.458e-005 3.8183 0.011905 0.00012057 0.0011786 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6497 0.616 0.18788 0.021197 20.1096 0.13112 0.00017251 0.75905 0.0097357 0.010755 0.0017146 0.9825 0.98783 3.7471e-006 1.4989e-005 0.16741 0.63356 0.74069 0.0015622 0.74318 0.35521 0.0020983 0.41625 1.5878 1.5838 16.0217 144.8843 0.00042803 -84.3746 0.18694
9.291 0.98816 5.458e-005 3.8183 0.011905 0.00012059 0.0011786 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6498 0.61605 0.18789 0.021198 20.113 0.13113 0.00017252 0.75905 0.009736 0.010755 0.0017119 0.98254 0.98791 3.7406e-006 1.4963e-005 0.16741 0.63465 0.74163 0.0015608 0.74463 0.35543 0.0020965 0.41626 1.59 1.5861 16.0218 144.8843 0.00042672 -84.3844 0.18794
9.292 0.98816 5.458e-005 3.8183 0.011905 0.0001206 0.0011786 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6499 0.61609 0.1879 0.021199 20.1164 0.13113 0.00017253 0.75904 0.0097363 0.010755 0.0017092 0.98258 0.98798 3.7343e-006 1.4938e-005 0.16742 0.63573 0.74257 0.0015595 0.74607 0.35564 0.0020948 0.41626 1.5922 1.5883 16.0218 144.8843 0.00042542 -84.3941 0.18894
9.293 0.98816 5.458e-005 3.8183 0.011905 0.00012061 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.65 0.61614 0.18792 0.0212 20.1197 0.13114 0.00017254 0.75904 0.0097367 0.010756 0.0017066 0.98262 0.98805 3.728e-006 1.4913e-005 0.16742 0.63681 0.7435 0.0015583 0.7475 0.35586 0.0020931 0.41627 1.5944 1.5905 16.0219 144.8843 0.00042413 -84.4038 0.18994
9.294 0.98816 5.458e-005 3.8183 0.011905 0.00012063 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.65 0.61618 0.18793 0.021201 20.1231 0.13114 0.00017255 0.75903 0.009737 0.010756 0.0017039 0.98265 0.98812 3.7217e-006 1.4887e-005 0.16742 0.63789 0.74443 0.001557 0.74893 0.35607 0.0020913 0.41627 1.5966 1.5927 16.022 144.8843 0.00042284 -84.4134 0.19094
9.295 0.98816 5.458e-005 3.8183 0.011905 0.00012064 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6501 0.61622 0.18794 0.021202 20.1265 0.13115 0.00017256 0.75902 0.0097373 0.010756 0.0017013 0.98269 0.98818 3.7155e-006 1.4862e-005 0.16742 0.63896 0.74535 0.0015557 0.75035 0.35629 0.0020897 0.41627 1.5988 1.5949 16.022 144.8843 0.00042157 -84.4229 0.19194
9.296 0.98816 5.458e-005 3.8183 0.011905 0.00012065 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6502 0.61627 0.18795 0.021203 20.1299 0.13115 0.00017257 0.75902 0.0097376 0.010757 0.0016986 0.98273 0.98825 3.7093e-006 1.4838e-005 0.16743 0.64003 0.74626 0.0015544 0.75176 0.35651 0.002088 0.41628 1.601 1.5971 16.0221 144.8843 0.00042029 -84.4323 0.19294
9.297 0.98816 5.458e-005 3.8183 0.011905 0.00012066 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6503 0.61631 0.18797 0.021204 20.1332 0.13116 0.00017258 0.75901 0.0097379 0.010757 0.001696 0.98277 0.98831 3.7031e-006 1.4813e-005 0.16743 0.64109 0.74717 0.0015532 0.75317 0.35672 0.0020863 0.41628 1.6032 1.5993 16.0222 144.8843 0.00041903 -84.4417 0.19394
9.298 0.98816 5.458e-005 3.8183 0.011905 0.00012068 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6504 0.61636 0.18798 0.021205 20.1366 0.13117 0.00017259 0.75901 0.0097383 0.010757 0.0016935 0.9828 0.98837 3.6971e-006 1.4789e-005 0.16743 0.64216 0.74807 0.0015519 0.75457 0.35694 0.0020847 0.41629 1.6054 1.6015 16.0222 144.8843 0.00041777 -84.451 0.19494
9.299 0.98816 5.458e-005 3.8183 0.011905 0.00012069 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6505 0.6164 0.18799 0.021206 20.14 0.13117 0.00017259 0.759 0.0097386 0.010758 0.0016909 0.98284 0.98842 3.6911e-006 1.4765e-005 0.16743 0.64322 0.74896 0.0015507 0.75596 0.35715 0.002083 0.41629 1.6076 1.6037 16.0223 144.8844 0.00041652 -84.4602 0.19594
9.3 0.98816 5.4579e-005 3.8183 0.011905 0.0001207 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6505 0.61644 0.18801 0.021207 20.1433 0.13118 0.0001726 0.75899 0.0097389 0.010758 0.0016883 0.98288 0.98848 3.6851e-006 1.4741e-005 0.16744 0.64427 0.74985 0.0015494 0.75735 0.35737 0.0020814 0.4163 1.6097 1.6059 16.0224 144.8844 0.00041527 -84.4693 0.19694
9.301 0.98816 5.4579e-005 3.8183 0.011905 0.00012072 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6506 0.61649 0.18802 0.021208 20.1467 0.13118 0.00017261 0.75899 0.0097392 0.010758 0.0016857 0.98291 0.98853 3.6791e-006 1.4717e-005 0.16744 0.64533 0.75074 0.0015482 0.75873 0.35758 0.0020798 0.4163 1.6119 1.6081 16.0224 144.8844 0.00041403 -84.4784 0.19794
9.302 0.98816 5.4579e-005 3.8183 0.011905 0.00012073 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6507 0.61653 0.18803 0.021209 20.1501 0.13119 0.00017262 0.75898 0.0097396 0.010759 0.0016831 0.98295 0.98858 3.6733e-006 1.4694e-005 0.16744 0.64638 0.75161 0.001547 0.7601 0.3578 0.0020782 0.41631 1.6141 1.6103 16.0225 144.8844 0.0004128 -84.4874 0.19894
9.303 0.98816 5.4579e-005 3.8183 0.011905 0.00012074 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6508 0.61658 0.18804 0.02121 20.1534 0.1312 0.00017263 0.75898 0.0097399 0.010759 0.0016806 0.98298 0.98863 3.6674e-006 1.467e-005 0.16744 0.64742 0.75248 0.0015457 0.76147 0.35801 0.0020766 0.41631 1.6163 1.6125 16.0225 144.8844 0.00041157 -84.4963 0.19994
9.304 0.98816 5.4579e-005 3.8183 0.011905 0.00012075 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6509 0.61662 0.18806 0.02121 20.1568 0.1312 0.00017264 0.75897 0.0097402 0.01076 0.0016781 0.98302 0.98868 3.6617e-006 1.4647e-005 0.16745 0.64847 0.75335 0.0015445 0.76283 0.35823 0.0020751 0.41632 1.6184 1.6146 16.0226 144.8844 0.00041035 -84.5052 0.20094
9.305 0.98816 5.4579e-005 3.8183 0.011905 0.00012077 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.651 0.61666 0.18807 0.021211 20.1602 0.13121 0.00017265 0.75897 0.0097405 0.01076 0.0016756 0.98305 0.98872 3.656e-006 1.4625e-005 0.16745 0.64951 0.75421 0.0015433 0.76418 0.35844 0.0020735 0.41633 1.6206 1.6168 16.0227 144.8844 0.00040913 -84.514 0.20194
9.306 0.98816 5.4579e-005 3.8183 0.011904 0.00012078 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.651 0.61671 0.18808 0.021212 20.1635 0.13121 0.00017266 0.75896 0.0097408 0.01076 0.0016732 0.98309 0.98876 3.6503e-006 1.4602e-005 0.16745 0.65054 0.75506 0.0015421 0.76553 0.35866 0.002072 0.41633 1.6227 1.619 16.0227 144.8844 0.00040793 -84.5227 0.20294
9.307 0.98816 5.4579e-005 3.8183 0.011904 0.00012079 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6511 0.61675 0.18809 0.021213 20.1669 0.13122 0.00017267 0.75895 0.0097412 0.010761 0.0016708 0.98312 0.98881 3.6448e-006 1.458e-005 0.16745 0.65158 0.75591 0.001541 0.76686 0.35888 0.0020704 0.41634 1.6249 1.6211 16.0228 144.8844 0.00040672 -84.5313 0.20394
9.308 0.98816 5.4579e-005 3.8183 0.011904 0.0001208 0.0011787 0.23352 0.00065931 0.23418 0.21609 0 0.032268 0.0389 0 1.6512 0.6168 0.18811 0.021214 20.1703 0.13122 0.00017268 0.75895 0.0097415 0.010761 0.0016684 0.98315 0.98885 3.6392e-006 1.4558e-005 0.16746 0.65261 0.75676 0.0015398 0.7682 0.35909 0.0020689 0.41634 1.627 1.6233 16.0228 144.8845 0.00040553 -84.5399 0.20494
9.309 0.98816 5.4579e-005 3.8183 0.011904 0.00012082 0.0011787 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6513 0.61684 0.18812 0.021215 20.1737 0.13123 0.00017268 0.75894 0.0097418 0.010761 0.001666 0.98319 0.98889 3.6338e-006 1.4536e-005 0.16746 0.65363 0.75759 0.0015387 0.76953 0.35931 0.0020674 0.41635 1.6291 1.6254 16.0229 144.8845 0.00040434 -84.5484 0.20594
9.31 0.98816 5.4579e-005 3.8183 0.011904 0.00012083 0.0011787 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6514 0.61688 0.18813 0.021216 20.177 0.13124 0.00017269 0.75894 0.0097421 0.010762 0.0016637 0.98322 0.98893 3.6284e-006 1.4514e-005 0.16746 0.65466 0.75843 0.0015375 0.77085 0.35952 0.002066 0.41635 1.6313 1.6276 16.0229 144.8845 0.00040316 -84.5569 0.20694
9.311 0.98816 5.4579e-005 3.8183 0.011904 0.00012084 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6514 0.61693 0.18815 0.021217 20.1804 0.13124 0.0001727 0.75893 0.0097425 0.010762 0.0016614 0.98325 0.98896 3.623e-006 1.4493e-005 0.16746 0.65568 0.75925 0.0015364 0.77216 0.35974 0.0020645 0.41636 1.6334 1.6297 16.023 144.8845 0.00040198 -84.5653 0.20794
9.312 0.98816 5.4578e-005 3.8183 0.011904 0.00012086 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6515 0.61697 0.18816 0.021218 20.1838 0.13125 0.00017271 0.75893 0.0097428 0.010762 0.0016592 0.98328 0.989 3.6177e-006 1.4471e-005 0.16747 0.6567 0.76007 0.0015353 0.77347 0.35995 0.002063 0.41637 1.6355 1.6318 16.0231 144.8845 0.00040081 -84.5736 0.20894
9.313 0.98816 5.4578e-005 3.8183 0.011904 0.00012087 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6516 0.61702 0.18817 0.021219 20.1872 0.13125 0.00017272 0.75892 0.0097431 0.010763 0.0016569 0.98331 0.98904 3.6124e-006 1.445e-005 0.16747 0.65771 0.76089 0.0015342 0.77477 0.36017 0.0020616 0.41637 1.6376 1.634 16.0231 144.8845 0.00039964 -84.5818 0.20994
9.314 0.98816 5.4578e-005 3.8183 0.011904 0.00012088 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6517 0.61706 0.18818 0.02122 20.1905 0.13126 0.00017273 0.75891 0.0097434 0.010763 0.0016547 0.98335 0.98907 3.6072e-006 1.4429e-005 0.16747 0.65872 0.7617 0.0015331 0.77606 0.36038 0.0020601 0.41638 1.6398 1.6361 16.0232 144.8845 0.00039848 -84.59 0.21094
9.315 0.98816 5.4578e-005 3.8183 0.011904 0.00012089 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6518 0.6171 0.1882 0.021221 20.1939 0.13126 0.00017274 0.75891 0.0097437 0.010763 0.0016524 0.98338 0.9891 3.602e-006 1.4409e-005 0.16747 0.65973 0.76251 0.0015321 0.77735 0.3606 0.0020587 0.41639 1.6419 1.6382 16.0232 144.8845 0.00039733 -84.5981 0.21194
9.316 0.98816 5.4578e-005 3.8183 0.011904 0.00012091 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6519 0.61715 0.18821 0.021222 20.1973 0.13127 0.00017275 0.7589 0.0097441 0.010764 0.0016502 0.98341 0.98914 3.5969e-006 1.4388e-005 0.16748 0.66074 0.76331 0.001531 0.77863 0.36081 0.0020573 0.41639 1.644 1.6403 16.0233 144.8846 0.00039618 -84.6062 0.21294
9.317 0.98816 5.4578e-005 3.8183 0.011904 0.00012092 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6519 0.61719 0.18822 0.021223 20.2007 0.13128 0.00017276 0.7589 0.0097444 0.010764 0.001648 0.98344 0.98917 3.5918e-006 1.4368e-005 0.16748 0.66174 0.7641 0.0015299 0.77991 0.36103 0.0020559 0.4164 1.6461 1.6424 16.0233 144.8846 0.00039504 -84.6142 0.21394
9.318 0.98816 5.4578e-005 3.8183 0.011904 0.00012093 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.652 0.61724 0.18823 0.021224 20.204 0.13128 0.00017276 0.75889 0.0097447 0.010764 0.0016458 0.98347 0.9892 3.5867e-006 1.4348e-005 0.16748 0.66274 0.76489 0.0015288 0.78117 0.36124 0.0020545 0.41641 1.6482 1.6446 16.0234 144.8846 0.0003939 -84.6221 0.21494
9.319 0.98816 5.4578e-005 3.8183 0.011904 0.00012094 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6521 0.61728 0.18825 0.021225 20.2074 0.13129 0.00017277 0.75888 0.009745 0.010765 0.0016437 0.9835 0.98923 3.5817e-006 1.4328e-005 0.16748 0.66374 0.76568 0.0015278 0.78244 0.36146 0.0020531 0.41641 1.6503 1.6467 16.0234 144.8846 0.00039277 -84.63 0.21594
9.32 0.98816 5.4578e-005 3.8183 0.011904 0.00012096 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6522 0.61732 0.18826 0.021226 20.2108 0.13129 0.00017278 0.75888 0.0097454 0.010765 0.0016415 0.98353 0.98926 3.5768e-006 1.4308e-005 0.16749 0.66473 0.76646 0.0015267 0.78369 0.36167 0.0020518 0.41642 1.6523 1.6488 16.0235 144.8846 0.00039164 -84.6378 0.21694
9.321 0.98816 5.4578e-005 3.8183 0.011904 0.00012097 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6523 0.61737 0.18827 0.021227 20.2142 0.1313 0.00017279 0.75887 0.0097457 0.010765 0.0016394 0.98356 0.98929 3.5719e-006 1.4288e-005 0.16749 0.66572 0.76724 0.0015257 0.78494 0.36189 0.0020504 0.41643 1.6544 1.6509 16.0235 144.8846 0.00039053 -84.6455 0.21794
9.322 0.98816 5.4578e-005 3.8183 0.011904 0.00012098 0.0011788 0.23352 0.00065931 0.23417 0.21609 0 0.032268 0.0389 0 1.6523 0.61741 0.18829 0.021228 20.2175 0.13131 0.0001728 0.75887 0.009746 0.010766 0.0016373 0.98359 0.98932 3.567e-006 1.4269e-005 0.16749 0.66671 0.76801 0.0015247 0.78618 0.3621 0.0020491 0.41643 1.6565 1.6529 16.0236 144.8846 0.00038941 -84.6532 0.21894
9.323 0.98816 5.4577e-005 3.8183 0.011904 0.000121 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6524 0.61746 0.1883 0.021229 20.2209 0.13131 0.00017281 0.75886 0.0097463 0.010766 0.0016352 0.98361 0.98934 3.5622e-006 1.4249e-005 0.16749 0.66769 0.76877 0.0015236 0.78742 0.36232 0.0020478 0.41644 1.6586 1.655 16.0237 144.8846 0.0003883 -84.6608 0.21994
9.324 0.98816 5.4577e-005 3.8183 0.011904 0.00012101 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6525 0.6175 0.18831 0.02123 20.2243 0.13132 0.00017282 0.75886 0.0097466 0.010766 0.0016331 0.98364 0.98937 3.5575e-006 1.423e-005 0.1675 0.66867 0.76953 0.0015226 0.78865 0.36253 0.0020464 0.41645 1.6606 1.6571 16.0237 144.8847 0.0003872 -84.6684 0.22094
9.325 0.98816 5.4577e-005 3.8183 0.011904 0.00012102 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6526 0.61754 0.18832 0.021231 20.2277 0.13132 0.00017283 0.75885 0.009747 0.010767 0.0016311 0.98367 0.9894 3.5527e-006 1.4211e-005 0.1675 0.66965 0.77029 0.0015216 0.78988 0.36275 0.0020451 0.41645 1.6627 1.6592 16.0238 144.8847 0.00038611 -84.6759 0.22194
9.326 0.98816 5.4577e-005 3.8183 0.011904 0.00012103 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6527 0.61759 0.18834 0.021232 20.231 0.13133 0.00017284 0.75884 0.0097473 0.010767 0.0016291 0.9837 0.98942 3.5481e-006 1.4193e-005 0.1675 0.67063 0.77104 0.0015206 0.79109 0.36296 0.0020438 0.41646 1.6648 1.6613 16.0238 144.8847 0.00038501 -84.6833 0.22294
9.327 0.98816 5.4577e-005 3.8183 0.011904 0.00012105 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6528 0.61763 0.18835 0.021233 20.2344 0.13133 0.00017284 0.75884 0.0097476 0.010767 0.0016271 0.98373 0.98945 3.5434e-006 1.4174e-005 0.1675 0.6716 0.77179 0.0015197 0.79231 0.36318 0.0020425 0.41647 1.6668 1.6633 16.0239 144.8847 0.00038393 -84.6907 0.22394
9.328 0.98816 5.4577e-005 3.8183 0.011904 0.00012106 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6528 0.61768 0.18836 0.021234 20.2378 0.13134 0.00017285 0.75883 0.0097479 0.010768 0.0016251 0.98375 0.98947 3.5388e-006 1.4156e-005 0.16751 0.67257 0.77253 0.0015187 0.79351 0.36339 0.0020413 0.41648 1.6689 1.6654 16.0239 144.8847 0.00038285 -84.698 0.22494
9.329 0.98816 5.4577e-005 3.8183 0.011904 0.00012107 0.0011788 0.23352 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6529 0.61772 0.18837 0.021235 20.2412 0.13135 0.00017286 0.75883 0.0097483 0.010768 0.0016232 0.98378 0.98949 3.5343e-006 1.4138e-005 0.16751 0.67353 0.77327 0.0015177 0.79471 0.36361 0.00204 0.41648 1.6709 1.6674 16.024 144.8847 0.00038177 -84.7053 0.22594
9.33 0.98816 5.4577e-005 3.8183 0.011904 0.00012109 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.653 0.61776 0.18839 0.021236 20.2446 0.13135 0.00017287 0.75882 0.0097486 0.010768 0.0016212 0.98381 0.98952 3.5298e-006 1.412e-005 0.16751 0.6745 0.774 0.0015168 0.79591 0.36382 0.0020388 0.41649 1.673 1.6695 16.024 144.8847 0.0003807 -84.7125 0.22694
9.331 0.98816 5.4577e-005 3.8183 0.011904 0.0001211 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6531 0.61781 0.1884 0.021237 20.2479 0.13136 0.00017288 0.75882 0.0097489 0.010769 0.0016193 0.98383 0.98954 3.5253e-006 1.4102e-005 0.16751 0.67546 0.77473 0.0015158 0.79709 0.36404 0.0020375 0.4165 1.675 1.6715 16.0241 144.8847 0.00037964 -84.7197 0.22794
9.332 0.98816 5.4577e-005 3.8183 0.011904 0.00012111 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6532 0.61785 0.18841 0.021238 20.2513 0.13136 0.00017289 0.75881 0.0097492 0.010769 0.0016174 0.98386 0.98956 3.5209e-006 1.4084e-005 0.16752 0.67641 0.77546 0.0015149 0.79827 0.36425 0.0020363 0.41651 1.677 1.6736 16.0241 144.8848 0.00037858 -84.7268 0.22894
9.333 0.98816 5.4577e-005 3.8183 0.011904 0.00012112 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6533 0.6179 0.18843 0.021239 20.2547 0.13137 0.0001729 0.7588 0.0097495 0.010769 0.0016155 0.98389 0.98959 3.5165e-006 1.4066e-005 0.16752 0.67737 0.77618 0.001514 0.79945 0.36447 0.0020351 0.41652 1.6791 1.6756 16.0242 144.8848 0.00037753 -84.7338 0.22994
9.334 0.98816 5.4577e-005 3.8183 0.011904 0.00012114 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6533 0.61794 0.18844 0.02124 20.2581 0.13137 0.00017291 0.7588 0.0097499 0.01077 0.0016136 0.98391 0.98961 3.5121e-006 1.4049e-005 0.16752 0.67832 0.77689 0.001513 0.80062 0.36468 0.0020339 0.41652 1.6811 1.6777 16.0242 144.8848 0.00037648 -84.7408 0.23094
9.335 0.98816 5.4576e-005 3.8183 0.011904 0.00012115 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6534 0.61798 0.18845 0.021241 20.2615 0.13138 0.00017292 0.75879 0.0097502 0.01077 0.0016118 0.98394 0.98963 3.5078e-006 1.4032e-005 0.16752 0.67927 0.7776 0.0015121 0.80178 0.3649 0.0020326 0.41653 1.6831 1.6797 16.0243 144.8848 0.00037544 -84.7478 0.23194
9.336 0.98816 5.4576e-005 3.8183 0.011904 0.00012116 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6535 0.61803 0.18846 0.021242 20.2648 0.13139 0.00017292 0.75879 0.0097505 0.01077 0.0016099 0.98396 0.98965 3.5036e-006 1.4015e-005 0.16753 0.68021 0.77831 0.0015112 0.80294 0.36511 0.0020315 0.41654 1.6851 1.6817 16.0243 144.8848 0.0003744 -84.7547 0.23294
9.337 0.98816 5.4576e-005 3.8183 0.011904 0.00012117 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6536 0.61807 0.18848 0.021243 20.2682 0.13139 0.00017293 0.75878 0.0097508 0.010771 0.0016081 0.98399 0.98967 3.4993e-006 1.3998e-005 0.16753 0.68116 0.77901 0.0015103 0.80409 0.36533 0.0020303 0.41655 1.6871 1.6837 16.0243 144.8848 0.00037337 -84.7615 0.23394
9.338 0.98816 5.4576e-005 3.8183 0.011904 0.00012119 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6537 0.61812 0.18849 0.021244 20.2716 0.1314 0.00017294 0.75878 0.0097511 0.010771 0.0016062 0.98401 0.98969 3.4951e-006 1.3981e-005 0.16753 0.6821 0.77971 0.0015094 0.80523 0.36554 0.0020291 0.41656 1.6891 1.6858 16.0244 144.8848 0.00037234 -84.7683 0.23494
9.339 0.98816 5.4576e-005 3.8183 0.011904 0.0001212 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6537 0.61816 0.1885 0.021245 20.275 0.1314 0.00017295 0.75877 0.0097515 0.010771 0.0016044 0.98404 0.98971 3.491e-006 1.3964e-005 0.16753 0.68303 0.78041 0.0015085 0.80637 0.36576 0.0020279 0.41657 1.6911 1.6878 16.0244 144.8849 0.00037132 -84.775 0.23594
9.34 0.98816 5.4576e-005 3.8183 0.011904 0.00012121 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032268 0.0389 0 1.6538 0.6182 0.18851 0.021246 20.2784 0.13141 0.00017296 0.75876 0.0097518 0.010772 0.0016026 0.98406 0.98973 3.4869e-006 1.3948e-005 0.16754 0.68397 0.7811 0.0015076 0.8075 0.36597 0.0020268 0.41657 1.6931 1.6898 16.0245 144.8849 0.0003703 -84.7817 0.23694
9.341 0.98816 5.4576e-005 3.8183 0.011904 0.00012123 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6539 0.61825 0.18853 0.021247 20.2817 0.13141 0.00017297 0.75876 0.0097521 0.010772 0.0016009 0.98409 0.98975 3.4828e-006 1.3931e-005 0.16754 0.6849 0.78179 0.0015067 0.80863 0.36619 0.0020257 0.41658 1.6951 1.6918 16.0245 144.8849 0.00036929 -84.7883 0.23794
9.342 0.98816 5.4576e-005 3.8183 0.011904 0.00012124 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.654 0.61829 0.18854 0.021248 20.2851 0.13142 0.00017298 0.75875 0.0097524 0.010772 0.0015991 0.98411 0.98977 3.4787e-006 1.3915e-005 0.16754 0.68583 0.78247 0.0015059 0.80975 0.3664 0.0020245 0.41659 1.6971 1.6938 16.0246 144.8849 0.00036828 -84.7949 0.23894
9.343 0.98816 5.4576e-005 3.8183 0.011904 0.00012125 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6541 0.61834 0.18855 0.021249 20.2885 0.13143 0.00017299 0.75875 0.0097527 0.010773 0.0015974 0.98414 0.98979 3.4747e-006 1.3899e-005 0.16754 0.68675 0.78315 0.001505 0.81087 0.36662 0.0020234 0.4166 1.6991 1.6958 16.0246 144.8849 0.00036728 -84.8014 0.23994
9.344 0.98816 5.4576e-005 3.8183 0.011904 0.00012126 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6542 0.61838 0.18857 0.02125 20.2919 0.13143 0.000173 0.75874 0.0097531 0.010773 0.0015957 0.98416 0.9898 3.4707e-006 1.3883e-005 0.16755 0.68767 0.78382 0.0015041 0.81198 0.36683 0.0020223 0.41661 1.7011 1.6978 16.0247 144.8849 0.00036628 -84.8079 0.24094
9.345 0.98816 5.4576e-005 3.8183 0.011904 0.00012128 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6542 0.61842 0.18858 0.02125 20.2953 0.13144 0.000173 0.75874 0.0097534 0.010773 0.001594 0.98418 0.98982 3.4668e-006 1.3868e-005 0.16755 0.68859 0.78449 0.0015033 0.81308 0.36705 0.0020212 0.41662 1.7031 1.6998 16.0247 144.8849 0.00036529 -84.8143 0.24194
9.346 0.98816 5.4576e-005 3.8183 0.011904 0.00012129 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6543 0.61847 0.18859 0.021251 20.2987 0.13144 0.00017301 0.75873 0.0097537 0.010774 0.0015923 0.98421 0.98984 3.4629e-006 1.3852e-005 0.16755 0.68951 0.78516 0.0015025 0.81418 0.36726 0.0020201 0.41663 1.705 1.7017 16.0247 144.885 0.0003643 -84.8207 0.24294
9.347 0.98816 5.4575e-005 3.8183 0.011904 0.0001213 0.0011789 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6544 0.61851 0.1886 0.021252 20.302 0.13145 0.00017302 0.75872 0.009754 0.010774 0.0015906 0.98423 0.98986 3.459e-006 1.3836e-005 0.16755 0.69042 0.78582 0.0015016 0.81527 0.36748 0.002019 0.41664 1.707 1.7037 16.0248 144.885 0.00036332 -84.827 0.24394
9.348 0.98816 5.4575e-005 3.8183 0.011904 0.00012131 0.001179 0.23351 0.00065931 0.23417 0.21608 0 0.032269 0.0389 0 1.6545 0.61856 0.18862 0.021253 20.3054 0.13145 0.00017303 0.75872 0.0097544 0.010774 0.0015889 0.98425 0.98987 3.4552e-006 1.3821e-005 0.16756 0.69133 0.78648 0.0015008 0.81635 0.36769 0.0020179 0.41664 1.7089 1.7057 16.0248 144.885 0.00036234 -84.8333 0.24494
9.349 0.98816 5.4575e-005 3.8183 0.011904 0.00012133 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6546 0.6186 0.18863 0.021254 20.3088 0.13146 0.00017304 0.75871 0.0097547 0.010775 0.0015873 0.98427 0.98989 3.4514e-006 1.3806e-005 0.16756 0.69224 0.78713 0.0015 0.81743 0.36791 0.0020168 0.41665 1.7109 1.7076 16.0249 144.885 0.00036137 -84.8395 0.24594
9.35 0.98816 5.4575e-005 3.8183 0.011904 0.00012134 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6546 0.61864 0.18864 0.021255 20.3122 0.13147 0.00017305 0.75871 0.009755 0.010775 0.0015857 0.9843 0.98991 3.4476e-006 1.3791e-005 0.16756 0.69315 0.78778 0.0014992 0.81851 0.36812 0.0020158 0.41666 1.7129 1.7096 16.0249 144.885 0.0003604 -84.8457 0.24694
9.351 0.98816 5.4575e-005 3.8183 0.011904 0.00012135 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6547 0.61869 0.18865 0.021256 20.3156 0.13147 0.00017306 0.7587 0.0097553 0.010775 0.0015841 0.98432 0.98992 3.4438e-006 1.3776e-005 0.16756 0.69405 0.78843 0.0014984 0.81958 0.36833 0.0020147 0.41667 1.7148 1.7116 16.025 144.885 0.00035944 -84.8518 0.24794
9.352 0.98816 5.4575e-005 3.8183 0.011904 0.00012137 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6548 0.61873 0.18867 0.021257 20.319 0.13148 0.00017307 0.7587 0.0097556 0.010776 0.0015825 0.98434 0.98994 3.4401e-006 1.3761e-005 0.16756 0.69495 0.78908 0.0014976 0.82064 0.36855 0.0020137 0.41668 1.7167 1.7135 16.025 144.885 0.00035848 -84.8579 0.24894
9.353 0.98816 5.4575e-005 3.8183 0.011904 0.00012138 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6549 0.61878 0.18868 0.021258 20.3224 0.13148 0.00017308 0.75869 0.009756 0.010776 0.0015809 0.98436 0.98996 3.4365e-006 1.3746e-005 0.16757 0.69585 0.78972 0.0014968 0.8217 0.36876 0.0020127 0.41669 1.7187 1.7155 16.025 144.8851 0.00035753 -84.8639 0.24994
9.354 0.98816 5.4575e-005 3.8183 0.011904 0.00012139 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.655 0.61882 0.18869 0.021259 20.3257 0.13149 0.00017308 0.75868 0.0097563 0.010776 0.0015793 0.98438 0.98997 3.4328e-006 1.3732e-005 0.16757 0.69674 0.79035 0.0014961 0.82275 0.36898 0.0020116 0.4167 1.7206 1.7174 16.0251 144.8851 0.00035658 -84.8699 0.25094
9.355 0.98816 5.4575e-005 3.8183 0.011904 0.0001214 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6551 0.61886 0.18871 0.02126 20.3291 0.1315 0.00017309 0.75868 0.0097566 0.010777 0.0015778 0.9844 0.98999 3.4292e-006 1.3717e-005 0.16757 0.69763 0.79098 0.0014953 0.82379 0.36919 0.0020106 0.41671 1.7225 1.7193 16.0251 144.8851 0.00035563 -84.8759 0.25194
9.356 0.98816 5.4575e-005 3.8183 0.011904 0.00012142 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6551 0.61891 0.18872 0.021261 20.3325 0.1315 0.0001731 0.75867 0.0097569 0.010777 0.0015762 0.98443 0.99 3.4256e-006 1.3703e-005 0.16757 0.69852 0.79161 0.0014945 0.82483 0.36941 0.0020096 0.41672 1.7245 1.7213 16.0252 144.8851 0.0003547 -84.8818 0.25294
9.357 0.98816 5.4575e-005 3.8183 0.011904 0.00012143 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6552 0.61895 0.18873 0.021262 20.3359 0.13151 0.00017311 0.75867 0.0097572 0.010777 0.0015747 0.98445 0.99002 3.4221e-006 1.3689e-005 0.16758 0.69941 0.79224 0.0014937 0.82587 0.36962 0.0020086 0.41673 1.7264 1.7232 16.0252 144.8851 0.00035376 -84.8876 0.25394
9.358 0.98816 5.4575e-005 3.8183 0.011904 0.00012144 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6553 0.619 0.18874 0.021263 20.3393 0.13151 0.00017312 0.75866 0.0097576 0.010778 0.0015731 0.98447 0.99003 3.4186e-006 1.3675e-005 0.16758 0.70029 0.79286 0.001493 0.8269 0.36983 0.0020076 0.41674 1.7283 1.7251 16.0252 144.8851 0.00035283 -84.8934 0.25494
9.359 0.98816 5.4574e-005 3.8183 0.011904 0.00012146 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6554 0.61904 0.18876 0.021264 20.3427 0.13152 0.00017313 0.75865 0.0097579 0.010778 0.0015716 0.98449 0.99005 3.4151e-006 1.3661e-005 0.16758 0.70117 0.79348 0.0014922 0.82792 0.37005 0.0020066 0.41675 1.7302 1.7271 16.0253 144.8851 0.0003519 -84.8992 0.25594
9.36 0.98816 5.4574e-005 3.8183 0.011904 0.00012147 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6555 0.61908 0.18877 0.021265 20.3461 0.13152 0.00017314 0.75865 0.0097582 0.010778 0.0015701 0.98451 0.99006 3.4116e-006 1.3647e-005 0.16758 0.70205 0.79409 0.0014915 0.82894 0.37026 0.0020057 0.41676 1.7321 1.729 16.0253 144.8852 0.00035098 -84.9049 0.25694
9.361 0.98816 5.4574e-005 3.8183 0.011903 0.00012148 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6555 0.61913 0.18878 0.021266 20.3495 0.13153 0.00017315 0.75864 0.0097585 0.010779 0.0015686 0.98453 0.99008 3.4082e-006 1.3633e-005 0.16759 0.70293 0.79471 0.0014907 0.82995 0.37048 0.0020047 0.41677 1.734 1.7309 16.0254 144.8852 0.00035007 -84.9106 0.25794
9.362 0.98816 5.4574e-005 3.8183 0.011903 0.00012149 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6556 0.61917 0.18879 0.021267 20.3528 0.13154 0.00017316 0.75864 0.0097588 0.010779 0.0015672 0.98455 0.99009 3.4048e-006 1.362e-005 0.16759 0.7038 0.79531 0.00149 0.83096 0.37069 0.0020037 0.41678 1.7359 1.7328 16.0254 144.8852 0.00034915 -84.9162 0.25894
9.363 0.98816 5.4574e-005 3.8183 0.011903 0.00012151 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6557 0.61921 0.18881 0.021268 20.3562 0.13154 0.00017316 0.75863 0.0097592 0.010779 0.0015657 0.98457 0.99011 3.4015e-006 1.3606e-005 0.16759 0.70467 0.79592 0.0014892 0.83196 0.37091 0.0020028 0.41679 1.7378 1.7347 16.0254 144.8852 0.00034825 -84.9218 0.25994
9.364 0.98816 5.4574e-005 3.8183 0.011903 0.00012152 0.001179 0.23351 0.00065931 0.23416 0.21608 0 0.032269 0.0389 0 1.6558 0.61926 0.18882 0.021269 20.3596 0.13155 0.00017317 0.75863 0.0097595 0.01078 0.0015643 0.98459 0.99012 3.3981e-006 1.3593e-005 0.16759 0.70554 0.79652 0.0014885 0.83296 0.37112 0.0020018 0.4168 1.7397 1.7366 16.0255 144.8852 0.00034734 -84.9273 0.26094
9.365 0.98816 5.4574e-005 3.8183 0.011903 0.00012153 0.001179 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6559 0.6193 0.18883 0.02127 20.363 0.13155 0.00017318 0.75862 0.0097598 0.01078 0.0015628 0.98461 0.99014 3.3948e-006 1.358e-005 0.1676 0.7064 0.79712 0.0014878 0.83395 0.37133 0.0020009 0.41681 1.7416 1.7385 16.0255 144.8852 0.00034644 -84.9328 0.26194
9.366 0.98816 5.4574e-005 3.8183 0.011903 0.00012154 0.0011791 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.656 0.61935 0.18885 0.021271 20.3664 0.13156 0.00017319 0.75861 0.0097601 0.01078 0.0015614 0.98463 0.99015 3.3915e-006 1.3566e-005 0.1676 0.70726 0.79771 0.0014871 0.83493 0.37155 0.002 0.41682 1.7435 1.7404 16.0256 144.8852 0.00034555 -84.9383 0.26294
9.367 0.98816 5.4574e-005 3.8183 0.011903 0.00012156 0.0011791 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.656 0.61939 0.18886 0.021272 20.3698 0.13156 0.0001732 0.75861 0.0097604 0.010781 0.00156 0.98465 0.99016 3.3883e-006 1.3553e-005 0.1676 0.70812 0.7983 0.0014864 0.83591 0.37176 0.001999 0.41683 1.7453 1.7423 16.0256 144.8853 0.00034466 -84.9437 0.26394
9.368 0.98816 5.4574e-005 3.8183 0.011903 0.00012157 0.0011791 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6561 0.61943 0.18887 0.021273 20.3732 0.13157 0.00017321 0.7586 0.0097608 0.010781 0.0015586 0.98466 0.99018 3.3851e-006 1.3541e-005 0.1676 0.70898 0.79889 0.0014857 0.83689 0.37197 0.0019981 0.41684 1.7472 1.7441 16.0256 144.8853 0.00034377 -84.9491 0.26494
9.369 0.98816 5.4574e-005 3.8183 0.011903 0.00012158 0.0011791 0.23351 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6562 0.61948 0.18888 0.021274 20.3766 0.13158 0.00017322 0.7586 0.0097611 0.010781 0.0015572 0.98468 0.99019 3.3819e-006 1.3528e-005 0.16761 0.70983 0.79948 0.001485 0.83785 0.37219 0.0019972 0.41685 1.7491 1.746 16.0257 144.8853 0.00034289 -84.9544 0.26594
9.37 0.98816 5.4573e-005 3.8183 0.011903 0.0001216 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6563 0.61952 0.1889 0.021275 20.38 0.13158 0.00017323 0.75859 0.0097614 0.010782 0.0015559 0.9847 0.9902 3.3787e-006 1.3515e-005 0.16761 0.71069 0.80006 0.0014843 0.83882 0.3724 0.0019963 0.41686 1.7509 1.7479 16.0257 144.8853 0.00034202 -84.9597 0.26694
9.371 0.98816 5.4573e-005 3.8183 0.011903 0.00012161 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6564 0.61957 0.18891 0.021276 20.3834 0.13159 0.00017324 0.75859 0.0097617 0.010782 0.0015545 0.98472 0.99022 3.3756e-006 1.3503e-005 0.16761 0.71153 0.80064 0.0014836 0.83978 0.37262 0.0019954 0.41687 1.7528 1.7498 16.0257 144.8853 0.00034114 -84.965 0.26794
9.372 0.98816 5.4573e-005 3.8183 0.011903 0.00012162 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6564 0.61961 0.18892 0.021277 20.3868 0.13159 0.00017324 0.75858 0.009762 0.010783 0.0015532 0.98474 0.99023 3.3724e-006 1.349e-005 0.16761 0.71238 0.80121 0.001483 0.84073 0.37283 0.0019945 0.41688 1.7546 1.7516 16.0258 144.8853 0.00034027 -84.9702 0.26894
9.373 0.98816 5.4573e-005 3.8183 0.011903 0.00012163 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6565 0.61965 0.18893 0.021278 20.3901 0.1316 0.00017325 0.75857 0.0097624 0.010783 0.0015518 0.98476 0.99024 3.3694e-006 1.3478e-005 0.16762 0.71322 0.80178 0.0014823 0.84168 0.37304 0.0019937 0.41689 1.7565 1.7535 16.0258 144.8854 0.00033941 -84.9754 0.26994
9.374 0.98816 5.4573e-005 3.8183 0.011903 0.00012165 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6566 0.6197 0.18895 0.021279 20.3935 0.1316 0.00017326 0.75857 0.0097627 0.010783 0.0015505 0.98477 0.99025 3.3663e-006 1.3465e-005 0.16762 0.71406 0.80235 0.0014816 0.84262 0.37326 0.0019928 0.4169 1.7583 1.7553 16.0258 144.8854 0.00033855 -84.9805 0.27094
9.375 0.98816 5.4573e-005 3.8183 0.011903 0.00012166 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6567 0.61974 0.18896 0.02128 20.3969 0.13161 0.00017327 0.75856 0.009763 0.010784 0.0015492 0.98479 0.99027 3.3633e-006 1.3453e-005 0.16762 0.7149 0.80292 0.001481 0.84356 0.37347 0.0019919 0.41691 1.7602 1.7572 16.0259 144.8854 0.00033769 -84.9856 0.27194
9.376 0.98816 5.4573e-005 3.8183 0.011903 0.00012167 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6568 0.61979 0.18897 0.021281 20.4003 0.13162 0.00017328 0.75856 0.0097633 0.010784 0.0015479 0.98481 0.99028 3.3603e-006 1.3441e-005 0.16762 0.71574 0.80348 0.0014803 0.84449 0.37369 0.0019911 0.41692 1.762 1.759 16.0259 144.8854 0.00033684 -84.9907 0.27294
9.377 0.98816 5.4573e-005 3.8183 0.011903 0.00012168 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6569 0.61983 0.18898 0.021282 20.4037 0.13162 0.00017329 0.75855 0.0097636 0.010784 0.0015466 0.98483 0.99029 3.3573e-006 1.3429e-005 0.16763 0.71657 0.80404 0.0014796 0.84542 0.3739 0.0019902 0.41693 1.7638 1.7609 16.0259 144.8854 0.00033599 -84.9957 0.27394
9.378 0.98816 5.4573e-005 3.8183 0.011903 0.0001217 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6569 0.61987 0.189 0.021283 20.4071 0.13163 0.0001733 0.75855 0.0097639 0.010785 0.0015453 0.98484 0.9903 3.3543e-006 1.3418e-005 0.16763 0.7174 0.8046 0.001479 0.84634 0.37411 0.0019894 0.41694 1.7656 1.7627 16.026 144.8854 0.00033515 -85.0007 0.27494
9.379 0.98816 5.4573e-005 3.8183 0.011903 0.00012171 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.657 0.61992 0.18901 0.021284 20.4105 0.13163 0.00017331 0.75854 0.0097643 0.010785 0.001544 0.98486 0.99031 3.3514e-006 1.3406e-005 0.16763 0.71823 0.80515 0.0014783 0.84726 0.37433 0.0019885 0.41695 1.7675 1.7645 16.026 144.8854 0.00033431 -85.0056 0.27594
9.38 0.98816 5.4573e-005 3.8183 0.011903 0.00012172 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6571 0.61996 0.18902 0.021285 20.4139 0.13164 0.00017332 0.75853 0.0097646 0.010785 0.0015427 0.98488 0.99033 3.3485e-006 1.3394e-005 0.16763 0.71906 0.8057 0.0014777 0.84817 0.37454 0.0019877 0.41696 1.7693 1.7664 16.026 144.8855 0.00033347 -85.0105 0.27694
9.381 0.98816 5.4573e-005 3.8183 0.011903 0.00012174 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6572 0.62001 0.18904 0.021285 20.4173 0.13164 0.00017332 0.75853 0.0097649 0.010786 0.0015415 0.9849 0.99034 3.3456e-006 1.3383e-005 0.16764 0.71988 0.80625 0.0014771 0.84907 0.37475 0.0019869 0.41698 1.7711 1.7682 16.0261 144.8855 0.00033264 -85.0154 0.27794
9.382 0.98816 5.4572e-005 3.8183 0.011903 0.00012175 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6573 0.62005 0.18905 0.021286 20.4207 0.13165 0.00017333 0.75852 0.0097652 0.010786 0.0015403 0.98491 0.99035 3.3427e-006 1.3371e-005 0.16764 0.7207 0.80679 0.0014765 0.84998 0.37497 0.0019861 0.41699 1.7729 1.77 16.0261 144.8855 0.00033182 -85.0202 0.27894
9.383 0.98816 5.4572e-005 3.8183 0.011903 0.00012176 0.0011791 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6574 0.62009 0.18906 0.021287 20.4241 0.13166 0.00017334 0.75852 0.0097655 0.010786 0.001539 0.98493 0.99036 3.3399e-006 1.336e-005 0.16764 0.72152 0.80733 0.0014758 0.85087 0.37518 0.0019853 0.417 1.7747 1.7718 16.0261 144.8855 0.00033099 -85.025 0.27994
9.384 0.98816 5.4572e-005 3.8183 0.011903 0.00012177 0.0011792 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6574 0.62014 0.18907 0.021288 20.4275 0.13166 0.00017335 0.75851 0.0097659 0.010787 0.0015378 0.98495 0.99037 3.3371e-006 1.3349e-005 0.16764 0.72233 0.80787 0.0014752 0.85176 0.37539 0.0019845 0.41701 1.7765 1.7736 16.0262 144.8855 0.00033017 -85.0297 0.28094
9.385 0.98816 5.4572e-005 3.8183 0.011903 0.00012179 0.0011792 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6575 0.62018 0.18909 0.021289 20.4309 0.13167 0.00017336 0.75851 0.0097662 0.010787 0.0015366 0.98496 0.99038 3.3343e-006 1.3337e-005 0.16765 0.72315 0.80841 0.0014746 0.85265 0.37561 0.0019837 0.41702 1.7783 1.7754 16.0262 144.8855 0.00032936 -85.0345 0.28194
9.386 0.98816 5.4572e-005 3.8183 0.011903 0.0001218 0.0011792 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6576 0.62023 0.1891 0.02129 20.4343 0.13167 0.00017337 0.7585 0.0097665 0.010787 0.0015354 0.98498 0.99039 3.3315e-006 1.3326e-005 0.16765 0.72396 0.80894 0.001474 0.85353 0.37582 0.0019829 0.41703 1.7801 1.7772 16.0262 144.8856 0.00032854 -85.0391 0.28294
9.387 0.98816 5.4572e-005 3.8183 0.011903 0.00012181 0.0011792 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6577 0.62027 0.18911 0.021291 20.4377 0.13168 0.00017338 0.75849 0.0097668 0.010788 0.0015342 0.98499 0.99041 3.3288e-006 1.3315e-005 0.16765 0.72476 0.80947 0.0014734 0.85441 0.37603 0.0019821 0.41704 1.7819 1.779 16.0263 144.8856 0.00032774 -85.0438 0.28394
9.388 0.98816 5.4572e-005 3.8183 0.011903 0.00012183 0.0011792 0.2335 0.00065931 0.23416 0.21607 0 0.032269 0.0389 0 1.6578 0.62031 0.18912 0.021292 20.4411 0.13168 0.00017339 0.75849 0.0097671 0.010788 0.001533 0.98501 0.99042 3.3261e-006 1.3305e-005 0.16765 0.72557 0.81 0.0014728 0.85528 0.37625 0.0019813 0.41705 1.7836 1.7808 16.0263 144.8856 0.00032693 -85.0484 0.28494
9.389 0.98816 5.4572e-005 3.8183 0.011903 0.00012184 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6578 0.62036 0.18914 0.021293 20.4445 0.13169 0.00017339 0.75848 0.0097675 0.010788 0.0015319 0.98503 0.99043 3.3234e-006 1.3294e-005 0.16766 0.72637 0.81053 0.0014722 0.85615 0.37646 0.0019805 0.41706 1.7854 1.7826 16.0263 144.8856 0.00032613 -85.053 0.28594
9.39 0.98816 5.4572e-005 3.8183 0.011903 0.00012185 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6579 0.6204 0.18915 0.021294 20.4479 0.1317 0.0001734 0.75848 0.0097678 0.010789 0.0015307 0.98504 0.99044 3.3207e-006 1.3283e-005 0.16766 0.72717 0.81105 0.0014717 0.85701 0.37667 0.0019798 0.41708 1.7872 1.7844 16.0263 144.8856 0.00032534 -85.0575 0.28694
9.391 0.98816 5.4572e-005 3.8183 0.011903 0.00012186 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.658 0.62045 0.18916 0.021295 20.4513 0.1317 0.00017341 0.75847 0.0097681 0.010789 0.0015296 0.98506 0.99045 3.3181e-006 1.3273e-005 0.16766 0.72797 0.81157 0.0014711 0.85787 0.37688 0.001979 0.41709 1.789 1.7861 16.0264 144.8856 0.00032454 -85.062 0.28794
9.392 0.98816 5.4572e-005 3.8183 0.011903 0.00012188 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6581 0.62049 0.18918 0.021296 20.4547 0.13171 0.00017342 0.75847 0.0097684 0.010789 0.0015284 0.98507 0.99046 3.3154e-006 1.3262e-005 0.16766 0.72876 0.81208 0.0014705 0.85872 0.3771 0.0019783 0.4171 1.7907 1.7879 16.0264 144.8857 0.00032376 -85.0665 0.28894
9.393 0.98816 5.4572e-005 3.8183 0.011903 0.00012189 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6582 0.62053 0.18919 0.021297 20.4581 0.13171 0.00017343 0.75846 0.0097687 0.01079 0.0015273 0.98509 0.99047 3.3128e-006 1.3252e-005 0.16766 0.72956 0.8126 0.0014699 0.85956 0.37731 0.0019775 0.41711 1.7925 1.7897 16.0264 144.8857 0.00032297 -85.071 0.28994
9.394 0.98816 5.4571e-005 3.8183 0.011903 0.0001219 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6583 0.62058 0.1892 0.021298 20.4615 0.13172 0.00017344 0.75845 0.009769 0.01079 0.0015262 0.9851 0.99048 3.3103e-006 1.3241e-005 0.16767 0.73035 0.81311 0.0014694 0.86041 0.37752 0.0019768 0.41712 1.7942 1.7914 16.0265 144.8857 0.00032219 -85.0754 0.29094
9.395 0.98816 5.4571e-005 3.8183 0.011903 0.00012191 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6583 0.62062 0.18921 0.021299 20.4649 0.13172 0.00017345 0.75845 0.0097694 0.01079 0.0015251 0.98512 0.99049 3.3077e-006 1.3231e-005 0.16767 0.73114 0.81362 0.0014688 0.86125 0.37774 0.001976 0.41713 1.796 1.7932 16.0265 144.8857 0.00032141 -85.0797 0.29194
9.396 0.98816 5.4571e-005 3.8183 0.011903 0.00012193 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6584 0.62067 0.18923 0.0213 20.4683 0.13173 0.00017346 0.75844 0.0097697 0.010791 0.001524 0.98513 0.9905 3.3052e-006 1.3221e-005 0.16767 0.73192 0.81412 0.0014683 0.86208 0.37795 0.0019753 0.41715 1.7977 1.795 16.0265 144.8857 0.00032064 -85.0841 0.29294
9.397 0.98816 5.4571e-005 3.8183 0.011903 0.00012194 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6585 0.62071 0.18924 0.021301 20.4717 0.13174 0.00017347 0.75844 0.00977 0.010791 0.0015229 0.98515 0.99051 3.3026e-006 1.3211e-005 0.16767 0.7327 0.81463 0.0014677 0.86291 0.37816 0.0019746 0.41716 1.7995 1.7967 16.0265 144.8857 0.00031987 -85.0884 0.29394
9.398 0.98816 5.4571e-005 3.8183 0.011903 0.00012195 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6586 0.62075 0.18925 0.021302 20.4751 0.13174 0.00017347 0.75843 0.0097703 0.010791 0.0015218 0.98516 0.99052 3.3001e-006 1.3201e-005 0.16768 0.73349 0.81513 0.0014672 0.86373 0.37837 0.0019739 0.41717 1.8012 1.7984 16.0266 144.8857 0.0003191 -85.0927 0.29494
9.399 0.98816 5.4571e-005 3.8183 0.011903 0.00012197 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6587 0.6208 0.18926 0.021303 20.4785 0.13175 0.00017348 0.75843 0.0097706 0.010792 0.0015207 0.98518 0.99053 3.2977e-006 1.3191e-005 0.16768 0.73426 0.81562 0.0014666 0.86455 0.37859 0.0019732 0.41718 1.8029 1.8002 16.0266 144.8858 0.00031834 -85.0969 0.29594
9.4 0.98816 5.4571e-005 3.8183 0.011903 0.00012198 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6587 0.62084 0.18928 0.021304 20.4819 0.13175 0.00017349 0.75842 0.009771 0.010792 0.0015196 0.98519 0.99054 3.2952e-006 1.3181e-005 0.16768 0.73504 0.81612 0.0014661 0.86536 0.3788 0.0019725 0.41719 1.8047 1.8019 16.0266 144.8858 0.00031758 -85.1011 0.29694
9.401 0.98816 5.4571e-005 3.8183 0.011903 0.00012199 0.0011792 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6588 0.62088 0.18929 0.021305 20.4853 0.13176 0.0001735 0.75841 0.0097713 0.010792 0.0015186 0.9852 0.99055 3.2928e-006 1.3171e-005 0.16768 0.73581 0.81661 0.0014655 0.86617 0.37901 0.0019718 0.4172 1.8064 1.8037 16.0267 144.8858 0.00031683 -85.1053 0.29794
9.402 0.98816 5.4571e-005 3.8183 0.011903 0.000122 0.0011793 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6589 0.62093 0.1893 0.021306 20.4887 0.13176 0.00017351 0.75841 0.0097716 0.010793 0.0015175 0.98522 0.99056 3.2904e-006 1.3162e-005 0.16769 0.73658 0.8171 0.001465 0.86698 0.37923 0.0019711 0.41722 1.8081 1.8054 16.0267 144.8858 0.00031607 -85.1094 0.29894
9.403 0.98816 5.4571e-005 3.8183 0.011903 0.00012202 0.0011793 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.659 0.62097 0.18931 0.021307 20.4921 0.13177 0.00017352 0.7584 0.0097719 0.010793 0.0015165 0.98523 0.99057 3.288e-006 1.3152e-005 0.16769 0.73735 0.81759 0.0014645 0.86778 0.37944 0.0019704 0.41723 1.8098 1.8071 16.0267 144.8858 0.00031533 -85.1135 0.29994
9.404 0.98816 5.4571e-005 3.8183 0.011903 0.00012203 0.0011793 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6591 0.62102 0.18933 0.021308 20.4955 0.13178 0.00017353 0.7584 0.0097722 0.010793 0.0015155 0.98525 0.99058 3.2856e-006 1.3143e-005 0.16769 0.73812 0.81808 0.001464 0.86857 0.37965 0.0019697 0.41724 1.8115 1.8088 16.0267 144.8858 0.00031458 -85.1176 0.30094
9.405 0.98816 5.4571e-005 3.8183 0.011903 0.00012204 0.0011793 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6592 0.62106 0.18934 0.021309 20.4989 0.13178 0.00017354 0.75839 0.0097725 0.010794 0.0015144 0.98526 0.99059 3.2832e-006 1.3133e-005 0.16769 0.73888 0.81856 0.0014634 0.86937 0.37986 0.001969 0.41725 1.8132 1.8105 16.0268 144.8859 0.00031384 -85.1217 0.30194
9.406 0.98816 5.457e-005 3.8183 0.011903 0.00012205 0.0011793 0.2335 0.00065931 0.23415 0.21607 0 0.032269 0.0389 0 1.6592 0.6211 0.18935 0.02131 20.5023 0.13179 0.00017355 0.75839 0.0097729 0.010794 0.0015134 0.98527 0.9906 3.2809e-006 1.3124e-005 0.1677 0.73965 0.81904 0.0014629 0.87015 0.38008 0.0019683 0.41726 1.8149 1.8122 16.0268 144.8859 0.0003131 -85.1257 0.30294
9.407 0.98816 5.457e-005 3.8183 0.011903 0.00012207 0.0011793 0.2335 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6593 0.62115 0.18937 0.021311 20.5057 0.13179 0.00017355 0.75838 0.0097732 0.010794 0.0015124 0.98529 0.99061 3.2786e-006 1.3114e-005 0.1677 0.7404 0.81952 0.0014624 0.87094 0.38029 0.0019677 0.41728 1.8166 1.814 16.0268 144.8859 0.00031237 -85.1297 0.30394
9.408 0.98816 5.457e-005 3.8183 0.011903 0.00012208 0.0011793 0.2335 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6594 0.62119 0.18938 0.021312 20.5091 0.1318 0.00017356 0.75837 0.0097735 0.010795 0.0015114 0.9853 0.99061 3.2763e-006 1.3105e-005 0.1677 0.74116 0.81999 0.0014619 0.87171 0.3805 0.001967 0.41729 1.8183 1.8157 16.0268 144.8859 0.00031164 -85.1337 0.30494
9.409 0.98816 5.457e-005 3.8183 0.011903 0.00012209 0.0011793 0.2335 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6595 0.62124 0.18939 0.021313 20.5125 0.1318 0.00017357 0.75837 0.0097738 0.010795 0.0015104 0.98531 0.99062 3.274e-006 1.3096e-005 0.1677 0.74192 0.82047 0.0014614 0.87249 0.38071 0.0019663 0.4173 1.82 1.8174 16.0269 144.8859 0.00031091 -85.1376 0.30594
9.41 0.98816 5.457e-005 3.8183 0.011903 0.00012211 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6596 0.62128 0.1894 0.021314 20.5159 0.13181 0.00017358 0.75836 0.0097741 0.010795 0.0015094 0.98533 0.99063 3.2717e-006 1.3087e-005 0.16771 0.74267 0.82094 0.0014609 0.87325 0.38092 0.0019657 0.41731 1.8217 1.819 16.0269 144.8859 0.00031019 -85.1415 0.30694
9.411 0.98816 5.457e-005 3.8183 0.011903 0.00012212 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6596 0.62132 0.18942 0.021315 20.5193 0.13182 0.00017359 0.75836 0.0097745 0.010796 0.0015085 0.98534 0.99064 3.2695e-006 1.3078e-005 0.16771 0.74342 0.82141 0.0014604 0.87402 0.38114 0.001965 0.41732 1.8234 1.8207 16.0269 144.886 0.00030947 -85.1454 0.30794
9.412 0.98816 5.457e-005 3.8183 0.011903 0.00012213 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6597 0.62137 0.18943 0.021316 20.5227 0.13182 0.0001736 0.75835 0.0097748 0.010796 0.0015075 0.98535 0.99065 3.2673e-006 1.3069e-005 0.16771 0.74417 0.82187 0.0014599 0.87478 0.38135 0.0019644 0.41734 1.825 1.8224 16.0269 144.886 0.00030875 -85.1492 0.30894
9.413 0.98816 5.457e-005 3.8183 0.011903 0.00012214 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6598 0.62141 0.18944 0.021316 20.5261 0.13183 0.00017361 0.75835 0.0097751 0.010796 0.0015065 0.98537 0.99066 3.2651e-006 1.306e-005 0.16771 0.74491 0.82234 0.0014594 0.87554 0.38156 0.0019638 0.41735 1.8267 1.8241 16.027 144.886 0.00030804 -85.153 0.30994
9.414 0.98816 5.457e-005 3.8183 0.011903 0.00012216 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6599 0.62146 0.18945 0.021317 20.5295 0.13183 0.00017362 0.75834 0.0097754 0.010797 0.0015056 0.98538 0.99067 3.2629e-006 1.3052e-005 0.16772 0.74565 0.8228 0.0014589 0.87629 0.38177 0.0019631 0.41736 1.8284 1.8258 16.027 144.886 0.00030733 -85.1568 0.31094
9.415 0.98816 5.457e-005 3.8183 0.011903 0.00012217 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.66 0.6215 0.18947 0.021318 20.5329 0.13184 0.00017362 0.75833 0.0097757 0.010797 0.0015047 0.98539 0.99068 3.2607e-006 1.3043e-005 0.16772 0.7464 0.82326 0.0014584 0.87703 0.38199 0.0019625 0.41737 1.83 1.8274 16.027 144.886 0.00030662 -85.1606 0.31194
9.416 0.98816 5.457e-005 3.8183 0.011902 0.00012218 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6601 0.62154 0.18948 0.021319 20.5363 0.13184 0.00017363 0.75833 0.009776 0.010797 0.0015037 0.9854 0.99068 3.2586e-006 1.3034e-005 0.16772 0.74713 0.82371 0.001458 0.87778 0.3822 0.0019619 0.41739 1.8317 1.8291 16.027 144.886 0.00030591 -85.1643 0.31294
9.417 0.98816 5.457e-005 3.8183 0.011902 0.0001222 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6601 0.62159 0.18949 0.02132 20.5397 0.13185 0.00017364 0.75832 0.0097764 0.010798 0.0015028 0.98542 0.99069 3.2564e-006 1.3026e-005 0.16772 0.74787 0.82417 0.0014575 0.87851 0.38241 0.0019613 0.4174 1.8334 1.8308 16.027 144.8861 0.00030521 -85.168 0.31394
9.418 0.98816 5.4569e-005 3.8183 0.011902 0.00012221 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6602 0.62163 0.1895 0.021321 20.5431 0.13186 0.00017365 0.75832 0.0097767 0.010798 0.0015019 0.98543 0.9907 3.2543e-006 1.3017e-005 0.16773 0.7486 0.82462 0.0014571 0.87925 0.38262 0.0019607 0.41741 1.835 1.8324 16.0271 144.8861 0.00030452 -85.1717 0.31494
9.419 0.98816 5.4569e-005 3.8183 0.011902 0.00012222 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6603 0.62168 0.18952 0.021322 20.5465 0.13186 0.00017366 0.75831 0.009777 0.010798 0.001501 0.98544 0.99071 3.2522e-006 1.3009e-005 0.16773 0.74934 0.82507 0.0014566 0.87998 0.38283 0.00196 0.41742 1.8366 1.8341 16.0271 144.8861 0.00030382 -85.1753 0.31594
9.42 0.98816 5.4569e-005 3.8183 0.011902 0.00012223 0.0011793 0.23349 0.00065931 0.23415 0.21606 0 0.032269 0.0389 0 1.6604 0.62172 0.18953 0.021323 20.55 0.13187 0.00017367 0.75831 0.0097773 0.010799 0.0015001 0.98545 0.99072 3.2501e-006 1.3001e-005 0.16773 0.75006 0.82552 0.0014561 0.8807 0.38304 0.0019594 0.41744 1.8383 1.8357 16.0271 144.8861 0.00030313 -85.1789 0.31694
9.421 0.98816 5.4569e-005 3.8183 0.011902 0.00012225 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.6605 0.62176 0.18954 0.021324 20.5534 0.13187 0.00017368 0.7583 0.0097776 0.010799 0.0014992 0.98546 0.99073 3.2481e-006 1.2992e-005 0.16773 0.75079 0.82596 0.0014557 0.88142 0.38326 0.0019588 0.41745 1.8399 1.8374 16.0271 144.8861 0.00030245 -85.1825 0.31794
9.422 0.98816 5.4569e-005 3.8183 0.011902 0.00012226 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.6605 0.62181 0.18956 0.021325 20.5568 0.13188 0.00017369 0.75829 0.0097779 0.010799 0.0014983 0.98548 0.99073 3.246e-006 1.2984e-005 0.16774 0.75152 0.82641 0.0014552 0.88214 0.38347 0.0019582 0.41746 1.8416 1.839 16.0272 144.8861 0.00030176 -85.1861 0.31894
9.423 0.98816 5.4569e-005 3.8183 0.011902 0.00012227 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.6606 0.62185 0.18957 0.021326 20.5602 0.13188 0.0001737 0.75829 0.0097783 0.0108 0.0014974 0.98549 0.99074 3.244e-006 1.2976e-005 0.16774 0.75224 0.82685 0.0014548 0.88285 0.38368 0.0019577 0.41747 1.8432 1.8406 16.0272 144.8862 0.00030108 -85.1896 0.31994
9.424 0.98816 5.4569e-005 3.8183 0.011902 0.00012228 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.6607 0.6219 0.18958 0.021327 20.5636 0.13189 0.0001737 0.75828 0.0097786 0.0108 0.0014965 0.9855 0.99075 3.242e-006 1.2968e-005 0.16774 0.75296 0.82729 0.0014543 0.88356 0.38389 0.0019571 0.41749 1.8448 1.8423 16.0272 144.8862 0.0003004 -85.1931 0.32094
9.425 0.98816 5.4569e-005 3.8183 0.011902 0.0001223 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.6608 0.62194 0.18959 0.021328 20.567 0.1319 0.00017371 0.75828 0.0097789 0.0108 0.0014956 0.98551 0.99076 3.24e-006 1.296e-005 0.16774 0.75368 0.82772 0.0014539 0.88427 0.3841 0.0019565 0.4175 1.8464 1.8439 16.0272 144.8862 0.00029973 -85.1966 0.32194
9.426 0.98816 5.4569e-005 3.8183 0.011902 0.00012231 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.6609 0.62198 0.18961 0.021329 20.5704 0.1319 0.00017372 0.75827 0.0097792 0.010801 0.0014948 0.98552 0.99076 3.238e-006 1.2952e-005 0.16774 0.75439 0.82816 0.0014534 0.88497 0.38431 0.0019559 0.41751 1.848 1.8455 16.0272 144.8862 0.00029906 -85.2001 0.32294
9.427 0.98816 5.4569e-005 3.8183 0.011902 0.00012232 0.0011794 0.23349 0.00065931 0.23415 0.21606 0 0.03227 0.0389 0 1.661 0.62203 0.18962 0.02133 20.5738 0.13191 0.00017373 0.75827 0.0097795 0.010801 0.0014939 0.98553 0.99077 3.236e-006 1.2944e-005 0.16775 0.75511 0.82859 0.001453 0.88567 0.38453 0.0019554 0.41753 1.8496 1.8472 16.0273 144.8862 0.00029839 -85.2035 0.32394
9.428 0.98816 5.4569e-005 3.8183 0.011902 0.00012234 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.661 0.62207 0.18963 0.021331 20.5772 0.13191 0.00017374 0.75826 0.0097798 0.010801 0.0014931 0.98554 0.99078 3.2341e-006 1.2936e-005 0.16775 0.75582 0.82902 0.0014525 0.88636 0.38474 0.0019548 0.41754 1.8513 1.8488 16.0273 144.8862 0.00029773 -85.2069 0.32494
9.429 0.98816 5.4568e-005 3.8183 0.011902 0.00012235 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6611 0.62211 0.18964 0.021332 20.5806 0.13192 0.00017375 0.75825 0.0097802 0.010802 0.0014922 0.98556 0.99079 3.2322e-006 1.2929e-005 0.16775 0.75653 0.82945 0.0014521 0.88705 0.38495 0.0019542 0.41755 1.8529 1.8504 16.0273 144.8863 0.00029706 -85.2103 0.32594
9.43 0.98816 5.4568e-005 3.8183 0.011902 0.00012236 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6612 0.62216 0.18966 0.021333 20.5841 0.13192 0.00017376 0.75825 0.0097805 0.010802 0.0014914 0.98557 0.9908 3.2302e-006 1.2921e-005 0.16775 0.75723 0.82987 0.0014517 0.88773 0.38516 0.0019537 0.41756 1.8545 1.852 16.0273 144.8863 0.0002964 -85.2136 0.32694
9.431 0.98816 5.4568e-005 3.8183 0.011902 0.00012237 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6613 0.6222 0.18967 0.021334 20.5875 0.13193 0.00017377 0.75824 0.0097808 0.010802 0.0014906 0.98558 0.9908 3.2283e-006 1.2913e-005 0.16776 0.75794 0.8303 0.0014513 0.88841 0.38537 0.0019531 0.41758 1.856 1.8536 16.0273 144.8863 0.00029575 -85.217 0.32794
9.432 0.98816 5.4568e-005 3.8183 0.011902 0.00012239 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6614 0.62225 0.18968 0.021335 20.5909 0.13194 0.00017377 0.75824 0.0097811 0.010803 0.0014898 0.98559 0.99081 3.2264e-006 1.2906e-005 0.16776 0.75864 0.83072 0.0014509 0.88909 0.38558 0.0019526 0.41759 1.8576 1.8552 16.0274 144.8863 0.0002951 -85.2203 0.32894
9.433 0.98816 5.4568e-005 3.8183 0.011902 0.0001224 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6614 0.62229 0.18969 0.021336 20.5943 0.13194 0.00017378 0.75823 0.0097814 0.010803 0.0014889 0.9856 0.99082 3.2246e-006 1.2898e-005 0.16776 0.75934 0.83114 0.0014505 0.88976 0.38579 0.001952 0.4176 1.8592 1.8568 16.0274 144.8863 0.00029445 -85.2235 0.32994
9.434 0.98816 5.4568e-005 3.8183 0.011902 0.00012241 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6615 0.62233 0.18971 0.021337 20.5977 0.13195 0.00017379 0.75823 0.0097817 0.010803 0.0014881 0.98561 0.99082 3.2227e-006 1.2891e-005 0.16776 0.76004 0.83156 0.0014501 0.89043 0.386 0.0019515 0.41762 1.8608 1.8584 16.0274 144.8863 0.0002938 -85.2268 0.33094
9.435 0.98816 5.4568e-005 3.8183 0.011902 0.00012242 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6616 0.62238 0.18972 0.021338 20.6011 0.13195 0.0001738 0.75822 0.0097821 0.010804 0.0014873 0.98562 0.99083 3.2209e-006 1.2884e-005 0.16777 0.76074 0.83198 0.0014497 0.89109 0.38622 0.0019509 0.41763 1.8624 1.8599 16.0274 144.8864 0.00029316 -85.23 0.33194
9.436 0.98816 5.4568e-005 3.8183 0.011902 0.00012244 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6617 0.62242 0.18973 0.021339 20.6045 0.13196 0.00017381 0.75821 0.0097824 0.010804 0.0014866 0.98563 0.99084 3.219e-006 1.2876e-005 0.16777 0.76143 0.83239 0.0014493 0.89175 0.38643 0.0019504 0.41764 1.864 1.8615 16.0274 144.8864 0.00029252 -85.2332 0.33294
9.437 0.98816 5.4568e-005 3.8183 0.011902 0.00012245 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6618 0.62247 0.18975 0.02134 20.6079 0.13196 0.00017382 0.75821 0.0097827 0.010804 0.0014858 0.98564 0.99085 3.2172e-006 1.2869e-005 0.16777 0.76212 0.8328 0.0014489 0.89241 0.38664 0.0019499 0.41766 1.8655 1.8631 16.0274 144.8864 0.00029188 -85.2364 0.33394
9.438 0.98816 5.4568e-005 3.8183 0.011902 0.00012246 0.0011794 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6619 0.62251 0.18976 0.021341 20.6113 0.13197 0.00017383 0.7582 0.009783 0.010805 0.001485 0.98565 0.99085 3.2154e-006 1.2862e-005 0.16777 0.76281 0.83321 0.0014485 0.89306 0.38685 0.0019494 0.41767 1.8671 1.8647 16.0275 144.8864 0.00029124 -85.2396 0.33494
9.439 0.98816 5.4568e-005 3.8183 0.011902 0.00012248 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6619 0.62255 0.18977 0.021342 20.6148 0.13198 0.00017384 0.7582 0.0097833 0.010805 0.0014842 0.98566 0.99086 3.2137e-006 1.2855e-005 0.16778 0.7635 0.83362 0.0014481 0.89371 0.38706 0.0019488 0.41768 1.8686 1.8662 16.0275 144.8864 0.00029061 -85.2427 0.33594
9.44 0.98816 5.4568e-005 3.8183 0.011902 0.00012249 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.662 0.6226 0.18978 0.021343 20.6182 0.13198 0.00017385 0.75819 0.0097836 0.010805 0.0014834 0.98567 0.99087 3.2119e-006 1.2848e-005 0.16778 0.76419 0.83402 0.0014477 0.89436 0.38727 0.0019483 0.4177 1.8702 1.8678 16.0275 144.8865 0.00028998 -85.2458 0.33694
9.441 0.98816 5.4567e-005 3.8183 0.011902 0.0001225 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6621 0.62264 0.1898 0.021344 20.6216 0.13199 0.00017385 0.75819 0.009784 0.010806 0.0014827 0.98568 0.99087 3.2101e-006 1.2841e-005 0.16778 0.76487 0.83443 0.0014472 0.895 0.38748 0.0019478 0.41771 1.8718 1.8694 16.0275 144.8865 0.00028936 -85.2489 0.33794
9.442 0.98816 5.4567e-005 3.8183 0.011902 0.00012251 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6622 0.62269 0.18981 0.021344 20.625 0.13199 0.00017386 0.75818 0.0097843 0.010806 0.0014819 0.98569 0.99088 3.2084e-006 1.2834e-005 0.16778 0.76555 0.83483 0.0014468 0.89563 0.38769 0.0019473 0.41772 1.8733 1.8709 16.0275 144.8865 0.00028873 -85.252 0.33894
9.443 0.98816 5.4567e-005 3.8183 0.011902 0.00012253 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6623 0.62273 0.18982 0.021345 20.6284 0.132 0.00017387 0.75818 0.0097846 0.010806 0.0014812 0.9857 0.99089 3.2067e-006 1.2827e-005 0.16779 0.76623 0.83523 0.0014464 0.89627 0.3879 0.0019468 0.41774 1.8748 1.8725 16.0275 144.8865 0.00028811 -85.255 0.33994
9.444 0.98816 5.4567e-005 3.8183 0.011902 0.00012254 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6623 0.62277 0.18983 0.021346 20.6318 0.132 0.00017388 0.75817 0.0097849 0.010807 0.0014804 0.98571 0.99089 3.205e-006 1.282e-005 0.16779 0.76691 0.83563 0.001446 0.8969 0.38811 0.0019463 0.41775 1.8764 1.874 16.0276 144.8865 0.0002875 -85.258 0.34094
9.445 0.98816 5.4567e-005 3.8183 0.011902 0.00012255 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6624 0.62282 0.18985 0.021347 20.6352 0.13201 0.00017389 0.75816 0.0097852 0.010807 0.0014797 0.98572 0.9909 3.2033e-006 1.2813e-005 0.16779 0.76758 0.83603 0.0014456 0.89752 0.38832 0.0019458 0.41776 1.8779 1.8756 16.0276 144.8865 0.00028688 -85.261 0.34194
9.446 0.98816 5.4567e-005 3.8183 0.011902 0.00012257 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6625 0.62286 0.18986 0.021348 20.6387 0.13202 0.0001739 0.75816 0.0097855 0.010807 0.0014789 0.98573 0.99091 3.2016e-006 1.2806e-005 0.16779 0.76825 0.83642 0.0014452 0.89815 0.38853 0.0019453 0.41778 1.8795 1.8771 16.0276 144.8866 0.00028627 -85.264 0.34294
9.447 0.98816 5.4567e-005 3.8183 0.011902 0.00012258 0.0011795 0.23349 0.00065931 0.23414 0.21606 0 0.03227 0.0389 0 1.6626 0.62291 0.18987 0.021349 20.6421 0.13202 0.00017391 0.75815 0.0097859 0.010808 0.0014782 0.98574 0.99091 3.1999e-006 1.28e-005 0.1678 0.76892 0.83681 0.0014449 0.89877 0.38874 0.0019448 0.41779 1.881 1.8786 16.0276 144.8866 0.00028566 -85.2669 0.34394
9.448 0.98816 5.4567e-005 3.8183 0.011902 0.00012259 0.0011795 0.23349 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6627 0.62295 0.18988 0.02135 20.6455 0.13203 0.00017392 0.75815 0.0097862 0.010808 0.0014775 0.98575 0.99092 3.1982e-006 1.2793e-005 0.1678 0.76959 0.8372 0.0014445 0.89938 0.38895 0.0019443 0.4178 1.8825 1.8802 16.0276 144.8866 0.00028506 -85.2699 0.34494
9.449 0.98816 5.4567e-005 3.8183 0.011902 0.0001226 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6628 0.62299 0.1899 0.021351 20.6489 0.13203 0.00017392 0.75814 0.0097865 0.010808 0.0014768 0.98576 0.99093 3.1966e-006 1.2787e-005 0.1678 0.77026 0.83759 0.0014442 0.89999 0.38916 0.0019439 0.41782 1.884 1.8817 16.0276 144.8866 0.00028445 -85.2728 0.34594
9.45 0.98816 5.4567e-005 3.8183 0.011902 0.00012262 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6628 0.62304 0.18991 0.021352 20.6523 0.13204 0.00017393 0.75814 0.0097868 0.010809 0.0014761 0.98577 0.99093 3.195e-006 1.278e-005 0.1678 0.77092 0.83798 0.0014438 0.9006 0.38937 0.0019434 0.41783 1.8855 1.8832 16.0277 144.8866 0.00028385 -85.2757 0.34694
9.451 0.98816 5.4567e-005 3.8183 0.011902 0.00012263 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6629 0.62308 0.18992 0.021353 20.6557 0.13204 0.00017394 0.75813 0.0097871 0.010809 0.0014754 0.98578 0.99094 3.1934e-006 1.2774e-005 0.16781 0.77159 0.83837 0.0014435 0.9012 0.38958 0.0019429 0.41784 1.887 1.8847 16.0277 144.8866 0.00028325 -85.2785 0.34794
9.452 0.98816 5.4567e-005 3.8183 0.011902 0.00012264 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.663 0.62312 0.18994 0.021354 20.6592 0.13205 0.00017395 0.75812 0.0097874 0.010809 0.0014747 0.98579 0.99094 3.1917e-006 1.2767e-005 0.16781 0.77225 0.83875 0.0014432 0.90181 0.3898 0.0019424 0.41786 1.8886 1.8863 16.0277 144.8867 0.00028266 -85.2814 0.34894
9.453 0.98816 5.4566e-005 3.8183 0.011902 0.00012265 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6631 0.62317 0.18995 0.021355 20.6626 0.13206 0.00017396 0.75812 0.0097878 0.01081 0.001474 0.9858 0.99095 3.1902e-006 1.2761e-005 0.16781 0.77291 0.83913 0.0014429 0.9024 0.39001 0.001942 0.41787 1.8901 1.8878 16.0277 144.8867 0.00028207 -85.2842 0.34994
9.454 0.98816 5.4566e-005 3.8183 0.011902 0.00012267 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6632 0.62321 0.18996 0.021356 20.666 0.13206 0.00017397 0.75811 0.0097881 0.01081 0.0014733 0.98581 0.99096 3.1886e-006 1.2754e-005 0.16781 0.77356 0.83951 0.0014425 0.903 0.39022 0.0019415 0.41788 1.8916 1.8893 16.0277 144.8867 0.00028148 -85.287 0.35094
9.455 0.98816 5.4566e-005 3.8183 0.011902 0.00012268 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6632 0.62326 0.18997 0.021357 20.6694 0.13207 0.00017398 0.75811 0.0097884 0.01081 0.0014726 0.98582 0.99096 3.187e-006 1.2748e-005 0.16781 0.77422 0.83989 0.0014422 0.90359 0.39043 0.0019411 0.4179 1.893 1.8908 16.0277 144.8867 0.00028089 -85.2898 0.35194
9.456 0.98816 5.4566e-005 3.8183 0.011902 0.00012269 0.0011795 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6633 0.6233 0.18999 0.021358 20.6728 0.13207 0.00017399 0.7581 0.0097887 0.010811 0.0014719 0.98583 0.99097 3.1854e-006 1.2742e-005 0.16782 0.77487 0.84027 0.0014418 0.90417 0.39064 0.0019406 0.41791 1.8945 1.8923 16.0277 144.8867 0.00028031 -85.2925 0.35294
9.457 0.98816 5.4566e-005 3.8183 0.011902 0.00012271 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6634 0.62334 0.19 0.021359 20.6763 0.13208 0.00017399 0.7581 0.009789 0.010811 0.0014713 0.98583 0.99097 3.1839e-006 1.2736e-005 0.16782 0.77552 0.84064 0.0014415 0.90476 0.39085 0.0019402 0.41792 1.896 1.8938 16.0278 144.8868 0.00027972 -85.2953 0.35394
9.458 0.98816 5.4566e-005 3.8183 0.011902 0.00012272 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6635 0.62339 0.19001 0.02136 20.6797 0.13208 0.000174 0.75809 0.0097893 0.010811 0.0014706 0.98584 0.99098 3.1824e-006 1.273e-005 0.16782 0.77617 0.84101 0.0014411 0.90533 0.39106 0.0019397 0.41794 1.8975 1.8953 16.0278 144.8868 0.00027915 -85.298 0.35494
9.459 0.98816 5.4566e-005 3.8183 0.011902 0.00012273 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6636 0.62343 0.19002 0.021361 20.6831 0.13209 0.00017401 0.75808 0.0097896 0.010812 0.0014699 0.98585 0.99099 3.1809e-006 1.2724e-005 0.16782 0.77681 0.84138 0.0014408 0.90591 0.39126 0.0019393 0.41795 1.899 1.8967 16.0278 144.8868 0.00027857 -85.3007 0.35594
9.46 0.98816 5.4566e-005 3.8183 0.011902 0.00012274 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6636 0.62348 0.19004 0.021362 20.6865 0.1321 0.00017402 0.75808 0.00979 0.010812 0.0014693 0.98586 0.99099 3.1794e-006 1.2717e-005 0.16783 0.77746 0.84175 0.0014404 0.90648 0.39147 0.0019388 0.41797 1.9005 1.8982 16.0278 144.8868 0.000278 -85.3034 0.35694
9.461 0.98816 5.4566e-005 3.8183 0.011902 0.00012276 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6637 0.62352 0.19005 0.021363 20.6899 0.1321 0.00017403 0.75807 0.0097903 0.010812 0.0014686 0.98587 0.991 3.1779e-006 1.2712e-005 0.16783 0.7781 0.84212 0.00144 0.90705 0.39168 0.0019384 0.41798 1.9019 1.8997 16.0278 144.8868 0.00027743 -85.306 0.35794
9.462 0.98816 5.4566e-005 3.8183 0.011902 0.00012277 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6638 0.62356 0.19006 0.021364 20.6934 0.13211 0.00017404 0.75807 0.0097906 0.010813 0.001468 0.98588 0.991 3.1764e-006 1.2706e-005 0.16783 0.77874 0.84249 0.0014396 0.90762 0.39189 0.0019379 0.41799 1.9034 1.9012 16.0278 144.8868 0.00027686 -85.3087 0.35894
9.463 0.98816 5.4566e-005 3.8183 0.011902 0.00012278 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6639 0.62361 0.19007 0.021365 20.6968 0.13211 0.00017405 0.75806 0.0097909 0.010813 0.0014673 0.98589 0.99101 3.1749e-006 1.27e-005 0.16783 0.77938 0.84285 0.0014393 0.90818 0.3921 0.0019375 0.41801 1.9049 1.9026 16.0278 144.8869 0.00027629 -85.3113 0.35994
9.464 0.98816 5.4566e-005 3.8183 0.011902 0.00012279 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.664 0.62365 0.19009 0.021366 20.7002 0.13212 0.00017406 0.75806 0.0097912 0.010813 0.0014667 0.98589 0.99101 3.1734e-006 1.2694e-005 0.16784 0.78001 0.84321 0.0014389 0.90874 0.39231 0.0019371 0.41802 1.9063 1.9041 16.0278 144.8869 0.00027573 -85.3139 0.36094
9.465 0.98816 5.4565e-005 3.8183 0.011902 0.00012281 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6641 0.6237 0.1901 0.021367 20.7036 0.13212 0.00017406 0.75805 0.0097915 0.010814 0.0014661 0.9859 0.99102 3.172e-006 1.2688e-005 0.16784 0.78065 0.84357 0.0014386 0.90929 0.39252 0.0019367 0.41803 1.9078 1.9056 16.0279 144.8869 0.00027517 -85.3164 0.36194
9.466 0.98816 5.4565e-005 3.8183 0.011902 0.00012282 0.0011796 0.23348 0.00065931 0.23414 0.21605 0 0.03227 0.0389 0 1.6641 0.62374 0.19011 0.021368 20.707 0.13213 0.00017407 0.75804 0.0097919 0.010814 0.0014654 0.98591 0.99103 3.1706e-006 1.2682e-005 0.16784 0.78128 0.84393 0.0014383 0.90985 0.39273 0.0019362 0.41805 1.9092 1.907 16.0279 144.8869 0.00027461 -85.319 0.36294
9.467 0.98816 5.4565e-005 3.8183 0.011902 0.00012283 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6642 0.62378 0.19012 0.021369 20.7105 0.13214 0.00017408 0.75804 0.0097922 0.010814 0.0014648 0.98592 0.99103 3.1691e-006 1.2677e-005 0.16784 0.78191 0.84429 0.001438 0.9104 0.39294 0.0019358 0.41806 1.9107 1.9085 16.0279 144.8869 0.00027405 -85.3215 0.36394
9.468 0.98816 5.4565e-005 3.8183 0.011902 0.00012285 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6643 0.62383 0.19014 0.02137 20.7139 0.13214 0.00017409 0.75803 0.0097925 0.010815 0.0014642 0.98593 0.99104 3.1677e-006 1.2671e-005 0.16785 0.78254 0.84465 0.0014377 0.91094 0.39315 0.0019354 0.41808 1.9121 1.9099 16.0279 144.8869 0.0002735 -85.3241 0.36494
9.469 0.98816 5.4565e-005 3.8183 0.011902 0.00012286 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6644 0.62387 0.19015 0.02137 20.7173 0.13215 0.0001741 0.75803 0.0097928 0.010815 0.0014636 0.98594 0.99104 3.1663e-006 1.2665e-005 0.16785 0.78317 0.845 0.0014374 0.91148 0.39336 0.001935 0.41809 1.9136 1.9114 16.0279 144.887 0.00027295 -85.3266 0.36594
9.47 0.98816 5.4565e-005 3.8183 0.011902 0.00012287 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6645 0.62391 0.19016 0.021371 20.7207 0.13215 0.00017411 0.75802 0.0097931 0.010815 0.001463 0.98594 0.99105 3.1649e-006 1.266e-005 0.16785 0.78379 0.84535 0.0014371 0.91202 0.39357 0.0019346 0.4181 1.915 1.9128 16.0279 144.887 0.0002724 -85.329 0.36694
9.471 0.98816 5.4565e-005 3.8183 0.011901 0.00012288 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6645 0.62396 0.19018 0.021372 20.7242 0.13216 0.00017412 0.75802 0.0097934 0.010816 0.0014624 0.98595 0.99105 3.1636e-006 1.2654e-005 0.16785 0.78441 0.84571 0.0014368 0.91256 0.39378 0.0019342 0.41812 1.9164 1.9143 16.0279 144.887 0.00027186 -85.3315 0.36794
9.472 0.98816 5.4565e-005 3.8183 0.011901 0.0001229 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6646 0.624 0.19019 0.021373 20.7276 0.13216 0.00017413 0.75801 0.0097937 0.010816 0.0014618 0.98596 0.99106 3.1622e-006 1.2649e-005 0.16786 0.78503 0.84605 0.0014365 0.91309 0.39399 0.0019338 0.41813 1.9178 1.9157 16.0279 144.887 0.00027131 -85.334 0.36894
9.473 0.98816 5.4565e-005 3.8183 0.011901 0.00012291 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6647 0.62405 0.1902 0.021374 20.731 0.13217 0.00017414 0.758 0.0097941 0.010816 0.0014612 0.98597 0.99106 3.1608e-006 1.2643e-005 0.16786 0.78565 0.8464 0.0014363 0.91362 0.3942 0.0019334 0.41815 1.9193 1.9171 16.0279 144.887 0.00027077 -85.3364 0.36994
9.474 0.98816 5.4565e-005 3.8183 0.011901 0.00012292 0.0011796 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6648 0.62409 0.19021 0.021375 20.7344 0.13218 0.00017414 0.758 0.0097944 0.010817 0.0014606 0.98597 0.99107 3.1595e-006 1.2638e-005 0.16786 0.78627 0.84675 0.001436 0.91415 0.39441 0.001933 0.41816 1.9207 1.9186 16.0279 144.8871 0.00027024 -85.3388 0.37094
9.475 0.98816 5.4565e-005 3.8183 0.011901 0.00012294 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6649 0.62413 0.19023 0.021376 20.7379 0.13218 0.00017415 0.75799 0.0097947 0.010817 0.00146 0.98598 0.99107 3.1581e-006 1.2633e-005 0.16786 0.78688 0.84709 0.0014357 0.91467 0.39461 0.0019326 0.41817 1.9221 1.92 16.028 144.8871 0.0002697 -85.3412 0.37194
9.476 0.98816 5.4564e-005 3.8183 0.011901 0.00012295 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.665 0.62418 0.19024 0.021377 20.7413 0.13219 0.00017416 0.75799 0.009795 0.010817 0.0014595 0.98599 0.99108 3.1568e-006 1.2627e-005 0.16787 0.7875 0.84744 0.0014354 0.91519 0.39482 0.0019322 0.41819 1.9235 1.9214 16.028 144.8871 0.00026917 -85.3436 0.37294
9.477 0.98816 5.4564e-005 3.8183 0.011901 0.00012296 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.665 0.62422 0.19025 0.021378 20.7447 0.13219 0.00017417 0.75798 0.0097953 0.010818 0.0014589 0.986 0.99108 3.1555e-006 1.2622e-005 0.16787 0.78811 0.84778 0.0014351 0.91571 0.39503 0.0019318 0.4182 1.9249 1.9228 16.028 144.8871 0.00026864 -85.3459 0.37394
9.478 0.98816 5.4564e-005 3.8183 0.011901 0.00012297 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6651 0.62427 0.19026 0.021379 20.7481 0.1322 0.00017418 0.75798 0.0097956 0.010818 0.0014583 0.98601 0.99109 3.1542e-006 1.2617e-005 0.16787 0.78872 0.84812 0.0014347 0.91622 0.39524 0.0019314 0.41822 1.9263 1.9242 16.028 144.8871 0.00026811 -85.3483 0.37494
9.479 0.98816 5.4564e-005 3.8183 0.011901 0.00012299 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6652 0.62431 0.19028 0.02138 20.7516 0.1322 0.00017419 0.75797 0.0097959 0.010818 0.0014577 0.98601 0.99109 3.1529e-006 1.2612e-005 0.16787 0.78933 0.84846 0.0014344 0.91673 0.39545 0.001931 0.41823 1.9277 1.9256 16.028 144.8871 0.00026758 -85.3506 0.37594
9.48 0.98816 5.4564e-005 3.8183 0.011901 0.000123 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6653 0.62435 0.19029 0.021381 20.755 0.13221 0.0001742 0.75796 0.0097963 0.010819 0.0014572 0.98602 0.9911 3.1516e-006 1.2606e-005 0.16788 0.78993 0.84879 0.0014341 0.91724 0.39566 0.0019307 0.41825 1.9291 1.927 16.028 144.8872 0.00026706 -85.3529 0.37694
9.481 0.98816 5.4564e-005 3.8183 0.011901 0.00012301 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6654 0.6244 0.1903 0.021382 20.7584 0.13221 0.00017421 0.75796 0.0097966 0.010819 0.0014566 0.98603 0.9911 3.1503e-006 1.2601e-005 0.16788 0.79053 0.84913 0.0014338 0.91774 0.39587 0.0019303 0.41826 1.9305 1.9284 16.028 144.8872 0.00026654 -85.3552 0.37794
9.482 0.98816 5.4564e-005 3.8183 0.011901 0.00012302 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6654 0.62444 0.19031 0.021383 20.7618 0.13222 0.00017421 0.75795 0.0097969 0.010819 0.0014561 0.98603 0.99111 3.1491e-006 1.2596e-005 0.16788 0.79114 0.84946 0.0014335 0.91824 0.39608 0.0019299 0.41827 1.9319 1.9298 16.028 144.8872 0.00026602 -85.3574 0.37894
9.483 0.98816 5.4564e-005 3.8183 0.011901 0.00012304 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6655 0.62449 0.19033 0.021384 20.7653 0.13223 0.00017422 0.75795 0.0097972 0.01082 0.0014555 0.98604 0.99111 3.1478e-006 1.2591e-005 0.16788 0.79174 0.84979 0.0014332 0.91874 0.39628 0.0019296 0.41829 1.9333 1.9312 16.028 144.8872 0.0002655 -85.3597 0.37994
9.484 0.98816 5.4564e-005 3.8183 0.011901 0.00012305 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6656 0.62453 0.19034 0.021385 20.7687 0.13223 0.00017423 0.75794 0.0097975 0.01082 0.001455 0.98605 0.99112 3.1466e-006 1.2586e-005 0.16788 0.79233 0.85013 0.0014329 0.91924 0.39649 0.0019292 0.4183 1.9347 1.9326 16.028 144.8872 0.00026499 -85.3619 0.38094
9.485 0.98816 5.4564e-005 3.8183 0.011901 0.00012306 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6657 0.62457 0.19035 0.021386 20.7721 0.13224 0.00017424 0.75794 0.0097978 0.01082 0.0014544 0.98606 0.99112 3.1453e-006 1.2581e-005 0.16789 0.79293 0.85045 0.0014326 0.91973 0.3967 0.0019288 0.41832 1.9361 1.934 16.028 144.8873 0.00026447 -85.3642 0.38194
9.486 0.98816 5.4564e-005 3.8183 0.011901 0.00012308 0.0011797 0.23348 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6658 0.62462 0.19036 0.021387 20.7756 0.13224 0.00017425 0.75793 0.0097981 0.010821 0.0014539 0.98606 0.99113 3.1441e-006 1.2576e-005 0.16789 0.79352 0.85078 0.0014323 0.92022 0.39691 0.0019285 0.41833 1.9374 1.9354 16.028 144.8873 0.00026396 -85.3664 0.38294
9.487 0.98816 5.4564e-005 3.8183 0.011901 0.00012309 0.0011797 0.23347 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6659 0.62466 0.19038 0.021388 20.779 0.13225 0.00017426 0.75793 0.0097985 0.010821 0.0014534 0.98607 0.99113 3.1429e-006 1.2572e-005 0.16789 0.79412 0.85111 0.0014321 0.9207 0.39712 0.0019281 0.41835 1.9388 1.9368 16.0281 144.8873 0.00026346 -85.3685 0.38394
9.488 0.98816 5.4563e-005 3.8183 0.011901 0.0001231 0.0011797 0.23347 0.00065931 0.23413 0.21605 0 0.03227 0.0389 0 1.6659 0.6247 0.19039 0.021389 20.7824 0.13225 0.00017427 0.75792 0.0097988 0.010821 0.0014529 0.98608 0.99114 3.1417e-006 1.2567e-005 0.16789 0.79471 0.85143 0.0014319 0.92119 0.39733 0.0019277 0.41836 1.9402 1.9381 16.0281 144.8873 0.00026295 -85.3707 0.38494
9.489 0.98816 5.4563e-005 3.8183 0.011901 0.00012311 0.0011797 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.666 0.62475 0.1904 0.02139 20.7858 0.13226 0.00017428 0.75791 0.0097991 0.010822 0.0014523 0.98608 0.99114 3.1405e-006 1.2562e-005 0.1679 0.7953 0.85176 0.0014316 0.92167 0.39753 0.0019274 0.41837 1.9415 1.9395 16.0281 144.8873 0.00026245 -85.3729 0.38594
9.49 0.98816 5.4563e-005 3.8183 0.011901 0.00012313 0.0011797 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6661 0.62479 0.19042 0.021391 20.7893 0.13227 0.00017428 0.75791 0.0097994 0.010822 0.0014518 0.98609 0.99114 3.1393e-006 1.2557e-005 0.1679 0.79588 0.85208 0.0014314 0.92214 0.39774 0.001927 0.41839 1.9429 1.9409 16.0281 144.8874 0.00026195 -85.375 0.38694
9.491 0.98816 5.4563e-005 3.8183 0.011901 0.00012314 0.0011797 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6662 0.62484 0.19043 0.021392 20.7927 0.13227 0.00017429 0.7579 0.0097997 0.010822 0.0014513 0.9861 0.99115 3.1381e-006 1.2552e-005 0.1679 0.79647 0.8524 0.0014312 0.92262 0.39795 0.0019267 0.4184 1.9442 1.9422 16.0281 144.8874 0.00026145 -85.3771 0.38794
9.492 0.98816 5.4563e-005 3.8183 0.011901 0.00012315 0.0011797 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6663 0.62488 0.19044 0.021393 20.7961 0.13228 0.0001743 0.7579 0.0098 0.010822 0.0014508 0.9861 0.99115 3.1369e-006 1.2548e-005 0.1679 0.79705 0.85272 0.001431 0.92309 0.39816 0.0019263 0.41842 1.9456 1.9436 16.0281 144.8874 0.00026095 -85.3792 0.38894
9.493 0.98816 5.4563e-005 3.8183 0.011901 0.00012316 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6663 0.62492 0.19045 0.021394 20.7996 0.13228 0.00017431 0.75789 0.0098003 0.010823 0.0014503 0.98611 0.99116 3.1358e-006 1.2543e-005 0.16791 0.79763 0.85304 0.0014307 0.92356 0.39837 0.001926 0.41843 1.9469 1.9449 16.0281 144.8874 0.00026046 -85.3813 0.38994
9.494 0.98816 5.4563e-005 3.8183 0.011901 0.00012318 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6664 0.62497 0.19047 0.021394 20.803 0.13229 0.00017432 0.75789 0.0098007 0.010823 0.0014498 0.98612 0.99116 3.1346e-006 1.2539e-005 0.16791 0.79821 0.85335 0.0014305 0.92402 0.39857 0.0019257 0.41845 1.9483 1.9463 16.0281 144.8874 0.00025997 -85.3834 0.39094
9.495 0.98816 5.4563e-005 3.8183 0.011901 0.00012319 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6665 0.62501 0.19048 0.021395 20.8064 0.13229 0.00017433 0.75788 0.009801 0.010823 0.0014493 0.98612 0.99117 3.1335e-006 1.2534e-005 0.16791 0.79879 0.85367 0.0014302 0.92449 0.39878 0.0019253 0.41846 1.9496 1.9476 16.0281 144.8874 0.00025948 -85.3855 0.39194
9.496 0.98816 5.4563e-005 3.8183 0.011901 0.0001232 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6666 0.62506 0.19049 0.021396 20.8099 0.1323 0.00017434 0.75787 0.0098013 0.010824 0.0014488 0.98613 0.99117 3.1324e-006 1.2529e-005 0.16791 0.79937 0.85398 0.0014299 0.92495 0.39899 0.001925 0.41848 1.951 1.949 16.0281 144.8875 0.00025899 -85.3875 0.39294
9.497 0.98816 5.4563e-005 3.8183 0.011901 0.00012322 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6667 0.6251 0.1905 0.021397 20.8133 0.13231 0.00017435 0.75787 0.0098016 0.010824 0.0014483 0.98614 0.99118 3.1312e-006 1.2525e-005 0.16792 0.79994 0.85429 0.0014296 0.9254 0.3992 0.0019247 0.41849 1.9523 1.9503 16.0281 144.8875 0.00025851 -85.3895 0.39394
9.498 0.98816 5.4563e-005 3.8183 0.011901 0.00012323 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.03227 0.0389 0 1.6668 0.62514 0.19052 0.021398 20.8167 0.13231 0.00017435 0.75786 0.0098019 0.010824 0.0014478 0.98614 0.99118 3.1301e-006 1.252e-005 0.16792 0.80051 0.8546 0.0014293 0.92586 0.3994 0.0019243 0.4185 1.9536 1.9517 16.0281 144.8875 0.00025802 -85.3916 0.39494
9.499 0.98816 5.4563e-005 3.8183 0.011901 0.00012324 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.6668 0.62519 0.19053 0.021399 20.8202 0.13232 0.00017436 0.75786 0.0098022 0.010825 0.0014473 0.98615 0.99118 3.129e-006 1.2516e-005 0.16792 0.80108 0.85491 0.001429 0.92631 0.39961 0.001924 0.41852 1.9549 1.953 16.0281 144.8875 0.00025754 -85.3936 0.39594
9.5 0.98816 5.4562e-005 3.8183 0.011901 0.00012325 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.6669 0.62523 0.19054 0.0214 20.8236 0.13232 0.00017437 0.75785 0.0098025 0.010825 0.0014468 0.98616 0.99119 3.1279e-006 1.2512e-005 0.16792 0.80165 0.85522 0.0014287 0.92676 0.39982 0.0019237 0.41853 1.9563 1.9543 16.0281 144.8875 0.00025706 -85.3955 0.39694
9.501 0.98816 5.4562e-005 3.8183 0.011901 0.00012327 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.667 0.62527 0.19055 0.021401 20.827 0.13233 0.00017438 0.75785 0.0098029 0.010825 0.0014464 0.98616 0.99119 3.1268e-006 1.2507e-005 0.16793 0.80222 0.85553 0.0014285 0.92721 0.40003 0.0019234 0.41855 1.9576 1.9556 16.0281 144.8876 0.00025659 -85.3975 0.39794
9.502 0.98816 5.4562e-005 3.8183 0.011901 0.00012328 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.6671 0.62532 0.19057 0.021402 20.8305 0.13233 0.00017439 0.75784 0.0098032 0.010826 0.0014459 0.98617 0.9912 3.1257e-006 1.2503e-005 0.16793 0.80278 0.85583 0.0014283 0.92765 0.40023 0.001923 0.41856 1.9589 1.957 16.0281 144.8876 0.00025611 -85.3995 0.39894
9.503 0.98816 5.4562e-005 3.8183 0.011901 0.00012329 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.6672 0.62536 0.19058 0.021403 20.8339 0.13234 0.0001744 0.75783 0.0098035 0.010826 0.0014454 0.98617 0.9912 3.1247e-006 1.2499e-005 0.16793 0.80335 0.85614 0.0014281 0.92809 0.40044 0.0019227 0.41858 1.9602 1.9583 16.0281 144.8876 0.00025564 -85.4014 0.39994
9.504 0.98816 5.4562e-005 3.8183 0.011901 0.0001233 0.0011798 0.23347 0.00065931 0.23413 0.21604 0 0.032271 0.0389 0 1.6672 0.62541 0.19059 0.021404 20.8373 0.13235 0.00017441 0.75783 0.0098038 0.010826 0.001445 0.98618 0.9912 3.1236e-006 1.2494e-005 0.16793 0.80391 0.85644 0.0014279 0.92853 0.40065 0.0019224 0.41859 1.9615 1.9596 16.0282 144.8876 0.00025517 -85.4033 0.40094
9.505 0.98816 5.4562e-005 3.8183 0.011901 0.00012332 0.0011798 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6673 0.62545 0.1906 0.021405 20.8408 0.13235 0.00017442 0.75782 0.0098041 0.010827 0.0014445 0.98619 0.99121 3.1225e-006 1.249e-005 0.16793 0.80447 0.85674 0.0014276 0.92896 0.40086 0.0019221 0.41861 1.9628 1.9609 16.0282 144.8876 0.0002547 -85.4052 0.40194
9.506 0.98816 5.4562e-005 3.8183 0.011901 0.00012333 0.0011798 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6674 0.62549 0.19062 0.021406 20.8442 0.13236 0.00017442 0.75782 0.0098044 0.010827 0.0014441 0.98619 0.99121 3.1215e-006 1.2486e-005 0.16794 0.80503 0.85704 0.0014273 0.9294 0.40106 0.0019218 0.41862 1.9641 1.9622 16.0282 144.8876 0.00025423 -85.4071 0.40294
9.507 0.98816 5.4562e-005 3.8183 0.011901 0.00012334 0.0011798 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6675 0.62554 0.19063 0.021407 20.8476 0.13236 0.00017443 0.75781 0.0098047 0.010827 0.0014436 0.9862 0.99122 3.1205e-006 1.2482e-005 0.16794 0.80558 0.85734 0.001427 0.92983 0.40127 0.0019215 0.41864 1.9654 1.9635 16.0282 144.8877 0.00025377 -85.409 0.40394
9.508 0.98816 5.4562e-005 3.8183 0.011901 0.00012336 0.0011798 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6676 0.62558 0.19064 0.021408 20.8511 0.13237 0.00017444 0.75781 0.009805 0.010828 0.0014431 0.9862 0.99122 3.1194e-006 1.2478e-005 0.16794 0.80614 0.85764 0.0014267 0.93025 0.40148 0.0019212 0.41865 1.9667 1.9648 16.0282 144.8877 0.00025331 -85.4109 0.40494
9.509 0.98816 5.4562e-005 3.8183 0.011901 0.00012337 0.0011798 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6676 0.62563 0.19065 0.021409 20.8545 0.13237 0.00017445 0.7578 0.0098054 0.010828 0.0014427 0.98621 0.99122 3.1184e-006 1.2474e-005 0.16794 0.80669 0.85793 0.0014264 0.93068 0.40168 0.0019209 0.41866 1.968 1.9661 16.0282 144.8877 0.00025285 -85.4128 0.40594
9.51 0.98816 5.4562e-005 3.8183 0.011901 0.00012338 0.0011798 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6677 0.62567 0.19067 0.02141 20.8579 0.13238 0.00017446 0.7578 0.0098057 0.010828 0.0014422 0.98622 0.99123 3.1174e-006 1.247e-005 0.16795 0.80724 0.85823 0.0014262 0.9311 0.40189 0.0019206 0.41868 1.9693 1.9674 16.0282 144.8877 0.00025239 -85.4146 0.40694
9.511 0.98816 5.4561e-005 3.8183 0.011901 0.00012339 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6678 0.62571 0.19068 0.021411 20.8614 0.13238 0.00017447 0.75779 0.009806 0.010829 0.0014418 0.98622 0.99123 3.1164e-006 1.2465e-005 0.16795 0.80779 0.85852 0.001426 0.93152 0.4021 0.0019203 0.41869 1.9706 1.9687 16.0282 144.8877 0.00025193 -85.4164 0.40794
9.512 0.98816 5.4561e-005 3.8183 0.011901 0.00012341 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6679 0.62576 0.19069 0.021412 20.8648 0.13239 0.00017448 0.75778 0.0098063 0.010829 0.0014414 0.98623 0.99124 3.1154e-006 1.2461e-005 0.16795 0.80834 0.85881 0.0014257 0.93194 0.40231 0.00192 0.41871 1.9719 1.97 16.0282 144.8878 0.00025148 -85.4182 0.40894
9.513 0.98816 5.4561e-005 3.8183 0.011901 0.00012342 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.668 0.6258 0.19071 0.021413 20.8682 0.1324 0.00017449 0.75778 0.0098066 0.010829 0.0014409 0.98623 0.99124 3.1144e-006 1.2458e-005 0.16795 0.80889 0.8591 0.0014255 0.93235 0.40251 0.0019197 0.41872 1.9731 1.9713 16.0282 144.8878 0.00025103 -85.42 0.40994
9.514 0.98816 5.4561e-005 3.8183 0.011901 0.00012343 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6681 0.62584 0.19072 0.021414 20.8717 0.1324 0.00017449 0.75777 0.0098069 0.01083 0.0014405 0.98624 0.99124 3.1134e-006 1.2454e-005 0.16796 0.80943 0.85939 0.0014253 0.93276 0.40272 0.0019194 0.41874 1.9744 1.9725 16.0282 144.8878 0.00025058 -85.4218 0.41094
9.515 0.98816 5.4561e-005 3.8183 0.011901 0.00012345 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6681 0.62589 0.19073 0.021415 20.8751 0.13241 0.0001745 0.75777 0.0098072 0.01083 0.0014401 0.98624 0.99125 3.1124e-006 1.245e-005 0.16796 0.80998 0.85968 0.0014252 0.93317 0.40293 0.0019191 0.41875 1.9757 1.9738 16.0282 144.8878 0.00025013 -85.4236 0.41194
9.516 0.98816 5.4561e-005 3.8183 0.011901 0.00012346 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6682 0.62593 0.19074 0.021416 20.8786 0.13241 0.00017451 0.75776 0.0098076 0.01083 0.0014397 0.98625 0.99125 3.1114e-006 1.2446e-005 0.16796 0.81052 0.85997 0.001425 0.93358 0.40313 0.0019188 0.41877 1.9769 1.9751 16.0282 144.8878 0.00024968 -85.4254 0.41294
9.517 0.98816 5.4561e-005 3.8183 0.011901 0.00012347 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6683 0.62598 0.19076 0.021417 20.882 0.13242 0.00017452 0.75776 0.0098079 0.010831 0.0014393 0.98626 0.99125 3.1105e-006 1.2442e-005 0.16796 0.81106 0.86025 0.0014249 0.93398 0.40334 0.0019185 0.41878 1.9782 1.9763 16.0282 144.8879 0.00024924 -85.4271 0.41394
9.518 0.98816 5.4561e-005 3.8183 0.011901 0.00012348 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6684 0.62602 0.19077 0.021417 20.8854 0.13242 0.00017453 0.75775 0.0098082 0.010831 0.0014388 0.98626 0.99126 3.1095e-006 1.2438e-005 0.16797 0.8116 0.86054 0.0014247 0.93439 0.40355 0.0019182 0.4188 1.9795 1.9776 16.0282 144.8879 0.0002488 -85.4289 0.41494
9.519 0.98816 5.4561e-005 3.8183 0.011901 0.0001235 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6685 0.62606 0.19078 0.021418 20.8889 0.13243 0.00017454 0.75774 0.0098085 0.010831 0.0014384 0.98627 0.99126 3.1086e-006 1.2434e-005 0.16797 0.81213 0.86082 0.0014245 0.93478 0.40375 0.001918 0.41881 1.9807 1.9789 16.0282 144.8879 0.00024836 -85.4306 0.41594
9.52 0.98816 5.4561e-005 3.8183 0.011901 0.00012351 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6685 0.62611 0.19079 0.021419 20.8923 0.13244 0.00017455 0.75774 0.0098088 0.010832 0.001438 0.98627 0.99126 3.1076e-006 1.2431e-005 0.16797 0.81267 0.8611 0.0014243 0.93518 0.40396 0.0019177 0.41883 1.982 1.9801 16.0282 144.8879 0.00024792 -85.4323 0.41694
9.521 0.98816 5.4561e-005 3.8183 0.011901 0.00012352 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6686 0.62615 0.19081 0.02142 20.8958 0.13244 0.00017456 0.75773 0.0098091 0.010832 0.0014376 0.98628 0.99127 3.1067e-006 1.2427e-005 0.16797 0.8132 0.86139 0.0014241 0.93558 0.40416 0.0019174 0.41884 1.9832 1.9814 16.0282 144.8879 0.00024748 -85.434 0.41794
9.522 0.98816 5.4561e-005 3.8183 0.011901 0.00012353 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6687 0.6262 0.19082 0.021421 20.8992 0.13245 0.00017456 0.75773 0.0098094 0.010832 0.0014372 0.98628 0.99127 3.1058e-006 1.2423e-005 0.16798 0.81373 0.86166 0.0014239 0.93597 0.40437 0.0019171 0.41886 1.9844 1.9826 16.0282 144.8879 0.00024705 -85.4357 0.41894
9.523 0.98816 5.456e-005 3.8183 0.011901 0.00012355 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6688 0.62624 0.19083 0.021422 20.9026 0.13245 0.00017457 0.75772 0.0098097 0.010833 0.0014368 0.98629 0.99127 3.1048e-006 1.2419e-005 0.16798 0.81426 0.86194 0.0014237 0.93636 0.40458 0.0019169 0.41887 1.9857 1.9839 16.0282 144.888 0.00024661 -85.4374 0.41994
9.524 0.98816 5.456e-005 3.8183 0.011901 0.00012356 0.0011799 0.23347 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6689 0.62628 0.19084 0.021423 20.9061 0.13246 0.00017458 0.75772 0.0098101 0.010833 0.0014364 0.98629 0.99128 3.1039e-006 1.2416e-005 0.16798 0.81479 0.86222 0.0014235 0.93674 0.40478 0.0019166 0.41889 1.9869 1.9851 16.0282 144.888 0.00024618 -85.439 0.42094
9.525 0.98816 5.456e-005 3.8183 0.0119 0.00012357 0.0011799 0.23346 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.669 0.62633 0.19086 0.021424 20.9095 0.13246 0.00017459 0.75771 0.0098104 0.010833 0.001436 0.9863 0.99128 3.103e-006 1.2412e-005 0.16798 0.81531 0.8625 0.0014232 0.93713 0.40499 0.0019163 0.4189 1.9882 1.9864 16.0282 144.888 0.00024576 -85.4407 0.42194
9.526 0.98816 5.456e-005 3.8183 0.0119 0.00012359 0.0011799 0.23346 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.669 0.62637 0.19087 0.021425 20.913 0.13247 0.0001746 0.75771 0.0098107 0.010834 0.0014356 0.9863 0.99128 3.1021e-006 1.2409e-005 0.16799 0.81584 0.86277 0.001423 0.93751 0.40519 0.001916 0.41892 1.9894 1.9876 16.0282 144.888 0.00024533 -85.4423 0.42294
9.527 0.98816 5.456e-005 3.8183 0.0119 0.0001236 0.0011799 0.23346 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6691 0.62641 0.19088 0.021426 20.9164 0.13248 0.00017461 0.7577 0.009811 0.010834 0.0014352 0.98631 0.99129 3.1012e-006 1.2405e-005 0.16799 0.81636 0.86304 0.0014227 0.93789 0.4054 0.0019158 0.41893 1.9906 1.9888 16.0282 144.888 0.0002449 -85.4439 0.42394
9.528 0.98816 5.456e-005 3.8183 0.0119 0.00012361 0.0011799 0.23346 0.00065931 0.23412 0.21604 0 0.032271 0.0389 0 1.6692 0.62646 0.19089 0.021427 20.9198 0.13248 0.00017462 0.75769 0.0098113 0.010834 0.0014348 0.98631 0.99129 3.1004e-006 1.2401e-005 0.16799 0.81688 0.86332 0.0014225 0.93827 0.40561 0.0019155 0.41895 1.9918 1.9901 16.0282 144.8881 0.00024448 -85.4455 0.42494
9.529 0.98816 5.456e-005 3.8183 0.0119 0.00012362 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6693 0.6265 0.19091 0.021428 20.9233 0.13249 0.00017463 0.75769 0.0098116 0.010835 0.0014344 0.98632 0.99129 3.0995e-006 1.2398e-005 0.16799 0.8174 0.86359 0.0014222 0.93864 0.40581 0.0019153 0.41896 1.9931 1.9913 16.0282 144.8881 0.00024406 -85.4471 0.42594
9.53 0.98816 5.456e-005 3.8183 0.0119 0.00012364 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6694 0.62655 0.19092 0.021429 20.9267 0.13249 0.00017463 0.75768 0.0098119 0.010835 0.0014341 0.98632 0.9913 3.0986e-006 1.2394e-005 0.16799 0.81792 0.86386 0.001422 0.93902 0.40602 0.001915 0.41898 1.9943 1.9925 16.0282 144.8881 0.00024364 -85.4487 0.42694
9.531 0.98816 5.456e-005 3.8183 0.0119 0.00012365 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6694 0.62659 0.19093 0.02143 20.9302 0.1325 0.00017464 0.75768 0.0098122 0.010835 0.0014337 0.98633 0.9913 3.0977e-006 1.2391e-005 0.168 0.81844 0.86413 0.0014218 0.93939 0.40622 0.0019147 0.41899 1.9955 1.9937 16.0282 144.8881 0.00024322 -85.4503 0.42794
9.532 0.98816 5.456e-005 3.8183 0.0119 0.00012366 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6695 0.62663 0.19094 0.021431 20.9336 0.1325 0.00017465 0.75767 0.0098126 0.010836 0.0014333 0.98633 0.9913 3.0969e-006 1.2388e-005 0.168 0.81895 0.8644 0.0014216 0.93976 0.40643 0.0019145 0.41901 1.9967 1.9949 16.0282 144.8881 0.00024281 -85.4519 0.42894
9.533 0.98816 5.456e-005 3.8183 0.0119 0.00012367 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6696 0.62668 0.19096 0.021432 20.9371 0.13251 0.00017466 0.75767 0.0098129 0.010836 0.0014329 0.98634 0.99131 3.096e-006 1.2384e-005 0.168 0.81947 0.86466 0.0014214 0.94012 0.40663 0.0019142 0.41902 1.9979 1.9962 16.0282 144.8882 0.00024239 -85.4534 0.42994
9.534 0.98816 5.456e-005 3.8183 0.0119 0.00012369 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6697 0.62672 0.19097 0.021433 20.9405 0.13251 0.00017467 0.75766 0.0098132 0.010836 0.0014326 0.98634 0.99131 3.0952e-006 1.2381e-005 0.168 0.81998 0.86493 0.0014213 0.94049 0.40684 0.001914 0.41904 1.9991 1.9974 16.0282 144.8882 0.00024198 -85.455 0.43094
9.535 0.98816 5.4559e-005 3.8183 0.0119 0.0001237 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6698 0.62677 0.19098 0.021434 20.9439 0.13252 0.00017468 0.75765 0.0098135 0.010837 0.0014322 0.98635 0.99131 3.0943e-006 1.2377e-005 0.16801 0.82049 0.86519 0.0014211 0.94085 0.40705 0.0019137 0.41905 2.0003 1.9986 16.0282 144.8882 0.00024157 -85.4565 0.43194
9.536 0.98816 5.4559e-005 3.8183 0.0119 0.00012371 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6698 0.62681 0.19099 0.021435 20.9474 0.13253 0.00017469 0.75765 0.0098138 0.010837 0.0014319 0.98635 0.99132 3.0935e-006 1.2374e-005 0.16801 0.821 0.86546 0.0014209 0.94121 0.40725 0.0019135 0.41907 2.0015 1.9998 16.0282 144.8882 0.00024116 -85.458 0.43294
9.537 0.98816 5.4559e-005 3.8183 0.0119 0.00012373 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6699 0.62685 0.19101 0.021436 20.9508 0.13253 0.0001747 0.75764 0.0098141 0.010837 0.0014315 0.98636 0.99132 3.0927e-006 1.2371e-005 0.16801 0.8215 0.86572 0.0014208 0.94156 0.40746 0.0019132 0.41908 2.0027 2.001 16.0282 144.8882 0.00024075 -85.4595 0.43394
9.538 0.98816 5.4559e-005 3.8183 0.0119 0.00012374 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.67 0.6269 0.19102 0.021437 20.9543 0.13254 0.0001747 0.75764 0.0098144 0.010838 0.0014311 0.98636 0.99132 3.0919e-006 1.2367e-005 0.16801 0.82201 0.86598 0.0014206 0.94192 0.40766 0.001913 0.4191 2.0039 2.0022 16.0282 144.8883 0.00024035 -85.461 0.43494
9.539 0.98816 5.4559e-005 3.8183 0.0119 0.00012375 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6701 0.62694 0.19103 0.021438 20.9577 0.13254 0.00017471 0.75763 0.0098147 0.010838 0.0014308 0.98637 0.99133 3.0911e-006 1.2364e-005 0.16802 0.82251 0.86624 0.0014204 0.94227 0.40787 0.0019128 0.41911 2.0051 2.0034 16.0282 144.8883 0.00023994 -85.4625 0.43594
9.54 0.98816 5.4559e-005 3.8183 0.0119 0.00012376 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6702 0.62698 0.19105 0.021439 20.9612 0.13255 0.00017472 0.75763 0.009815 0.010838 0.0014304 0.98637 0.99133 3.0902e-006 1.2361e-005 0.16802 0.82302 0.8665 0.0014203 0.94262 0.40807 0.0019125 0.41913 2.0063 2.0046 16.0282 144.8883 0.00023954 -85.464 0.43694
9.541 0.98816 5.4559e-005 3.8183 0.0119 0.00012378 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6703 0.62703 0.19106 0.021439 20.9646 0.13255 0.00017473 0.75762 0.0098154 0.010839 0.0014301 0.98638 0.99133 3.0894e-006 1.2358e-005 0.16802 0.82352 0.86676 0.0014201 0.94297 0.40828 0.0019123 0.41914 2.0074 2.0057 16.0282 144.8883 0.00023914 -85.4655 0.43794
9.542 0.98816 5.4559e-005 3.8183 0.0119 0.00012379 0.00118 0.23346 0.00065931 0.23412 0.21603 0 0.032271 0.0389 0 1.6703 0.62707 0.19107 0.02144 20.9681 0.13256 0.00017474 0.75761 0.0098157 0.010839 0.0014297 0.98638 0.99134 3.0887e-006 1.2355e-005 0.16802 0.82402 0.86701 0.0014199 0.94332 0.40848 0.001912 0.41916 2.0086 2.0069 16.0282 144.8883 0.00023874 -85.4669 0.43894
9.543 0.98816 5.4559e-005 3.8183 0.0119 0.0001238 0.00118 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6704 0.62712 0.19108 0.021441 20.9715 0.13257 0.00017475 0.75761 0.009816 0.010839 0.0014294 0.98638 0.99134 3.0879e-006 1.2351e-005 0.16803 0.82451 0.86727 0.0014198 0.94366 0.40869 0.0019118 0.41917 2.0098 2.0081 16.0282 144.8883 0.00023835 -85.4684 0.43994
9.544 0.98816 5.4559e-005 3.8183 0.0119 0.00012381 0.00118 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6705 0.62716 0.1911 0.021442 20.975 0.13257 0.00017476 0.7576 0.0098163 0.01084 0.0014291 0.98639 0.99134 3.0871e-006 1.2348e-005 0.16803 0.82501 0.86752 0.0014196 0.944 0.40889 0.0019116 0.41919 2.011 2.0093 16.0282 144.8884 0.00023795 -85.4698 0.44094
9.545 0.98816 5.4559e-005 3.8183 0.0119 0.00012383 0.00118 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6706 0.6272 0.19111 0.021443 20.9784 0.13258 0.00017477 0.7576 0.0098166 0.01084 0.0014287 0.98639 0.99134 3.0863e-006 1.2345e-005 0.16803 0.8255 0.86778 0.0014194 0.94434 0.4091 0.0019113 0.4192 2.0121 2.0105 16.0282 144.8884 0.00023756 -85.4712 0.44194
9.546 0.98816 5.4559e-005 3.8183 0.0119 0.00012384 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6707 0.62725 0.19112 0.021444 20.9818 0.13258 0.00017477 0.75759 0.0098169 0.01084 0.0014284 0.9864 0.99135 3.0855e-006 1.2342e-005 0.16803 0.826 0.86803 0.0014192 0.94468 0.4093 0.0019111 0.41922 2.0133 2.0116 16.0282 144.8884 0.00023717 -85.4726 0.44294
9.547 0.98816 5.4558e-005 3.8183 0.0119 0.00012385 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6707 0.62729 0.19113 0.021445 20.9853 0.13259 0.00017478 0.75759 0.0098172 0.010841 0.001428 0.9864 0.99135 3.0848e-006 1.2339e-005 0.16804 0.82649 0.86828 0.001419 0.94501 0.40951 0.0019109 0.41923 2.0145 2.0128 16.0282 144.8884 0.00023678 -85.474 0.44394
9.548 0.98816 5.4558e-005 3.8183 0.0119 0.00012387 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6708 0.62734 0.19115 0.021446 20.9887 0.13259 0.00017479 0.75758 0.0098175 0.010841 0.0014277 0.98641 0.99135 3.084e-006 1.2336e-005 0.16804 0.82698 0.86853 0.0014188 0.94535 0.40971 0.0019107 0.41925 2.0156 2.014 16.0282 144.8884 0.00023639 -85.4754 0.44494
9.549 0.98816 5.4558e-005 3.8183 0.0119 0.00012388 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6709 0.62738 0.19116 0.021447 20.9922 0.1326 0.0001748 0.75758 0.0098179 0.010841 0.0014274 0.98641 0.99136 3.0833e-006 1.2333e-005 0.16804 0.82747 0.86878 0.0014187 0.94568 0.40992 0.0019104 0.41926 2.0168 2.0151 16.0282 144.8885 0.000236 -85.4768 0.44594
9.55 0.98816 5.4558e-005 3.8183 0.0119 0.00012389 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.671 0.62742 0.19117 0.021448 20.9956 0.1326 0.00017481 0.75757 0.0098182 0.010842 0.0014271 0.98641 0.99136 3.0825e-006 1.233e-005 0.16804 0.82795 0.86903 0.0014185 0.94601 0.41012 0.0019102 0.41928 2.0179 2.0163 16.0282 144.8885 0.00023562 -85.4782 0.44694
9.551 0.98816 5.4558e-005 3.8183 0.0119 0.0001239 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6711 0.62747 0.19118 0.021449 20.9991 0.13261 0.00017482 0.75756 0.0098185 0.010842 0.0014267 0.98642 0.99136 3.0818e-006 1.2327e-005 0.16804 0.82844 0.86927 0.0014183 0.94634 0.41032 0.00191 0.41929 2.0191 2.0174 16.0282 144.8885 0.00023524 -85.4795 0.44794
9.552 0.98816 5.4558e-005 3.8183 0.0119 0.00012392 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6712 0.62751 0.1912 0.02145 21.0025 0.13262 0.00017483 0.75756 0.0098188 0.010842 0.0014264 0.98642 0.99136 3.081e-006 1.2324e-005 0.16805 0.82892 0.86952 0.0014181 0.94666 0.41053 0.0019098 0.41931 2.0202 2.0186 16.0282 144.8885 0.00023485 -85.4809 0.44894
9.553 0.98816 5.4558e-005 3.8183 0.0119 0.00012393 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6712 0.62755 0.19121 0.021451 21.006 0.13262 0.00017484 0.75755 0.0098191 0.010843 0.0014261 0.98643 0.99137 3.0803e-006 1.2321e-005 0.16805 0.82941 0.86976 0.001418 0.94698 0.41073 0.0019096 0.41932 2.0214 2.0197 16.0282 144.8885 0.00023447 -85.4822 0.44994
9.554 0.98816 5.4558e-005 3.8183 0.0119 0.00012394 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6713 0.6276 0.19122 0.021452 21.0094 0.13263 0.00017484 0.75755 0.0098194 0.010843 0.0014258 0.98643 0.99137 3.0796e-006 1.2318e-005 0.16805 0.82989 0.87001 0.0014178 0.9473 0.41094 0.0019093 0.41934 2.0225 2.0209 16.0282 144.8886 0.0002341 -85.4836 0.45094
9.555 0.98816 5.4558e-005 3.8183 0.0119 0.00012396 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6714 0.62764 0.19123 0.021453 21.0129 0.13263 0.00017485 0.75754 0.0098197 0.010843 0.0014255 0.98644 0.99137 3.0788e-006 1.2315e-005 0.16805 0.83037 0.87025 0.0014176 0.94762 0.41114 0.0019091 0.41935 2.0236 2.022 16.0282 144.8886 0.00023372 -85.4849 0.45194
9.556 0.98816 5.4558e-005 3.8183 0.0119 0.00012397 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6715 0.62769 0.19125 0.021454 21.0163 0.13264 0.00017486 0.75754 0.00982 0.010844 0.0014251 0.98644 0.99137 3.0781e-006 1.2313e-005 0.16806 0.83084 0.87049 0.0014175 0.94794 0.41135 0.0019089 0.41937 2.0248 2.0231 16.0282 144.8886 0.00023334 -85.4862 0.45294
9.557 0.98816 5.4558e-005 3.8183 0.0119 0.00012398 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6716 0.62773 0.19126 0.021455 21.0198 0.13264 0.00017487 0.75753 0.0098203 0.010844 0.0014248 0.98644 0.99138 3.0774e-006 1.231e-005 0.16806 0.83132 0.87073 0.0014173 0.94826 0.41155 0.0019087 0.41938 2.0259 2.0243 16.0281 144.8886 0.00023297 -85.4875 0.45394
9.558 0.98816 5.4557e-005 3.8183 0.0119 0.00012399 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6716 0.62777 0.19127 0.021456 21.0232 0.13265 0.00017488 0.75752 0.0098207 0.010844 0.0014245 0.98645 0.99138 3.0767e-006 1.2307e-005 0.16806 0.8318 0.87097 0.0014172 0.94857 0.41175 0.0019085 0.4194 2.027 2.0254 16.0281 144.8886 0.0002326 -85.4888 0.45494
9.559 0.98816 5.4557e-005 3.8183 0.0119 0.00012401 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6717 0.62782 0.19128 0.021457 21.0267 0.13266 0.00017489 0.75752 0.009821 0.010845 0.0014242 0.98645 0.99138 3.076e-006 1.2304e-005 0.16806 0.83227 0.87121 0.001417 0.94888 0.41196 0.0019083 0.41941 2.0281 2.0265 16.0281 144.8887 0.00023223 -85.4901 0.45594
9.56 0.98816 5.4557e-005 3.8183 0.0119 0.00012402 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6718 0.62786 0.1913 0.021458 21.0301 0.13266 0.0001749 0.75751 0.0098213 0.010845 0.0014239 0.98646 0.99139 3.0753e-006 1.2301e-005 0.16807 0.83274 0.87145 0.0014168 0.94919 0.41216 0.0019081 0.41943 2.0293 2.0277 16.0281 144.8887 0.00023186 -85.4913 0.45694
9.561 0.98816 5.4557e-005 3.8183 0.0119 0.00012403 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6719 0.62791 0.19131 0.021459 21.0336 0.13267 0.0001749 0.75751 0.0098216 0.010845 0.0014236 0.98646 0.99139 3.0746e-006 1.2299e-005 0.16807 0.83321 0.87169 0.0014167 0.9495 0.41237 0.0019079 0.41944 2.0304 2.0288 16.0281 144.8887 0.00023149 -85.4926 0.45794
9.562 0.98816 5.4557e-005 3.8183 0.0119 0.00012404 0.0011801 0.23346 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.672 0.62795 0.19132 0.02146 21.037 0.13267 0.00017491 0.7575 0.0098219 0.010845 0.0014233 0.98646 0.99139 3.074e-006 1.2296e-005 0.16807 0.83368 0.87192 0.0014165 0.9498 0.41257 0.0019077 0.41946 2.0315 2.0299 16.0281 144.8887 0.00023113 -85.4939 0.45894
9.563 0.98816 5.4557e-005 3.8183 0.0119 0.00012406 0.0011801 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.672 0.62799 0.19133 0.02146 21.0405 0.13268 0.00017492 0.7575 0.0098222 0.010846 0.001423 0.98647 0.99139 3.0733e-006 1.2293e-005 0.16807 0.83415 0.87216 0.0014164 0.9501 0.41277 0.0019075 0.41947 2.0326 2.031 16.0281 144.8887 0.00023076 -85.4951 0.45994
9.564 0.98816 5.4557e-005 3.8183 0.0119 0.00012407 0.0011802 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6721 0.62804 0.19135 0.021461 21.044 0.13268 0.00017493 0.75749 0.0098225 0.010846 0.0014227 0.98647 0.9914 3.0726e-006 1.229e-005 0.16808 0.83461 0.87239 0.0014162 0.95041 0.41298 0.0019073 0.41949 2.0337 2.0321 16.0281 144.8888 0.0002304 -85.4963 0.46094
9.565 0.98816 5.4557e-005 3.8183 0.0119 0.00012408 0.0011802 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6722 0.62808 0.19136 0.021462 21.0474 0.13269 0.00017494 0.75749 0.0098228 0.010846 0.0014224 0.98648 0.9914 3.0719e-006 1.2288e-005 0.16808 0.83508 0.87262 0.0014161 0.95071 0.41318 0.0019071 0.41951 2.0348 2.0332 16.0281 144.8888 0.00023004 -85.4976 0.46194
9.566 0.98816 5.4557e-005 3.8183 0.0119 0.0001241 0.0011802 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6723 0.62812 0.19137 0.021463 21.0509 0.13269 0.00017495 0.75748 0.0098231 0.010847 0.0014222 0.98648 0.9914 3.0713e-006 1.2285e-005 0.16808 0.83554 0.87286 0.0014159 0.951 0.41338 0.0019069 0.41952 2.0359 2.0343 16.0281 144.8888 0.00022968 -85.4988 0.46294
9.567 0.98816 5.4557e-005 3.8183 0.0119 0.00012411 0.0011802 0.23345 0.00065931 0.23411 0.21603 0 0.032271 0.0389 0 1.6724 0.62817 0.19138 0.021464 21.0543 0.1327 0.00017496 0.75747 0.0098234 0.010847 0.0014219 0.98648 0.9914 3.0706e-006 1.2282e-005 0.16808 0.836 0.87309 0.0014158 0.9513 0.41359 0.0019067 0.41954 2.037 2.0355 16.0281 144.8888 0.00022932 -85.5 0.46394
9.568 0.98816 5.4557e-005 3.8183 0.0119 0.00012412 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6725 0.62821 0.1914 0.021465 21.0578 0.13271 0.00017497 0.75747 0.0098238 0.010847 0.0014216 0.98649 0.99141 3.07e-006 1.228e-005 0.16808 0.83647 0.87332 0.0014156 0.95159 0.41379 0.0019065 0.41955 2.0381 2.0366 16.0281 144.8888 0.00022897 -85.5012 0.46494
9.569 0.98816 5.4557e-005 3.8183 0.0119 0.00012413 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6725 0.62826 0.19141 0.021466 21.0612 0.13271 0.00017497 0.75746 0.0098241 0.010848 0.0014213 0.98649 0.99141 3.0693e-006 1.2277e-005 0.16809 0.83692 0.87355 0.0014155 0.95189 0.41399 0.0019063 0.41957 2.0392 2.0376 16.0281 144.8888 0.00022861 -85.5024 0.46594
9.57 0.98816 5.4556e-005 3.8183 0.0119 0.00012415 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6726 0.6283 0.19142 0.021467 21.0647 0.13272 0.00017498 0.75746 0.0098244 0.010848 0.001421 0.98649 0.99141 3.0687e-006 1.2275e-005 0.16809 0.83738 0.87377 0.0014153 0.95218 0.4142 0.0019061 0.41958 2.0403 2.0387 16.0281 144.8889 0.00022826 -85.5036 0.46694
9.571 0.98816 5.4556e-005 3.8183 0.0119 0.00012416 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6727 0.62834 0.19144 0.021468 21.0681 0.13272 0.00017499 0.75745 0.0098247 0.010848 0.0014207 0.9865 0.99141 3.068e-006 1.2272e-005 0.16809 0.83784 0.874 0.0014152 0.95246 0.4144 0.0019059 0.4196 2.0414 2.0398 16.0281 144.8889 0.00022791 -85.5047 0.46794
9.572 0.98816 5.4556e-005 3.8183 0.0119 0.00012417 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6728 0.62839 0.19145 0.021469 21.0716 0.13273 0.000175 0.75745 0.009825 0.010849 0.0014205 0.9865 0.99142 3.0674e-006 1.227e-005 0.16809 0.83829 0.87423 0.001415 0.95275 0.4146 0.0019057 0.41961 2.0425 2.0409 16.0281 144.8889 0.00022756 -85.5059 0.46894
9.573 0.98816 5.4556e-005 3.8183 0.0119 0.00012418 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6729 0.62843 0.19146 0.02147 21.075 0.13273 0.00017501 0.75744 0.0098253 0.010849 0.0014202 0.9865 0.99142 3.0668e-006 1.2267e-005 0.1681 0.83875 0.87445 0.0014149 0.95304 0.41481 0.0019055 0.41963 2.0435 2.042 16.0281 144.8889 0.00022721 -85.5071 0.46994
9.574 0.98816 5.4556e-005 3.8183 0.0119 0.0001242 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032271 0.0389 0 1.6729 0.62847 0.19147 0.021471 21.0785 0.13274 0.00017502 0.75744 0.0098256 0.010849 0.0014199 0.98651 0.99142 3.0662e-006 1.2265e-005 0.1681 0.8392 0.87468 0.0014148 0.95332 0.41501 0.0019053 0.41964 2.0446 2.0431 16.0281 144.8889 0.00022686 -85.5082 0.47094
9.575 0.98816 5.4556e-005 3.8183 0.0119 0.00012421 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.673 0.62852 0.19149 0.021472 21.082 0.13275 0.00017503 0.75743 0.0098259 0.01085 0.0014196 0.98651 0.99142 3.0655e-006 1.2262e-005 0.1681 0.83965 0.8749 0.0014146 0.9536 0.41521 0.0019052 0.41966 2.0457 2.0442 16.0281 144.889 0.00022652 -85.5094 0.47194
9.576 0.98816 5.4556e-005 3.8183 0.0119 0.00012422 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.6731 0.62856 0.1915 0.021473 21.0854 0.13275 0.00017504 0.75742 0.0098262 0.01085 0.0014194 0.98651 0.99142 3.0649e-006 1.226e-005 0.1681 0.8401 0.87512 0.0014145 0.95388 0.41542 0.001905 0.41967 2.0468 2.0452 16.028 144.889 0.00022617 -85.5105 0.47294
9.577 0.98816 5.4556e-005 3.8183 0.0119 0.00012424 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.6732 0.62861 0.19151 0.021474 21.0889 0.13276 0.00017504 0.75742 0.0098265 0.01085 0.0014191 0.98652 0.99143 3.0643e-006 1.2257e-005 0.16811 0.84054 0.87534 0.0014143 0.95416 0.41562 0.0019048 0.41969 2.0478 2.0463 16.028 144.889 0.00022583 -85.5116 0.47394
9.578 0.98816 5.4556e-005 3.8183 0.0119 0.00012425 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.6733 0.62865 0.19152 0.021475 21.0923 0.13276 0.00017505 0.75741 0.0098269 0.010851 0.0014189 0.98652 0.99143 3.0637e-006 1.2255e-005 0.16811 0.84099 0.87556 0.0014142 0.95443 0.41582 0.0019046 0.4197 2.0489 2.0474 16.028 144.889 0.00022549 -85.5127 0.47494
9.579 0.98816 5.4556e-005 3.8183 0.0119 0.00012426 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.6733 0.62869 0.19154 0.021476 21.0958 0.13277 0.00017506 0.75741 0.0098272 0.010851 0.0014186 0.98653 0.99143 3.0631e-006 1.2252e-005 0.16811 0.84144 0.87578 0.0014141 0.95471 0.41602 0.0019044 0.41972 2.05 2.0485 16.028 144.889 0.00022515 -85.5138 0.47594
9.58 0.98816 5.4556e-005 3.8183 0.011899 0.00012427 0.0011802 0.23345 0.00065931 0.23411 0.21602 0 0.032272 0.0389 0 1.6734 0.62874 0.19155 0.021477 21.0992 0.13277 0.00017507 0.7574 0.0098275 0.010851 0.0014183 0.98653 0.99143 3.0625e-006 1.225e-005 0.16811 0.84188 0.876 0.001414 0.95498 0.41623 0.0019043 0.41974 2.051 2.0495 16.028 144.8891 0.00022481 -85.5149 0.47694
9.581 0.98816 5.4556e-005 3.8183 0.011899 0.00012429 0.0011802 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6735 0.62878 0.19156 0.021478 21.1027 0.13278 0.00017508 0.7574 0.0098278 0.010852 0.0014181 0.98653 0.99144 3.0619e-006 1.2248e-005 0.16812 0.84232 0.87622 0.0014138 0.95525 0.41643 0.0019041 0.41975 2.0521 2.0506 16.028 144.8891 0.00022447 -85.516 0.47794
9.582 0.98816 5.4555e-005 3.8183 0.011899 0.0001243 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6736 0.62883 0.19157 0.021479 21.1062 0.13278 0.00017509 0.75739 0.0098281 0.010852 0.0014178 0.98654 0.99144 3.0613e-006 1.2245e-005 0.16812 0.84276 0.87644 0.0014137 0.95552 0.41663 0.0019039 0.41977 2.0531 2.0516 16.028 144.8891 0.00022413 -85.5171 0.47894
9.583 0.98816 5.4555e-005 3.8183 0.011899 0.00012431 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6737 0.62887 0.19159 0.021479 21.1096 0.13279 0.0001751 0.75738 0.0098284 0.010852 0.0014176 0.98654 0.99144 3.0608e-006 1.2243e-005 0.16812 0.8432 0.87665 0.0014136 0.95579 0.41683 0.0019037 0.41978 2.0542 2.0527 16.028 144.8891 0.0002238 -85.5182 0.47994
9.584 0.98816 5.4555e-005 3.8183 0.011899 0.00012432 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6738 0.62891 0.1916 0.02148 21.1131 0.1328 0.0001751 0.75738 0.0098287 0.010853 0.0014173 0.98654 0.99144 3.0602e-006 1.2241e-005 0.16812 0.84364 0.87687 0.0014134 0.95605 0.41704 0.0019036 0.4198 2.0552 2.0538 16.028 144.8891 0.00022347 -85.5193 0.48094
9.585 0.98816 5.4555e-005 3.8183 0.011899 0.00012434 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6738 0.62896 0.19161 0.021481 21.1165 0.1328 0.00017511 0.75737 0.009829 0.010853 0.0014171 0.98655 0.99144 3.0596e-006 1.2238e-005 0.16813 0.84408 0.87708 0.0014133 0.95632 0.41724 0.0019034 0.41981 2.0563 2.0548 16.028 144.8892 0.00022314 -85.5203 0.48194
9.586 0.98816 5.4555e-005 3.8183 0.011899 0.00012435 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6739 0.629 0.19162 0.021482 21.12 0.13281 0.00017512 0.75737 0.0098293 0.010853 0.0014168 0.98655 0.99145 3.059e-006 1.2236e-005 0.16813 0.84451 0.8773 0.0014132 0.95658 0.41744 0.0019032 0.41983 2.0573 2.0559 16.028 144.8892 0.00022281 -85.5214 0.48294
9.587 0.98816 5.4555e-005 3.8183 0.011899 0.00012436 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.674 0.62904 0.19164 0.021483 21.1235 0.13281 0.00017513 0.75736 0.0098296 0.010854 0.0014166 0.98655 0.99145 3.0585e-006 1.2234e-005 0.16813 0.84495 0.87751 0.001413 0.95684 0.41764 0.001903 0.41984 2.0584 2.0569 16.028 144.8892 0.00022248 -85.5224 0.48394
9.588 0.98816 5.4555e-005 3.8183 0.011899 0.00012438 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6741 0.62909 0.19165 0.021484 21.1269 0.13282 0.00017514 0.75736 0.00983 0.010854 0.0014163 0.98655 0.99145 3.0579e-006 1.2232e-005 0.16813 0.84538 0.87772 0.0014129 0.9571 0.41785 0.0019029 0.41986 2.0594 2.0579 16.028 144.8892 0.00022215 -85.5234 0.48494
9.589 0.98816 5.4555e-005 3.8183 0.011899 0.00012439 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6742 0.62913 0.19166 0.021485 21.1304 0.13282 0.00017515 0.75735 0.0098303 0.010854 0.0014161 0.98656 0.99145 3.0574e-006 1.2229e-005 0.16813 0.84581 0.87793 0.0014128 0.95736 0.41805 0.0019027 0.41987 2.0604 2.059 16.028 144.8892 0.00022182 -85.5245 0.48594
9.59 0.98816 5.4555e-005 3.8183 0.011899 0.0001244 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6742 0.62918 0.19167 0.021486 21.1338 0.13283 0.00017516 0.75735 0.0098306 0.010855 0.0014158 0.98656 0.99145 3.0568e-006 1.2227e-005 0.16814 0.84624 0.87814 0.0014126 0.95761 0.41825 0.0019025 0.41989 2.0615 2.06 16.0279 144.8893 0.0002215 -85.5255 0.48694
9.591 0.98816 5.4555e-005 3.8183 0.011899 0.00012441 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6743 0.62922 0.19169 0.021487 21.1373 0.13284 0.00017517 0.75734 0.0098309 0.010855 0.0014156 0.98656 0.99146 3.0562e-006 1.2225e-005 0.16814 0.84667 0.87835 0.0014125 0.95787 0.41845 0.0019024 0.4199 2.0625 2.061 16.0279 144.8893 0.00022118 -85.5265 0.48794
9.592 0.98816 5.4555e-005 3.8183 0.011899 0.00012443 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6744 0.62926 0.1917 0.021488 21.1408 0.13284 0.00017517 0.75733 0.0098312 0.010855 0.0014154 0.98657 0.99146 3.0557e-006 1.2223e-005 0.16814 0.84709 0.87856 0.0014124 0.95812 0.41865 0.0019022 0.41992 2.0635 2.0621 16.0279 144.8893 0.00022085 -85.5275 0.48894
9.593 0.98816 5.4554e-005 3.8183 0.011899 0.00012444 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6745 0.62931 0.19171 0.021489 21.1442 0.13285 0.00017518 0.75733 0.0098315 0.010856 0.0014151 0.98657 0.99146 3.0552e-006 1.2221e-005 0.16814 0.84752 0.87877 0.0014123 0.95837 0.41886 0.0019021 0.41993 2.0645 2.0631 16.0279 144.8893 0.00022053 -85.5285 0.48994
9.594 0.98816 5.4554e-005 3.8183 0.011899 0.00012445 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6746 0.62935 0.19172 0.02149 21.1477 0.13285 0.00017519 0.75732 0.0098318 0.010856 0.0014149 0.98657 0.99146 3.0546e-006 1.2218e-005 0.16815 0.84794 0.87897 0.0014121 0.95862 0.41906 0.0019019 0.41995 2.0656 2.0641 16.0279 144.8893 0.00022021 -85.5295 0.49094
9.595 0.98816 5.4554e-005 3.8183 0.011899 0.00012447 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6746 0.62939 0.19174 0.021491 21.1512 0.13286 0.0001752 0.75732 0.0098321 0.010856 0.0014147 0.98658 0.99146 3.0541e-006 1.2216e-005 0.16815 0.84837 0.87918 0.001412 0.95887 0.41926 0.0019017 0.41997 2.0666 2.0651 16.0279 144.8894 0.0002199 -85.5305 0.49194
9.596 0.98816 5.4554e-005 3.8183 0.011899 0.00012448 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6747 0.62944 0.19175 0.021492 21.1546 0.13286 0.00017521 0.75731 0.0098324 0.010857 0.0014144 0.98658 0.99147 3.0536e-006 1.2214e-005 0.16815 0.84879 0.87938 0.0014119 0.95911 0.41946 0.0019016 0.41998 2.0676 2.0662 16.0279 144.8894 0.00021958 -85.5315 0.49294
9.597 0.98816 5.4554e-005 3.8183 0.011899 0.00012449 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6748 0.62948 0.19176 0.021493 21.1581 0.13287 0.00017522 0.75731 0.0098327 0.010857 0.0014142 0.98658 0.99147 3.053e-006 1.2212e-005 0.16815 0.84921 0.87959 0.0014118 0.95936 0.41966 0.0019014 0.42 2.0686 2.0672 16.0279 144.8894 0.00021926 -85.5324 0.49394
9.598 0.98816 5.4554e-005 3.8183 0.011899 0.0001245 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6749 0.62953 0.19177 0.021494 21.1615 0.13287 0.00017523 0.7573 0.0098331 0.010857 0.001414 0.98659 0.99147 3.0525e-006 1.221e-005 0.16816 0.84963 0.87979 0.0014117 0.9596 0.41986 0.0019013 0.42001 2.0696 2.0682 16.0279 144.8894 0.00021895 -85.5334 0.49494
9.599 0.98816 5.4554e-005 3.8183 0.011899 0.00012452 0.0011803 0.23345 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.675 0.62957 0.19179 0.021495 21.165 0.13288 0.00017524 0.7573 0.0098334 0.010858 0.0014137 0.98659 0.99147 3.052e-006 1.2208e-005 0.16816 0.85005 0.87999 0.0014115 0.95984 0.42007 0.0019011 0.42003 2.0706 2.0692 16.0279 144.8894 0.00021864 -85.5344 0.49594
9.6 0.98816 5.4554e-005 3.8183 0.011899 0.00012453 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6751 0.62961 0.1918 0.021496 21.1685 0.13289 0.00017524 0.75729 0.0098337 0.010858 0.0014135 0.98659 0.99147 3.0515e-006 1.2206e-005 0.16816 0.85046 0.88019 0.0014114 0.96008 0.42027 0.001901 0.42004 2.0716 2.0702 16.0279 144.8895 0.00021833 -85.5353 0.49694
9.601 0.98816 5.4554e-005 3.8183 0.011899 0.00012454 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6751 0.62966 0.19181 0.021497 21.1719 0.13289 0.00017525 0.75728 0.009834 0.010858 0.0014133 0.98659 0.99148 3.051e-006 1.2204e-005 0.16816 0.85088 0.8804 0.0014113 0.96032 0.42047 0.0019008 0.42006 2.0726 2.0712 16.0278 144.8895 0.00021802 -85.5362 0.49794
9.602 0.98816 5.4554e-005 3.8183 0.011899 0.00012455 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6752 0.6297 0.19182 0.021498 21.1754 0.1329 0.00017526 0.75728 0.0098343 0.010859 0.0014131 0.9866 0.99148 3.0505e-006 1.2202e-005 0.16817 0.85129 0.8806 0.0014112 0.96056 0.42067 0.0019007 0.42007 2.0736 2.0722 16.0278 144.8895 0.00021771 -85.5372 0.49894
9.603 0.98816 5.4554e-005 3.8183 0.011899 0.00012457 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6753 0.62974 0.19184 0.021498 21.1789 0.1329 0.00017527 0.75727 0.0098346 0.010859 0.0014129 0.9866 0.99148 3.05e-006 1.22e-005 0.16817 0.85171 0.88079 0.0014111 0.96079 0.42087 0.0019005 0.42009 2.0746 2.0732 16.0278 144.8895 0.0002174 -85.5381 0.49994
9.604 0.98816 5.4554e-005 3.8183 0.011899 0.00012458 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6754 0.62979 0.19185 0.021499 21.1823 0.13291 0.00017528 0.75727 0.0098349 0.010859 0.0014126 0.9866 0.99148 3.0495e-006 1.2198e-005 0.16817 0.85212 0.88099 0.001411 0.96103 0.42107 0.0019004 0.4201 2.0756 2.0742 16.0278 144.8895 0.00021709 -85.539 0.50094
9.605 0.98816 5.4553e-005 3.8183 0.011899 0.00012459 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6755 0.62983 0.19186 0.0215 21.1858 0.13291 0.00017529 0.75726 0.0098352 0.010859 0.0014124 0.98661 0.99148 3.049e-006 1.2196e-005 0.16817 0.85253 0.88119 0.0014108 0.96126 0.42127 0.0019002 0.42012 2.0766 2.0752 16.0278 144.8896 0.00021679 -85.5399 0.50194
9.606 0.98816 5.4553e-005 3.8183 0.011899 0.00012461 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6755 0.62988 0.19187 0.021501 21.1893 0.13292 0.0001753 0.75726 0.0098355 0.01086 0.0014122 0.98661 0.99149 3.0485e-006 1.2194e-005 0.16817 0.85294 0.88139 0.0014107 0.96149 0.42147 0.0019001 0.42014 2.0776 2.0762 16.0278 144.8896 0.00021648 -85.5409 0.50294
9.607 0.98816 5.4553e-005 3.8183 0.011899 0.00012462 0.0011804 0.23344 0.00065931 0.2341 0.21602 0 0.032272 0.0389 0 1.6756 0.62992 0.19189 0.021502 21.1927 0.13292 0.0001753 0.75725 0.0098358 0.01086 0.001412 0.98661 0.99149 3.048e-006 1.2192e-005 0.16818 0.85335 0.88158 0.0014106 0.96172 0.42168 0.0018999 0.42015 2.0786 2.0772 16.0278 144.8896 0.00021618 -85.5418 0.50394
9.608 0.98816 5.4553e-005 3.8183 0.011899 0.00012463 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6757 0.62996 0.1919 0.021503 21.1962 0.13293 0.00017531 0.75724 0.0098361 0.01086 0.0014118 0.98661 0.99149 3.0475e-006 1.219e-005 0.16818 0.85375 0.88178 0.0014105 0.96195 0.42188 0.0018998 0.42017 2.0796 2.0782 16.0278 144.8896 0.00021588 -85.5427 0.50494
9.609 0.98816 5.4553e-005 3.8183 0.011899 0.00012464 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6758 0.63001 0.19191 0.021504 21.1997 0.13294 0.00017532 0.75724 0.0098364 0.010861 0.0014116 0.98662 0.99149 3.0471e-006 1.2188e-005 0.16818 0.85416 0.88197 0.0014104 0.96218 0.42208 0.0018996 0.42018 2.0805 2.0792 16.0278 144.8896 0.00021558 -85.5435 0.50594
9.61 0.98816 5.4553e-005 3.8183 0.011899 0.00012466 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6759 0.63005 0.19192 0.021505 21.2031 0.13294 0.00017533 0.75723 0.0098368 0.010861 0.0014114 0.98662 0.99149 3.0466e-006 1.2186e-005 0.16818 0.85456 0.88217 0.0014103 0.9624 0.42228 0.0018995 0.4202 2.0815 2.0801 16.0278 144.8897 0.00021528 -85.5444 0.50694
9.611 0.98816 5.4553e-005 3.8183 0.011899 0.00012467 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6759 0.63009 0.19194 0.021506 21.2066 0.13295 0.00017534 0.75723 0.0098371 0.010861 0.0014112 0.98662 0.99149 3.0461e-006 1.2184e-005 0.16819 0.85496 0.88236 0.0014102 0.96263 0.42248 0.0018993 0.42021 2.0825 2.0811 16.0277 144.8897 0.00021498 -85.5453 0.50794
9.612 0.98816 5.4553e-005 3.8183 0.011899 0.00012468 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.676 0.63014 0.19195 0.021507 21.2101 0.13295 0.00017535 0.75722 0.0098374 0.010862 0.001411 0.98662 0.9915 3.0456e-006 1.2182e-005 0.16819 0.85536 0.88255 0.0014101 0.96285 0.42268 0.0018992 0.42023 2.0835 2.0821 16.0277 144.8897 0.00021469 -85.5462 0.50894
9.613 0.98816 5.4553e-005 3.8183 0.011899 0.00012469 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6761 0.63018 0.19196 0.021508 21.2135 0.13296 0.00017536 0.75722 0.0098377 0.010862 0.0014108 0.98663 0.9915 3.0451e-006 1.2181e-005 0.16819 0.85576 0.88274 0.0014099 0.96307 0.42288 0.0018991 0.42024 2.0844 2.0831 16.0277 144.8897 0.00021439 -85.547 0.50994
9.614 0.98816 5.4553e-005 3.8183 0.011899 0.00012471 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6762 0.63023 0.19198 0.021509 21.217 0.13296 0.00017537 0.75721 0.009838 0.010862 0.0014105 0.98663 0.9915 3.0447e-006 1.2179e-005 0.16819 0.85616 0.88293 0.0014098 0.96329 0.42308 0.0018989 0.42026 2.0854 2.084 16.0277 144.8897 0.0002141 -85.5479 0.51094
9.615 0.98816 5.4553e-005 3.8183 0.011899 0.00012472 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6763 0.63027 0.19199 0.02151 21.2205 0.13297 0.00017537 0.75721 0.0098383 0.010863 0.0014103 0.98663 0.9915 3.0442e-006 1.2177e-005 0.1682 0.85656 0.88312 0.0014097 0.96351 0.42328 0.0018988 0.42027 2.0863 2.085 16.0277 144.8898 0.00021381 -85.5487 0.51194
9.616 0.98816 5.4553e-005 3.8183 0.011899 0.00012473 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6764 0.63031 0.192 0.021511 21.224 0.13298 0.00017538 0.7572 0.0098386 0.010863 0.0014102 0.98663 0.9915 3.0438e-006 1.2175e-005 0.1682 0.85696 0.88331 0.0014096 0.96372 0.42348 0.0018987 0.42029 2.0873 2.086 16.0277 144.8898 0.00021352 -85.5496 0.51294
9.617 0.98816 5.4552e-005 3.8183 0.011899 0.00012475 0.0011804 0.23344 0.00065931 0.2341 0.21601 0 0.032272 0.0389 0 1.6764 0.63036 0.19201 0.021512 21.2274 0.13298 0.00017539 0.75719 0.0098389 0.010863 0.00141 0.98664 0.9915 3.0433e-006 1.2173e-005 0.1682 0.85735 0.8835 0.0014095 0.96394 0.42368 0.0018985 0.42031 2.0883 2.0869 16.0277 144.8898 0.00021323 -85.5504 0.51394
9.618 0.98816 5.4552e-005 3.8183 0.011899 0.00012476 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6765 0.6304 0.19203 0.021513 21.2309 0.13299 0.0001754 0.75719 0.0098392 0.010864 0.0014098 0.98664 0.99151 3.0429e-006 1.2171e-005 0.1682 0.85775 0.88369 0.0014094 0.96415 0.42388 0.0018984 0.42032 2.0892 2.0879 16.0277 144.8898 0.00021294 -85.5513 0.51494
9.619 0.98816 5.4552e-005 3.8183 0.011899 0.00012477 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6766 0.63045 0.19204 0.021514 21.2344 0.13299 0.00017541 0.75718 0.0098395 0.010864 0.0014096 0.98664 0.99151 3.0424e-006 1.217e-005 0.16821 0.85814 0.88387 0.0014093 0.96437 0.42408 0.0018983 0.42034 2.0902 2.0888 16.0277 144.8898 0.00021265 -85.5521 0.51594
9.62 0.98816 5.4552e-005 3.8183 0.011899 0.00012478 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6767 0.63049 0.19205 0.021515 21.2378 0.133 0.00017542 0.75718 0.0098398 0.010864 0.0014094 0.98665 0.99151 3.042e-006 1.2168e-005 0.16821 0.85853 0.88406 0.0014092 0.96458 0.42428 0.0018981 0.42035 2.0911 2.0898 16.0276 144.8899 0.00021236 -85.5529 0.51694
9.621 0.98816 5.4552e-005 3.8183 0.011899 0.0001248 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6768 0.63053 0.19206 0.021516 21.2413 0.133 0.00017543 0.75717 0.0098401 0.010865 0.0014092 0.98665 0.99151 3.0415e-006 1.2166e-005 0.16821 0.85892 0.88424 0.0014091 0.96479 0.42448 0.001898 0.42037 2.0921 2.0908 16.0276 144.8899 0.00021208 -85.5537 0.51794
9.622 0.98816 5.4552e-005 3.8183 0.011899 0.00012481 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6768 0.63058 0.19208 0.021517 21.2448 0.13301 0.00017543 0.75717 0.0098405 0.010865 0.001409 0.98665 0.99151 3.0411e-006 1.2164e-005 0.16821 0.85931 0.88443 0.001409 0.965 0.42468 0.0018979 0.42038 2.093 2.0917 16.0276 144.8899 0.00021179 -85.5545 0.51894
9.623 0.98816 5.4552e-005 3.8183 0.011899 0.00012482 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6769 0.63062 0.19209 0.021517 21.2482 0.13301 0.00017544 0.75716 0.0098408 0.010865 0.0014088 0.98665 0.99151 3.0407e-006 1.2163e-005 0.16821 0.8597 0.88461 0.0014089 0.9652 0.42488 0.0018977 0.4204 2.094 2.0926 16.0276 144.8899 0.00021151 -85.5553 0.51994
9.624 0.98816 5.4552e-005 3.8183 0.011899 0.00012483 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.677 0.63066 0.1921 0.021518 21.2517 0.13302 0.00017545 0.75716 0.0098411 0.010866 0.0014086 0.98665 0.99152 3.0403e-006 1.2161e-005 0.16822 0.86008 0.88479 0.0014088 0.96541 0.42508 0.0018976 0.42041 2.0949 2.0936 16.0276 144.8899 0.00021123 -85.5561 0.52094
9.625 0.98816 5.4552e-005 3.8183 0.011899 0.00012485 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6771 0.63071 0.19211 0.021519 21.2552 0.13303 0.00017546 0.75715 0.0098414 0.010866 0.0014084 0.98666 0.99152 3.0398e-006 1.2159e-005 0.16822 0.86047 0.88498 0.0014087 0.96561 0.42528 0.0018975 0.42043 2.0958 2.0945 16.0276 144.89 0.00021095 -85.5569 0.52194
9.626 0.98816 5.4552e-005 3.8183 0.011899 0.00012486 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6772 0.63075 0.19213 0.02152 21.2587 0.13303 0.00017547 0.75714 0.0098417 0.010866 0.0014082 0.98666 0.99152 3.0394e-006 1.2158e-005 0.16822 0.86085 0.88516 0.0014086 0.96582 0.42548 0.0018973 0.42045 2.0968 2.0955 16.0276 144.89 0.00021067 -85.5577 0.52294
9.627 0.98816 5.4552e-005 3.8183 0.011899 0.00012487 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6772 0.6308 0.19214 0.021521 21.2621 0.13304 0.00017548 0.75714 0.009842 0.010867 0.0014081 0.98666 0.99152 3.039e-006 1.2156e-005 0.16822 0.86124 0.88534 0.0014086 0.96602 0.42568 0.0018972 0.42046 2.0977 2.0964 16.0276 144.89 0.00021039 -85.5585 0.52394
9.628 0.98816 5.4552e-005 3.8183 0.011899 0.00012489 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6773 0.63084 0.19215 0.021522 21.2656 0.13304 0.00017549 0.75713 0.0098423 0.010867 0.0014079 0.98666 0.99152 3.0386e-006 1.2154e-005 0.16823 0.86162 0.88552 0.0014085 0.96622 0.42588 0.0018971 0.42048 2.0986 2.0973 16.0275 144.89 0.00021011 -85.5592 0.52494
9.629 0.98816 5.4551e-005 3.8183 0.011899 0.0001249 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6774 0.63088 0.19216 0.021523 21.2691 0.13305 0.0001755 0.75713 0.0098426 0.010867 0.0014077 0.98667 0.99152 3.0382e-006 1.2153e-005 0.16823 0.862 0.8857 0.0014084 0.96642 0.42608 0.001897 0.42049 2.0996 2.0983 16.0275 144.89 0.00020983 -85.56 0.52594
9.63 0.98816 5.4551e-005 3.8183 0.011899 0.00012491 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6775 0.63093 0.19218 0.021524 21.2726 0.13305 0.0001755 0.75712 0.0098429 0.010868 0.0014075 0.98667 0.99153 3.0378e-006 1.2151e-005 0.16823 0.86238 0.88588 0.0014083 0.96662 0.42628 0.0018969 0.42051 2.1005 2.0992 16.0275 144.89 0.00020956 -85.5608 0.52694
9.631 0.98816 5.4551e-005 3.8183 0.011899 0.00012492 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6776 0.63097 0.19219 0.021525 21.276 0.13306 0.00017551 0.75712 0.0098432 0.010868 0.0014073 0.98667 0.99153 3.0374e-006 1.215e-005 0.16823 0.86276 0.88605 0.0014082 0.96682 0.42648 0.0018967 0.42052 2.1014 2.1001 16.0275 144.8901 0.00020928 -85.5615 0.52794
9.632 0.98816 5.4551e-005 3.8183 0.011899 0.00012494 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6777 0.63101 0.1922 0.021526 21.2795 0.13306 0.00017552 0.75711 0.0098435 0.010868 0.0014072 0.98667 0.99153 3.037e-006 1.2148e-005 0.16824 0.86313 0.88623 0.0014081 0.96701 0.42668 0.0018966 0.42054 2.1023 2.1011 16.0275 144.8901 0.00020901 -85.5623 0.52894
9.633 0.98816 5.4551e-005 3.8183 0.011899 0.00012495 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6777 0.63106 0.19221 0.021527 21.283 0.13307 0.00017553 0.75711 0.0098438 0.010869 0.001407 0.98668 0.99153 3.0366e-006 1.2146e-005 0.16824 0.86351 0.88641 0.001408 0.96721 0.42688 0.0018965 0.42055 2.1032 2.102 16.0275 144.8901 0.00020874 -85.563 0.52994
9.634 0.98816 5.4551e-005 3.8183 0.011898 0.00012496 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6778 0.6311 0.19223 0.021528 21.2865 0.13308 0.00017554 0.7571 0.0098442 0.010869 0.0014068 0.98668 0.99153 3.0362e-006 1.2145e-005 0.16824 0.86389 0.88658 0.0014079 0.9674 0.42708 0.0018964 0.42057 2.1042 2.1029 16.0275 144.8901 0.00020847 -85.5638 0.53094
9.635 0.98816 5.4551e-005 3.8183 0.011898 0.00012498 0.0011805 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6779 0.63115 0.19224 0.021529 21.2899 0.13308 0.00017555 0.75709 0.0098445 0.010869 0.0014066 0.98668 0.99153 3.0358e-006 1.2143e-005 0.16824 0.86426 0.88676 0.0014078 0.96759 0.42728 0.0018963 0.42058 2.1051 2.1038 16.0275 144.8901 0.0002082 -85.5645 0.53194
9.636 0.98816 5.4551e-005 3.8183 0.011898 0.00012499 0.0011806 0.23344 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.678 0.63119 0.19225 0.02153 21.2934 0.13309 0.00017556 0.75709 0.0098448 0.01087 0.0014065 0.98668 0.99153 3.0354e-006 1.2141e-005 0.16825 0.86463 0.88693 0.0014077 0.96778 0.42747 0.0018961 0.4206 2.106 2.1047 16.0274 144.8902 0.00020793 -85.5652 0.53294
9.637 0.98816 5.4551e-005 3.8183 0.011898 0.000125 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6781 0.63123 0.19226 0.021531 21.2969 0.13309 0.00017556 0.75708 0.0098451 0.01087 0.0014063 0.98668 0.99154 3.035e-006 1.214e-005 0.16825 0.865 0.88711 0.0014076 0.96797 0.42767 0.001896 0.42062 2.1069 2.1056 16.0274 144.8902 0.00020766 -85.566 0.53394
9.638 0.98816 5.4551e-005 3.8183 0.011898 0.00012501 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6781 0.63128 0.19228 0.021532 21.3004 0.1331 0.00017557 0.75708 0.0098454 0.01087 0.0014061 0.98669 0.99154 3.0346e-006 1.2138e-005 0.16825 0.86537 0.88728 0.0014075 0.96816 0.42787 0.0018959 0.42063 2.1078 2.1065 16.0274 144.8902 0.0002074 -85.5667 0.53494
9.639 0.98816 5.4551e-005 3.8183 0.011898 0.00012503 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6782 0.63132 0.19229 0.021533 21.3038 0.1331 0.00017558 0.75707 0.0098457 0.010871 0.001406 0.98669 0.99154 3.0342e-006 1.2137e-005 0.16825 0.86574 0.88745 0.0014075 0.96835 0.42807 0.0018958 0.42065 2.1087 2.1075 16.0274 144.8902 0.00020713 -85.5674 0.53594
9.64 0.98816 5.455e-005 3.8183 0.011898 0.00012504 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6783 0.63136 0.1923 0.021534 21.3073 0.13311 0.00017559 0.75707 0.009846 0.010871 0.0014058 0.98669 0.99154 3.0338e-006 1.2135e-005 0.16825 0.86611 0.88762 0.0014074 0.96853 0.42827 0.0018957 0.42066 2.1096 2.1084 16.0274 144.8902 0.00020687 -85.5681 0.53694
9.641 0.98816 5.455e-005 3.8183 0.011898 0.00012505 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6784 0.63141 0.19231 0.021534 21.3108 0.13311 0.0001756 0.75706 0.0098463 0.010871 0.0014056 0.98669 0.99154 3.0335e-006 1.2134e-005 0.16826 0.86648 0.88779 0.0014073 0.96872 0.42847 0.0018956 0.42068 2.1105 2.1093 16.0274 144.8903 0.0002066 -85.5688 0.53794
9.642 0.98816 5.455e-005 3.8183 0.011898 0.00012506 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6785 0.63145 0.19233 0.021535 21.3143 0.13312 0.00017561 0.75706 0.0098466 0.010871 0.0014055 0.9867 0.99154 3.0331e-006 1.2132e-005 0.16826 0.86684 0.88796 0.0014072 0.9689 0.42867 0.0018954 0.42069 2.1114 2.1102 16.0274 144.8903 0.00020634 -85.5695 0.53894
9.643 0.98816 5.455e-005 3.8183 0.011898 0.00012508 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6785 0.6315 0.19234 0.021536 21.3178 0.13313 0.00017562 0.75705 0.0098469 0.010872 0.0014053 0.9867 0.99154 3.0327e-006 1.2131e-005 0.16826 0.86721 0.88813 0.0014071 0.96908 0.42887 0.0018953 0.42071 2.1123 2.1111 16.0273 144.8903 0.00020608 -85.5702 0.53994
9.644 0.98816 5.455e-005 3.8183 0.011898 0.00012509 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6786 0.63154 0.19235 0.021537 21.3212 0.13313 0.00017563 0.75704 0.0098472 0.010872 0.0014052 0.9867 0.99155 3.0324e-006 1.2129e-005 0.16826 0.86757 0.8883 0.001407 0.96927 0.42907 0.0018952 0.42072 2.1132 2.1119 16.0273 144.8903 0.00020582 -85.5709 0.54094
9.645 0.98816 5.455e-005 3.8183 0.011898 0.0001251 0.0011806 0.23343 0.00065931 0.23409 0.21601 0 0.032272 0.0389 0 1.6787 0.63158 0.19236 0.021538 21.3247 0.13314 0.00017563 0.75704 0.0098475 0.010872 0.001405 0.9867 0.99155 3.032e-006 1.2128e-005 0.16827 0.86793 0.88847 0.0014069 0.96945 0.42926 0.0018951 0.42074 2.1141 2.1128 16.0273 144.8903 0.00020556 -85.5716 0.54194
9.646 0.98816 5.455e-005 3.8183 0.011898 0.00012512 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032272 0.0389 0 1.6788 0.63163 0.19238 0.021539 21.3282 0.13314 0.00017564 0.75703 0.0098478 0.010873 0.0014048 0.9867 0.99155 3.0316e-006 1.2126e-005 0.16827 0.86829 0.88864 0.0014068 0.96963 0.42946 0.001895 0.42076 2.115 2.1137 16.0273 144.8904 0.0002053 -85.5722 0.54294
9.647 0.98816 5.455e-005 3.8183 0.011898 0.00012513 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032272 0.0389 0 1.6789 0.63167 0.19239 0.02154 21.3317 0.13315 0.00017565 0.75703 0.0098481 0.010873 0.0014047 0.98671 0.99155 3.0312e-006 1.2125e-005 0.16827 0.86865 0.8888 0.0014068 0.9698 0.42966 0.0018949 0.42077 2.1158 2.1146 16.0273 144.8904 0.00020505 -85.5729 0.54394
9.648 0.98816 5.455e-005 3.8183 0.011898 0.00012514 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032272 0.0389 0 1.679 0.63171 0.1924 0.021541 21.3351 0.13315 0.00017566 0.75702 0.0098485 0.010873 0.0014045 0.98671 0.99155 3.0309e-006 1.2123e-005 0.16827 0.86901 0.88897 0.0014067 0.96998 0.42986 0.0018948 0.42079 2.1167 2.1155 16.0273 144.8904 0.00020479 -85.5736 0.54494
9.649 0.98816 5.455e-005 3.8183 0.011898 0.00012515 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.679 0.63176 0.19241 0.021542 21.3386 0.13316 0.00017567 0.75702 0.0098488 0.010874 0.0014044 0.98671 0.99155 3.0305e-006 1.2122e-005 0.16828 0.86937 0.88914 0.0014066 0.97016 0.43006 0.0018947 0.4208 2.1176 2.1164 16.0273 144.8904 0.00020454 -85.5742 0.54594
9.65 0.98816 5.455e-005 3.8183 0.011898 0.00012517 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.6791 0.6318 0.19243 0.021543 21.3421 0.13316 0.00017568 0.75701 0.0098491 0.010874 0.0014042 0.98671 0.99155 3.0302e-006 1.2121e-005 0.16828 0.86972 0.8893 0.0014065 0.97033 0.43026 0.0018946 0.42082 2.1185 2.1173 16.0272 144.8904 0.00020428 -85.5749 0.54694
9.651 0.98816 5.455e-005 3.8183 0.011898 0.00012518 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.6792 0.63185 0.19244 0.021544 21.3456 0.13317 0.00017569 0.75701 0.0098494 0.010874 0.0014041 0.98671 0.99155 3.0298e-006 1.2119e-005 0.16828 0.87008 0.88947 0.0014065 0.9705 0.43045 0.0018945 0.42083 2.1193 2.1181 16.0272 144.8905 0.00020403 -85.5756 0.54794
9.652 0.98816 5.4549e-005 3.8183 0.011898 0.00012519 0.0011806 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.6793 0.63189 0.19245 0.021545 21.3491 0.13318 0.00017569 0.757 0.0098497 0.010875 0.0014039 0.98672 0.99156 3.0295e-006 1.2118e-005 0.16828 0.87043 0.88963 0.0014064 0.97068 0.43065 0.0018944 0.42085 2.1202 2.119 16.0272 144.8905 0.00020378 -85.5762 0.54894
9.653 0.98816 5.4549e-005 3.8183 0.011898 0.0001252 0.0011807 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.6794 0.63193 0.19246 0.021546 21.3525 0.13318 0.0001757 0.75699 0.00985 0.010875 0.0014038 0.98672 0.99156 3.0292e-006 1.2117e-005 0.16828 0.87079 0.88979 0.0014063 0.97085 0.43085 0.0018943 0.42086 2.1211 2.1199 16.0272 144.8905 0.00020353 -85.5768 0.54994
9.654 0.98816 5.4549e-005 3.8183 0.011898 0.00012522 0.0011807 0.23343 0.00065931 0.23409 0.216 0 0.032273 0.0389 0 1.6794 0.63198 0.19248 0.021547 21.356 0.13319 0.00017571 0.75699 0.0098503 0.010875 0.0014036 0.98672 0.99156 3.0288e-006 1.2115e-005 0.16829 0.87114 0.88995 0.0014062 0.97102 0.43105 0.0018942 0.42088 2.122 2.1208 16.0272 144.8905 0.00020328 -85.5775 0.55094
9.655 0.98816 5.4549e-005 3.8183 0.011898 0.00012523 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6795 0.63202 0.19249 0.021548 21.3595 0.13319 0.00017572 0.75698 0.0098506 0.010876 0.0014035 0.98672 0.99156 3.0285e-006 1.2114e-005 0.16829 0.87149 0.89012 0.0014061 0.97119 0.43125 0.0018941 0.4209 2.1228 2.1216 16.0272 144.8905 0.00020303 -85.5781 0.55194
9.656 0.98816 5.4549e-005 3.8183 0.011898 0.00012524 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6796 0.63206 0.1925 0.021549 21.363 0.1332 0.00017573 0.75698 0.0098509 0.010876 0.0014033 0.98672 0.99156 3.0281e-006 1.2112e-005 0.16829 0.87184 0.89028 0.001406 0.97135 0.43144 0.001894 0.42091 2.1237 2.1225 16.0272 144.8906 0.00020278 -85.5788 0.55294
9.657 0.98816 5.4549e-005 3.8183 0.011898 0.00012526 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6797 0.63211 0.19251 0.02155 21.3665 0.1332 0.00017574 0.75697 0.0098512 0.010876 0.0014032 0.98673 0.99156 3.0277e-006 1.2111e-005 0.16829 0.87219 0.89044 0.0014059 0.97152 0.43164 0.0018939 0.42093 2.1245 2.1234 16.0271 144.8906 0.00020254 -85.5794 0.55394
9.658 0.98816 5.4549e-005 3.8183 0.011898 0.00012527 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6798 0.63215 0.19253 0.021551 21.37 0.13321 0.00017575 0.75697 0.0098515 0.010877 0.001403 0.98673 0.99156 3.0274e-006 1.211e-005 0.1683 0.87254 0.8906 0.0014058 0.97169 0.43184 0.0018938 0.42094 2.1254 2.1242 16.0271 144.8906 0.00020229 -85.58 0.55494
9.659 0.98816 5.4549e-005 3.8183 0.011898 0.00012528 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6798 0.6322 0.19254 0.021551 21.3734 0.13322 0.00017575 0.75696 0.0098518 0.010877 0.0014029 0.98673 0.99156 3.0271e-006 1.2108e-005 0.1683 0.87288 0.89076 0.0014058 0.97185 0.43204 0.0018937 0.42096 2.1263 2.1251 16.0271 144.8906 0.00020205 -85.5806 0.55594
9.66 0.98816 5.4549e-005 3.8183 0.011898 0.00012529 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6799 0.63224 0.19255 0.021552 21.3769 0.13322 0.00017576 0.75696 0.0098521 0.010877 0.0014027 0.98673 0.99157 3.0268e-006 1.2107e-005 0.1683 0.87323 0.89091 0.0014058 0.97202 0.43223 0.0018936 0.42097 2.1271 2.1259 16.0271 144.8906 0.0002018 -85.5812 0.55694
9.661 0.98816 5.4549e-005 3.8183 0.011898 0.00012531 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.68 0.63228 0.19256 0.021553 21.3804 0.13323 0.00017577 0.75695 0.0098524 0.010878 0.0014026 0.98673 0.99157 3.0265e-006 1.2106e-005 0.1683 0.87357 0.89107 0.0014058 0.97218 0.43243 0.0018935 0.42099 2.128 2.1268 16.0271 144.8907 0.00020156 -85.5818 0.55794
9.662 0.98816 5.4549e-005 3.8183 0.011898 0.00012532 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6801 0.63233 0.19258 0.021554 21.3839 0.13323 0.00017578 0.75694 0.0098527 0.010878 0.0014024 0.98673 0.99157 3.0263e-006 1.2105e-005 0.16831 0.87392 0.89123 0.0014058 0.97234 0.43263 0.0018934 0.421 2.1288 2.1276 16.0271 144.8907 0.00020132 -85.5824 0.55894
9.663 0.98816 5.4549e-005 3.8183 0.011898 0.00012533 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6802 0.63237 0.19259 0.021555 21.3874 0.13324 0.00017579 0.75694 0.009853 0.010878 0.0014023 0.98674 0.99157 3.026e-006 1.2104e-005 0.16831 0.87426 0.89139 0.0014057 0.9725 0.43283 0.0018933 0.42102 2.1297 2.1285 16.027 144.8907 0.00020108 -85.583 0.55994
9.664 0.98816 5.4548e-005 3.8183 0.011898 0.00012534 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6802 0.63241 0.1926 0.021556 21.3909 0.13324 0.0001758 0.75693 0.0098534 0.010879 0.0014022 0.98674 0.99157 3.0256e-006 1.2102e-005 0.16831 0.8746 0.89154 0.0014057 0.97266 0.43302 0.0018932 0.42103 2.1305 2.1293 16.027 144.8907 0.00020084 -85.5836 0.56094
9.665 0.98816 5.4548e-005 3.8183 0.011898 0.00012536 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6803 0.63246 0.19261 0.021557 21.3943 0.13325 0.00017581 0.75693 0.0098537 0.010879 0.001402 0.98674 0.99157 3.0253e-006 1.2101e-005 0.16831 0.87494 0.8917 0.0014056 0.97282 0.43322 0.0018931 0.42105 2.1313 2.1302 16.027 144.8907 0.0002006 -85.5842 0.56194
9.666 0.98816 5.4548e-005 3.8183 0.011898 0.00012537 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6804 0.6325 0.19263 0.021558 21.3978 0.13325 0.00017581 0.75692 0.009854 0.010879 0.0014019 0.98674 0.99157 3.025e-006 1.21e-005 0.16832 0.87528 0.89185 0.0014055 0.97298 0.43342 0.001893 0.42107 2.1322 2.131 16.027 144.8908 0.00020036 -85.5848 0.56294
9.667 0.98816 5.4548e-005 3.8183 0.011898 0.00012538 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6805 0.63255 0.19264 0.021559 21.4013 0.13326 0.00017582 0.75692 0.0098543 0.01088 0.0014018 0.98674 0.99157 3.0246e-006 1.2098e-005 0.16832 0.87562 0.89201 0.0014054 0.97313 0.43361 0.0018929 0.42108 2.133 2.1319 16.027 144.8908 0.00020012 -85.5854 0.56394
9.668 0.98816 5.4548e-005 3.8183 0.011898 0.0001254 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6806 0.63259 0.19265 0.02156 21.4048 0.13327 0.00017583 0.75691 0.0098546 0.01088 0.0014016 0.98675 0.99158 3.0243e-006 1.2097e-005 0.16832 0.87596 0.89216 0.0014053 0.97329 0.43381 0.0018928 0.4211 2.1339 2.1327 16.027 144.8908 0.00019989 -85.586 0.56494
9.669 0.98816 5.4548e-005 3.8183 0.011898 0.00012541 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6807 0.63263 0.19266 0.021561 21.4083 0.13327 0.00017584 0.75691 0.0098549 0.01088 0.0014015 0.98675 0.99158 3.024e-006 1.2096e-005 0.16832 0.87629 0.89231 0.0014052 0.97344 0.43401 0.0018927 0.42111 2.1347 2.1336 16.0269 144.8908 0.00019965 -85.5865 0.56594
9.67 0.98816 5.4548e-005 3.8183 0.011898 0.00012542 0.0011807 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6807 0.63268 0.19268 0.021562 21.4118 0.13328 0.00017585 0.7569 0.0098552 0.01088 0.0014014 0.98675 0.99158 3.0237e-006 1.2095e-005 0.16832 0.87663 0.89247 0.0014051 0.9736 0.43421 0.0018926 0.42113 2.1355 2.1344 16.0269 144.8908 0.00019942 -85.5871 0.56694
9.671 0.98816 5.4548e-005 3.8183 0.011898 0.00012543 0.0011808 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6808 0.63272 0.19269 0.021563 21.4153 0.13328 0.00017586 0.75689 0.0098555 0.010881 0.0014012 0.98675 0.99158 3.0234e-006 1.2093e-005 0.16833 0.87696 0.89262 0.001405 0.97375 0.4344 0.0018925 0.42114 2.1364 2.1352 16.0269 144.8909 0.00019918 -85.5877 0.56794
9.672 0.98816 5.4548e-005 3.8183 0.011898 0.00012545 0.0011808 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6809 0.63276 0.1927 0.021564 21.4187 0.13329 0.00017587 0.75689 0.0098558 0.010881 0.0014011 0.98675 0.99158 3.023e-006 1.2092e-005 0.16833 0.87729 0.89277 0.0014049 0.9739 0.4346 0.0018924 0.42116 2.1372 2.1361 16.0269 144.8909 0.00019895 -85.5882 0.56894
9.673 0.98816 5.4548e-005 3.8183 0.011898 0.00012546 0.0011808 0.23343 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.681 0.63281 0.19271 0.021565 21.4222 0.13329 0.00017588 0.75688 0.0098561 0.010881 0.001401 0.98675 0.99158 3.0227e-006 1.2091e-005 0.16833 0.87762 0.89292 0.0014048 0.97405 0.4348 0.0018923 0.42117 2.138 2.1369 16.0269 144.8909 0.00019872 -85.5888 0.56994
9.674 0.98816 5.4548e-005 3.8183 0.011898 0.00012547 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6811 0.63285 0.19273 0.021566 21.4257 0.1333 0.00017588 0.75688 0.0098564 0.010882 0.0014008 0.98676 0.99158 3.0224e-006 1.209e-005 0.16833 0.87796 0.89307 0.0014047 0.9742 0.43499 0.0018923 0.42119 2.1388 2.1377 16.0269 144.8909 0.00019849 -85.5893 0.57094
9.675 0.98816 5.4547e-005 3.8183 0.011898 0.00012548 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6811 0.6329 0.19274 0.021567 21.4292 0.1333 0.00017589 0.75687 0.0098567 0.010882 0.0014007 0.98676 0.99158 3.0221e-006 1.2089e-005 0.16834 0.87829 0.89322 0.0014046 0.97435 0.43519 0.0018922 0.42121 2.1397 2.1385 16.0268 144.891 0.00019826 -85.5899 0.57194
9.676 0.98816 5.4547e-005 3.8183 0.011898 0.0001255 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6812 0.63294 0.19275 0.021568 21.4327 0.13331 0.0001759 0.75687 0.009857 0.010882 0.0014006 0.98676 0.99158 3.0218e-006 1.2087e-005 0.16834 0.87861 0.89337 0.0014045 0.9745 0.43539 0.0018921 0.42122 2.1405 2.1394 16.0268 144.891 0.00019803 -85.5904 0.57294
9.677 0.98816 5.4547e-005 3.8183 0.011898 0.00012551 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6813 0.63298 0.19276 0.021568 21.4362 0.13332 0.00017591 0.75686 0.0098573 0.010883 0.0014005 0.98676 0.99159 3.0216e-006 1.2086e-005 0.16834 0.87894 0.89352 0.0014045 0.97464 0.43558 0.001892 0.42124 2.1413 2.1402 16.0268 144.891 0.0001978 -85.591 0.57394
9.678 0.98816 5.4547e-005 3.8183 0.011898 0.00012552 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6814 0.63303 0.19278 0.021569 21.4397 0.13332 0.00017592 0.75686 0.0098576 0.010883 0.0014003 0.98676 0.99159 3.0213e-006 1.2085e-005 0.16834 0.87927 0.89366 0.0014044 0.97479 0.43578 0.0018919 0.42125 2.1421 2.141 16.0268 144.891 0.00019758 -85.5915 0.57494
9.679 0.98816 5.4547e-005 3.8183 0.011898 0.00012554 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6815 0.63307 0.19279 0.02157 21.4432 0.13333 0.00017593 0.75685 0.0098579 0.010883 0.0014002 0.98676 0.99159 3.021e-006 1.2084e-005 0.16835 0.87959 0.89381 0.0014043 0.97493 0.43597 0.0018918 0.42127 2.1429 2.1418 16.0268 144.891 0.00019735 -85.592 0.57594
9.68 0.98816 5.4547e-005 3.8183 0.011898 0.00012555 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6815 0.63311 0.1928 0.021571 21.4467 0.13333 0.00017594 0.75684 0.0098582 0.010884 0.0014001 0.98677 0.99159 3.0207e-006 1.2083e-005 0.16835 0.87992 0.89396 0.0014043 0.97508 0.43617 0.0018917 0.42128 2.1437 2.1426 16.0268 144.8911 0.00019713 -85.5926 0.57694
9.681 0.98816 5.4547e-005 3.8183 0.011898 0.00012556 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6816 0.63316 0.19281 0.021572 21.4501 0.13334 0.00017594 0.75684 0.0098586 0.010884 0.0014 0.98677 0.99159 3.0205e-006 1.2082e-005 0.16835 0.88024 0.8941 0.0014043 0.97522 0.43637 0.0018917 0.4213 2.1445 2.1434 16.0267 144.8911 0.0001969 -85.5931 0.57794
9.682 0.98816 5.4547e-005 3.8183 0.011898 0.00012557 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6817 0.6332 0.19283 0.021573 21.4536 0.13334 0.00017595 0.75683 0.0098589 0.010884 0.0013998 0.98677 0.99159 3.0202e-006 1.2081e-005 0.16835 0.88057 0.89425 0.0014042 0.97536 0.43656 0.0018916 0.42131 2.1453 2.1442 16.0267 144.8911 0.00019668 -85.5936 0.57894
9.683 0.98816 5.4547e-005 3.8183 0.011898 0.00012559 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6818 0.63325 0.19284 0.021574 21.4571 0.13335 0.00017596 0.75683 0.0098592 0.010885 0.0013997 0.98677 0.99159 3.0199e-006 1.208e-005 0.16835 0.88089 0.89439 0.0014042 0.9755 0.43676 0.0018915 0.42133 2.1461 2.145 16.0267 144.8911 0.00019646 -85.5941 0.57994
9.684 0.98816 5.4547e-005 3.8183 0.011898 0.0001256 0.0011808 0.23342 0.00065931 0.23408 0.216 0 0.032273 0.0389 0 1.6819 0.63329 0.19285 0.021575 21.4606 0.13335 0.00017597 0.75682 0.0098595 0.010885 0.0013996 0.98677 0.99159 3.0196e-006 1.2078e-005 0.16836 0.88121 0.89454 0.0014041 0.97564 0.43695 0.0018914 0.42134 2.1469 2.1458 16.0267 144.8911 0.00019624 -85.5946 0.58094
9.685 0.98816 5.4547e-005 3.8183 0.011898 0.00012561 0.0011808 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.6819 0.63333 0.19286 0.021576 21.4641 0.13336 0.00017598 0.75682 0.0098598 0.010885 0.0013995 0.98677 0.99159 3.0194e-006 1.2077e-005 0.16836 0.88153 0.89468 0.0014041 0.97578 0.43715 0.0018913 0.42136 2.1477 2.1467 16.0267 144.8912 0.00019601 -85.5951 0.58194
9.686 0.98816 5.4547e-005 3.8183 0.011898 0.00012563 0.0011808 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.682 0.63338 0.19288 0.021577 21.4676 0.13337 0.00017599 0.75681 0.0098601 0.010886 0.0013994 0.98677 0.99159 3.0191e-006 1.2076e-005 0.16836 0.88185 0.89482 0.001404 0.97592 0.43735 0.0018912 0.42138 2.1485 2.1475 16.0267 144.8912 0.00019579 -85.5957 0.58294
9.687 0.98816 5.4546e-005 3.8183 0.011898 0.00012564 0.0011808 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.6821 0.63342 0.19289 0.021578 21.4711 0.13337 0.000176 0.75681 0.0098604 0.010886 0.0013992 0.98678 0.9916 3.0188e-006 1.2075e-005 0.16836 0.88216 0.89497 0.001404 0.97606 0.43754 0.0018912 0.42139 2.1493 2.1482 16.0266 144.8912 0.00019558 -85.5962 0.58394
9.688 0.98816 5.4546e-005 3.8183 0.011897 0.00012565 0.0011808 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.6822 0.63346 0.1929 0.021579 21.4746 0.13338 0.000176 0.7568 0.0098607 0.010886 0.0013991 0.98678 0.9916 3.0186e-006 1.2074e-005 0.16837 0.88248 0.89511 0.0014039 0.9762 0.43774 0.0018911 0.42141 2.1501 2.149 16.0266 144.8912 0.00019536 -85.5967 0.58494
9.689 0.98816 5.4546e-005 3.8183 0.011897 0.00012566 0.0011809 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.6823 0.63351 0.19291 0.02158 21.4781 0.13338 0.00017601 0.75679 0.009861 0.010887 0.001399 0.98678 0.9916 3.0183e-006 1.2073e-005 0.16837 0.8828 0.89525 0.0014038 0.97633 0.43793 0.001891 0.42142 2.1509 2.1498 16.0266 144.8912 0.00019514 -85.5971 0.58594
9.69 0.98816 5.4546e-005 3.8183 0.011897 0.00012568 0.0011809 0.23342 0.00065931 0.23408 0.21599 0 0.032273 0.0389 0 1.6824 0.63355 0.19293 0.021581 21.4816 0.13339 0.00017602 0.75679 0.0098613 0.010887 0.0013989 0.98678 0.9916 3.018e-006 1.2072e-005 0.16837 0.88311 0.89539 0.0014038 0.97647 0.43813 0.0018909 0.42144 2.1517 2.1506 16.0266 144.8913 0.00019492 -85.5976 0.58694
9.691 0.98816 5.4546e-005 3.8183 0.011897 0.00012569 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6824 0.63359 0.19294 0.021582 21.4851 0.13339 0.00017603 0.75678 0.0098616 0.010887 0.0013988 0.98678 0.9916 3.0178e-006 1.2071e-005 0.16837 0.88342 0.89553 0.0014037 0.9766 0.43832 0.0018908 0.42145 2.1525 2.1514 16.0266 144.8913 0.00019471 -85.5981 0.58794
9.692 0.98816 5.4546e-005 3.8183 0.011897 0.0001257 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6825 0.63364 0.19295 0.021583 21.4886 0.1334 0.00017604 0.75678 0.0098619 0.010888 0.0013987 0.98678 0.9916 3.0175e-006 1.207e-005 0.16838 0.88374 0.89567 0.0014036 0.97673 0.43852 0.0018908 0.42147 2.1533 2.1522 16.0265 144.8913 0.00019449 -85.5986 0.58894
9.693 0.98816 5.4546e-005 3.8183 0.011897 0.00012571 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6826 0.63368 0.19296 0.021584 21.4921 0.1334 0.00017605 0.75677 0.0098622 0.010888 0.0013986 0.98679 0.9916 3.0172e-006 1.2069e-005 0.16838 0.88405 0.89581 0.0014036 0.97687 0.43872 0.0018907 0.42148 2.1541 2.153 16.0265 144.8913 0.00019428 -85.5991 0.58994
9.694 0.98816 5.4546e-005 3.8183 0.011897 0.00012573 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6827 0.63373 0.19298 0.021584 21.4955 0.13341 0.00017606 0.75677 0.0098625 0.010888 0.0013984 0.98679 0.9916 3.017e-006 1.2068e-005 0.16838 0.88436 0.89595 0.0014035 0.977 0.43891 0.0018906 0.4215 2.1548 2.1538 16.0265 144.8913 0.00019407 -85.5996 0.59094
9.695 0.98816 5.4546e-005 3.8183 0.011897 0.00012574 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6828 0.63377 0.19299 0.021585 21.499 0.13342 0.00017606 0.75676 0.0098628 0.010889 0.0013983 0.98679 0.9916 3.0167e-006 1.2067e-005 0.16838 0.88467 0.89609 0.0014034 0.97713 0.43911 0.0018905 0.42152 2.1556 2.1546 16.0265 144.8914 0.00019386 -85.6 0.59194
9.696 0.98816 5.4546e-005 3.8183 0.011897 0.00012575 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6828 0.63381 0.193 0.021586 21.5025 0.13342 0.00017607 0.75676 0.0098631 0.010889 0.0013982 0.98679 0.9916 3.0165e-006 1.2066e-005 0.16839 0.88498 0.89623 0.0014034 0.97726 0.4393 0.0018905 0.42153 2.1564 2.1553 16.0265 144.8914 0.00019364 -85.6005 0.59294
9.697 0.98816 5.4546e-005 3.8183 0.011897 0.00012577 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6829 0.63386 0.19301 0.021587 21.506 0.13343 0.00017608 0.75675 0.0098634 0.010889 0.0013981 0.98679 0.9916 3.0162e-006 1.2065e-005 0.16839 0.88529 0.89636 0.0014033 0.97739 0.4395 0.0018904 0.42155 2.1572 2.1561 16.0265 144.8914 0.00019343 -85.601 0.59394
9.698 0.98816 5.4546e-005 3.8183 0.011897 0.00012578 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.683 0.6339 0.19303 0.021588 21.5095 0.13343 0.00017609 0.75674 0.0098637 0.010889 0.001398 0.98679 0.99161 3.016e-006 1.2064e-005 0.16839 0.88559 0.8965 0.0014032 0.97752 0.43969 0.0018903 0.42156 2.1579 2.1569 16.0264 144.8914 0.00019322 -85.6014 0.59494
9.699 0.98816 5.4545e-005 3.8183 0.011897 0.00012579 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6831 0.63394 0.19304 0.021589 21.513 0.13344 0.0001761 0.75674 0.009864 0.01089 0.0013979 0.98679 0.99161 3.0157e-006 1.2063e-005 0.16839 0.8859 0.89664 0.0014032 0.97764 0.43989 0.0018902 0.42158 2.1587 2.1577 16.0264 144.8914 0.00019302 -85.6019 0.59594
9.7 0.98816 5.4545e-005 3.8183 0.011897 0.0001258 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6832 0.63399 0.19305 0.02159 21.5165 0.13344 0.00017611 0.75673 0.0098643 0.01089 0.0013978 0.9868 0.99161 3.0155e-006 1.2062e-005 0.16839 0.8862 0.89677 0.0014031 0.97777 0.44008 0.0018902 0.42159 2.1595 2.1584 16.0264 144.8915 0.00019281 -85.6024 0.59694
9.701 0.98816 5.4545e-005 3.8183 0.011897 0.00012582 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6832 0.63403 0.19306 0.021591 21.52 0.13345 0.00017612 0.75673 0.0098647 0.01089 0.0013977 0.9868 0.99161 3.0153e-006 1.2061e-005 0.1684 0.88651 0.89691 0.0014031 0.9779 0.44028 0.0018901 0.42161 2.1603 2.1592 16.0264 144.8915 0.0001926 -85.6028 0.59794
9.702 0.98816 5.4545e-005 3.8183 0.011897 0.00012583 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6833 0.63408 0.19308 0.021592 21.5235 0.13345 0.00017613 0.75672 0.009865 0.010891 0.0013976 0.9868 0.99161 3.015e-006 1.206e-005 0.1684 0.88681 0.89704 0.001403 0.97802 0.44047 0.00189 0.42162 2.161 2.16 16.0264 144.8915 0.00019239 -85.6033 0.59894
9.703 0.98816 5.4545e-005 3.8183 0.011897 0.00012584 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6834 0.63412 0.19309 0.021593 21.527 0.13346 0.00017613 0.75672 0.0098653 0.010891 0.0013975 0.9868 0.99161 3.0148e-006 1.2059e-005 0.1684 0.88711 0.89717 0.001403 0.97814 0.44067 0.0018899 0.42164 2.1618 2.1607 16.0263 144.8915 0.00019219 -85.6037 0.59994
9.704 0.98816 5.4545e-005 3.8183 0.011897 0.00012585 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6835 0.63416 0.1931 0.021594 21.5305 0.13346 0.00017614 0.75671 0.0098656 0.010891 0.0013974 0.9868 0.99161 3.0145e-006 1.2058e-005 0.1684 0.88741 0.89731 0.0014029 0.97827 0.44086 0.0018899 0.42165 2.1625 2.1615 16.0263 144.8915 0.00019198 -85.6042 0.60094
9.705 0.98816 5.4545e-005 3.8183 0.011897 0.00012587 0.0011809 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6836 0.63421 0.19311 0.021595 21.534 0.13347 0.00017615 0.75671 0.0098659 0.010892 0.0013973 0.9868 0.99161 3.0143e-006 1.2057e-005 0.16841 0.88771 0.89744 0.0014029 0.97839 0.44106 0.0018898 0.42167 2.1633 2.1623 16.0263 144.8916 0.00019178 -85.6046 0.60194
9.706 0.98816 5.4545e-005 3.8183 0.011897 0.00012588 0.001181 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6836 0.63425 0.19313 0.021596 21.5375 0.13348 0.00017616 0.7567 0.0098662 0.010892 0.0013972 0.9868 0.99161 3.0141e-006 1.2056e-005 0.16841 0.88801 0.89757 0.0014028 0.97851 0.44125 0.0018897 0.42169 2.1641 2.163 16.0263 144.8916 0.00019158 -85.605 0.60294
9.707 0.98816 5.4545e-005 3.8183 0.011897 0.00012589 0.001181 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6837 0.63429 0.19314 0.021597 21.541 0.13348 0.00017617 0.75669 0.0098665 0.010892 0.0013971 0.9868 0.99161 3.0138e-006 1.2055e-005 0.16841 0.88831 0.89771 0.0014028 0.97863 0.44144 0.0018897 0.4217 2.1648 2.1638 16.0263 144.8916 0.00019137 -85.6055 0.60394
9.708 0.98816 5.4545e-005 3.8183 0.011897 0.00012591 0.001181 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6838 0.63434 0.19315 0.021598 21.5445 0.13349 0.00017618 0.75669 0.0098668 0.010893 0.001397 0.98681 0.99161 3.0136e-006 1.2054e-005 0.16841 0.88861 0.89784 0.0014027 0.97875 0.44164 0.0018896 0.42172 2.1656 2.1645 16.0262 144.8916 0.00019117 -85.6059 0.60494
9.709 0.98816 5.4545e-005 3.8183 0.011897 0.00012592 0.001181 0.23342 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6839 0.63438 0.19316 0.021599 21.548 0.13349 0.00017619 0.75668 0.0098671 0.010893 0.0013969 0.98681 0.99162 3.0134e-006 1.2053e-005 0.16842 0.88891 0.89797 0.0014027 0.97887 0.44183 0.0018895 0.42173 2.1663 2.1653 16.0262 144.8916 0.00019097 -85.6063 0.60594
9.71 0.98816 5.4544e-005 3.8183 0.011897 0.00012593 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.684 0.63443 0.19318 0.021599 21.5515 0.1335 0.00017619 0.75668 0.0098674 0.010893 0.0013968 0.98681 0.99162 3.0132e-006 1.2053e-005 0.16842 0.8892 0.8981 0.0014026 0.97899 0.44203 0.0018895 0.42175 2.1671 2.1661 16.0262 144.8917 0.00019077 -85.6067 0.60694
9.711 0.98816 5.4544e-005 3.8183 0.011897 0.00012594 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6841 0.63447 0.19319 0.0216 21.555 0.1335 0.0001762 0.75667 0.0098677 0.010894 0.0013967 0.98681 0.99162 3.0129e-006 1.2052e-005 0.16842 0.8895 0.89823 0.0014026 0.97911 0.44222 0.0018894 0.42176 2.1678 2.1668 16.0262 144.8917 0.00019057 -85.6072 0.60794
9.712 0.98816 5.4544e-005 3.8183 0.011897 0.00012596 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6841 0.63451 0.1932 0.021601 21.5585 0.13351 0.00017621 0.75667 0.009868 0.010894 0.0013966 0.98681 0.99162 3.0127e-006 1.2051e-005 0.16842 0.88979 0.89836 0.0014025 0.97923 0.44242 0.0018893 0.42178 2.1686 2.1676 16.0262 144.8917 0.00019037 -85.6076 0.60894
9.713 0.98816 5.4544e-005 3.8183 0.011897 0.00012597 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6842 0.63456 0.19321 0.021602 21.562 0.13351 0.00017622 0.75666 0.0098683 0.010894 0.0013965 0.98681 0.99162 3.0125e-006 1.205e-005 0.16842 0.89008 0.89849 0.0014024 0.97934 0.44261 0.0018893 0.42179 2.1693 2.1683 16.0261 144.8917 0.00019018 -85.608 0.60994
9.714 0.98816 5.4544e-005 3.8183 0.011897 0.00012598 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6843 0.6346 0.19323 0.021603 21.5655 0.13352 0.00017623 0.75666 0.0098686 0.010895 0.0013964 0.98681 0.99162 3.0123e-006 1.2049e-005 0.16843 0.89037 0.89862 0.0014024 0.97946 0.4428 0.0018892 0.42181 2.17 2.169 16.0261 144.8917 0.00018998 -85.6084 0.61094
9.715 0.98816 5.4544e-005 3.8183 0.011897 0.00012599 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6844 0.63464 0.19324 0.021604 21.569 0.13353 0.00017624 0.75665 0.0098689 0.010895 0.0013963 0.98681 0.99162 3.0121e-006 1.2048e-005 0.16843 0.89067 0.89874 0.0014023 0.97957 0.443 0.0018891 0.42182 2.1708 2.1698 16.0261 144.8918 0.00018978 -85.6088 0.61194
9.716 0.98816 5.4544e-005 3.8183 0.011897 0.00012601 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6845 0.63469 0.19325 0.021605 21.5725 0.13353 0.00017625 0.75664 0.0098692 0.010895 0.0013962 0.98682 0.99162 3.0118e-006 1.2047e-005 0.16843 0.89096 0.89887 0.0014023 0.97969 0.44319 0.0018891 0.42184 2.1715 2.1705 16.0261 144.8918 0.00018959 -85.6092 0.61294
9.717 0.98816 5.4544e-005 3.8183 0.011897 0.00012602 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6845 0.63473 0.19326 0.021606 21.576 0.13354 0.00017625 0.75664 0.0098695 0.010896 0.0013961 0.98682 0.99162 3.0116e-006 1.2046e-005 0.16843 0.89124 0.899 0.0014022 0.9798 0.44339 0.001889 0.42186 2.1723 2.1713 16.0261 144.8918 0.00018939 -85.6096 0.61394
9.718 0.98816 5.4544e-005 3.8183 0.011897 0.00012603 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6846 0.63478 0.19328 0.021607 21.5795 0.13354 0.00017626 0.75663 0.0098698 0.010896 0.001396 0.98682 0.99162 3.0114e-006 1.2046e-005 0.16844 0.89153 0.89912 0.0014022 0.97991 0.44358 0.0018889 0.42187 2.173 2.172 16.026 144.8918 0.0001892 -85.61 0.61494
9.719 0.98816 5.4544e-005 3.8183 0.011897 0.00012605 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6847 0.63482 0.19329 0.021608 21.583 0.13355 0.00017627 0.75663 0.0098701 0.010896 0.0013959 0.98682 0.99162 3.0112e-006 1.2045e-005 0.16844 0.89182 0.89925 0.0014022 0.98002 0.44377 0.0018889 0.42189 2.1737 2.1727 16.026 144.8918 0.00018901 -85.6104 0.61594
9.72 0.98816 5.4544e-005 3.8183 0.011897 0.00012606 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6848 0.63486 0.1933 0.021609 21.5865 0.13355 0.00017628 0.75662 0.0098704 0.010897 0.0013958 0.98682 0.99162 3.011e-006 1.2044e-005 0.16844 0.89211 0.89938 0.0014021 0.98014 0.44397 0.0018888 0.4219 2.1745 2.1735 16.026 144.8919 0.00018881 -85.6108 0.61694
9.721 0.98816 5.4544e-005 3.8183 0.011897 0.00012607 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032273 0.0389 0 1.6849 0.63491 0.19331 0.02161 21.59 0.13356 0.00017629 0.75662 0.0098707 0.010897 0.0013957 0.98682 0.99163 3.0108e-006 1.2043e-005 0.16844 0.89239 0.8995 0.0014021 0.98025 0.44416 0.0018887 0.42192 2.1752 2.1742 16.026 144.8919 0.00018862 -85.6112 0.61794
9.722 0.98816 5.4543e-005 3.8183 0.011897 0.00012608 0.001181 0.23341 0.00065931 0.23407 0.21599 0 0.032274 0.0389 0 1.6849 0.63495 0.19333 0.021611 21.5935 0.13356 0.0001763 0.75661 0.009871 0.010897 0.0013956 0.98682 0.99163 3.0106e-006 1.2042e-005 0.16845 0.89268 0.89963 0.001402 0.98036 0.44435 0.0018887 0.42193 2.1759 2.1749 16.026 144.8919 0.00018843 -85.6116 0.61894
9.723 0.98816 5.4543e-005 3.8183 0.011897 0.0001261 0.001181 0.23341 0.00065931 0.23407 0.21598 0 0.032274 0.0389 0 1.685 0.63499 0.19334 0.021612 21.597 0.13357 0.00017631 0.75661 0.0098713 0.010897 0.0013955 0.98682 0.99163 3.0104e-006 1.2041e-005 0.16845 0.89296 0.89975 0.001402 0.98046 0.44455 0.0018886 0.42195 2.1766 2.1757 16.0259 144.8919 0.00018824 -85.612 0.61994
9.724 0.98816 5.4543e-005 3.8183 0.011897 0.00012611 0.0011811 0.23341 0.00065931 0.23407 0.21598 0 0.032274 0.0389 0 1.6851 0.63504 0.19335 0.021613 21.6005 0.13358 0.00017631 0.7566 0.0098716 0.010898 0.0013955 0.98683 0.99163 3.0102e-006 1.2041e-005 0.16845 0.89324 0.89987 0.0014019 0.98057 0.44474 0.0018886 0.42196 2.1774 2.1764 16.0259 144.8919 0.00018805 -85.6124 0.62094
9.725 0.98816 5.4543e-005 3.8183 0.011897 0.00012612 0.0011811 0.23341 0.00065931 0.23407 0.21598 0 0.032274 0.0389 0 1.6852 0.63508 0.19336 0.021614 21.604 0.13358 0.00017632 0.7566 0.009872 0.010898 0.0013954 0.98683 0.99163 3.01e-006 1.204e-005 0.16845 0.89353 0.9 0.0014019 0.98068 0.44493 0.0018885 0.42198 2.1781 2.1771 16.0259 144.892 0.00018786 -85.6128 0.62194
9.726 0.98816 5.4543e-005 3.8183 0.011897 0.00012613 0.0011811 0.23341 0.00065931 0.23407 0.21598 0 0.032274 0.0389 0 1.6853 0.63512 0.19338 0.021615 21.6075 0.13359 0.00017633 0.75659 0.0098723 0.010898 0.0013953 0.98683 0.99163 3.0098e-006 1.2039e-005 0.16845 0.89381 0.90012 0.0014018 0.98079 0.44513 0.0018884 0.42199 2.1788 2.1778 16.0259 144.892 0.00018767 -85.6131 0.62294
9.727 0.98816 5.4543e-005 3.8183 0.011897 0.00012615 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6853 0.63517 0.19339 0.021615 21.611 0.13359 0.00017634 0.75658 0.0098726 0.010899 0.0013952 0.98683 0.99163 3.0096e-006 1.2038e-005 0.16846 0.89409 0.90024 0.0014018 0.98089 0.44532 0.0018884 0.42201 2.1795 2.1786 16.0259 144.892 0.00018749 -85.6135 0.62394
9.728 0.98816 5.4543e-005 3.8183 0.011897 0.00012616 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6854 0.63521 0.1934 0.021616 21.6145 0.1336 0.00017635 0.75658 0.0098729 0.010899 0.0013951 0.98683 0.99163 3.0094e-006 1.2037e-005 0.16846 0.89437 0.90036 0.0014017 0.981 0.44551 0.0018883 0.42202 2.1802 2.1793 16.0258 144.892 0.0001873 -85.6139 0.62494
9.729 0.98816 5.4543e-005 3.8183 0.011897 0.00012617 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6855 0.63526 0.19341 0.021617 21.618 0.1336 0.00017636 0.75657 0.0098732 0.010899 0.001395 0.98683 0.99163 3.0092e-006 1.2037e-005 0.16846 0.89465 0.90048 0.0014017 0.9811 0.44571 0.0018883 0.42204 2.181 2.18 16.0258 144.892 0.00018711 -85.6142 0.62594
9.73 0.98816 5.4543e-005 3.8183 0.011897 0.00012619 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6856 0.6353 0.19343 0.021618 21.6215 0.13361 0.00017637 0.75657 0.0098735 0.0109 0.0013949 0.98683 0.99163 3.009e-006 1.2036e-005 0.16846 0.89492 0.90061 0.0014017 0.98121 0.4459 0.0018882 0.42206 2.1817 2.1807 16.0258 144.8921 0.00018693 -85.6146 0.62694
9.731 0.98816 5.4543e-005 3.8183 0.011897 0.0001262 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6857 0.63534 0.19344 0.021619 21.625 0.13361 0.00017637 0.75656 0.0098738 0.0109 0.0013948 0.98683 0.99163 3.0088e-006 1.2035e-005 0.16847 0.8952 0.90073 0.0014016 0.98131 0.44609 0.0018881 0.42207 2.1824 2.1814 16.0258 144.8921 0.00018675 -85.615 0.62794
9.732 0.98816 5.4543e-005 3.8183 0.011897 0.00012621 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6858 0.63539 0.19345 0.02162 21.6286 0.13362 0.00017638 0.75656 0.0098741 0.0109 0.0013948 0.98683 0.99163 3.0086e-006 1.2034e-005 0.16847 0.89548 0.90085 0.0014016 0.98142 0.44629 0.0018881 0.42209 2.1831 2.1821 16.0258 144.8921 0.00018656 -85.6153 0.62894
9.733 0.98816 5.4543e-005 3.8183 0.011897 0.00012622 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6858 0.63543 0.19346 0.021621 21.6321 0.13363 0.00017639 0.75655 0.0098744 0.010901 0.0013947 0.98684 0.99163 3.0084e-006 1.2033e-005 0.16847 0.89575 0.90097 0.0014015 0.98152 0.44648 0.001888 0.4221 2.1838 2.1828 16.0257 144.8921 0.00018638 -85.6157 0.62994
9.734 0.98816 5.4542e-005 3.8183 0.011897 0.00012624 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6859 0.63547 0.19348 0.021622 21.6356 0.13363 0.0001764 0.75655 0.0098747 0.010901 0.0013946 0.98684 0.99163 3.0082e-006 1.2033e-005 0.16847 0.89603 0.90108 0.0014015 0.98162 0.44667 0.001888 0.42212 2.1845 2.1835 16.0257 144.8921 0.0001862 -85.6161 0.63094
9.735 0.98816 5.4542e-005 3.8183 0.011897 0.00012625 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.686 0.63552 0.19349 0.021623 21.6391 0.13364 0.00017641 0.75654 0.009875 0.010901 0.0013945 0.98684 0.99164 3.008e-006 1.2032e-005 0.16848 0.8963 0.9012 0.0014015 0.98172 0.44686 0.0018879 0.42213 2.1852 2.1843 16.0257 144.8922 0.00018601 -85.6164 0.63194
9.736 0.98816 5.4542e-005 3.8183 0.011897 0.00012626 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6861 0.63556 0.1935 0.021624 21.6426 0.13364 0.00017642 0.75653 0.0098753 0.010902 0.0013944 0.98684 0.99164 3.0078e-006 1.2031e-005 0.16848 0.89657 0.90132 0.0014014 0.98182 0.44706 0.0018878 0.42215 2.1859 2.185 16.0257 144.8922 0.00018583 -85.6168 0.63294
9.737 0.98816 5.4542e-005 3.8183 0.011897 0.00012627 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6862 0.63561 0.19351 0.021625 21.6461 0.13365 0.00017643 0.75653 0.0098756 0.010902 0.0013944 0.98684 0.99164 3.0076e-006 1.203e-005 0.16848 0.89684 0.90144 0.0014014 0.98192 0.44725 0.0018878 0.42216 2.1866 2.1857 16.0256 144.8922 0.00018565 -85.6171 0.63394
9.738 0.98816 5.4542e-005 3.8183 0.011897 0.00012629 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6862 0.63565 0.19353 0.021626 21.6496 0.13365 0.00017643 0.75652 0.0098759 0.010902 0.0013943 0.98684 0.99164 3.0075e-006 1.203e-005 0.16848 0.89711 0.90156 0.0014013 0.98202 0.44744 0.0018877 0.42218 2.1873 2.1864 16.0256 144.8922 0.00018547 -85.6174 0.63494
9.739 0.98816 5.4542e-005 3.8183 0.011897 0.0001263 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6863 0.63569 0.19354 0.021627 21.6531 0.13366 0.00017644 0.75652 0.0098762 0.010903 0.0013942 0.98684 0.99164 3.0073e-006 1.2029e-005 0.16848 0.89738 0.90167 0.0014013 0.98212 0.44763 0.0018877 0.42219 2.188 2.1871 16.0256 144.8922 0.0001853 -85.6178 0.63594
9.74 0.98816 5.4542e-005 3.8183 0.011897 0.00012631 0.0011811 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6864 0.63574 0.19355 0.021628 21.6566 0.13366 0.00017645 0.75651 0.0098765 0.010903 0.0013941 0.98684 0.99164 3.0071e-006 1.2028e-005 0.16849 0.89765 0.90179 0.0014012 0.98221 0.44783 0.0018876 0.42221 2.1887 2.1878 16.0256 144.8923 0.00018512 -85.6181 0.63694
9.741 0.98816 5.4542e-005 3.8183 0.011897 0.00012633 0.0011812 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6865 0.63578 0.19356 0.021629 21.6601 0.13367 0.00017646 0.75651 0.0098768 0.010903 0.001394 0.98684 0.99164 3.0069e-006 1.2028e-005 0.16849 0.89792 0.9019 0.0014012 0.98231 0.44802 0.0018876 0.42222 2.1894 2.1885 16.0256 144.8923 0.00018494 -85.6185 0.63794
9.742 0.98816 5.4542e-005 3.8183 0.011897 0.00012634 0.0011812 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6866 0.63582 0.19358 0.021629 21.6636 0.13367 0.00017647 0.7565 0.0098771 0.010904 0.001394 0.98684 0.99164 3.0067e-006 1.2027e-005 0.16849 0.89819 0.90202 0.0014011 0.98241 0.44821 0.0018875 0.42224 2.1901 2.1892 16.0255 144.8923 0.00018476 -85.6188 0.63894
9.743 0.98816 5.4542e-005 3.8183 0.011896 0.00012635 0.0011812 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6866 0.63587 0.19359 0.02163 21.6671 0.13368 0.00017648 0.7565 0.0098774 0.010904 0.0013939 0.98685 0.99164 3.0066e-006 1.2026e-005 0.16849 0.89846 0.90214 0.0014011 0.9825 0.4484 0.0018875 0.42226 2.1908 2.1898 16.0255 144.8923 0.00018459 -85.6191 0.63994
9.744 0.98816 5.4542e-005 3.8183 0.011896 0.00012636 0.0011812 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6867 0.63591 0.1936 0.021631 21.6706 0.13369 0.00017649 0.75649 0.0098777 0.010904 0.0013938 0.98685 0.99164 3.0064e-006 1.2025e-005 0.1685 0.89872 0.90225 0.0014011 0.9826 0.44859 0.0018874 0.42227 2.1915 2.1905 16.0255 144.8923 0.00018441 -85.6195 0.64094
9.745 0.98816 5.4541e-005 3.8183 0.011896 0.00012638 0.0011812 0.23341 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6868 0.63595 0.19361 0.021632 21.6742 0.13369 0.00017649 0.75648 0.009878 0.010904 0.0013937 0.98685 0.99164 3.0062e-006 1.2025e-005 0.1685 0.89899 0.90236 0.001401 0.98269 0.44879 0.0018874 0.42229 2.1921 2.1912 16.0255 144.8924 0.00018424 -85.6198 0.64194
9.746 0.98816 5.4541e-005 3.8183 0.011896 0.00012639 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6869 0.636 0.19362 0.021633 21.6777 0.1337 0.0001765 0.75648 0.0098783 0.010905 0.0013937 0.98685 0.99164 3.006e-006 1.2024e-005 0.1685 0.89925 0.90248 0.001401 0.98279 0.44898 0.0018873 0.4223 2.1928 2.1919 16.0254 144.8924 0.00018406 -85.6201 0.64294
9.747 0.98816 5.4541e-005 3.8183 0.011896 0.0001264 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.687 0.63604 0.19364 0.021634 21.6812 0.1337 0.00017651 0.75647 0.0098786 0.010905 0.0013936 0.98685 0.99164 3.0059e-006 1.2023e-005 0.1685 0.89951 0.90259 0.0014009 0.98288 0.44917 0.0018873 0.42232 2.1935 2.1926 16.0254 144.8924 0.00018389 -85.6204 0.64394
9.748 0.98816 5.4541e-005 3.8183 0.011896 0.00012642 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.687 0.63609 0.19365 0.021635 21.6847 0.13371 0.00017652 0.75647 0.0098789 0.010905 0.0013935 0.98685 0.99164 3.0057e-006 1.2023e-005 0.16851 0.89978 0.9027 0.0014009 0.98297 0.44936 0.0018872 0.42233 2.1942 2.1933 16.0254 144.8924 0.00018372 -85.6208 0.64494
9.749 0.98816 5.4541e-005 3.8183 0.011896 0.00012643 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6871 0.63613 0.19366 0.021636 21.6882 0.13371 0.00017653 0.75646 0.0098792 0.010906 0.0013934 0.98685 0.99164 3.0055e-006 1.2022e-005 0.16851 0.90004 0.90282 0.0014009 0.98307 0.44955 0.0018872 0.42235 2.1949 2.194 16.0254 144.8925 0.00018354 -85.6211 0.64594
9.75 0.98816 5.4541e-005 3.8183 0.011896 0.00012644 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6872 0.63617 0.19367 0.021637 21.6917 0.13372 0.00017654 0.75646 0.0098795 0.010906 0.0013934 0.98685 0.99165 3.0054e-006 1.2021e-005 0.16851 0.9003 0.90293 0.0014008 0.98316 0.44975 0.0018871 0.42236 2.1955 2.1946 16.0254 144.8925 0.00018337 -85.6214 0.64694
9.751 0.98816 5.4541e-005 3.8183 0.011896 0.00012645 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6873 0.63622 0.19369 0.021638 21.6952 0.13372 0.00017655 0.75645 0.0098798 0.010906 0.0013933 0.98685 0.99165 3.0052e-006 1.2021e-005 0.16851 0.90056 0.90304 0.0014008 0.98325 0.44994 0.0018871 0.42238 2.1962 2.1953 16.0253 144.8925 0.0001832 -85.6217 0.64794
9.752 0.98816 5.4541e-005 3.8183 0.011896 0.00012647 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6874 0.63626 0.1937 0.021639 21.6987 0.13373 0.00017655 0.75645 0.0098801 0.010907 0.0013932 0.98685 0.99165 3.005e-006 1.202e-005 0.16851 0.90082 0.90315 0.0014007 0.98334 0.45013 0.001887 0.42239 2.1969 2.196 16.0253 144.8925 0.00018303 -85.622 0.64894
9.753 0.98816 5.4541e-005 3.8183 0.011896 0.00012648 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6874 0.6363 0.19371 0.02164 21.7022 0.13374 0.00017656 0.75644 0.0098804 0.010907 0.0013931 0.98686 0.99165 3.0048e-006 1.2019e-005 0.16852 0.90108 0.90326 0.0014007 0.98343 0.45032 0.001887 0.42241 2.1976 2.1967 16.0253 144.8925 0.00018286 -85.6223 0.64994
9.754 0.98816 5.4541e-005 3.8183 0.011896 0.00012649 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6875 0.63635 0.19372 0.021641 21.7058 0.13374 0.00017657 0.75644 0.0098807 0.010907 0.0013931 0.98686 0.99165 3.0047e-006 1.2019e-005 0.16852 0.90133 0.90337 0.0014007 0.98352 0.45051 0.0018869 0.42242 2.1982 2.1973 16.0253 144.8926 0.00018269 -85.6226 0.65094
9.755 0.98816 5.4541e-005 3.8183 0.011896 0.0001265 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6876 0.63639 0.19374 0.021642 21.7093 0.13375 0.00017658 0.75643 0.009881 0.010908 0.001393 0.98686 0.99165 3.0045e-006 1.2018e-005 0.16852 0.90159 0.90348 0.0014006 0.98361 0.4507 0.0018869 0.42244 2.1989 2.198 16.0252 144.8926 0.00018253 -85.6229 0.65194
9.756 0.98816 5.4541e-005 3.8183 0.011896 0.00012652 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6877 0.63644 0.19375 0.021643 21.7128 0.13375 0.00017659 0.75642 0.0098813 0.010908 0.0013929 0.98686 0.99165 3.0044e-006 1.2017e-005 0.16852 0.90185 0.90359 0.0014006 0.98369 0.45089 0.0018868 0.42245 2.1996 2.1987 16.0252 144.8926 0.00018236 -85.6232 0.65294
9.757 0.98816 5.454e-005 3.8183 0.011896 0.00012653 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6878 0.63648 0.19376 0.021644 21.7163 0.13376 0.0001766 0.75642 0.0098816 0.010908 0.0013929 0.98686 0.99165 3.0042e-006 1.2017e-005 0.16853 0.9021 0.9037 0.0014006 0.98378 0.45109 0.0018868 0.42247 2.2002 2.1994 16.0252 144.8926 0.00018219 -85.6235 0.65394
9.758 0.98816 5.454e-005 3.8183 0.011896 0.00012654 0.0011812 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6879 0.63652 0.19377 0.021644 21.7198 0.13376 0.00017661 0.75641 0.0098819 0.010909 0.0013928 0.98686 0.99165 3.0041e-006 1.2016e-005 0.16853 0.90236 0.90381 0.0014005 0.98387 0.45128 0.0018867 0.42248 2.2009 2.2 16.0252 144.8926 0.00018202 -85.6238 0.65494
9.759 0.98816 5.454e-005 3.8183 0.011896 0.00012656 0.0011813 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.6879 0.63657 0.19379 0.021645 21.7233 0.13377 0.00017661 0.75641 0.0098822 0.010909 0.0013927 0.98686 0.99165 3.0039e-006 1.2016e-005 0.16853 0.90261 0.90392 0.0014005 0.98396 0.45147 0.0018867 0.4225 2.2016 2.2007 16.0251 144.8927 0.00018186 -85.6241 0.65594
9.76 0.98816 5.454e-005 3.8183 0.011896 0.00012657 0.0011813 0.2334 0.00065931 0.23406 0.21598 0 0.032274 0.0389 0 1.688 0.63661 0.1938 0.021646 21.7268 0.13377 0.00017662 0.7564 0.0098825 0.010909 0.0013927 0.98686 0.99165 3.0038e-006 1.2015e-005 0.16853 0.90286 0.90402 0.0014005 0.98404 0.45166 0.0018866 0.42252 2.2022 2.2014 16.0251 144.8927 0.00018169 -85.6244 0.65694
9.761 0.98816 5.454e-005 3.8183 0.011896 0.00012658 0.0011813 0.2334 0.00065931 0.23406 0.21597 0 0.032274 0.0389 0 1.6881 0.63665 0.19381 0.021647 21.7304 0.13378 0.00017663 0.7564 0.0098828 0.01091 0.0013926 0.98686 0.99165 3.0036e-006 1.2014e-005 0.16854 0.90312 0.90413 0.0014004 0.98413 0.45185 0.0018866 0.42253 2.2029 2.202 16.0251 144.8927 0.00018153 -85.6247 0.65794
9.762 0.98816 5.454e-005 3.8183 0.011896 0.00012659 0.0011813 0.2334 0.00065931 0.23406 0.21597 0 0.032274 0.0389 0 1.6882 0.6367 0.19382 0.021648 21.7339 0.13379 0.00017664 0.75639 0.0098832 0.01091 0.0013925 0.98686 0.99165 3.0034e-006 1.2014e-005 0.16854 0.90337 0.90424 0.0014004 0.98421 0.45204 0.0018865 0.42255 2.2036 2.2027 16.0251 144.8927 0.00018137 -85.625 0.65894
9.763 0.98816 5.454e-005 3.8183 0.011896 0.00012661 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6883 0.63674 0.19384 0.021649 21.7374 0.13379 0.00017665 0.75639 0.0098835 0.01091 0.0013925 0.98686 0.99165 3.0033e-006 1.2013e-005 0.16854 0.90362 0.90435 0.0014004 0.9843 0.45223 0.0018865 0.42256 2.2042 2.2033 16.0251 144.8927 0.0001812 -85.6253 0.65994
9.764 0.98816 5.454e-005 3.8183 0.011896 0.00012662 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6883 0.63678 0.19385 0.02165 21.7409 0.1338 0.00017666 0.75638 0.0098838 0.010911 0.0013924 0.98687 0.99165 3.0031e-006 1.2012e-005 0.16854 0.90387 0.90445 0.0014003 0.98438 0.45242 0.0018864 0.42258 2.2049 2.204 16.025 144.8928 0.00018104 -85.6256 0.66094
9.765 0.98816 5.454e-005 3.8183 0.011896 0.00012663 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6884 0.63683 0.19386 0.021651 21.7444 0.1338 0.00017667 0.75637 0.0098841 0.010911 0.0013923 0.98687 0.99165 3.003e-006 1.2012e-005 0.16854 0.90412 0.90456 0.0014003 0.98446 0.45261 0.0018864 0.42259 2.2055 2.2046 16.025 144.8928 0.00018088 -85.6259 0.66194
9.766 0.98816 5.454e-005 3.8183 0.011896 0.00012664 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6885 0.63687 0.19387 0.021652 21.7479 0.13381 0.00017667 0.75637 0.0098844 0.010911 0.0013923 0.98687 0.99165 3.0028e-006 1.2011e-005 0.16855 0.90436 0.90466 0.0014002 0.98454 0.4528 0.0018863 0.42261 2.2062 2.2053 16.025 144.8928 0.00018072 -85.6262 0.66294
9.767 0.98816 5.454e-005 3.8183 0.011896 0.00012666 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6886 0.63692 0.19389 0.021653 21.7515 0.13381 0.00017668 0.75636 0.0098847 0.010911 0.0013922 0.98687 0.99165 3.0027e-006 1.2011e-005 0.16855 0.90461 0.90477 0.0014002 0.98463 0.45299 0.0018863 0.42262 2.2068 2.206 16.025 144.8928 0.00018056 -85.6264 0.66394
9.768 0.98816 5.454e-005 3.8183 0.011896 0.00012667 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6887 0.63696 0.1939 0.021654 21.755 0.13382 0.00017669 0.75636 0.009885 0.010912 0.0013921 0.98687 0.99166 3.0025e-006 1.201e-005 0.16855 0.90486 0.90487 0.0014002 0.98471 0.45318 0.0018863 0.42264 2.2075 2.2066 16.0249 144.8928 0.0001804 -85.6267 0.66494
9.769 0.98816 5.4539e-005 3.8183 0.011896 0.00012668 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6887 0.637 0.19391 0.021655 21.7585 0.13382 0.0001767 0.75635 0.0098853 0.010912 0.0013921 0.98687 0.99166 3.0024e-006 1.2009e-005 0.16855 0.9051 0.90498 0.0014001 0.98479 0.45338 0.0018862 0.42265 2.2081 2.2073 16.0249 144.8929 0.00018024 -85.627 0.66594
9.77 0.98816 5.4539e-005 3.8183 0.011896 0.0001267 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6888 0.63705 0.19392 0.021656 21.762 0.13383 0.00017671 0.75635 0.0098856 0.010912 0.001392 0.98687 0.99166 3.0022e-006 1.2009e-005 0.16856 0.90535 0.90508 0.0014001 0.98487 0.45357 0.0018862 0.42267 2.2088 2.2079 16.0249 144.8929 0.00018008 -85.6273 0.66694
9.771 0.98816 5.4539e-005 3.8183 0.011896 0.00012671 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6889 0.63709 0.19394 0.021657 21.7655 0.13383 0.00017672 0.75634 0.0098859 0.010913 0.0013919 0.98687 0.99166 3.0021e-006 1.2008e-005 0.16856 0.90559 0.90518 0.0014001 0.98495 0.45376 0.0018861 0.42268 2.2094 2.2086 16.0249 144.8929 0.00017992 -85.6275 0.66794
9.772 0.98816 5.4539e-005 3.8183 0.011896 0.00012672 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.689 0.63713 0.19395 0.021658 21.769 0.13384 0.00017672 0.75634 0.0098862 0.010913 0.0013919 0.98687 0.99166 3.002e-006 1.2008e-005 0.16856 0.90584 0.90529 0.0014 0.98503 0.45395 0.0018861 0.4227 2.2101 2.2092 16.0248 144.8929 0.00017976 -85.6278 0.66894
9.773 0.98816 5.4539e-005 3.8183 0.011896 0.00012673 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6891 0.63718 0.19396 0.021658 21.7726 0.13385 0.00017673 0.75633 0.0098865 0.010913 0.0013918 0.98687 0.99166 3.0018e-006 1.2007e-005 0.16856 0.90608 0.90539 0.0014 0.98511 0.45414 0.001886 0.42271 2.2107 2.2098 16.0248 144.8929 0.0001796 -85.6281 0.66994
9.774 0.98816 5.4539e-005 3.8183 0.011896 0.00012675 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6891 0.63722 0.19397 0.021659 21.7761 0.13385 0.00017674 0.75633 0.0098868 0.010914 0.0013917 0.98687 0.99166 3.0017e-006 1.2007e-005 0.16857 0.90632 0.90549 0.0014 0.98519 0.45433 0.001886 0.42273 2.2113 2.2105 16.0248 144.893 0.00017945 -85.6283 0.67094
9.775 0.98816 5.4539e-005 3.8183 0.011896 0.00012676 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6892 0.63726 0.19399 0.02166 21.7796 0.13386 0.00017675 0.75632 0.0098871 0.010914 0.0013917 0.98687 0.99166 3.0015e-006 1.2006e-005 0.16857 0.90656 0.90559 0.0013999 0.98526 0.45452 0.001886 0.42274 2.212 2.2111 16.0248 144.893 0.00017929 -85.6286 0.67194
9.776 0.98816 5.4539e-005 3.8183 0.011896 0.00012677 0.0011813 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6893 0.63731 0.194 0.021661 21.7831 0.13386 0.00017676 0.75631 0.0098874 0.010914 0.0013916 0.98687 0.99166 3.0014e-006 1.2005e-005 0.16857 0.9068 0.9057 0.0013999 0.98534 0.45471 0.0018859 0.42276 2.2126 2.2118 16.0247 144.893 0.00017914 -85.6289 0.67294
9.777 0.98816 5.4539e-005 3.8183 0.011896 0.00012678 0.0011814 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6894 0.63735 0.19401 0.021662 21.7866 0.13387 0.00017677 0.75631 0.0098877 0.010915 0.0013916 0.98688 0.99166 3.0013e-006 1.2005e-005 0.16857 0.90704 0.9058 0.0013999 0.98542 0.4549 0.0018859 0.42277 2.2132 2.2124 16.0247 144.893 0.00017898 -85.6291 0.67394
9.778 0.98817 5.4539e-005 3.8183 0.011896 0.0001268 0.0011814 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6895 0.6374 0.19402 0.021663 21.7902 0.13387 0.00017678 0.7563 0.009888 0.010915 0.0013915 0.98688 0.99166 3.0011e-006 1.2004e-005 0.16857 0.90728 0.9059 0.0013998 0.98549 0.45509 0.0018858 0.42279 2.2139 2.213 16.0247 144.893 0.00017883 -85.6294 0.67494
9.779 0.98817 5.4539e-005 3.8183 0.011896 0.00012681 0.0011814 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6895 0.63744 0.19404 0.021664 21.7937 0.13388 0.00017678 0.7563 0.0098883 0.010915 0.0013914 0.98688 0.99166 3.001e-006 1.2004e-005 0.16858 0.90752 0.906 0.0013998 0.98557 0.45528 0.0018858 0.42281 2.2145 2.2137 16.0247 144.8931 0.00017867 -85.6296 0.67594
9.78 0.98817 5.4538e-005 3.8183 0.011896 0.00012682 0.0011814 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6896 0.63748 0.19405 0.021665 21.7972 0.13388 0.00017679 0.75629 0.0098886 0.010916 0.0013914 0.98688 0.99166 3.0009e-006 1.2003e-005 0.16858 0.90776 0.9061 0.0013998 0.98565 0.45547 0.0018857 0.42282 2.2151 2.2143 16.0247 144.8931 0.00017852 -85.6299 0.67694
9.781 0.98817 5.4538e-005 3.8183 0.011896 0.00012684 0.0011814 0.2334 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6897 0.63753 0.19406 0.021666 21.8007 0.13389 0.0001768 0.75629 0.0098889 0.010916 0.0013913 0.98688 0.99166 3.0007e-006 1.2003e-005 0.16858 0.90799 0.9062 0.0013997 0.98572 0.45566 0.0018857 0.42284 2.2158 2.2149 16.0246 144.8931 0.00017837 -85.6301 0.67794
9.782 0.98817 5.4538e-005 3.8183 0.011896 0.00012685 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6898 0.63757 0.19407 0.021667 21.8042 0.1339 0.00017681 0.75628 0.0098892 0.010916 0.0013913 0.98688 0.99166 3.0006e-006 1.2002e-005 0.16858 0.90823 0.9063 0.0013997 0.9858 0.45584 0.0018857 0.42285 2.2164 2.2156 16.0246 144.8931 0.00017822 -85.6304 0.67894
9.783 0.98817 5.4538e-005 3.8183 0.011896 0.00012686 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6899 0.63761 0.19409 0.021668 21.8078 0.1339 0.00017682 0.75628 0.0098895 0.010917 0.0013912 0.98688 0.99166 3.0005e-006 1.2002e-005 0.16859 0.90847 0.9064 0.0013997 0.98587 0.45603 0.0018856 0.42287 2.217 2.2162 16.0246 144.8931 0.00017807 -85.6306 0.67994
9.784 0.98817 5.4538e-005 3.8183 0.011896 0.00012687 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.69 0.63766 0.1941 0.021669 21.8113 0.13391 0.00017683 0.75627 0.0098898 0.010917 0.0013912 0.98688 0.99166 3.0003e-006 1.2001e-005 0.16859 0.9087 0.9065 0.0013996 0.98594 0.45622 0.0018856 0.42288 2.2176 2.2168 16.0246 144.8932 0.00017791 -85.6309 0.68094
9.785 0.98817 5.4538e-005 3.8183 0.011896 0.00012689 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.69 0.6377 0.19411 0.02167 21.8148 0.13391 0.00017684 0.75627 0.0098901 0.010917 0.0013911 0.98688 0.99166 3.0002e-006 1.2001e-005 0.16859 0.90893 0.90659 0.0013996 0.98602 0.45641 0.0018855 0.4229 2.2183 2.2174 16.0245 144.8932 0.00017776 -85.6311 0.68194
9.786 0.98817 5.4538e-005 3.8183 0.011896 0.0001269 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6901 0.63774 0.19412 0.021671 21.8183 0.13392 0.00017684 0.75626 0.0098904 0.010917 0.001391 0.98688 0.99166 3.0001e-006 1.2e-005 0.16859 0.90917 0.90669 0.0013996 0.98609 0.4566 0.0018855 0.42291 2.2189 2.2181 16.0245 144.8932 0.00017761 -85.6314 0.68294
9.787 0.98817 5.4538e-005 3.8183 0.011896 0.00012691 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6902 0.63779 0.19414 0.021672 21.8219 0.13392 0.00017685 0.75625 0.0098907 0.010918 0.001391 0.98688 0.99167 2.9999e-006 1.2e-005 0.1686 0.9094 0.90679 0.0013996 0.98616 0.45679 0.0018855 0.42293 2.2195 2.2187 16.0245 144.8932 0.00017747 -85.6316 0.68394
9.788 0.98817 5.4538e-005 3.8183 0.011896 0.00012692 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6903 0.63783 0.19415 0.021672 21.8254 0.13393 0.00017686 0.75625 0.009891 0.010918 0.0013909 0.98688 0.99167 2.9998e-006 1.1999e-005 0.1686 0.90963 0.90689 0.0013995 0.98623 0.45698 0.0018854 0.42294 2.2201 2.2193 16.0245 144.8932 0.00017732 -85.6318 0.68494
9.789 0.98817 5.4538e-005 3.8183 0.011896 0.00012694 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6904 0.63788 0.19416 0.021673 21.8289 0.13393 0.00017687 0.75624 0.0098913 0.010918 0.0013909 0.98688 0.99167 2.9997e-006 1.1999e-005 0.1686 0.90986 0.90698 0.0013995 0.9863 0.45717 0.0018854 0.42296 2.2207 2.2199 16.0244 144.8933 0.00017717 -85.6321 0.68594
9.79 0.98817 5.4538e-005 3.8183 0.011896 0.00012695 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6904 0.63792 0.19417 0.021674 21.8324 0.13394 0.00017688 0.75624 0.0098916 0.010919 0.0013908 0.98689 0.99167 2.9996e-006 1.1998e-005 0.1686 0.91009 0.90708 0.0013995 0.98637 0.45736 0.0018854 0.42297 2.2214 2.2205 16.0244 144.8933 0.00017702 -85.6323 0.68694
9.791 0.98817 5.4538e-005 3.8183 0.011896 0.00012696 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6905 0.63796 0.19418 0.021675 21.836 0.13394 0.00017689 0.75623 0.0098919 0.010919 0.0013908 0.98689 0.99167 2.9994e-006 1.1998e-005 0.1686 0.91032 0.90718 0.0013994 0.98644 0.45755 0.0018853 0.42299 2.222 2.2212 16.0244 144.8933 0.00017688 -85.6325 0.68794
9.792 0.98817 5.4537e-005 3.8183 0.011896 0.00012698 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6906 0.63801 0.1942 0.021676 21.8395 0.13395 0.0001769 0.75623 0.0098922 0.010919 0.0013907 0.98689 0.99167 2.9993e-006 1.1997e-005 0.16861 0.91055 0.90727 0.0013994 0.98651 0.45774 0.0018853 0.423 2.2226 2.2218 16.0244 144.8933 0.00017673 -85.6328 0.68894
9.793 0.98817 5.4537e-005 3.8183 0.011896 0.00012699 0.0011814 0.23339 0.00065931 0.23405 0.21597 0 0.032274 0.0389 0 1.6907 0.63805 0.19421 0.021677 21.843 0.13396 0.0001769 0.75622 0.0098925 0.01092 0.0013907 0.98689 0.99167 2.9992e-006 1.1997e-005 0.16861 0.91078 0.90737 0.0013994 0.98658 0.45793 0.0018852 0.42302 2.2232 2.2224 16.0243 144.8933 0.00017658 -85.633 0.68994
9.794 0.98817 5.4537e-005 3.8183 0.011896 0.000127 0.0011815 0.23339 0.00065931 0.23405 0.21597 0 0.032275 0.0389 0 1.6908 0.63809 0.19422 0.021678 21.8465 0.13396 0.00017691 0.75622 0.0098928 0.01092 0.0013906 0.98689 0.99167 2.9991e-006 1.1996e-005 0.16861 0.91101 0.90746 0.0013994 0.98665 0.45812 0.0018852 0.42303 2.2238 2.223 16.0243 144.8934 0.00017644 -85.6332 0.69094
9.795 0.98817 5.4537e-005 3.8183 0.011896 0.00012701 0.0011815 0.23339 0.00065931 0.23405 0.21597 0 0.032275 0.0389 0 1.6908 0.63814 0.19423 0.021679 21.8501 0.13397 0.00017692 0.75621 0.0098931 0.01092 0.0013906 0.98689 0.99167 2.9989e-006 1.1996e-005 0.16861 0.91123 0.90756 0.0013993 0.98672 0.4583 0.0018852 0.42305 2.2244 2.2236 16.0243 144.8934 0.00017629 -85.6335 0.69194
9.796 0.98817 5.4537e-005 3.8183 0.011896 0.00012703 0.0011815 0.23339 0.00065931 0.23405 0.21597 0 0.032275 0.0389 0 1.6909 0.63818 0.19425 0.02168 21.8536 0.13397 0.00017693 0.7562 0.0098934 0.010921 0.0013905 0.98689 0.99167 2.9988e-006 1.1995e-005 0.16862 0.91146 0.90765 0.0013993 0.98679 0.45849 0.0018851 0.42306 2.225 2.2242 16.0243 144.8934 0.00017615 -85.6337 0.69294
9.797 0.98817 5.4537e-005 3.8183 0.011895 0.00012704 0.0011815 0.23339 0.00065931 0.23405 0.21597 0 0.032275 0.0389 0 1.691 0.63823 0.19426 0.021681 21.8571 0.13398 0.00017694 0.7562 0.0098937 0.010921 0.0013904 0.98689 0.99167 2.9987e-006 1.1995e-005 0.16862 0.91168 0.90774 0.0013993 0.98686 0.45868 0.0018851 0.42308 2.2256 2.2248 16.0242 144.8934 0.00017601 -85.6339 0.69394
9.798 0.98817 5.4537e-005 3.8183 0.011895 0.00012705 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6911 0.63827 0.19427 0.021682 21.8606 0.13398 0.00017695 0.75619 0.009894 0.010921 0.0013904 0.98689 0.99167 2.9986e-006 1.1994e-005 0.16862 0.91191 0.90784 0.0013993 0.98692 0.45887 0.0018851 0.42309 2.2262 2.2254 16.0242 144.8935 0.00017586 -85.6341 0.69494
9.799 0.98817 5.4537e-005 3.8183 0.011895 0.00012706 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6912 0.63831 0.19428 0.021683 21.8642 0.13399 0.00017696 0.75619 0.0098943 0.010922 0.0013903 0.98689 0.99167 2.9985e-006 1.1994e-005 0.16862 0.91213 0.90793 0.0013992 0.98699 0.45906 0.001885 0.42311 2.2268 2.226 16.0242 144.8935 0.00017572 -85.6343 0.69594
9.8 0.98817 5.4537e-005 3.8183 0.011895 0.00012708 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6912 0.63836 0.1943 0.021684 21.8677 0.13399 0.00017696 0.75618 0.0098946 0.010922 0.0013903 0.98689 0.99167 2.9984e-006 1.1993e-005 0.16863 0.91236 0.90802 0.0013992 0.98706 0.45925 0.001885 0.42312 2.2274 2.2266 16.0242 144.8935 0.00017558 -85.6346 0.69694
9.801 0.98817 5.4537e-005 3.8183 0.011895 0.00012709 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6913 0.6384 0.19431 0.021685 21.8712 0.134 0.00017697 0.75618 0.0098949 0.010922 0.0013903 0.98689 0.99167 2.9982e-006 1.1993e-005 0.16863 0.91258 0.90812 0.0013992 0.98712 0.45944 0.001885 0.42314 2.228 2.2272 16.0241 144.8935 0.00017544 -85.6348 0.69794
9.802 0.98817 5.4537e-005 3.8183 0.011895 0.0001271 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6914 0.63844 0.19432 0.021685 21.8747 0.134 0.00017698 0.75617 0.0098952 0.010923 0.0013902 0.98689 0.99167 2.9981e-006 1.1992e-005 0.16863 0.9128 0.90821 0.0013991 0.98719 0.45962 0.0018849 0.42315 2.2286 2.2278 16.0241 144.8935 0.0001753 -85.635 0.69894
9.803 0.98817 5.4537e-005 3.8183 0.011895 0.00012712 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6915 0.63849 0.19433 0.021686 21.8783 0.13401 0.00017699 0.75617 0.0098955 0.010923 0.0013902 0.98689 0.99167 2.998e-006 1.1992e-005 0.16863 0.91302 0.9083 0.0013991 0.98725 0.45981 0.0018849 0.42317 2.2292 2.2284 16.0241 144.8936 0.00017516 -85.6352 0.69994
9.804 0.98817 5.4536e-005 3.8183 0.011895 0.00012713 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6916 0.63853 0.19435 0.021687 21.8818 0.13402 0.000177 0.75616 0.0098958 0.010923 0.0013901 0.98689 0.99167 2.9979e-006 1.1992e-005 0.16863 0.91324 0.90839 0.0013991 0.98732 0.46 0.0018849 0.42318 2.2298 2.229 16.024 144.8936 0.00017502 -85.6354 0.70094
9.805 0.98817 5.4536e-005 3.8183 0.011895 0.00012714 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6916 0.63857 0.19436 0.021688 21.8853 0.13402 0.00017701 0.75616 0.0098961 0.010923 0.0013901 0.9869 0.99167 2.9978e-006 1.1991e-005 0.16864 0.91346 0.90848 0.0013991 0.98738 0.46019 0.0018848 0.4232 2.2304 2.2296 16.024 144.8936 0.00017488 -85.6356 0.70194
9.806 0.98817 5.4536e-005 3.8183 0.011895 0.00012715 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6917 0.63862 0.19437 0.021689 21.8889 0.13403 0.00017701 0.75615 0.0098964 0.010924 0.00139 0.9869 0.99167 2.9977e-006 1.1991e-005 0.16864 0.91368 0.90857 0.001399 0.98744 0.46038 0.0018848 0.42321 2.231 2.2302 16.024 144.8936 0.00017474 -85.6358 0.70294
9.807 0.98817 5.4536e-005 3.8183 0.011895 0.00012717 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6918 0.63866 0.19438 0.02169 21.8924 0.13403 0.00017702 0.75614 0.0098967 0.010924 0.00139 0.9869 0.99167 2.9976e-006 1.199e-005 0.16864 0.9139 0.90866 0.001399 0.98751 0.46056 0.0018848 0.42323 2.2316 2.2308 16.024 144.8936 0.0001746 -85.636 0.70394
9.808 0.98817 5.4536e-005 3.8183 0.011895 0.00012718 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6919 0.63871 0.1944 0.021691 21.8959 0.13404 0.00017703 0.75614 0.009897 0.010924 0.0013899 0.9869 0.99167 2.9975e-006 1.199e-005 0.16864 0.91412 0.90875 0.001399 0.98757 0.46075 0.0018847 0.42324 2.2322 2.2314 16.0239 144.8937 0.00017446 -85.6363 0.70494
9.809 0.98817 5.4536e-005 3.8183 0.011895 0.00012719 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.692 0.63875 0.19441 0.021692 21.8994 0.13404 0.00017704 0.75613 0.0098973 0.010925 0.0013899 0.9869 0.99167 2.9974e-006 1.1989e-005 0.16865 0.91433 0.90884 0.001399 0.98763 0.46094 0.0018847 0.42326 2.2328 2.232 16.0239 144.8937 0.00017432 -85.6365 0.70594
9.81 0.98817 5.4536e-005 3.8183 0.011895 0.0001272 0.0011815 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.692 0.63879 0.19442 0.021693 21.903 0.13405 0.00017705 0.75613 0.0098976 0.010925 0.0013898 0.9869 0.99167 2.9973e-006 1.1989e-005 0.16865 0.91455 0.90893 0.0013989 0.98769 0.46113 0.0018847 0.42327 2.2334 2.2326 16.0239 144.8937 0.00017419 -85.6367 0.70694
9.811 0.98817 5.4536e-005 3.8183 0.011895 0.00012722 0.0011816 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6921 0.63884 0.19443 0.021694 21.9065 0.13405 0.00017706 0.75612 0.0098979 0.010925 0.0013898 0.9869 0.99168 2.9971e-006 1.1988e-005 0.16865 0.91476 0.90902 0.0013989 0.98776 0.46132 0.0018846 0.42329 2.234 2.2332 16.0239 144.8937 0.00017405 -85.6369 0.70794
9.812 0.98817 5.4536e-005 3.8183 0.011895 0.00012723 0.0011816 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6922 0.63888 0.19445 0.021695 21.91 0.13406 0.00017707 0.75612 0.0098982 0.010926 0.0013897 0.9869 0.99168 2.997e-006 1.1988e-005 0.16865 0.91498 0.90911 0.0013989 0.98782 0.4615 0.0018846 0.4233 2.2345 2.2338 16.0238 144.8937 0.00017391 -85.6371 0.70894
9.813 0.98817 5.4536e-005 3.8183 0.011895 0.00012724 0.0011816 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6923 0.63892 0.19446 0.021696 21.9136 0.13407 0.00017707 0.75611 0.0098985 0.010926 0.0013897 0.9869 0.99168 2.9969e-006 1.1988e-005 0.16865 0.91519 0.9092 0.0013989 0.98788 0.46169 0.0018846 0.42332 2.2351 2.2344 16.0238 144.8938 0.00017378 -85.6373 0.70994
9.814 0.98817 5.4536e-005 3.8183 0.011895 0.00012726 0.0011816 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6924 0.63897 0.19447 0.021697 21.9171 0.13407 0.00017708 0.75611 0.0098988 0.010926 0.0013896 0.9869 0.99168 2.9968e-006 1.1987e-005 0.16866 0.91541 0.90929 0.0013988 0.98794 0.46188 0.0018845 0.42333 2.2357 2.2349 16.0238 144.8938 0.00017364 -85.6375 0.71094
9.815 0.98817 5.4535e-005 3.8183 0.011895 0.00012727 0.0011816 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6925 0.63901 0.19448 0.021698 21.9206 0.13408 0.00017709 0.7561 0.0098991 0.010927 0.0013896 0.9869 0.99168 2.9967e-006 1.1987e-005 0.16866 0.91562 0.90938 0.0013988 0.988 0.46207 0.0018845 0.42335 2.2363 2.2355 16.0238 144.8938 0.00017351 -85.6376 0.71194
9.816 0.98817 5.4535e-005 3.8183 0.011895 0.00012728 0.0011816 0.23339 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6925 0.63905 0.1945 0.021699 21.9242 0.13408 0.0001771 0.7561 0.0098994 0.010927 0.0013895 0.9869 0.99168 2.9966e-006 1.1986e-005 0.16866 0.91583 0.90946 0.0013988 0.98806 0.46225 0.0018845 0.42336 2.2369 2.2361 16.0237 144.8938 0.00017338 -85.6378 0.71294
9.817 0.98817 5.4535e-005 3.8183 0.011895 0.00012729 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6926 0.6391 0.19451 0.021699 21.9277 0.13409 0.00017711 0.75609 0.0098997 0.010927 0.0013895 0.9869 0.99168 2.9965e-006 1.1986e-005 0.16866 0.91604 0.90955 0.0013988 0.98812 0.46244 0.0018844 0.42338 2.2374 2.2367 16.0237 144.8938 0.00017324 -85.638 0.71394
9.818 0.98817 5.4535e-005 3.8183 0.011895 0.00012731 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6927 0.63914 0.19452 0.0217 21.9312 0.13409 0.00017712 0.75608 0.0099 0.010928 0.0013895 0.9869 0.99168 2.9964e-006 1.1986e-005 0.16867 0.91625 0.90964 0.0013988 0.98818 0.46263 0.0018844 0.42339 2.238 2.2373 16.0237 144.8939 0.00017311 -85.6382 0.71494
9.819 0.98817 5.4535e-005 3.8183 0.011895 0.00012732 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6928 0.63918 0.19453 0.021701 21.9348 0.1341 0.00017713 0.75608 0.0099003 0.010928 0.0013894 0.9869 0.99168 2.9963e-006 1.1985e-005 0.16867 0.91646 0.90972 0.0013987 0.98823 0.46281 0.0018844 0.42341 2.2386 2.2378 16.0237 144.8939 0.00017298 -85.6384 0.71594
9.82 0.98817 5.4535e-005 3.8183 0.011895 0.00012733 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6929 0.63923 0.19454 0.021702 21.9383 0.1341 0.00017713 0.75607 0.0099006 0.010928 0.0013894 0.9869 0.99168 2.9962e-006 1.1985e-005 0.16867 0.91667 0.90981 0.0013987 0.98829 0.463 0.0018843 0.42342 2.2392 2.2384 16.0236 144.8939 0.00017285 -85.6386 0.71694
9.821 0.98817 5.4535e-005 3.8183 0.011895 0.00012735 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6929 0.63927 0.19456 0.021703 21.9418 0.13411 0.00017714 0.75607 0.0099009 0.010928 0.0013893 0.9869 0.99168 2.9961e-006 1.1984e-005 0.16867 0.91688 0.9099 0.0013987 0.98835 0.46319 0.0018843 0.42344 2.2397 2.239 16.0236 144.8939 0.00017271 -85.6388 0.71794
9.822 0.98817 5.4535e-005 3.8183 0.011895 0.00012736 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.693 0.63932 0.19457 0.021704 21.9454 0.13411 0.00017715 0.75606 0.0099012 0.010929 0.0013893 0.98691 0.99168 2.996e-006 1.1984e-005 0.16868 0.91709 0.90998 0.0013987 0.98841 0.46338 0.0018843 0.42345 2.2403 2.2396 16.0236 144.8939 0.00017258 -85.639 0.71894
9.823 0.98817 5.4535e-005 3.8183 0.011895 0.00012737 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6931 0.63936 0.19458 0.021705 21.9489 0.13412 0.00017716 0.75606 0.0099015 0.010929 0.0013892 0.98691 0.99168 2.9959e-006 1.1984e-005 0.16868 0.9173 0.91007 0.0013987 0.98846 0.46356 0.0018843 0.42347 2.2409 2.2401 16.0236 144.894 0.00017245 -85.6392 0.71994
9.824 0.98817 5.4535e-005 3.8183 0.011895 0.00012738 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6932 0.6394 0.19459 0.021706 21.9524 0.13413 0.00017717 0.75605 0.0099018 0.010929 0.0013892 0.98691 0.99168 2.9958e-006 1.1983e-005 0.16868 0.91751 0.91015 0.0013986 0.98852 0.46375 0.0018842 0.42348 2.2414 2.2407 16.0235 144.894 0.00017232 -85.6393 0.72094
9.825 0.98817 5.4535e-005 3.8183 0.011895 0.0001274 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6933 0.63945 0.19461 0.021707 21.956 0.13413 0.00017718 0.75605 0.0099021 0.01093 0.0013891 0.98691 0.99168 2.9957e-006 1.1983e-005 0.16868 0.91771 0.91024 0.0013986 0.98858 0.46394 0.0018842 0.4235 2.242 2.2413 16.0235 144.894 0.00017219 -85.6395 0.72194
9.826 0.98817 5.4535e-005 3.8183 0.011895 0.00012741 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6933 0.63949 0.19462 0.021708 21.9595 0.13414 0.00017719 0.75604 0.0099024 0.01093 0.0013891 0.98691 0.99168 2.9956e-006 1.1982e-005 0.16868 0.91792 0.91032 0.0013986 0.98863 0.46412 0.0018842 0.42351 2.2426 2.2418 16.0235 144.894 0.00017206 -85.6397 0.72294
9.827 0.98817 5.4534e-005 3.8183 0.011895 0.00012742 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6934 0.63953 0.19463 0.021709 21.963 0.13414 0.00017719 0.75604 0.0099027 0.01093 0.0013891 0.98691 0.99168 2.9955e-006 1.1982e-005 0.16869 0.91812 0.91041 0.0013986 0.98869 0.46431 0.0018841 0.42353 2.2431 2.2424 16.0234 144.894 0.00017194 -85.6399 0.72394
9.828 0.98817 5.4534e-005 3.8183 0.011895 0.00012743 0.0011816 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6935 0.63958 0.19464 0.02171 21.9666 0.13415 0.0001772 0.75603 0.009903 0.010931 0.001389 0.98691 0.99168 2.9954e-006 1.1982e-005 0.16869 0.91833 0.91049 0.0013985 0.98874 0.4645 0.0018841 0.42354 2.2437 2.243 16.0234 144.8941 0.00017181 -85.6401 0.72494
9.829 0.98817 5.4534e-005 3.8183 0.011895 0.00012745 0.0011817 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6936 0.63962 0.19466 0.021711 21.9701 0.13415 0.00017721 0.75602 0.0099033 0.010931 0.001389 0.98691 0.99168 2.9954e-006 1.1981e-005 0.16869 0.91853 0.91057 0.0013985 0.9888 0.46468 0.0018841 0.42356 2.2443 2.2435 16.0234 144.8941 0.00017168 -85.6402 0.72594
9.83 0.98817 5.4534e-005 3.8183 0.011895 0.00012746 0.0011817 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6937 0.63966 0.19467 0.021712 21.9736 0.13416 0.00017722 0.75602 0.0099036 0.010931 0.0013889 0.98691 0.99168 2.9953e-006 1.1981e-005 0.16869 0.91873 0.91066 0.0013985 0.98885 0.46487 0.0018841 0.42357 2.2448 2.2441 16.0234 144.8941 0.00017155 -85.6404 0.72694
9.831 0.98817 5.4534e-005 3.8183 0.011895 0.00012747 0.0011817 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6937 0.63971 0.19468 0.021712 21.9772 0.13416 0.00017723 0.75601 0.0099039 0.010932 0.0013889 0.98691 0.99168 2.9952e-006 1.1981e-005 0.1687 0.91894 0.91074 0.0013985 0.98891 0.46506 0.001884 0.42359 2.2454 2.2447 16.0233 144.8941 0.00017143 -85.6406 0.72794
9.832 0.98817 5.4534e-005 3.8183 0.011895 0.00012749 0.0011817 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6938 0.63975 0.19469 0.021713 21.9807 0.13417 0.00017724 0.75601 0.0099042 0.010932 0.0013889 0.98691 0.99168 2.9951e-006 1.198e-005 0.1687 0.91914 0.91082 0.0013985 0.98896 0.46524 0.001884 0.4236 2.246 2.2452 16.0233 144.8941 0.0001713 -85.6407 0.72894
9.833 0.98817 5.4534e-005 3.8183 0.011895 0.0001275 0.0011817 0.23338 0.00065931 0.23404 0.21596 0 0.032275 0.0389 0 1.6939 0.6398 0.19471 0.021714 21.9843 0.13417 0.00017724 0.756 0.0099045 0.010932 0.0013888 0.98691 0.99168 2.995e-006 1.198e-005 0.1687 0.91934 0.9109 0.0013984 0.98901 0.46543 0.001884 0.42362 2.2465 2.2458 16.0233 144.8942 0.00017118 -85.6409 0.72994
9.834 0.98817 5.4534e-005 3.8183 0.011895 0.00012751 0.0011817 0.23338 0.00065931 0.23403 0.21596 0 0.032275 0.0389 0 1.694 0.63984 0.19472 0.021715 21.9878 0.13418 0.00017725 0.756 0.0099048 0.010933 0.0013888 0.98691 0.99168 2.9949e-006 1.198e-005 0.1687 0.91954 0.91099 0.0013984 0.98907 0.46562 0.0018839 0.42363 2.2471 2.2463 16.0233 144.8942 0.00017105 -85.6411 0.73094
9.835 0.98817 5.4534e-005 3.8183 0.011895 0.00012752 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6941 0.63988 0.19473 0.021716 21.9913 0.13419 0.00017726 0.75599 0.0099051 0.010933 0.0013887 0.98691 0.99168 2.9948e-006 1.1979e-005 0.1687 0.91974 0.91107 0.0013984 0.98912 0.4658 0.0018839 0.42365 2.2476 2.2469 16.0232 144.8942 0.00017093 -85.6413 0.73194
9.836 0.98817 5.4534e-005 3.8183 0.011895 0.00012754 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6941 0.63993 0.19474 0.021717 21.9949 0.13419 0.00017727 0.75599 0.0099054 0.010933 0.0013887 0.98691 0.99168 2.9947e-006 1.1979e-005 0.16871 0.91994 0.91115 0.0013984 0.98917 0.46599 0.0018839 0.42366 2.2482 2.2474 16.0232 144.8942 0.0001708 -85.6414 0.73294
9.837 0.98817 5.4534e-005 3.8183 0.011895 0.00012755 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6942 0.63997 0.19476 0.021718 21.9984 0.1342 0.00017728 0.75598 0.0099057 0.010934 0.0013887 0.98691 0.99168 2.9946e-006 1.1978e-005 0.16871 0.92014 0.91123 0.0013984 0.98922 0.46617 0.0018839 0.42368 2.2487 2.248 16.0232 144.8943 0.00017068 -85.6416 0.73394
9.838 0.98817 5.4533e-005 3.8183 0.011895 0.00012756 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6943 0.64001 0.19477 0.021719 22.0019 0.1342 0.00017729 0.75598 0.009906 0.010934 0.0013886 0.98691 0.99168 2.9946e-006 1.1978e-005 0.16871 0.92034 0.91131 0.0013983 0.98928 0.46636 0.0018838 0.42369 2.2493 2.2486 16.0231 144.8943 0.00017055 -85.6417 0.73494
9.839 0.98817 5.4533e-005 3.8183 0.011895 0.00012757 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6944 0.64006 0.19478 0.02172 22.0055 0.13421 0.0001773 0.75597 0.0099063 0.010934 0.0013886 0.98691 0.99169 2.9945e-006 1.1978e-005 0.16871 0.92053 0.91139 0.0013983 0.98933 0.46655 0.0018838 0.42371 2.2498 2.2491 16.0231 144.8943 0.00017043 -85.6419 0.73594
9.84 0.98817 5.4533e-005 3.8183 0.011895 0.00012759 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6945 0.6401 0.19479 0.021721 22.009 0.13421 0.0001773 0.75596 0.0099066 0.010934 0.0013886 0.98691 0.99169 2.9944e-006 1.1977e-005 0.16872 0.92073 0.91147 0.0013983 0.98938 0.46673 0.0018838 0.42372 2.2504 2.2497 16.0231 144.8943 0.00017031 -85.6421 0.73694
9.841 0.98817 5.4533e-005 3.8183 0.011895 0.0001276 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6945 0.64014 0.19481 0.021722 22.0126 0.13422 0.00017731 0.75596 0.0099069 0.010935 0.0013885 0.98691 0.99169 2.9943e-006 1.1977e-005 0.16872 0.92093 0.91155 0.0013983 0.98943 0.46692 0.0018838 0.42374 2.2509 2.2502 16.0231 144.8943 0.00017019 -85.6422 0.73794
9.842 0.98817 5.4533e-005 3.8183 0.011895 0.00012761 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6946 0.64019 0.19482 0.021723 22.0161 0.13422 0.00017732 0.75595 0.0099072 0.010935 0.0013885 0.98692 0.99169 2.9942e-006 1.1977e-005 0.16872 0.92112 0.91163 0.0013982 0.98948 0.4671 0.0018837 0.42375 2.2515 2.2508 16.023 144.8944 0.00017006 -85.6424 0.73894
9.843 0.98817 5.4533e-005 3.8183 0.011895 0.00012763 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6947 0.64023 0.19483 0.021724 22.0196 0.13423 0.00017733 0.75595 0.0099075 0.010935 0.0013884 0.98692 0.99169 2.9941e-006 1.1976e-005 0.16872 0.92132 0.91171 0.0013982 0.98953 0.46729 0.0018837 0.42377 2.252 2.2513 16.023 144.8944 0.00016994 -85.6425 0.73994
9.844 0.98817 5.4533e-005 3.8183 0.011895 0.00012764 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6948 0.64028 0.19484 0.021724 22.0232 0.13423 0.00017734 0.75594 0.0099078 0.010936 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.16873 0.92151 0.91179 0.0013982 0.98958 0.46747 0.0018837 0.42378 2.2526 2.2518 16.023 144.8944 0.00016982 -85.6427 0.74094
9.845 0.98817 5.4533e-005 3.8183 0.011895 0.00012765 0.0011817 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6949 0.64032 0.19485 0.021725 22.0267 0.13424 0.00017735 0.75594 0.0099081 0.010936 0.0013884 0.98692 0.99169 2.994e-006 1.1976e-005 0.16873 0.92171 0.91187 0.0013982 0.98963 0.46766 0.0018837 0.4238 2.2531 2.2524 16.023 144.8944 0.0001697 -85.6429 0.74194
9.846 0.98817 5.4533e-005 3.8183 0.011895 0.00012766 0.0011818 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6949 0.64036 0.19487 0.021726 22.0303 0.13425 0.00017735 0.75593 0.0099084 0.010936 0.0013883 0.98692 0.99169 2.9939e-006 1.1975e-005 0.16873 0.9219 0.91195 0.0013982 0.98968 0.46785 0.0018836 0.42381 2.2536 2.2529 16.0229 144.8944 0.00016958 -85.643 0.74294
9.847 0.98817 5.4533e-005 3.8183 0.011895 0.00012768 0.0011818 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.695 0.64041 0.19488 0.021727 22.0338 0.13425 0.00017736 0.75593 0.0099087 0.010937 0.0013883 0.98692 0.99169 2.9938e-006 1.1975e-005 0.16873 0.92209 0.91202 0.0013982 0.98973 0.46803 0.0018836 0.42383 2.2542 2.2535 16.0229 144.8945 0.00016946 -85.6432 0.74394
9.848 0.98817 5.4533e-005 3.8183 0.011895 0.00012769 0.0011818 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6951 0.64045 0.19489 0.021728 22.0374 0.13426 0.00017737 0.75592 0.009909 0.010937 0.0013883 0.98692 0.99169 2.9937e-006 1.1975e-005 0.16873 0.92228 0.9121 0.0013982 0.98978 0.46822 0.0018836 0.42384 2.2547 2.254 16.0229 144.8945 0.00016934 -85.6433 0.74494
9.849 0.98817 5.4533e-005 3.8183 0.011895 0.0001277 0.0011818 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6952 0.64049 0.1949 0.021729 22.0409 0.13426 0.00017738 0.75592 0.0099093 0.010937 0.0013882 0.98692 0.99169 2.9937e-006 1.1975e-005 0.16874 0.92248 0.91218 0.0013981 0.98982 0.4684 0.0018836 0.42386 2.2553 2.2546 16.0228 144.8945 0.00016923 -85.6435 0.74594
9.85 0.98817 5.4532e-005 3.8183 0.011895 0.00012771 0.0011818 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6953 0.64054 0.19492 0.02173 22.0444 0.13427 0.00017739 0.75591 0.0099096 0.010938 0.0013882 0.98692 0.99169 2.9936e-006 1.1974e-005 0.16874 0.92267 0.91226 0.0013981 0.98987 0.46859 0.0018835 0.42387 2.2558 2.2551 16.0228 144.8945 0.00016911 -85.6436 0.74694
9.851 0.98817 5.4532e-005 3.8183 0.011894 0.00012773 0.0011818 0.23338 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6954 0.64058 0.19493 0.021731 22.048 0.13427 0.0001774 0.7559 0.0099098 0.010938 0.0013882 0.98692 0.99169 2.9935e-006 1.1974e-005 0.16874 0.92286 0.91233 0.0013981 0.98992 0.46877 0.0018835 0.42389 2.2563 2.2556 16.0228 144.8945 0.00016899 -85.6438 0.74794
9.852 0.98817 5.4532e-005 3.8183 0.011894 0.00012774 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6954 0.64062 0.19494 0.021732 22.0515 0.13428 0.00017741 0.7559 0.0099101 0.010938 0.0013881 0.98692 0.99169 2.9934e-006 1.1974e-005 0.16874 0.92305 0.91241 0.0013981 0.98997 0.46896 0.0018835 0.4239 2.2569 2.2562 16.0228 144.8946 0.00016887 -85.6439 0.74894
9.853 0.98817 5.4532e-005 3.8183 0.011894 0.00012775 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6955 0.64067 0.19495 0.021733 22.0551 0.13428 0.00017741 0.75589 0.0099104 0.010939 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.16875 0.92324 0.91249 0.0013981 0.99001 0.46914 0.0018835 0.42392 2.2574 2.2567 16.0227 144.8946 0.00016876 -85.6441 0.74994
9.854 0.98817 5.4532e-005 3.8183 0.011894 0.00012777 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6956 0.64071 0.19497 0.021734 22.0586 0.13429 0.00017742 0.75589 0.0099107 0.010939 0.0013881 0.98692 0.99169 2.9933e-006 1.1973e-005 0.16875 0.92342 0.91256 0.001398 0.99006 0.46933 0.0018835 0.42393 2.2579 2.2572 16.0227 144.8946 0.00016864 -85.6442 0.75094
9.855 0.98817 5.4532e-005 3.8183 0.011894 0.00012778 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6957 0.64075 0.19498 0.021735 22.0622 0.13429 0.00017743 0.75588 0.009911 0.010939 0.001388 0.98692 0.99169 2.9932e-006 1.1973e-005 0.16875 0.92361 0.91264 0.001398 0.99011 0.46951 0.0018834 0.42395 2.2585 2.2578 16.0227 144.8946 0.00016852 -85.6443 0.75194
9.856 0.98817 5.4532e-005 3.8183 0.011894 0.00012779 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6958 0.6408 0.19499 0.021736 22.0657 0.1343 0.00017744 0.75588 0.0099113 0.010939 0.001388 0.98692 0.99169 2.9931e-006 1.1972e-005 0.16875 0.9238 0.91271 0.001398 0.99015 0.4697 0.0018834 0.42396 2.259 2.2583 16.0226 144.8946 0.00016841 -85.6445 0.75294
9.857 0.98817 5.4532e-005 3.8183 0.011894 0.0001278 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6958 0.64084 0.195 0.021737 22.0692 0.13431 0.00017745 0.75587 0.0099116 0.01094 0.001388 0.98692 0.99169 2.993e-006 1.1972e-005 0.16875 0.92399 0.91279 0.001398 0.9902 0.46988 0.0018834 0.42398 2.2595 2.2588 16.0226 144.8947 0.00016829 -85.6446 0.75394
9.858 0.98817 5.4532e-005 3.8183 0.011894 0.00012782 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6959 0.64089 0.19502 0.021737 22.0728 0.13431 0.00017746 0.75587 0.0099119 0.01094 0.0013879 0.98692 0.99169 2.993e-006 1.1972e-005 0.16876 0.92417 0.91286 0.001398 0.99024 0.47007 0.0018834 0.42399 2.26 2.2594 16.0226 144.8947 0.00016818 -85.6448 0.75494
9.859 0.98817 5.4532e-005 3.8183 0.011894 0.00012783 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.696 0.64093 0.19503 0.021738 22.0763 0.13432 0.00017747 0.75586 0.0099122 0.01094 0.0013879 0.98692 0.99169 2.9929e-006 1.1971e-005 0.16876 0.92436 0.91294 0.0013979 0.99029 0.47025 0.0018833 0.42401 2.2606 2.2599 16.0226 144.8947 0.00016806 -85.6449 0.75594
9.86 0.98817 5.4532e-005 3.8183 0.011894 0.00012784 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6961 0.64097 0.19504 0.021739 22.0799 0.13432 0.00017747 0.75586 0.0099125 0.010941 0.0013879 0.98692 0.99169 2.9928e-006 1.1971e-005 0.16876 0.92454 0.91301 0.0013979 0.99033 0.47044 0.0018833 0.42402 2.2611 2.2604 16.0225 144.8947 0.00016795 -85.6451 0.75694
9.861 0.98817 5.4532e-005 3.8183 0.011894 0.00012785 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6962 0.64102 0.19505 0.02174 22.0834 0.13433 0.00017748 0.75585 0.0099128 0.010941 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.16876 0.92473 0.91309 0.0013979 0.99038 0.47062 0.0018833 0.42404 2.2616 2.2609 16.0225 144.8947 0.00016784 -85.6452 0.75794
9.862 0.98817 5.4531e-005 3.8183 0.011894 0.00012787 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6962 0.64106 0.19507 0.021741 22.087 0.13433 0.00017749 0.75584 0.0099131 0.010941 0.0013878 0.98692 0.99169 2.9927e-006 1.1971e-005 0.16877 0.92491 0.91316 0.0013979 0.99042 0.4708 0.0018833 0.42405 2.2621 2.2615 16.0225 144.8948 0.00016772 -85.6453 0.75894
9.863 0.98817 5.4531e-005 3.8183 0.011894 0.00012788 0.0011818 0.23337 0.00065931 0.23403 0.21595 0 0.032275 0.0389 0 1.6963 0.6411 0.19508 0.021742 22.0905 0.13434 0.0001775 0.75584 0.0099134 0.010942 0.0013878 0.98692 0.99169 2.9926e-006 1.197e-005 0.16877 0.92509 0.91324 0.0013979 0.99047 0.47099 0.0018832 0.42407 2.2627 2.262 16.0224 144.8948 0.00016761 -85.6455 0.75994
9.864 0.98817 5.4531e-005 3.8183 0.011894 0.00012789 0.0011819 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.6964 0.64115 0.19509 0.021743 22.0941 0.13434 0.00017751 0.75583 0.0099137 0.010942 0.0013877 0.98692 0.99169 2.9925e-006 1.197e-005 0.16877 0.92528 0.91331 0.0013979 0.99051 0.47117 0.0018832 0.42408 2.2632 2.2625 16.0224 144.8948 0.0001675 -85.6456 0.76094
9.865 0.98817 5.4531e-005 3.8183 0.011894 0.00012791 0.0011819 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.6965 0.64119 0.1951 0.021744 22.0976 0.13435 0.00017752 0.75583 0.009914 0.010942 0.0013877 0.98693 0.99169 2.9924e-006 1.197e-005 0.16877 0.92546 0.91338 0.0013978 0.99055 0.47136 0.0018832 0.42409 2.2637 2.263 16.0224 144.8948 0.00016739 -85.6457 0.76194
9.866 0.98817 5.4531e-005 3.8183 0.011894 0.00012792 0.0011819 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.6966 0.64123 0.19512 0.021745 22.1012 0.13435 0.00017752 0.75582 0.0099143 0.010943 0.0013877 0.98693 0.99169 2.9924e-006 1.1969e-005 0.16878 0.92564 0.91346 0.0013978 0.9906 0.47154 0.0018832 0.42411 2.2642 2.2635 16.0224 144.8948 0.00016727 -85.6459 0.76294
9.867 0.98817 5.4531e-005 3.8183 0.011894 0.00012793 0.0011819 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.6966 0.64128 0.19513 0.021746 22.1047 0.13436 0.00017753 0.75582 0.0099146 0.010943 0.0013876 0.98693 0.99169 2.9923e-006 1.1969e-005 0.16878 0.92582 0.91353 0.0013978 0.99064 0.47173 0.0018832 0.42412 2.2647 2.2641 16.0223 144.8949 0.00016716 -85.646 0.76394
9.868 0.98817 5.4531e-005 3.8183 0.011894 0.00012794 0.0011819 0.23337 0.00065931 0.23403 0.21595 0 0.032276 0.0389 0 1.6967 0.64132 0.19514 0.021747 22.1083 0.13437 0.00017754 0.75581 0.0099149 0.010943 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.16878 0.926 0.9136 0.0013978 0.99068 0.47191 0.0018831 0.42414 2.2652 2.2646 16.0223 144.8949 0.00016705 -85.6461 0.76494
9.869 0.98817 5.4531e-005 3.8183 0.011894 0.00012796 0.0011819 0.23337 0.00065931 0.23402 0.21595 0 0.032276 0.0389 0 1.6968 0.64137 0.19515 0.021748 22.1118 0.13437 0.00017755 0.75581 0.0099152 0.010944 0.0013876 0.98693 0.99169 2.9922e-006 1.1969e-005 0.16878 0.92618 0.91367 0.0013978 0.99072 0.47209 0.0018831 0.42415 2.2658 2.2651 16.0223 144.8949 0.00016694 -85.6462 0.76594
9.87 0.98817 5.4531e-005 3.8183 0.011894 0.00012797 0.0011819 0.23337 0.00065931 0.23402 0.21595 0 0.032276 0.0389 0 1.6969 0.64141 0.19516 0.021749 22.1154 0.13438 0.00017756 0.7558 0.0099155 0.010944 0.0013876 0.98693 0.99169 2.9921e-006 1.1968e-005 0.16878 0.92636 0.91374 0.0013977 0.99076 0.47228 0.0018831 0.42417 2.2663 2.2656 16.0222 144.8949 0.00016683 -85.6464 0.76694
9.871 0.98817 5.4531e-005 3.8183 0.011894 0.00012798 0.0011819 0.23337 0.00065931 0.23402 0.21595 0 0.032276 0.0389 0 1.697 0.64145 0.19518 0.021749 22.1189 0.13438 0.00017757 0.7558 0.0099158 0.010944 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16879 0.92654 0.91382 0.0013977 0.99081 0.47246 0.0018831 0.42418 2.2668 2.2661 16.0222 144.895 0.00016672 -85.6465 0.76794
9.872 0.98817 5.4531e-005 3.8183 0.011894 0.00012799 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.697 0.6415 0.19519 0.02175 22.1225 0.13439 0.00017758 0.75579 0.0099161 0.010944 0.0013875 0.98693 0.99169 2.992e-006 1.1968e-005 0.16879 0.92672 0.91389 0.0013977 0.99085 0.47265 0.0018831 0.4242 2.2673 2.2666 16.0222 144.895 0.00016661 -85.6466 0.76894
9.873 0.98817 5.453e-005 3.8183 0.011894 0.00012801 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6971 0.64154 0.1952 0.021751 22.126 0.13439 0.00017758 0.75578 0.0099164 0.010945 0.0013875 0.98693 0.99169 2.9919e-006 1.1968e-005 0.16879 0.92689 0.91396 0.0013977 0.99089 0.47283 0.001883 0.42421 2.2678 2.2671 16.0222 144.895 0.00016651 -85.6468 0.76994
9.874 0.98817 5.453e-005 3.8183 0.011894 0.00012802 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6972 0.64158 0.19521 0.021752 22.1296 0.1344 0.00017759 0.75578 0.0099167 0.010945 0.0013874 0.98693 0.99169 2.9918e-006 1.1967e-005 0.16879 0.92707 0.91403 0.0013977 0.99093 0.47301 0.001883 0.42423 2.2683 2.2677 16.0221 144.895 0.0001664 -85.6469 0.77094
9.875 0.98817 5.453e-005 3.8183 0.011894 0.00012803 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6973 0.64163 0.19523 0.021753 22.1331 0.1344 0.0001776 0.75577 0.009917 0.010945 0.0013874 0.98693 0.9917 2.9918e-006 1.1967e-005 0.1688 0.92725 0.9141 0.0013977 0.99097 0.4732 0.001883 0.42424 2.2688 2.2682 16.0221 144.895 0.00016629 -85.647 0.77194
9.876 0.98817 5.453e-005 3.8183 0.011894 0.00012805 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6974 0.64167 0.19524 0.021754 22.1367 0.13441 0.00017761 0.75577 0.0099173 0.010946 0.0013874 0.98693 0.9917 2.9917e-006 1.1967e-005 0.1688 0.92742 0.91417 0.0013977 0.99101 0.47338 0.001883 0.42426 2.2693 2.2687 16.0221 144.8951 0.00016618 -85.6471 0.77294
9.877 0.98817 5.453e-005 3.8183 0.011894 0.00012806 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6974 0.64171 0.19525 0.021755 22.1402 0.13441 0.00017762 0.75576 0.0099176 0.010946 0.0013874 0.98693 0.9917 2.9916e-006 1.1966e-005 0.1688 0.9276 0.91424 0.0013976 0.99105 0.47356 0.001883 0.42427 2.2698 2.2692 16.022 144.8951 0.00016607 -85.6472 0.77394
9.878 0.98817 5.453e-005 3.8183 0.011894 0.00012807 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6975 0.64176 0.19526 0.021756 22.1438 0.13442 0.00017763 0.75576 0.0099179 0.010946 0.0013873 0.98693 0.9917 2.9916e-006 1.1966e-005 0.1688 0.92777 0.91431 0.0013976 0.99109 0.47375 0.0018829 0.42429 2.2703 2.2697 16.022 144.8951 0.00016597 -85.6474 0.77494
9.879 0.98817 5.453e-005 3.8183 0.011894 0.00012808 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6976 0.6418 0.19528 0.021757 22.1473 0.13443 0.00017763 0.75575 0.0099182 0.010947 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.1688 0.92795 0.91438 0.0013976 0.99113 0.47393 0.0018829 0.4243 2.2708 2.2702 16.022 144.8951 0.00016586 -85.6475 0.77594
9.88 0.98817 5.453e-005 3.8183 0.011894 0.0001281 0.0011819 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6977 0.64184 0.19529 0.021758 22.1509 0.13443 0.00017764 0.75575 0.0099185 0.010947 0.0013873 0.98693 0.9917 2.9915e-006 1.1966e-005 0.16881 0.92812 0.91445 0.0013976 0.99117 0.47411 0.0018829 0.42432 2.2714 2.2707 16.022 144.8951 0.00016576 -85.6476 0.77694
9.881 0.98817 5.453e-005 3.8183 0.011894 0.00012811 0.001182 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6978 0.64189 0.1953 0.021759 22.1544 0.13444 0.00017765 0.75574 0.0099188 0.010947 0.0013872 0.98693 0.9917 2.9914e-006 1.1965e-005 0.16881 0.9283 0.91452 0.0013976 0.99121 0.4743 0.0018829 0.42433 2.2719 2.2712 16.0219 144.8952 0.00016565 -85.6477 0.77794
9.882 0.98817 5.453e-005 3.8183 0.011894 0.00012812 0.001182 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6978 0.64193 0.19531 0.02176 22.158 0.13444 0.00017766 0.75574 0.0099191 0.010948 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16881 0.92847 0.91459 0.0013976 0.99125 0.47448 0.0018829 0.42434 2.2724 2.2717 16.0219 144.8952 0.00016554 -85.6478 0.77894
9.883 0.98817 5.453e-005 3.8183 0.011894 0.00012813 0.001182 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6979 0.64198 0.19533 0.021761 22.1615 0.13445 0.00017767 0.75573 0.0099194 0.010948 0.0013872 0.98693 0.9917 2.9913e-006 1.1965e-005 0.16881 0.92864 0.91466 0.0013976 0.99129 0.47466 0.0018829 0.42436 2.2729 2.2722 16.0219 144.8952 0.00016544 -85.648 0.77994
9.884 0.98817 5.453e-005 3.8183 0.011894 0.00012815 0.001182 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.698 0.64202 0.19534 0.021761 22.1651 0.13445 0.00017768 0.75573 0.0099197 0.010948 0.0013872 0.98693 0.9917 2.9912e-006 1.1965e-005 0.16882 0.92881 0.91472 0.0013976 0.99132 0.47485 0.0018828 0.42437 2.2734 2.2727 16.0218 144.8952 0.00016534 -85.6481 0.78094
9.885 0.98817 5.4529e-005 3.8183 0.011894 0.00012816 0.001182 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6981 0.64206 0.19535 0.021762 22.1686 0.13446 0.00017769 0.75572 0.00992 0.010949 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.16882 0.92898 0.91479 0.0013975 0.99136 0.47503 0.0018828 0.42439 2.2738 2.2732 16.0218 144.8952 0.00016523 -85.6482 0.78194
9.886 0.98817 5.4529e-005 3.8183 0.011894 0.00012817 0.001182 0.23337 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6982 0.64211 0.19536 0.021763 22.1722 0.13446 0.00017769 0.75571 0.0099203 0.010949 0.0013871 0.98693 0.9917 2.9911e-006 1.1964e-005 0.16882 0.92915 0.91486 0.0013975 0.9914 0.47521 0.0018828 0.4244 2.2743 2.2737 16.0218 144.8953 0.00016513 -85.6483 0.78294
9.887 0.98817 5.4529e-005 3.8183 0.011894 0.00012819 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6982 0.64215 0.19537 0.021764 22.1757 0.13447 0.0001777 0.75571 0.0099206 0.010949 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16882 0.92932 0.91493 0.0013975 0.99144 0.4754 0.0018828 0.42442 2.2748 2.2742 16.0218 144.8953 0.00016502 -85.6484 0.78394
9.888 0.98817 5.4529e-005 3.8183 0.011894 0.0001282 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6983 0.64219 0.19539 0.021765 22.1793 0.13447 0.00017771 0.7557 0.0099208 0.010949 0.0013871 0.98693 0.9917 2.991e-006 1.1964e-005 0.16883 0.92949 0.91499 0.0013975 0.99148 0.47558 0.0018828 0.42443 2.2753 2.2747 16.0217 144.8953 0.00016492 -85.6485 0.78494
9.889 0.98817 5.4529e-005 3.8183 0.011894 0.00012821 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6984 0.64224 0.1954 0.021766 22.1828 0.13448 0.00017772 0.7557 0.0099211 0.01095 0.001387 0.98693 0.9917 2.9909e-006 1.1964e-005 0.16883 0.92966 0.91506 0.0013975 0.99151 0.47576 0.0018827 0.42445 2.2758 2.2752 16.0217 144.8953 0.00016482 -85.6486 0.78594
9.89 0.98817 5.4529e-005 3.8183 0.011894 0.00012822 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6985 0.64228 0.19541 0.021767 22.1864 0.13449 0.00017773 0.75569 0.0099214 0.01095 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.16883 0.92983 0.91513 0.0013975 0.99155 0.47594 0.0018827 0.42446 2.2763 2.2757 16.0217 144.8953 0.00016472 -85.6487 0.78694
9.891 0.98817 5.4529e-005 3.8183 0.011894 0.00012824 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6986 0.64232 0.19542 0.021768 22.19 0.13449 0.00017774 0.75569 0.0099217 0.01095 0.001387 0.98693 0.9917 2.9908e-006 1.1963e-005 0.16883 0.93 0.9152 0.0013975 0.99159 0.47613 0.0018827 0.42448 2.2768 2.2762 16.0216 144.8954 0.00016461 -85.6488 0.78794
9.892 0.98817 5.4529e-005 3.8183 0.011894 0.00012825 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6986 0.64237 0.19544 0.021769 22.1935 0.1345 0.00017774 0.75568 0.009922 0.010951 0.001387 0.98694 0.9917 2.9907e-006 1.1963e-005 0.16883 0.93017 0.91526 0.0013974 0.99162 0.47631 0.0018827 0.42449 2.2773 2.2767 16.0216 144.8954 0.00016451 -85.649 0.78894
9.893 0.98817 5.4529e-005 3.8183 0.011894 0.00012826 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6987 0.64241 0.19545 0.02177 22.1971 0.1345 0.00017775 0.75568 0.0099223 0.010951 0.0013869 0.98694 0.9917 2.9907e-006 1.1963e-005 0.16884 0.93033 0.91533 0.0013974 0.99166 0.47649 0.0018827 0.42451 2.2778 2.2772 16.0216 144.8954 0.00016441 -85.6491 0.78994
9.894 0.98817 5.4529e-005 3.8183 0.011894 0.00012827 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6988 0.64245 0.19546 0.021771 22.2006 0.13451 0.00017776 0.75567 0.0099226 0.010951 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16884 0.9305 0.91539 0.0013974 0.99169 0.47667 0.0018827 0.42452 2.2783 2.2776 16.0215 144.8954 0.00016431 -85.6492 0.79094
9.895 0.98817 5.4529e-005 3.8183 0.011894 0.00012829 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6989 0.6425 0.19547 0.021772 22.2042 0.13451 0.00017777 0.75567 0.0099229 0.010952 0.0013869 0.98694 0.9917 2.9906e-006 1.1962e-005 0.16884 0.93066 0.91546 0.0013974 0.99173 0.47686 0.0018826 0.42454 2.2788 2.2781 16.0215 144.8954 0.00016421 -85.6493 0.79194
9.896 0.98817 5.4529e-005 3.8183 0.011894 0.0001283 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.699 0.64254 0.19549 0.021773 22.2077 0.13452 0.00017778 0.75566 0.0099232 0.010952 0.0013869 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16884 0.93083 0.91552 0.0013974 0.99177 0.47704 0.0018826 0.42455 2.2792 2.2786 16.0215 144.8955 0.00016411 -85.6494 0.79294
9.897 0.98817 5.4528e-005 3.8183 0.011894 0.00012831 0.001182 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6991 0.64259 0.1955 0.021773 22.2113 0.13452 0.00017779 0.75565 0.0099235 0.010952 0.0013868 0.98694 0.9917 2.9905e-006 1.1962e-005 0.16885 0.93099 0.91559 0.0013974 0.9918 0.47722 0.0018826 0.42456 2.2797 2.2791 16.0215 144.8955 0.00016401 -85.6495 0.79394
9.898 0.98817 5.4528e-005 3.8183 0.011894 0.00012833 0.0011821 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6991 0.64263 0.19551 0.021774 22.2149 0.13453 0.0001778 0.75565 0.0099238 0.010953 0.0013868 0.98694 0.9917 2.9904e-006 1.1962e-005 0.16885 0.93116 0.91565 0.0013974 0.99184 0.4774 0.0018826 0.42458 2.2802 2.2796 16.0214 144.8955 0.00016391 -85.6496 0.79494
9.899 0.98817 5.4528e-005 3.8183 0.011894 0.00012834 0.0011821 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6992 0.64267 0.19552 0.021775 22.2184 0.13453 0.0001778 0.75564 0.0099241 0.010953 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16885 0.93132 0.91572 0.0013973 0.99187 0.47759 0.0018826 0.42459 2.2807 2.2801 16.0214 144.8955 0.00016381 -85.6497 0.79594
9.9 0.98817 5.4528e-005 3.8184 0.011894 0.00012835 0.0011821 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6993 0.64272 0.19554 0.021776 22.222 0.13454 0.00017781 0.75564 0.0099244 0.010953 0.0013868 0.98694 0.9917 2.9903e-006 1.1961e-005 0.16885 0.93149 0.91578 0.0013973 0.9919 0.47777 0.0018826 0.42461 2.2812 2.2806 16.0214 144.8955 0.00016371 -85.6498 0.79694
9.901 0.98817 5.4528e-005 3.8184 0.011894 0.00012836 0.0011821 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6994 0.64276 0.19555 0.021777 22.2255 0.13454 0.00017782 0.75563 0.0099247 0.010953 0.0013868 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16885 0.93165 0.91585 0.0013973 0.99194 0.47795 0.0018825 0.42462 2.2817 2.281 16.0213 144.8956 0.00016362 -85.6499 0.79794
9.902 0.98817 5.4528e-005 3.8184 0.011894 0.00012838 0.0011821 0.23336 0.00065931 0.23402 0.21594 0 0.032276 0.0389 0 1.6995 0.6428 0.19556 0.021778 22.2291 0.13455 0.00017783 0.75563 0.009925 0.010954 0.0013867 0.98694 0.9917 2.9902e-006 1.1961e-005 0.16886 0.93181 0.91591 0.0013973 0.99197 0.47813 0.0018825 0.42464 2.2821 2.2815 16.0213 144.8956 0.00016352 -85.65 0.79894
9.903 0.98817 5.4528e-005 3.8184 0.011894 0.00012839 0.0011821 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.6995 0.64285 0.19557 0.021779 22.2326 0.13456 0.00017784 0.75562 0.0099253 0.010954 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.16886 0.93197 0.91598 0.0013973 0.99201 0.47831 0.0018825 0.42465 2.2826 2.282 16.0213 144.8956 0.00016342 -85.6501 0.79994
9.904 0.98817 5.4528e-005 3.8184 0.011894 0.0001284 0.0011821 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.6996 0.64289 0.19559 0.02178 22.2362 0.13456 0.00017785 0.75562 0.0099256 0.010954 0.0013867 0.98694 0.9917 2.9901e-006 1.196e-005 0.16886 0.93213 0.91604 0.0013973 0.99204 0.47849 0.0018825 0.42467 2.2831 2.2825 16.0212 144.8956 0.00016332 -85.6502 0.80094
9.905 0.98817 5.4528e-005 3.8184 0.011893 0.00012841 0.0011821 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.6997 0.64293 0.1956 0.021781 22.2398 0.13457 0.00017785 0.75561 0.0099259 0.010955 0.0013867 0.98694 0.9917 2.99e-006 1.196e-005 0.16886 0.93229 0.9161 0.0013973 0.99207 0.47868 0.0018825 0.42468 2.2836 2.283 16.0212 144.8957 0.00016323 -85.6503 0.80194
9.906 0.98817 5.4528e-005 3.8184 0.011893 0.00012843 0.0011821 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.6998 0.64298 0.19561 0.021782 22.2433 0.13457 0.00017786 0.75561 0.0099262 0.010955 0.0013866 0.98694 0.9917 2.99e-006 1.196e-005 0.16887 0.93245 0.91617 0.0013973 0.99211 0.47886 0.0018825 0.4247 2.2841 2.2834 16.0212 144.8957 0.00016313 -85.6504 0.80294
9.907 0.98817 5.4528e-005 3.8184 0.011893 0.00012844 0.0011821 0.23336 0.00065931 0.23401 0.21594 0 0.032276 0.0389 0 1.6999 0.64302 0.19562 0.021783 22.2469 0.13458 0.00017787 0.7556 0.0099265 0.010955 0.0013866 0.98694 0.9917 2.9899e-006 1.196e-005 0.16887 0.93261 0.91623 0.0013973 0.99214 0.47904 0.0018824 0.42471 2.2845 2.2839 16.0212 144.8957 0.00016303 -85.6505 0.80394
9.908 0.98817 5.4527e-005 3.8184 0.011893 0.00012845 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.6999 0.64306 0.19563 0.021784 22.2504 0.13458 0.00017788 0.7556 0.0099268 0.010956 0.0013866 0.98694 0.9917 2.9899e-006 1.1959e-005 0.16887 0.93277 0.91629 0.0013972 0.99217 0.47922 0.0018824 0.42472 2.285 2.2844 16.0211 144.8957 0.00016294 -85.6506 0.80494
9.909 0.98817 5.4527e-005 3.8184 0.011893 0.00012847 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7 0.64311 0.19565 0.021785 22.254 0.13459 0.00017789 0.75559 0.0099271 0.010956 0.0013866 0.98694 0.9917 2.9898e-006 1.1959e-005 0.16887 0.93293 0.91635 0.0013972 0.99221 0.4794 0.0018824 0.42474 2.2855 2.2849 16.0211 144.8957 0.00016284 -85.6507 0.80594
9.91 0.98817 5.4527e-005 3.8184 0.011893 0.00012848 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7001 0.64315 0.19566 0.021785 22.2576 0.13459 0.0001779 0.75558 0.0099274 0.010956 0.0013865 0.98694 0.9917 2.9898e-006 1.1959e-005 0.16887 0.93309 0.91642 0.0013972 0.99224 0.47958 0.0018824 0.42475 2.2859 2.2853 16.0211 144.8958 0.00016275 -85.6508 0.80694
9.911 0.98817 5.4527e-005 3.8184 0.011893 0.00012849 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7002 0.6432 0.19567 0.021786 22.2611 0.1346 0.0001779 0.75558 0.0099277 0.010957 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.16888 0.93325 0.91648 0.0013972 0.99227 0.47977 0.0018824 0.42477 2.2864 2.2858 16.021 144.8958 0.00016265 -85.6508 0.80794
9.912 0.98817 5.4527e-005 3.8184 0.011893 0.0001285 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7003 0.64324 0.19568 0.021787 22.2647 0.1346 0.00017791 0.75557 0.009928 0.010957 0.0013865 0.98694 0.9917 2.9897e-006 1.1959e-005 0.16888 0.9334 0.91654 0.0013972 0.9923 0.47995 0.0018824 0.42478 2.2869 2.2863 16.021 144.8958 0.00016256 -85.6509 0.80894
9.913 0.98817 5.4527e-005 3.8184 0.011893 0.00012852 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7003 0.64328 0.1957 0.021788 22.2683 0.13461 0.00017792 0.75557 0.0099282 0.010957 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16888 0.93356 0.9166 0.0013972 0.99233 0.48013 0.0018824 0.4248 2.2874 2.2868 16.021 144.8958 0.00016246 -85.651 0.80994
9.914 0.98817 5.4527e-005 3.8184 0.011893 0.00012853 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7004 0.64333 0.19571 0.021789 22.2718 0.13462 0.00017793 0.75556 0.0099285 0.010958 0.0013865 0.98694 0.9917 2.9896e-006 1.1958e-005 0.16888 0.93372 0.91666 0.0013972 0.99236 0.48031 0.0018823 0.42481 2.2878 2.2872 16.0209 144.8958 0.00016237 -85.6511 0.81094
9.915 0.98817 5.4527e-005 3.8184 0.011893 0.00012854 0.0011821 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7005 0.64337 0.19572 0.02179 22.2754 0.13462 0.00017794 0.75556 0.0099288 0.010958 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16889 0.93387 0.91672 0.0013972 0.9924 0.48049 0.0018823 0.42483 2.2883 2.2877 16.0209 144.8959 0.00016228 -85.6512 0.81194
9.916 0.98817 5.4527e-005 3.8184 0.011893 0.00012855 0.0011822 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7006 0.64341 0.19573 0.021791 22.2789 0.13463 0.00017795 0.75555 0.0099291 0.010958 0.0013864 0.98694 0.9917 2.9895e-006 1.1958e-005 0.16889 0.93403 0.91679 0.0013972 0.99243 0.48067 0.0018823 0.42484 2.2888 2.2882 16.0209 144.8959 0.00016218 -85.6513 0.81294
9.917 0.98817 5.4527e-005 3.8184 0.011893 0.00012857 0.0011822 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7007 0.64346 0.19575 0.021792 22.2825 0.13463 0.00017796 0.75555 0.0099294 0.010958 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.16889 0.93418 0.91685 0.0013972 0.99246 0.48085 0.0018823 0.42486 2.2892 2.2886 16.0209 144.8959 0.00016209 -85.6514 0.81394
9.918 0.98817 5.4527e-005 3.8184 0.011893 0.00012858 0.0011822 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7007 0.6435 0.19576 0.021793 22.2861 0.13464 0.00017796 0.75554 0.0099297 0.010959 0.0013864 0.98694 0.9917 2.9894e-006 1.1958e-005 0.16889 0.93434 0.91691 0.0013971 0.99249 0.48103 0.0018823 0.42487 2.2897 2.2891 16.0208 144.8959 0.000162 -85.6515 0.81494
9.919 0.98817 5.4527e-005 3.8184 0.011893 0.00012859 0.0011822 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7008 0.64354 0.19577 0.021794 22.2896 0.13464 0.00017797 0.75554 0.00993 0.010959 0.0013864 0.98694 0.9917 2.9894e-006 1.1957e-005 0.16889 0.93449 0.91697 0.0013971 0.99252 0.48121 0.0018823 0.42488 2.2902 2.2896 16.0208 144.8959 0.00016191 -85.6516 0.81594
9.92 0.98817 5.4526e-005 3.8184 0.011893 0.00012861 0.0011822 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7009 0.64359 0.19578 0.021795 22.2932 0.13465 0.00017798 0.75553 0.0099303 0.010959 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.1689 0.93464 0.91703 0.0013971 0.99255 0.48139 0.0018823 0.4249 2.2906 2.29 16.0208 144.896 0.00016181 -85.6516 0.81694
9.921 0.98817 5.4526e-005 3.8184 0.011893 0.00012862 0.0011822 0.23336 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.701 0.64363 0.1958 0.021796 22.2968 0.13465 0.00017799 0.75552 0.0099306 0.01096 0.0013863 0.98694 0.9917 2.9893e-006 1.1957e-005 0.1689 0.9348 0.91709 0.0013971 0.99258 0.48158 0.0018822 0.42491 2.2911 2.2905 16.0207 144.896 0.00016172 -85.6517 0.81794
9.922 0.98817 5.4526e-005 3.8184 0.011893 0.00012863 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7011 0.64367 0.19581 0.021796 22.3003 0.13466 0.000178 0.75552 0.0099309 0.01096 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.1689 0.93495 0.91715 0.0013971 0.99261 0.48176 0.0018822 0.42493 2.2915 2.2909 16.0207 144.896 0.00016163 -85.6518 0.81894
9.923 0.98817 5.4526e-005 3.8184 0.011893 0.00012864 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7011 0.64372 0.19582 0.021797 22.3039 0.13466 0.00017801 0.75551 0.0099312 0.01096 0.0013863 0.98694 0.9917 2.9892e-006 1.1957e-005 0.1689 0.9351 0.91721 0.0013971 0.99264 0.48194 0.0018822 0.42494 2.292 2.2914 16.0207 144.896 0.00016154 -85.6519 0.81994
9.924 0.98817 5.4526e-005 3.8184 0.011893 0.00012866 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7012 0.64376 0.19583 0.021798 22.3075 0.13467 0.00017801 0.75551 0.0099315 0.010961 0.0013863 0.98694 0.9917 2.9891e-006 1.1956e-005 0.16891 0.93525 0.91726 0.0013971 0.99267 0.48212 0.0018822 0.42496 2.2925 2.2919 16.0206 144.896 0.00016145 -85.652 0.82094
9.925 0.98817 5.4526e-005 3.8184 0.011893 0.00012867 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7013 0.6438 0.19584 0.021799 22.311 0.13467 0.00017802 0.7555 0.0099318 0.010961 0.0013862 0.98694 0.99171 2.9891e-006 1.1956e-005 0.16891 0.9354 0.91732 0.0013971 0.9927 0.4823 0.0018822 0.42497 2.2929 2.2923 16.0206 144.8961 0.00016136 -85.6521 0.82194
9.926 0.98817 5.4526e-005 3.8184 0.011893 0.00012868 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7014 0.64385 0.19586 0.0218 22.3146 0.13468 0.00017803 0.7555 0.0099321 0.010961 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16891 0.93555 0.91738 0.0013971 0.99273 0.48248 0.0018822 0.42499 2.2934 2.2928 16.0206 144.8961 0.00016127 -85.6522 0.82294
9.927 0.98817 5.4526e-005 3.8184 0.011893 0.00012869 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7015 0.64389 0.19587 0.021801 22.3182 0.13469 0.00017804 0.75549 0.0099324 0.010962 0.0013862 0.98694 0.99171 2.989e-006 1.1956e-005 0.16891 0.9357 0.91744 0.001397 0.99276 0.48266 0.0018822 0.425 2.2938 2.2932 16.0205 144.8961 0.00016118 -85.6522 0.82394
9.928 0.98817 5.4526e-005 3.8184 0.011893 0.00012871 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7015 0.64394 0.19588 0.021802 22.3217 0.13469 0.00017805 0.75549 0.0099327 0.010962 0.0013862 0.98695 0.99171 2.989e-006 1.1956e-005 0.16892 0.93585 0.9175 0.001397 0.99278 0.48284 0.0018822 0.42501 2.2943 2.2937 16.0205 144.8961 0.00016109 -85.6523 0.82494
9.929 0.98817 5.4526e-005 3.8184 0.011893 0.00012872 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7016 0.64398 0.19589 0.021803 22.3253 0.1347 0.00017806 0.75548 0.009933 0.010962 0.0013862 0.98695 0.99171 2.9889e-006 1.1956e-005 0.16892 0.936 0.91756 0.001397 0.99281 0.48302 0.0018821 0.42503 2.2947 2.2942 16.0205 144.8961 0.000161 -85.6524 0.82594
9.93 0.98817 5.4526e-005 3.8184 0.011893 0.00012873 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7017 0.64402 0.19591 0.021804 22.3289 0.1347 0.00017806 0.75548 0.0099333 0.010962 0.0013861 0.98695 0.99171 2.9889e-006 1.1955e-005 0.16892 0.93615 0.91762 0.001397 0.99284 0.4832 0.0018821 0.42504 2.2952 2.2946 16.0205 144.8962 0.00016091 -85.6525 0.82694
9.931 0.98817 5.4525e-005 3.8184 0.011893 0.00012875 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7018 0.64407 0.19592 0.021805 22.3324 0.13471 0.00017807 0.75547 0.0099336 0.010963 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16892 0.9363 0.91767 0.001397 0.99287 0.48338 0.0018821 0.42506 2.2956 2.2951 16.0204 144.8962 0.00016083 -85.6526 0.82794
9.932 0.98817 5.4525e-005 3.8184 0.011893 0.00012876 0.0011822 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7019 0.64411 0.19593 0.021806 22.336 0.13471 0.00017808 0.75547 0.0099339 0.010963 0.0013861 0.98695 0.99171 2.9888e-006 1.1955e-005 0.16892 0.93645 0.91773 0.001397 0.9929 0.48356 0.0018821 0.42507 2.2961 2.2955 16.0204 144.8962 0.00016074 -85.6526 0.82894
9.933 0.98817 5.4525e-005 3.8184 0.011893 0.00012877 0.0011823 0.23335 0.00065931 0.23401 0.21593 0 0.032276 0.0389 0 1.7019 0.64415 0.19594 0.021807 22.3396 0.13472 0.00017809 0.75546 0.0099342 0.010963 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16893 0.93659 0.91779 0.001397 0.99293 0.48374 0.0018821 0.42509 2.2965 2.296 16.0204 144.8962 0.00016065 -85.6527 0.82994
9.934 0.98817 5.4525e-005 3.8184 0.011893 0.00012878 0.0011823 0.23335 0.00065931 0.23401 0.21593 0 0.032277 0.0389 0 1.702 0.6442 0.19596 0.021808 22.3431 0.13472 0.0001781 0.75545 0.0099344 0.010964 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16893 0.93674 0.91785 0.001397 0.99295 0.48392 0.0018821 0.4251 2.297 2.2964 16.0203 144.8962 0.00016056 -85.6528 0.83094
9.935 0.98817 5.4525e-005 3.8184 0.011893 0.0001288 0.0011823 0.23335 0.00065931 0.23401 0.21593 0 0.032277 0.0389 0 1.7021 0.64424 0.19597 0.021808 22.3467 0.13473 0.00017811 0.75545 0.0099347 0.010964 0.0013861 0.98695 0.99171 2.9887e-006 1.1955e-005 0.16893 0.93689 0.9179 0.001397 0.99298 0.4841 0.0018821 0.42511 2.2974 2.2969 16.0203 144.8963 0.00016047 -85.6529 0.83194
9.936 0.98817 5.4525e-005 3.8184 0.011893 0.00012881 0.0011823 0.23335 0.00065931 0.23401 0.21593 0 0.032277 0.0389 0 1.7022 0.64428 0.19598 0.021809 22.3503 0.13473 0.00017812 0.75544 0.009935 0.010964 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16893 0.93703 0.91796 0.001397 0.99301 0.48428 0.0018821 0.42513 2.2979 2.2973 16.0203 144.8963 0.00016039 -85.6529 0.83294
9.937 0.98817 5.4525e-005 3.8184 0.011893 0.00012882 0.0011823 0.23335 0.00065931 0.23401 0.21593 0 0.032277 0.0389 0 1.7023 0.64433 0.19599 0.02181 22.3538 0.13474 0.00017812 0.75544 0.0099353 0.010965 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16894 0.93718 0.91802 0.001397 0.99303 0.48446 0.001882 0.42514 2.2983 2.2978 16.0202 144.8963 0.0001603 -85.653 0.83394
9.938 0.98817 5.4525e-005 3.8184 0.011893 0.00012884 0.0011823 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.7023 0.64437 0.196 0.021811 22.3574 0.13475 0.00017813 0.75543 0.0099356 0.010965 0.001386 0.98695 0.99171 2.9886e-006 1.1954e-005 0.16894 0.93732 0.91807 0.001397 0.99306 0.48464 0.001882 0.42516 2.2988 2.2982 16.0202 144.8963 0.00016022 -85.6531 0.83494
9.939 0.98817 5.4525e-005 3.8184 0.011893 0.00012885 0.0011823 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.7024 0.64441 0.19602 0.021812 22.361 0.13475 0.00017814 0.75543 0.0099359 0.010965 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16894 0.93747 0.91813 0.0013969 0.99309 0.48482 0.001882 0.42517 2.2992 2.2987 16.0202 144.8964 0.00016013 -85.6532 0.83594
9.94 0.98817 5.4525e-005 3.8184 0.011893 0.00012886 0.0011823 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.7025 0.64446 0.19603 0.021813 22.3645 0.13476 0.00017815 0.75542 0.0099362 0.010966 0.001386 0.98695 0.99171 2.9885e-006 1.1954e-005 0.16894 0.93761 0.91818 0.0013969 0.99312 0.485 0.001882 0.42519 2.2997 2.2991 16.0201 144.8964 0.00016004 -85.6532 0.83694
9.941 0.98817 5.4525e-005 3.8184 0.011893 0.00012887 0.0011823 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.7026 0.6445 0.19604 0.021814 22.3681 0.13476 0.00017816 0.75542 0.0099365 0.010966 0.001386 0.98695 0.99171 2.9884e-006 1.1954e-005 0.16894 0.93775 0.91824 0.0013969 0.99314 0.48518 0.001882 0.4252 2.3001 2.2995 16.0201 144.8964 0.00015996 -85.6533 0.83794
9.942 0.98817 5.4525e-005 3.8184 0.011893 0.00012889 0.0011823 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.7027 0.64455 0.19605 0.021815 22.3717 0.13477 0.00017817 0.75541 0.0099368 0.010966 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.16895 0.9379 0.9183 0.0013969 0.99317 0.48536 0.001882 0.42522 2.3006 2.3 16.0201 144.8964 0.00015987 -85.6534 0.83894
9.943 0.98817 5.4524e-005 3.8184 0.011893 0.0001289 0.0011823 0.23335 0.00065931 0.234 0.21593 0 0.032277 0.0389 0 1.7027 0.64459 0.19607 0.021816 22.3753 0.13477 0.00017817 0.75541 0.0099371 0.010966 0.0013859 0.98695 0.99171 2.9884e-006 1.1953e-005 0.16895 0.93804 0.91835 0.0013969 0.99319 0.48554 0.001882 0.42523 2.301 2.3004 16.02 144.8964 0.00015979 -85.6534 0.83994
9.944 0.98817 5.4524e-005 3.8184 0.011893 0.00012891 0.0011823 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7028 0.64463 0.19608 0.021817 22.3788 0.13478 0.00017818 0.7554 0.0099374 0.010967 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16895 0.93818 0.91841 0.0013969 0.99322 0.48572 0.001882 0.42524 2.3014 2.3009 16.02 144.8965 0.0001597 -85.6535 0.84094
9.945 0.98817 5.4524e-005 3.8184 0.011893 0.00012892 0.0011823 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7029 0.64468 0.19609 0.021818 22.3824 0.13478 0.00017819 0.7554 0.0099377 0.010967 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16895 0.93832 0.91846 0.0013969 0.99325 0.48589 0.0018819 0.42526 2.3019 2.3013 16.02 144.8965 0.00015962 -85.6536 0.84194
9.946 0.98817 5.4524e-005 3.8184 0.011893 0.00012894 0.0011823 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.703 0.64472 0.1961 0.021819 22.386 0.13479 0.0001782 0.75539 0.009938 0.010967 0.0013859 0.98695 0.99171 2.9883e-006 1.1953e-005 0.16896 0.93847 0.91852 0.0013969 0.99327 0.48607 0.0018819 0.42527 2.3023 2.3018 16.02 144.8965 0.00015954 -85.6537 0.84294
9.947 0.98817 5.4524e-005 3.8184 0.011893 0.00012895 0.0011823 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7031 0.64476 0.19612 0.021819 22.3896 0.13479 0.00017821 0.75538 0.0099383 0.010968 0.0013859 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16896 0.93861 0.91857 0.0013969 0.9933 0.48625 0.0018819 0.42529 2.3028 2.3022 16.0199 144.8965 0.00015945 -85.6537 0.84394
9.948 0.98817 5.4524e-005 3.8184 0.011893 0.00012896 0.0011823 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7031 0.64481 0.19613 0.02182 22.3931 0.1348 0.00017822 0.75538 0.0099386 0.010968 0.0013858 0.98695 0.99171 2.9882e-006 1.1953e-005 0.16896 0.93875 0.91862 0.0013969 0.99332 0.48643 0.0018819 0.4253 2.3032 2.3026 16.0199 144.8965 0.00015937 -85.6538 0.84494
9.949 0.98817 5.4524e-005 3.8184 0.011893 0.00012898 0.0011823 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7032 0.64485 0.19614 0.021821 22.3967 0.1348 0.00017822 0.75537 0.0099389 0.010968 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16896 0.93889 0.91868 0.0013968 0.99335 0.48661 0.0018819 0.42532 2.3036 2.3031 16.0199 144.8966 0.00015929 -85.6539 0.84594
9.95 0.98817 5.4524e-005 3.8184 0.011893 0.00012899 0.0011824 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7033 0.64489 0.19615 0.021822 22.4003 0.13481 0.00017823 0.75537 0.0099392 0.010969 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16896 0.93903 0.91873 0.0013968 0.99337 0.48679 0.0018819 0.42533 2.3041 2.3035 16.0198 144.8966 0.0001592 -85.6539 0.84694
9.951 0.98817 5.4524e-005 3.8184 0.011893 0.000129 0.0011824 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7034 0.64494 0.19617 0.021823 22.4038 0.13482 0.00017824 0.75536 0.0099394 0.010969 0.0013858 0.98695 0.99171 2.9881e-006 1.1952e-005 0.16897 0.93917 0.91879 0.0013968 0.9934 0.48697 0.0018819 0.42534 2.3045 2.3039 16.0198 144.8966 0.00015912 -85.654 0.84794
9.952 0.98817 5.4524e-005 3.8184 0.011893 0.00012901 0.0011824 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7035 0.64498 0.19618 0.021824 22.4074 0.13482 0.00017825 0.75536 0.0099397 0.010969 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16897 0.9393 0.91884 0.0013968 0.99342 0.48715 0.0018819 0.42536 2.3049 2.3044 16.0198 144.8966 0.00015904 -85.6541 0.84894
9.953 0.98817 5.4524e-005 3.8184 0.011893 0.00012903 0.0011824 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7035 0.64502 0.19619 0.021825 22.411 0.13483 0.00017826 0.75535 0.00994 0.01097 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16897 0.93944 0.91889 0.0013968 0.99345 0.48733 0.0018819 0.42537 2.3054 2.3048 16.0197 144.8966 0.00015896 -85.6541 0.84994
9.954 0.98817 5.4524e-005 3.8184 0.011893 0.00012904 0.0011824 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7036 0.64507 0.1962 0.021826 22.4146 0.13483 0.00017827 0.75535 0.0099403 0.01097 0.0013858 0.98695 0.99171 2.988e-006 1.1952e-005 0.16897 0.93958 0.91895 0.0013968 0.99347 0.4875 0.0018819 0.42539 2.3058 2.3052 16.0197 144.8967 0.00015888 -85.6542 0.85094
9.955 0.98817 5.4523e-005 3.8184 0.011893 0.00012905 0.0011824 0.23335 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7037 0.64511 0.19621 0.021827 22.4181 0.13484 0.00017828 0.75534 0.0099406 0.01097 0.0013857 0.98695 0.99171 2.9879e-006 1.1952e-005 0.16898 0.93972 0.919 0.0013968 0.99349 0.48768 0.0018818 0.4254 2.3062 2.3057 16.0197 144.8967 0.0001588 -85.6543 0.85194
9.956 0.98817 5.4523e-005 3.8184 0.011893 0.00012906 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7038 0.64515 0.19623 0.021828 22.4217 0.13484 0.00017828 0.75534 0.0099409 0.01097 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.16898 0.93985 0.91905 0.0013968 0.99352 0.48786 0.0018818 0.42542 2.3067 2.3061 16.0196 144.8967 0.00015872 -85.6543 0.85294
9.957 0.98817 5.4523e-005 3.8184 0.011893 0.00012908 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7039 0.6452 0.19624 0.021829 22.4253 0.13485 0.00017829 0.75533 0.0099412 0.010971 0.0013857 0.98695 0.99171 2.9879e-006 1.1951e-005 0.16898 0.93999 0.91911 0.0013968 0.99354 0.48804 0.0018818 0.42543 2.3071 2.3065 16.0196 144.8967 0.00015863 -85.6544 0.85394
9.958 0.98817 5.4523e-005 3.8184 0.011893 0.00012909 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7039 0.64524 0.19625 0.02183 22.4289 0.13485 0.0001783 0.75533 0.0099415 0.010971 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16898 0.94013 0.91916 0.0013968 0.99357 0.48822 0.0018818 0.42544 2.3075 2.307 16.0196 144.8967 0.00015855 -85.6544 0.85494
9.959 0.98817 5.4523e-005 3.8184 0.011892 0.0001291 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.704 0.64529 0.19626 0.02183 22.4324 0.13486 0.00017831 0.75532 0.0099418 0.010971 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16898 0.94026 0.91921 0.0013967 0.99359 0.4884 0.0018818 0.42546 2.308 2.3074 16.0195 144.8968 0.00015847 -85.6545 0.85594
9.96 0.98817 5.4523e-005 3.8184 0.011892 0.00012912 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7041 0.64533 0.19628 0.021831 22.436 0.13486 0.00017832 0.75531 0.0099421 0.010972 0.0013857 0.98695 0.99171 2.9878e-006 1.1951e-005 0.16899 0.9404 0.91926 0.0013967 0.99361 0.48858 0.0018818 0.42547 2.3084 2.3078 16.0195 144.8968 0.00015839 -85.6546 0.85694
9.961 0.98817 5.4523e-005 3.8184 0.011892 0.00012913 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7042 0.64537 0.19629 0.021832 22.4396 0.13487 0.00017833 0.75531 0.0099424 0.010972 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16899 0.94053 0.91931 0.0013967 0.99364 0.48875 0.0018818 0.42549 2.3088 2.3083 16.0195 144.8968 0.00015832 -85.6546 0.85794
9.962 0.98817 5.4523e-005 3.8184 0.011892 0.00012914 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7043 0.64542 0.1963 0.021833 22.4432 0.13487 0.00017833 0.7553 0.0099427 0.010972 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16899 0.94067 0.91937 0.0013967 0.99366 0.48893 0.0018818 0.4255 2.3092 2.3087 16.0194 144.8968 0.00015824 -85.6547 0.85894
9.963 0.98817 5.4523e-005 3.8184 0.011892 0.00012915 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7043 0.64546 0.19631 0.021834 22.4468 0.13488 0.00017834 0.7553 0.009943 0.010973 0.0013856 0.98695 0.99171 2.9877e-006 1.1951e-005 0.16899 0.9408 0.91942 0.0013967 0.99368 0.48911 0.0018818 0.42551 2.3097 2.3091 16.0194 144.8968 0.00015816 -85.6548 0.85994
9.964 0.98817 5.4523e-005 3.8184 0.011892 0.00012917 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7044 0.6455 0.19633 0.021835 22.4503 0.13489 0.00017835 0.75529 0.0099433 0.010973 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.169 0.94093 0.91947 0.0013967 0.9937 0.48929 0.0018818 0.42553 2.3101 2.3095 16.0194 144.8969 0.00015808 -85.6548 0.86094
9.965 0.98817 5.4523e-005 3.8184 0.011892 0.00012918 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7045 0.64555 0.19634 0.021836 22.4539 0.13489 0.00017836 0.75529 0.0099436 0.010973 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.169 0.94107 0.91952 0.0013967 0.99373 0.48947 0.0018817 0.42554 2.3105 2.31 16.0193 144.8969 0.000158 -85.6549 0.86194
9.966 0.98817 5.4522e-005 3.8184 0.011892 0.00012919 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7046 0.64559 0.19635 0.021837 22.4575 0.1349 0.00017837 0.75528 0.0099438 0.010974 0.0013856 0.98695 0.99171 2.9876e-006 1.195e-005 0.169 0.9412 0.91957 0.0013967 0.99375 0.48964 0.0018817 0.42556 2.3109 2.3104 16.0193 144.8969 0.00015792 -85.6549 0.86294
9.967 0.98817 5.4522e-005 3.8184 0.011892 0.0001292 0.0011824 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7047 0.64563 0.19636 0.021838 22.4611 0.1349 0.00017838 0.75528 0.0099441 0.010974 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.169 0.94133 0.91962 0.0013967 0.99377 0.48982 0.0018817 0.42557 2.3113 2.3108 16.0193 144.8969 0.00015784 -85.655 0.86394
9.968 0.98817 5.4522e-005 3.8184 0.011892 0.00012922 0.0011825 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7047 0.64568 0.19637 0.021839 22.4646 0.13491 0.00017838 0.75527 0.0099444 0.010974 0.0013856 0.98695 0.99171 2.9875e-006 1.195e-005 0.169 0.94146 0.91967 0.0013967 0.99379 0.49 0.0018817 0.42559 2.3118 2.3112 16.0193 144.897 0.00015777 -85.655 0.86494
9.969 0.98817 5.4522e-005 3.8184 0.011892 0.00012923 0.0011825 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7048 0.64572 0.19639 0.02184 22.4682 0.13491 0.00017839 0.75527 0.0099447 0.010974 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.16901 0.9416 0.91972 0.0013967 0.99382 0.49018 0.0018817 0.4256 2.3122 2.3117 16.0192 144.897 0.00015769 -85.6551 0.86594
9.97 0.98817 5.4522e-005 3.8184 0.011892 0.00012924 0.0011825 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.7049 0.64576 0.1964 0.021841 22.4718 0.13492 0.0001784 0.75526 0.009945 0.010975 0.0013855 0.98695 0.99171 2.9875e-006 1.195e-005 0.16901 0.94173 0.91977 0.0013967 0.99384 0.49035 0.0018817 0.42561 2.3126 2.3121 16.0192 144.897 0.00015761 -85.6552 0.86694
9.971 0.98817 5.4522e-005 3.8184 0.011892 0.00012926 0.0011825 0.23334 0.00065931 0.234 0.21592 0 0.032277 0.0389 0 1.705 0.64581 0.19641 0.021841 22.4754 0.13492 0.00017841 0.75526 0.0099453 0.010975 0.0013855 0.98695 0.99171 2.9874e-006 1.195e-005 0.16901 0.94186 0.91982 0.0013967 0.99386 0.49053 0.0018817 0.42563 2.313 2.3125 16.0192 144.897 0.00015754 -85.6552 0.86794
9.972 0.98817 5.4522e-005 3.8184 0.011892 0.00012927 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7051 0.64585 0.19642 0.021842 22.479 0.13493 0.00017842 0.75525 0.0099456 0.010975 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.16901 0.94199 0.91987 0.0013967 0.99388 0.49071 0.0018817 0.42564 2.3134 2.3129 16.0191 144.897 0.00015746 -85.6553 0.86894
9.973 0.98817 5.4522e-005 3.8184 0.011892 0.00012928 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7051 0.64589 0.19644 0.021843 22.4825 0.13493 0.00017843 0.75524 0.0099459 0.010976 0.0013855 0.98695 0.99171 2.9874e-006 1.1949e-005 0.16902 0.94212 0.91992 0.0013967 0.9939 0.49089 0.0018817 0.42566 2.3139 2.3133 16.0191 144.8971 0.00015738 -85.6553 0.86994
9.974 0.98817 5.4522e-005 3.8184 0.011892 0.00012929 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7052 0.64594 0.19645 0.021844 22.4861 0.13494 0.00017843 0.75524 0.0099462 0.010976 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16902 0.94225 0.91997 0.0013967 0.99392 0.49106 0.0018817 0.42567 2.3143 2.3137 16.0191 144.8971 0.00015731 -85.6554 0.87094
9.975 0.98817 5.4522e-005 3.8184 0.011892 0.00012931 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7053 0.64598 0.19646 0.021845 22.4897 0.13494 0.00017844 0.75523 0.0099465 0.010976 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16902 0.94238 0.92002 0.0013967 0.99394 0.49124 0.0018817 0.42568 2.3147 2.3142 16.019 144.8971 0.00015723 -85.6554 0.87194
9.976 0.98817 5.4522e-005 3.8184 0.011892 0.00012932 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7054 0.64602 0.19647 0.021846 22.4933 0.13495 0.00017845 0.75523 0.0099468 0.010977 0.0013855 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16902 0.94251 0.92007 0.0013966 0.99397 0.49142 0.0018816 0.4257 2.3151 2.3146 16.019 144.8971 0.00015716 -85.6555 0.87294
9.977 0.98817 5.4522e-005 3.8184 0.011892 0.00012933 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7055 0.64607 0.19649 0.021847 22.4969 0.13496 0.00017846 0.75522 0.0099471 0.010977 0.0013854 0.98695 0.99171 2.9873e-006 1.1949e-005 0.16902 0.94263 0.92012 0.0013966 0.99399 0.4916 0.0018816 0.42571 2.3155 2.315 16.019 144.8971 0.00015708 -85.6555 0.87394
9.978 0.98817 5.4521e-005 3.8184 0.011892 0.00012934 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7055 0.64611 0.1965 0.021848 22.5005 0.13496 0.00017847 0.75522 0.0099474 0.010977 0.0013854 0.98695 0.99171 2.9872e-006 1.1949e-005 0.16903 0.94276 0.92017 0.0013966 0.99401 0.49177 0.0018816 0.42573 2.3159 2.3154 16.0189 144.8972 0.00015701 -85.6556 0.87494
9.979 0.98817 5.4521e-005 3.8184 0.011892 0.00012936 0.0011825 0.23334 0.00065931 0.23399 0.21592 0 0.032277 0.0389 0 1.7056 0.64616 0.19651 0.021849 22.504 0.13497 0.00017848 0.75521 0.0099477 0.010978 0.0013854 0.98696 0.99171 2.9872e-006 1.1949e-005 0.16903 0.94289 0.92022 0.0013966 0.99403 0.49195 0.0018816 0.42574 2.3163 2.3158 16.0189 144.8972 0.00015693 -85.6556 0.87594
9.98 0.98817 5.4521e-005 3.8184 0.011892 0.00012937 0.0011825 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7057 0.6462 0.19652 0.02185 22.5076 0.13497 0.00017848 0.75521 0.009948 0.010978 0.0013854 0.98696 0.99171 2.9872e-006 1.1949e-005 0.16903 0.94302 0.92027 0.0013966 0.99405 0.49213 0.0018816 0.42576 2.3168 2.3162 16.0189 144.8972 0.00015686 -85.6557 0.87694
9.981 0.98817 5.4521e-005 3.8184 0.011892 0.00012938 0.0011825 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7058 0.64624 0.19653 0.021851 22.5112 0.13498 0.00017849 0.7552 0.0099482 0.010978 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16903 0.94314 0.92032 0.0013966 0.99407 0.49231 0.0018816 0.42577 2.3172 2.3166 16.0188 144.8972 0.00015678 -85.6557 0.87794
9.982 0.98817 5.4521e-005 3.8184 0.011892 0.0001294 0.0011825 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7059 0.64629 0.19655 0.021852 22.5148 0.13498 0.0001785 0.7552 0.0099485 0.010978 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16904 0.94327 0.92036 0.0013966 0.99409 0.49248 0.0018816 0.42578 2.3176 2.3171 16.0188 144.8972 0.00015671 -85.6558 0.87894
9.983 0.98817 5.4521e-005 3.8184 0.011892 0.00012941 0.0011825 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7059 0.64633 0.19656 0.021852 22.5184 0.13499 0.00017851 0.75519 0.0099488 0.010979 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16904 0.94339 0.92041 0.0013966 0.99411 0.49266 0.0018816 0.4258 2.318 2.3175 16.0188 144.8973 0.00015664 -85.6559 0.87994
9.984 0.98817 5.4521e-005 3.8184 0.011892 0.00012942 0.0011825 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.706 0.64637 0.19657 0.021853 22.522 0.13499 0.00017852 0.75519 0.0099491 0.010979 0.0013854 0.98696 0.99171 2.9871e-006 1.1948e-005 0.16904 0.94352 0.92046 0.0013966 0.99413 0.49284 0.0018816 0.42581 2.3184 2.3179 16.0187 144.8973 0.00015656 -85.6559 0.88094
9.985 0.98817 5.4521e-005 3.8184 0.011892 0.00012943 0.0011826 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7061 0.64642 0.19658 0.021854 22.5255 0.135 0.00017853 0.75518 0.0099494 0.010979 0.0013854 0.98696 0.99171 2.987e-006 1.1948e-005 0.16904 0.94365 0.92051 0.0013966 0.99415 0.49301 0.0018816 0.42583 2.3188 2.3183 16.0187 144.8973 0.00015649 -85.656 0.88194
9.986 0.98817 5.4521e-005 3.8184 0.011892 0.00012945 0.0011826 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7062 0.64646 0.1966 0.021855 22.5291 0.135 0.00017854 0.75517 0.0099497 0.01098 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16904 0.94377 0.92055 0.0013966 0.99417 0.49319 0.0018816 0.42584 2.3192 2.3187 16.0187 144.8973 0.00015642 -85.656 0.88294
9.987 0.98817 5.4521e-005 3.8184 0.011892 0.00012946 0.0011826 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7063 0.6465 0.19661 0.021856 22.5327 0.13501 0.00017854 0.75517 0.00995 0.01098 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16905 0.94389 0.9206 0.0013966 0.99419 0.49337 0.0018816 0.42585 2.3196 2.3191 16.0186 144.8973 0.00015634 -85.656 0.88394
9.988 0.98817 5.4521e-005 3.8184 0.011892 0.00012947 0.0011826 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7063 0.64655 0.19662 0.021857 22.5363 0.13501 0.00017855 0.75516 0.0099503 0.01098 0.0013853 0.98696 0.99171 2.987e-006 1.1948e-005 0.16905 0.94402 0.92065 0.0013966 0.99421 0.49354 0.0018815 0.42587 2.32 2.3195 16.0186 144.8974 0.00015627 -85.6561 0.88494
9.989 0.98817 5.452e-005 3.8184 0.011892 0.00012948 0.0011826 0.23334 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7064 0.64659 0.19663 0.021858 22.5399 0.13502 0.00017856 0.75516 0.0099506 0.010981 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16905 0.94414 0.9207 0.0013966 0.99423 0.49372 0.0018815 0.42588 2.3204 2.3199 16.0186 144.8974 0.0001562 -85.6561 0.88594
9.99 0.98817 5.452e-005 3.8184 0.011892 0.0001295 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7065 0.64663 0.19665 0.021859 22.5435 0.13503 0.00017857 0.75515 0.0099509 0.010981 0.0013853 0.98696 0.99171 2.9869e-006 1.1948e-005 0.16905 0.94426 0.92074 0.0013965 0.99425 0.4939 0.0018815 0.4259 2.3208 2.3203 16.0185 144.8974 0.00015613 -85.6562 0.88694
9.991 0.98817 5.452e-005 3.8184 0.011892 0.00012951 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7066 0.64668 0.19666 0.02186 22.5471 0.13503 0.00017858 0.75515 0.0099512 0.010981 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16906 0.94439 0.92079 0.0013965 0.99426 0.49407 0.0018815 0.42591 2.3212 2.3207 16.0185 144.8974 0.00015606 -85.6562 0.88794
9.992 0.98817 5.452e-005 3.8184 0.011892 0.00012952 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7067 0.64672 0.19667 0.021861 22.5506 0.13504 0.00017859 0.75514 0.0099515 0.010982 0.0013853 0.98696 0.99171 2.9869e-006 1.1947e-005 0.16906 0.94451 0.92084 0.0013965 0.99428 0.49425 0.0018815 0.42592 2.3216 2.3211 16.0185 144.8974 0.00015598 -85.6563 0.88894
9.993 0.98817 5.452e-005 3.8184 0.011892 0.00012954 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7067 0.64676 0.19668 0.021862 22.5542 0.13504 0.00017859 0.75514 0.0099518 0.010982 0.0013853 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16906 0.94463 0.92088 0.0013965 0.9943 0.49442 0.0018815 0.42594 2.322 2.3215 16.0184 144.8975 0.00015591 -85.6563 0.88994
9.994 0.98817 5.452e-005 3.8184 0.011892 0.00012955 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7068 0.64681 0.19669 0.021862 22.5578 0.13505 0.0001786 0.75513 0.009952 0.010982 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16906 0.94475 0.92093 0.0013965 0.99432 0.4946 0.0018815 0.42595 2.3224 2.3219 16.0184 144.8975 0.00015584 -85.6564 0.89094
9.995 0.98817 5.452e-005 3.8184 0.011892 0.00012956 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7069 0.64685 0.19671 0.021863 22.5614 0.13505 0.00017861 0.75513 0.0099523 0.010982 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16906 0.94487 0.92098 0.0013965 0.99434 0.49478 0.0018815 0.42597 2.3228 2.3223 16.0184 144.8975 0.00015577 -85.6564 0.89194
9.996 0.98817 5.452e-005 3.8184 0.011892 0.00012957 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.707 0.64689 0.19672 0.021864 22.565 0.13506 0.00017862 0.75512 0.0099526 0.010983 0.0013852 0.98696 0.99171 2.9868e-006 1.1947e-005 0.16907 0.945 0.92102 0.0013965 0.99436 0.49495 0.0018815 0.42598 2.3232 2.3227 16.0183 144.8975 0.0001557 -85.6565 0.89294
9.997 0.98817 5.452e-005 3.8184 0.011892 0.00012959 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7071 0.64694 0.19673 0.021865 22.5686 0.13506 0.00017863 0.75512 0.0099529 0.010983 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16907 0.94512 0.92107 0.0013965 0.99438 0.49513 0.0018815 0.42599 2.3236 2.3231 16.0183 144.8975 0.00015563 -85.6565 0.89394
9.998 0.98817 5.452e-005 3.8184 0.011892 0.0001296 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7071 0.64698 0.19674 0.021866 22.5722 0.13507 0.00017864 0.75511 0.0099532 0.010983 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16907 0.94524 0.92111 0.0013965 0.99439 0.4953 0.0018815 0.42601 2.324 2.3235 16.0183 144.8976 0.00015556 -85.6566 0.89494
9.999 0.98817 5.452e-005 3.8184 0.011892 0.00012961 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7072 0.64703 0.19676 0.021867 22.5758 0.13507 0.00017864 0.75511 0.0099535 0.010984 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16907 0.94536 0.92116 0.0013965 0.99441 0.49548 0.0018815 0.42602 2.3244 2.3239 16.0182 144.8976 0.00015549 -85.6566 0.89594
10 0.98817 5.452e-005 3.8184 0.011892 0.00012962 0.0011826 0.23333 0.00065931 0.23399 0.21591 0 0.032277 0.0389 0 1.7073 0.64707 0.19677 0.021868 22.5793 0.13508 0.00017865 0.7551 0.0099538 0.010984 0.0013852 0.98696 0.99171 2.9867e-006 1.1947e-005 0.16908 0.94547 0.9212 0.0013965 0.99443 0.49566 0.0018815 0.42604 2.3248 2.3243 16.0182 144.8976 0.00015542 -85.6566 0.89694
